VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO PAD_DVDD
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN PAD_DVDD 0 0 ;
  SIZE 100 BY 123 ;
  SYMMETRY X Y R90 ;
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER TOP_M ;
        RECT 52.5 120 96 123 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 4 120 47.5 123 ;
    END
    PORT
      LAYER M3 ;
        RECT 0 34 100 64 ;
      LAYER M4 ;
        RECT 0 34 100 64 ;
      LAYER TOP_V ;
        RECT 82.87 33.16 83.23 33.52 ;
        RECT 82.87 31.59 83.23 31.95 ;
        RECT 82.87 23.49 83.23 23.85 ;
        RECT 82.87 21.92 83.23 22.28 ;
        RECT 82.87 20.35 83.23 20.71 ;
        RECT 82.87 12.25 83.23 12.61 ;
        RECT 82.87 10.68 83.23 11.04 ;
        RECT 82.87 9.11 83.23 9.47 ;
        RECT 83.68 90.93 84.04 91.29 ;
        RECT 83.68 89.36 84.04 89.72 ;
        RECT 83.68 87.79 84.04 88.15 ;
        RECT 83.68 79.69 84.04 80.05 ;
        RECT 83.68 78.12 84.04 78.48 ;
        RECT 83.68 76.55 84.04 76.91 ;
        RECT 83.68 68.45 84.04 68.81 ;
        RECT 83.68 66.88 84.04 67.24 ;
        RECT 83.68 65.31 84.04 65.67 ;
        RECT 83.68 57.21 84.04 57.57 ;
        RECT 83.68 55.64 84.04 56 ;
        RECT 83.68 54.07 84.04 54.43 ;
        RECT 83.68 45.97 84.04 46.33 ;
        RECT 83.68 44.4 84.04 44.76 ;
        RECT 83.68 42.83 84.04 43.19 ;
        RECT 83.68 34.73 84.04 35.09 ;
        RECT 83.68 33.16 84.04 33.52 ;
        RECT 83.68 31.59 84.04 31.95 ;
        RECT 83.68 23.49 84.04 23.85 ;
        RECT 83.68 21.92 84.04 22.28 ;
        RECT 83.68 20.35 84.04 20.71 ;
        RECT 83.68 12.25 84.04 12.61 ;
        RECT 83.68 10.68 84.04 11.04 ;
        RECT 83.68 9.11 84.04 9.47 ;
        RECT 83.74 85.3 84.1 85.66 ;
        RECT 83.74 84.49 84.1 84.85 ;
        RECT 83.74 83.68 84.1 84.04 ;
        RECT 83.74 82.87 84.1 83.23 ;
        RECT 83.74 82.06 84.1 82.42 ;
        RECT 83.74 74.06 84.1 74.42 ;
        RECT 83.74 73.25 84.1 73.61 ;
        RECT 83.74 72.44 84.1 72.8 ;
        RECT 83.74 71.63 84.1 71.99 ;
        RECT 83.74 70.82 84.1 71.18 ;
        RECT 83.74 62.82 84.1 63.18 ;
        RECT 83.74 62.01 84.1 62.37 ;
        RECT 83.74 61.2 84.1 61.56 ;
        RECT 83.74 60.39 84.1 60.75 ;
        RECT 83.74 59.58 84.1 59.94 ;
        RECT 83.74 51.58 84.1 51.94 ;
        RECT 83.74 50.77 84.1 51.13 ;
        RECT 83.74 49.96 84.1 50.32 ;
        RECT 83.74 49.15 84.1 49.51 ;
        RECT 83.74 48.34 84.1 48.7 ;
        RECT 83.74 40.34 84.1 40.7 ;
        RECT 83.74 39.53 84.1 39.89 ;
        RECT 83.74 38.72 84.1 39.08 ;
        RECT 83.74 37.91 84.1 38.27 ;
        RECT 83.74 37.1 84.1 37.46 ;
        RECT 83.74 29.1 84.1 29.46 ;
        RECT 83.74 28.29 84.1 28.65 ;
        RECT 83.74 27.48 84.1 27.84 ;
        RECT 83.74 26.67 84.1 27.03 ;
        RECT 83.74 25.86 84.1 26.22 ;
        RECT 83.74 17.86 84.1 18.22 ;
        RECT 83.74 17.05 84.1 17.41 ;
        RECT 83.74 16.24 84.1 16.6 ;
        RECT 83.74 15.43 84.1 15.79 ;
        RECT 83.74 14.62 84.1 14.98 ;
        RECT 84.49 90.93 84.85 91.29 ;
        RECT 84.49 89.36 84.85 89.72 ;
        RECT 84.49 87.79 84.85 88.15 ;
        RECT 84.49 79.69 84.85 80.05 ;
        RECT 84.49 78.12 84.85 78.48 ;
        RECT 84.49 76.55 84.85 76.91 ;
        RECT 84.49 68.45 84.85 68.81 ;
        RECT 84.49 66.88 84.85 67.24 ;
        RECT 84.49 65.31 84.85 65.67 ;
        RECT 84.49 57.21 84.85 57.57 ;
        RECT 84.49 55.64 84.85 56 ;
        RECT 84.49 54.07 84.85 54.43 ;
        RECT 84.49 45.97 84.85 46.33 ;
        RECT 84.49 44.4 84.85 44.76 ;
        RECT 84.49 42.83 84.85 43.19 ;
        RECT 84.49 34.73 84.85 35.09 ;
        RECT 84.49 33.16 84.85 33.52 ;
        RECT 84.49 31.59 84.85 31.95 ;
        RECT 84.49 23.49 84.85 23.85 ;
        RECT 84.49 21.92 84.85 22.28 ;
        RECT 84.49 20.35 84.85 20.71 ;
        RECT 84.49 12.25 84.85 12.61 ;
        RECT 84.49 10.68 84.85 11.04 ;
        RECT 84.49 9.11 84.85 9.47 ;
        RECT 85.3 90.93 85.66 91.29 ;
        RECT 85.3 89.36 85.66 89.72 ;
        RECT 85.3 87.79 85.66 88.15 ;
        RECT 85.3 79.69 85.66 80.05 ;
        RECT 85.3 78.12 85.66 78.48 ;
        RECT 85.3 76.55 85.66 76.91 ;
        RECT 85.3 68.45 85.66 68.81 ;
        RECT 85.3 66.88 85.66 67.24 ;
        RECT 85.3 65.31 85.66 65.67 ;
        RECT 85.3 57.21 85.66 57.57 ;
        RECT 85.3 55.64 85.66 56 ;
        RECT 85.3 54.07 85.66 54.43 ;
        RECT 85.3 45.97 85.66 46.33 ;
        RECT 85.3 44.4 85.66 44.76 ;
        RECT 85.3 42.83 85.66 43.19 ;
        RECT 85.3 34.73 85.66 35.09 ;
        RECT 85.3 33.16 85.66 33.52 ;
        RECT 85.3 31.59 85.66 31.95 ;
        RECT 85.3 23.49 85.66 23.85 ;
        RECT 85.3 21.92 85.66 22.28 ;
        RECT 85.3 20.35 85.66 20.71 ;
        RECT 85.3 12.25 85.66 12.61 ;
        RECT 85.3 10.68 85.66 11.04 ;
        RECT 85.3 9.11 85.66 9.47 ;
        RECT 85.31 85.3 85.67 85.66 ;
        RECT 85.31 84.49 85.67 84.85 ;
        RECT 85.31 83.68 85.67 84.04 ;
        RECT 85.31 82.87 85.67 83.23 ;
        RECT 85.31 82.06 85.67 82.42 ;
        RECT 85.31 74.06 85.67 74.42 ;
        RECT 85.31 73.25 85.67 73.61 ;
        RECT 85.31 72.44 85.67 72.8 ;
        RECT 85.31 71.63 85.67 71.99 ;
        RECT 85.31 70.82 85.67 71.18 ;
        RECT 85.31 62.82 85.67 63.18 ;
        RECT 85.31 62.01 85.67 62.37 ;
        RECT 85.31 61.2 85.67 61.56 ;
        RECT 85.31 60.39 85.67 60.75 ;
        RECT 85.31 59.58 85.67 59.94 ;
        RECT 85.31 51.58 85.67 51.94 ;
        RECT 85.31 50.77 85.67 51.13 ;
        RECT 85.31 49.96 85.67 50.32 ;
        RECT 85.31 49.15 85.67 49.51 ;
        RECT 85.31 48.34 85.67 48.7 ;
        RECT 85.31 40.34 85.67 40.7 ;
        RECT 85.31 39.53 85.67 39.89 ;
        RECT 85.31 38.72 85.67 39.08 ;
        RECT 85.31 37.91 85.67 38.27 ;
        RECT 85.31 37.1 85.67 37.46 ;
        RECT 85.31 29.1 85.67 29.46 ;
        RECT 85.31 28.29 85.67 28.65 ;
        RECT 85.31 27.48 85.67 27.84 ;
        RECT 85.31 26.67 85.67 27.03 ;
        RECT 85.31 25.86 85.67 26.22 ;
        RECT 85.31 17.86 85.67 18.22 ;
        RECT 85.31 17.05 85.67 17.41 ;
        RECT 85.31 16.24 85.67 16.6 ;
        RECT 85.31 15.43 85.67 15.79 ;
        RECT 85.31 14.62 85.67 14.98 ;
        RECT 87.73 90.92 88.09 91.28 ;
        RECT 87.73 90.11 88.09 90.47 ;
        RECT 87.73 89.3 88.09 89.66 ;
        RECT 87.73 88.49 88.09 88.85 ;
        RECT 87.73 87.68 88.09 88.04 ;
        RECT 87.73 79.68 88.09 80.04 ;
        RECT 87.73 78.87 88.09 79.23 ;
        RECT 87.73 78.06 88.09 78.42 ;
        RECT 87.73 77.25 88.09 77.61 ;
        RECT 87.73 76.44 88.09 76.8 ;
        RECT 87.73 68.44 88.09 68.8 ;
        RECT 87.73 67.63 88.09 67.99 ;
        RECT 87.73 66.82 88.09 67.18 ;
        RECT 87.73 66.01 88.09 66.37 ;
        RECT 87.73 65.2 88.09 65.56 ;
        RECT 87.73 57.2 88.09 57.56 ;
        RECT 87.73 56.39 88.09 56.75 ;
        RECT 87.73 55.58 88.09 55.94 ;
        RECT 87.73 54.77 88.09 55.13 ;
        RECT 87.73 53.96 88.09 54.32 ;
        RECT 87.73 45.96 88.09 46.32 ;
        RECT 87.73 45.15 88.09 45.51 ;
        RECT 87.73 44.34 88.09 44.7 ;
        RECT 87.73 43.53 88.09 43.89 ;
        RECT 87.73 42.72 88.09 43.08 ;
        RECT 87.73 34.72 88.09 35.08 ;
        RECT 87.73 33.91 88.09 34.27 ;
        RECT 87.73 33.1 88.09 33.46 ;
        RECT 87.73 32.29 88.09 32.65 ;
        RECT 87.73 31.48 88.09 31.84 ;
        RECT 87.73 23.48 88.09 23.84 ;
        RECT 87.73 22.67 88.09 23.03 ;
        RECT 87.73 21.86 88.09 22.22 ;
        RECT 87.73 21.05 88.09 21.41 ;
        RECT 87.73 20.24 88.09 20.6 ;
        RECT 87.73 12.24 88.09 12.6 ;
        RECT 87.73 11.43 88.09 11.79 ;
        RECT 87.73 10.62 88.09 10.98 ;
        RECT 87.73 9.81 88.09 10.17 ;
        RECT 87.73 9 88.09 9.36 ;
        RECT 87.74 85.31 88.1 85.67 ;
        RECT 87.74 83.74 88.1 84.1 ;
        RECT 87.74 82.17 88.1 82.53 ;
        RECT 87.74 74.07 88.1 74.43 ;
        RECT 87.74 72.5 88.1 72.86 ;
        RECT 87.74 70.93 88.1 71.29 ;
        RECT 87.74 62.83 88.1 63.19 ;
        RECT 87.74 61.26 88.1 61.62 ;
        RECT 87.74 59.69 88.1 60.05 ;
        RECT 87.74 51.59 88.1 51.95 ;
        RECT 87.74 50.02 88.1 50.38 ;
        RECT 87.74 48.45 88.1 48.81 ;
        RECT 87.74 40.35 88.1 40.71 ;
        RECT 87.74 38.78 88.1 39.14 ;
        RECT 87.74 37.21 88.1 37.57 ;
        RECT 87.74 29.11 88.1 29.47 ;
        RECT 87.74 27.54 88.1 27.9 ;
        RECT 87.74 25.97 88.1 26.33 ;
        RECT 87.74 17.87 88.1 18.23 ;
        RECT 87.74 16.3 88.1 16.66 ;
        RECT 87.74 14.73 88.1 15.09 ;
        RECT 88.55 85.31 88.91 85.67 ;
        RECT 88.55 83.74 88.91 84.1 ;
        RECT 88.55 82.17 88.91 82.53 ;
        RECT 88.55 74.07 88.91 74.43 ;
        RECT 88.55 72.5 88.91 72.86 ;
        RECT 88.55 70.93 88.91 71.29 ;
        RECT 88.55 62.83 88.91 63.19 ;
        RECT 88.55 61.26 88.91 61.62 ;
        RECT 88.55 59.69 88.91 60.05 ;
        RECT 88.55 51.59 88.91 51.95 ;
        RECT 88.55 50.02 88.91 50.38 ;
        RECT 88.55 48.45 88.91 48.81 ;
        RECT 88.55 40.35 88.91 40.71 ;
        RECT 88.55 38.78 88.91 39.14 ;
        RECT 88.55 37.21 88.91 37.57 ;
        RECT 88.55 29.11 88.91 29.47 ;
        RECT 88.55 27.54 88.91 27.9 ;
        RECT 88.55 25.97 88.91 26.33 ;
        RECT 88.55 17.87 88.91 18.23 ;
        RECT 88.55 16.3 88.91 16.66 ;
        RECT 88.55 14.73 88.91 15.09 ;
        RECT 89.3 90.92 89.66 91.28 ;
        RECT 89.3 90.11 89.66 90.47 ;
        RECT 89.3 89.3 89.66 89.66 ;
        RECT 89.3 88.49 89.66 88.85 ;
        RECT 89.3 87.68 89.66 88.04 ;
        RECT 89.3 79.68 89.66 80.04 ;
        RECT 89.3 78.87 89.66 79.23 ;
        RECT 89.3 78.06 89.66 78.42 ;
        RECT 89.3 77.25 89.66 77.61 ;
        RECT 89.3 76.44 89.66 76.8 ;
        RECT 89.3 68.44 89.66 68.8 ;
        RECT 89.3 67.63 89.66 67.99 ;
        RECT 89.3 66.82 89.66 67.18 ;
        RECT 89.3 66.01 89.66 66.37 ;
        RECT 89.3 65.2 89.66 65.56 ;
        RECT 89.3 57.2 89.66 57.56 ;
        RECT 89.3 56.39 89.66 56.75 ;
        RECT 89.3 55.58 89.66 55.94 ;
        RECT 89.3 54.77 89.66 55.13 ;
        RECT 89.3 53.96 89.66 54.32 ;
        RECT 89.3 45.96 89.66 46.32 ;
        RECT 89.3 45.15 89.66 45.51 ;
        RECT 89.3 44.34 89.66 44.7 ;
        RECT 89.3 43.53 89.66 43.89 ;
        RECT 89.3 42.72 89.66 43.08 ;
        RECT 89.3 34.72 89.66 35.08 ;
        RECT 89.3 33.91 89.66 34.27 ;
        RECT 89.3 33.1 89.66 33.46 ;
        RECT 89.3 32.29 89.66 32.65 ;
        RECT 89.3 31.48 89.66 31.84 ;
        RECT 89.3 23.48 89.66 23.84 ;
        RECT 89.3 22.67 89.66 23.03 ;
        RECT 89.3 21.86 89.66 22.22 ;
        RECT 89.3 21.05 89.66 21.41 ;
        RECT 89.3 20.24 89.66 20.6 ;
        RECT 89.3 12.24 89.66 12.6 ;
        RECT 89.3 11.43 89.66 11.79 ;
        RECT 89.3 10.62 89.66 10.98 ;
        RECT 89.3 9.81 89.66 10.17 ;
        RECT 89.3 9 89.66 9.36 ;
        RECT 89.36 85.31 89.72 85.67 ;
        RECT 89.36 83.74 89.72 84.1 ;
        RECT 89.36 82.17 89.72 82.53 ;
        RECT 89.36 74.07 89.72 74.43 ;
        RECT 89.36 72.5 89.72 72.86 ;
        RECT 89.36 70.93 89.72 71.29 ;
        RECT 89.36 62.83 89.72 63.19 ;
        RECT 89.36 61.26 89.72 61.62 ;
        RECT 89.36 59.69 89.72 60.05 ;
        RECT 89.36 51.59 89.72 51.95 ;
        RECT 89.36 50.02 89.72 50.38 ;
        RECT 89.36 48.45 89.72 48.81 ;
        RECT 89.36 40.35 89.72 40.71 ;
        RECT 89.36 38.78 89.72 39.14 ;
        RECT 89.36 37.21 89.72 37.57 ;
        RECT 89.36 29.11 89.72 29.47 ;
        RECT 89.36 27.54 89.72 27.9 ;
        RECT 89.36 25.97 89.72 26.33 ;
        RECT 89.36 17.87 89.72 18.23 ;
        RECT 89.36 16.3 89.72 16.66 ;
        RECT 89.36 14.73 89.72 15.09 ;
        RECT 90.17 85.31 90.53 85.67 ;
        RECT 90.17 83.74 90.53 84.1 ;
        RECT 90.17 82.17 90.53 82.53 ;
        RECT 90.17 74.07 90.53 74.43 ;
        RECT 90.17 72.5 90.53 72.86 ;
        RECT 90.17 70.93 90.53 71.29 ;
        RECT 90.17 62.83 90.53 63.19 ;
        RECT 90.17 61.26 90.53 61.62 ;
        RECT 90.17 59.69 90.53 60.05 ;
        RECT 90.17 51.59 90.53 51.95 ;
        RECT 90.17 50.02 90.53 50.38 ;
        RECT 90.17 48.45 90.53 48.81 ;
        RECT 90.17 40.35 90.53 40.71 ;
        RECT 90.17 38.78 90.53 39.14 ;
        RECT 90.17 37.21 90.53 37.57 ;
        RECT 90.17 29.11 90.53 29.47 ;
        RECT 90.17 27.54 90.53 27.9 ;
        RECT 90.17 25.97 90.53 26.33 ;
        RECT 90.17 17.87 90.53 18.23 ;
        RECT 90.17 16.3 90.53 16.66 ;
        RECT 90.17 14.73 90.53 15.09 ;
        RECT 90.87 90.92 91.23 91.28 ;
        RECT 90.87 90.11 91.23 90.47 ;
        RECT 90.87 89.3 91.23 89.66 ;
        RECT 90.87 88.49 91.23 88.85 ;
        RECT 90.87 87.68 91.23 88.04 ;
        RECT 90.87 79.68 91.23 80.04 ;
        RECT 90.87 78.87 91.23 79.23 ;
        RECT 90.87 78.06 91.23 78.42 ;
        RECT 90.87 77.25 91.23 77.61 ;
        RECT 90.87 76.44 91.23 76.8 ;
        RECT 90.87 68.44 91.23 68.8 ;
        RECT 90.87 67.63 91.23 67.99 ;
        RECT 90.87 66.82 91.23 67.18 ;
        RECT 90.87 66.01 91.23 66.37 ;
        RECT 90.87 65.2 91.23 65.56 ;
        RECT 90.87 57.2 91.23 57.56 ;
        RECT 90.87 56.39 91.23 56.75 ;
        RECT 90.87 55.58 91.23 55.94 ;
        RECT 90.87 54.77 91.23 55.13 ;
        RECT 90.87 53.96 91.23 54.32 ;
        RECT 90.87 45.96 91.23 46.32 ;
        RECT 90.87 45.15 91.23 45.51 ;
        RECT 90.87 44.34 91.23 44.7 ;
        RECT 90.87 43.53 91.23 43.89 ;
        RECT 90.87 42.72 91.23 43.08 ;
        RECT 90.87 34.72 91.23 35.08 ;
        RECT 90.87 33.91 91.23 34.27 ;
        RECT 90.87 33.1 91.23 33.46 ;
        RECT 90.87 32.29 91.23 32.65 ;
        RECT 90.87 31.48 91.23 31.84 ;
        RECT 90.87 23.48 91.23 23.84 ;
        RECT 90.87 22.67 91.23 23.03 ;
        RECT 90.87 21.86 91.23 22.22 ;
        RECT 90.87 21.05 91.23 21.41 ;
        RECT 90.87 20.24 91.23 20.6 ;
        RECT 90.87 12.24 91.23 12.6 ;
        RECT 90.87 11.43 91.23 11.79 ;
        RECT 90.87 10.62 91.23 10.98 ;
        RECT 90.87 9.81 91.23 10.17 ;
        RECT 90.87 9 91.23 9.36 ;
        RECT 90.98 85.31 91.34 85.67 ;
        RECT 90.98 83.74 91.34 84.1 ;
        RECT 90.98 82.17 91.34 82.53 ;
        RECT 90.98 74.07 91.34 74.43 ;
        RECT 90.98 72.5 91.34 72.86 ;
        RECT 90.98 70.93 91.34 71.29 ;
        RECT 90.98 62.83 91.34 63.19 ;
        RECT 90.98 61.26 91.34 61.62 ;
        RECT 90.98 59.69 91.34 60.05 ;
        RECT 90.98 51.59 91.34 51.95 ;
        RECT 90.98 50.02 91.34 50.38 ;
        RECT 90.98 48.45 91.34 48.81 ;
        RECT 90.98 40.35 91.34 40.71 ;
        RECT 90.98 38.78 91.34 39.14 ;
        RECT 90.98 37.21 91.34 37.57 ;
        RECT 90.98 29.11 91.34 29.47 ;
        RECT 90.98 27.54 91.34 27.9 ;
        RECT 90.98 25.97 91.34 26.33 ;
        RECT 90.98 17.87 91.34 18.23 ;
        RECT 90.98 16.3 91.34 16.66 ;
        RECT 90.98 14.73 91.34 15.09 ;
        RECT 57.15 11.43 57.51 11.79 ;
        RECT 57.15 10.62 57.51 10.98 ;
        RECT 57.15 9.81 57.51 10.17 ;
        RECT 57.15 9 57.51 9.36 ;
        RECT 57.26 85.31 57.62 85.67 ;
        RECT 57.26 83.74 57.62 84.1 ;
        RECT 57.26 82.17 57.62 82.53 ;
        RECT 57.26 74.07 57.62 74.43 ;
        RECT 57.26 72.5 57.62 72.86 ;
        RECT 57.26 70.93 57.62 71.29 ;
        RECT 57.26 62.83 57.62 63.19 ;
        RECT 57.26 61.26 57.62 61.62 ;
        RECT 57.26 59.69 57.62 60.05 ;
        RECT 57.26 51.59 57.62 51.95 ;
        RECT 57.26 50.02 57.62 50.38 ;
        RECT 57.26 48.45 57.62 48.81 ;
        RECT 57.26 40.35 57.62 40.71 ;
        RECT 57.26 38.78 57.62 39.14 ;
        RECT 57.26 37.21 57.62 37.57 ;
        RECT 57.26 29.11 57.62 29.47 ;
        RECT 57.26 27.54 57.62 27.9 ;
        RECT 57.26 25.97 57.62 26.33 ;
        RECT 57.26 17.87 57.62 18.23 ;
        RECT 57.26 16.3 57.62 16.66 ;
        RECT 57.26 14.73 57.62 15.09 ;
        RECT 59.58 90.93 59.94 91.29 ;
        RECT 59.58 89.36 59.94 89.72 ;
        RECT 59.58 87.79 59.94 88.15 ;
        RECT 59.58 79.69 59.94 80.05 ;
        RECT 59.58 78.12 59.94 78.48 ;
        RECT 59.58 76.55 59.94 76.91 ;
        RECT 59.58 68.45 59.94 68.81 ;
        RECT 59.58 66.88 59.94 67.24 ;
        RECT 59.58 65.31 59.94 65.67 ;
        RECT 59.58 57.21 59.94 57.57 ;
        RECT 59.58 55.64 59.94 56 ;
        RECT 59.58 54.07 59.94 54.43 ;
        RECT 59.58 45.97 59.94 46.33 ;
        RECT 59.58 44.4 59.94 44.76 ;
        RECT 59.58 42.83 59.94 43.19 ;
        RECT 59.58 34.73 59.94 35.09 ;
        RECT 59.58 33.16 59.94 33.52 ;
        RECT 59.58 31.59 59.94 31.95 ;
        RECT 59.58 23.49 59.94 23.85 ;
        RECT 59.58 21.92 59.94 22.28 ;
        RECT 59.58 20.35 59.94 20.71 ;
        RECT 59.58 12.25 59.94 12.61 ;
        RECT 59.58 10.68 59.94 11.04 ;
        RECT 59.58 9.11 59.94 9.47 ;
        RECT 59.69 85.3 60.05 85.66 ;
        RECT 59.69 84.49 60.05 84.85 ;
        RECT 59.69 83.68 60.05 84.04 ;
        RECT 59.69 82.87 60.05 83.23 ;
        RECT 59.69 82.06 60.05 82.42 ;
        RECT 59.69 74.06 60.05 74.42 ;
        RECT 59.69 73.25 60.05 73.61 ;
        RECT 59.69 72.44 60.05 72.8 ;
        RECT 59.69 71.63 60.05 71.99 ;
        RECT 59.69 70.82 60.05 71.18 ;
        RECT 59.69 62.82 60.05 63.18 ;
        RECT 59.69 62.01 60.05 62.37 ;
        RECT 59.69 61.2 60.05 61.56 ;
        RECT 59.69 60.39 60.05 60.75 ;
        RECT 59.69 59.58 60.05 59.94 ;
        RECT 59.69 51.58 60.05 51.94 ;
        RECT 59.69 50.77 60.05 51.13 ;
        RECT 59.69 49.96 60.05 50.32 ;
        RECT 59.69 49.15 60.05 49.51 ;
        RECT 59.69 48.34 60.05 48.7 ;
        RECT 59.69 40.34 60.05 40.7 ;
        RECT 59.69 39.53 60.05 39.89 ;
        RECT 59.69 38.72 60.05 39.08 ;
        RECT 59.69 37.91 60.05 38.27 ;
        RECT 59.69 37.1 60.05 37.46 ;
        RECT 59.69 29.1 60.05 29.46 ;
        RECT 59.69 28.29 60.05 28.65 ;
        RECT 59.69 27.48 60.05 27.84 ;
        RECT 59.69 26.67 60.05 27.03 ;
        RECT 59.69 25.86 60.05 26.22 ;
        RECT 59.69 17.86 60.05 18.22 ;
        RECT 59.69 17.05 60.05 17.41 ;
        RECT 59.69 16.24 60.05 16.6 ;
        RECT 59.69 15.43 60.05 15.79 ;
        RECT 59.69 14.62 60.05 14.98 ;
        RECT 60.39 90.93 60.75 91.29 ;
        RECT 60.39 89.36 60.75 89.72 ;
        RECT 60.39 87.79 60.75 88.15 ;
        RECT 60.39 79.69 60.75 80.05 ;
        RECT 60.39 78.12 60.75 78.48 ;
        RECT 60.39 76.55 60.75 76.91 ;
        RECT 60.39 68.45 60.75 68.81 ;
        RECT 60.39 66.88 60.75 67.24 ;
        RECT 60.39 65.31 60.75 65.67 ;
        RECT 60.39 57.21 60.75 57.57 ;
        RECT 60.39 55.64 60.75 56 ;
        RECT 60.39 54.07 60.75 54.43 ;
        RECT 60.39 45.97 60.75 46.33 ;
        RECT 60.39 44.4 60.75 44.76 ;
        RECT 60.39 42.83 60.75 43.19 ;
        RECT 60.39 34.73 60.75 35.09 ;
        RECT 60.39 33.16 60.75 33.52 ;
        RECT 60.39 31.59 60.75 31.95 ;
        RECT 60.39 23.49 60.75 23.85 ;
        RECT 60.39 21.92 60.75 22.28 ;
        RECT 60.39 20.35 60.75 20.71 ;
        RECT 60.39 12.25 60.75 12.61 ;
        RECT 60.39 10.68 60.75 11.04 ;
        RECT 60.39 9.11 60.75 9.47 ;
        RECT 61.2 90.93 61.56 91.29 ;
        RECT 61.2 89.36 61.56 89.72 ;
        RECT 61.2 87.79 61.56 88.15 ;
        RECT 61.2 79.69 61.56 80.05 ;
        RECT 61.2 78.12 61.56 78.48 ;
        RECT 61.2 76.55 61.56 76.91 ;
        RECT 61.2 68.45 61.56 68.81 ;
        RECT 61.2 66.88 61.56 67.24 ;
        RECT 61.2 65.31 61.56 65.67 ;
        RECT 61.2 57.21 61.56 57.57 ;
        RECT 61.2 55.64 61.56 56 ;
        RECT 61.2 54.07 61.56 54.43 ;
        RECT 61.2 45.97 61.56 46.33 ;
        RECT 61.2 44.4 61.56 44.76 ;
        RECT 61.2 42.83 61.56 43.19 ;
        RECT 61.2 34.73 61.56 35.09 ;
        RECT 61.2 33.16 61.56 33.52 ;
        RECT 61.2 31.59 61.56 31.95 ;
        RECT 61.2 23.49 61.56 23.85 ;
        RECT 61.2 21.92 61.56 22.28 ;
        RECT 61.2 20.35 61.56 20.71 ;
        RECT 61.2 12.25 61.56 12.61 ;
        RECT 61.2 10.68 61.56 11.04 ;
        RECT 61.2 9.11 61.56 9.47 ;
        RECT 61.26 85.3 61.62 85.66 ;
        RECT 61.26 84.49 61.62 84.85 ;
        RECT 61.26 83.68 61.62 84.04 ;
        RECT 61.26 82.87 61.62 83.23 ;
        RECT 61.26 82.06 61.62 82.42 ;
        RECT 61.26 74.06 61.62 74.42 ;
        RECT 61.26 73.25 61.62 73.61 ;
        RECT 61.26 72.44 61.62 72.8 ;
        RECT 61.26 71.63 61.62 71.99 ;
        RECT 61.26 70.82 61.62 71.18 ;
        RECT 61.26 62.82 61.62 63.18 ;
        RECT 61.26 62.01 61.62 62.37 ;
        RECT 61.26 61.2 61.62 61.56 ;
        RECT 61.26 60.39 61.62 60.75 ;
        RECT 61.26 59.58 61.62 59.94 ;
        RECT 61.26 51.58 61.62 51.94 ;
        RECT 61.26 50.77 61.62 51.13 ;
        RECT 61.26 49.96 61.62 50.32 ;
        RECT 61.26 49.15 61.62 49.51 ;
        RECT 61.26 48.34 61.62 48.7 ;
        RECT 61.26 40.34 61.62 40.7 ;
        RECT 61.26 39.53 61.62 39.89 ;
        RECT 61.26 38.72 61.62 39.08 ;
        RECT 61.26 37.91 61.62 38.27 ;
        RECT 61.26 37.1 61.62 37.46 ;
        RECT 61.26 29.1 61.62 29.46 ;
        RECT 61.26 28.29 61.62 28.65 ;
        RECT 61.26 27.48 61.62 27.84 ;
        RECT 61.26 26.67 61.62 27.03 ;
        RECT 61.26 25.86 61.62 26.22 ;
        RECT 61.26 17.86 61.62 18.22 ;
        RECT 61.26 17.05 61.62 17.41 ;
        RECT 61.26 16.24 61.62 16.6 ;
        RECT 61.26 15.43 61.62 15.79 ;
        RECT 61.26 14.62 61.62 14.98 ;
        RECT 62.01 90.93 62.37 91.29 ;
        RECT 62.01 89.36 62.37 89.72 ;
        RECT 62.01 87.79 62.37 88.15 ;
        RECT 62.01 79.69 62.37 80.05 ;
        RECT 62.01 78.12 62.37 78.48 ;
        RECT 62.01 76.55 62.37 76.91 ;
        RECT 62.01 68.45 62.37 68.81 ;
        RECT 62.01 66.88 62.37 67.24 ;
        RECT 62.01 65.31 62.37 65.67 ;
        RECT 62.01 57.21 62.37 57.57 ;
        RECT 62.01 55.64 62.37 56 ;
        RECT 62.01 54.07 62.37 54.43 ;
        RECT 62.01 45.97 62.37 46.33 ;
        RECT 62.01 44.4 62.37 44.76 ;
        RECT 62.01 42.83 62.37 43.19 ;
        RECT 62.01 34.73 62.37 35.09 ;
        RECT 62.01 33.16 62.37 33.52 ;
        RECT 62.01 31.59 62.37 31.95 ;
        RECT 62.01 23.49 62.37 23.85 ;
        RECT 62.01 21.92 62.37 22.28 ;
        RECT 62.01 20.35 62.37 20.71 ;
        RECT 62.01 12.25 62.37 12.61 ;
        RECT 62.01 10.68 62.37 11.04 ;
        RECT 62.01 9.11 62.37 9.47 ;
        RECT 62.82 90.93 63.18 91.29 ;
        RECT 62.82 89.36 63.18 89.72 ;
        RECT 62.82 87.79 63.18 88.15 ;
        RECT 62.82 79.69 63.18 80.05 ;
        RECT 62.82 78.12 63.18 78.48 ;
        RECT 62.82 76.55 63.18 76.91 ;
        RECT 62.82 68.45 63.18 68.81 ;
        RECT 62.82 66.88 63.18 67.24 ;
        RECT 62.82 65.31 63.18 65.67 ;
        RECT 62.82 57.21 63.18 57.57 ;
        RECT 62.82 55.64 63.18 56 ;
        RECT 62.82 54.07 63.18 54.43 ;
        RECT 62.82 45.97 63.18 46.33 ;
        RECT 62.82 44.4 63.18 44.76 ;
        RECT 62.82 42.83 63.18 43.19 ;
        RECT 62.82 34.73 63.18 35.09 ;
        RECT 62.82 33.16 63.18 33.52 ;
        RECT 62.82 31.59 63.18 31.95 ;
        RECT 62.82 23.49 63.18 23.85 ;
        RECT 62.82 21.92 63.18 22.28 ;
        RECT 62.82 20.35 63.18 20.71 ;
        RECT 62.82 12.25 63.18 12.61 ;
        RECT 62.82 10.68 63.18 11.04 ;
        RECT 62.82 9.11 63.18 9.47 ;
        RECT 62.83 85.3 63.19 85.66 ;
        RECT 62.83 84.49 63.19 84.85 ;
        RECT 62.83 83.68 63.19 84.04 ;
        RECT 62.83 82.87 63.19 83.23 ;
        RECT 62.83 82.06 63.19 82.42 ;
        RECT 62.83 74.06 63.19 74.42 ;
        RECT 62.83 73.25 63.19 73.61 ;
        RECT 62.83 72.44 63.19 72.8 ;
        RECT 62.83 71.63 63.19 71.99 ;
        RECT 62.83 70.82 63.19 71.18 ;
        RECT 62.83 62.82 63.19 63.18 ;
        RECT 62.83 62.01 63.19 62.37 ;
        RECT 62.83 61.2 63.19 61.56 ;
        RECT 62.83 60.39 63.19 60.75 ;
        RECT 62.83 59.58 63.19 59.94 ;
        RECT 62.83 51.58 63.19 51.94 ;
        RECT 62.83 50.77 63.19 51.13 ;
        RECT 62.83 49.96 63.19 50.32 ;
        RECT 62.83 49.15 63.19 49.51 ;
        RECT 62.83 48.34 63.19 48.7 ;
        RECT 62.83 40.34 63.19 40.7 ;
        RECT 62.83 39.53 63.19 39.89 ;
        RECT 62.83 38.72 63.19 39.08 ;
        RECT 62.83 37.91 63.19 38.27 ;
        RECT 62.83 37.1 63.19 37.46 ;
        RECT 62.83 29.1 63.19 29.46 ;
        RECT 62.83 28.29 63.19 28.65 ;
        RECT 62.83 27.48 63.19 27.84 ;
        RECT 62.83 26.67 63.19 27.03 ;
        RECT 62.83 25.86 63.19 26.22 ;
        RECT 62.83 17.86 63.19 18.22 ;
        RECT 62.83 17.05 63.19 17.41 ;
        RECT 62.83 16.24 63.19 16.6 ;
        RECT 62.83 15.43 63.19 15.79 ;
        RECT 62.83 14.62 63.19 14.98 ;
        RECT 65.25 90.92 65.61 91.28 ;
        RECT 65.25 90.11 65.61 90.47 ;
        RECT 65.25 89.3 65.61 89.66 ;
        RECT 65.25 88.49 65.61 88.85 ;
        RECT 65.25 87.68 65.61 88.04 ;
        RECT 65.25 79.68 65.61 80.04 ;
        RECT 65.25 78.87 65.61 79.23 ;
        RECT 65.25 78.06 65.61 78.42 ;
        RECT 65.25 77.25 65.61 77.61 ;
        RECT 65.25 76.44 65.61 76.8 ;
        RECT 65.25 68.44 65.61 68.8 ;
        RECT 65.25 67.63 65.61 67.99 ;
        RECT 65.25 66.82 65.61 67.18 ;
        RECT 65.25 66.01 65.61 66.37 ;
        RECT 65.25 65.2 65.61 65.56 ;
        RECT 65.25 57.2 65.61 57.56 ;
        RECT 65.25 56.39 65.61 56.75 ;
        RECT 65.25 55.58 65.61 55.94 ;
        RECT 65.25 54.77 65.61 55.13 ;
        RECT 65.25 53.96 65.61 54.32 ;
        RECT 65.25 45.96 65.61 46.32 ;
        RECT 65.25 45.15 65.61 45.51 ;
        RECT 65.25 44.34 65.61 44.7 ;
        RECT 65.25 43.53 65.61 43.89 ;
        RECT 65.25 42.72 65.61 43.08 ;
        RECT 65.25 34.72 65.61 35.08 ;
        RECT 65.25 33.91 65.61 34.27 ;
        RECT 65.25 33.1 65.61 33.46 ;
        RECT 65.25 32.29 65.61 32.65 ;
        RECT 65.25 31.48 65.61 31.84 ;
        RECT 65.25 23.48 65.61 23.84 ;
        RECT 65.25 22.67 65.61 23.03 ;
        RECT 65.25 21.86 65.61 22.22 ;
        RECT 65.25 21.05 65.61 21.41 ;
        RECT 65.25 20.24 65.61 20.6 ;
        RECT 65.25 12.24 65.61 12.6 ;
        RECT 65.25 11.43 65.61 11.79 ;
        RECT 65.25 10.62 65.61 10.98 ;
        RECT 65.25 9.81 65.61 10.17 ;
        RECT 65.25 9 65.61 9.36 ;
        RECT 65.26 85.31 65.62 85.67 ;
        RECT 65.26 83.74 65.62 84.1 ;
        RECT 65.26 82.17 65.62 82.53 ;
        RECT 65.26 74.07 65.62 74.43 ;
        RECT 65.26 72.5 65.62 72.86 ;
        RECT 65.26 70.93 65.62 71.29 ;
        RECT 65.26 62.83 65.62 63.19 ;
        RECT 65.26 61.26 65.62 61.62 ;
        RECT 65.26 59.69 65.62 60.05 ;
        RECT 65.26 51.59 65.62 51.95 ;
        RECT 65.26 50.02 65.62 50.38 ;
        RECT 65.26 48.45 65.62 48.81 ;
        RECT 65.26 40.35 65.62 40.71 ;
        RECT 65.26 38.78 65.62 39.14 ;
        RECT 65.26 37.21 65.62 37.57 ;
        RECT 65.26 29.11 65.62 29.47 ;
        RECT 65.26 27.54 65.62 27.9 ;
        RECT 65.26 25.97 65.62 26.33 ;
        RECT 65.26 17.87 65.62 18.23 ;
        RECT 65.26 16.3 65.62 16.66 ;
        RECT 65.26 14.73 65.62 15.09 ;
        RECT 66.07 85.31 66.43 85.67 ;
        RECT 66.07 83.74 66.43 84.1 ;
        RECT 66.07 82.17 66.43 82.53 ;
        RECT 66.07 74.07 66.43 74.43 ;
        RECT 66.07 72.5 66.43 72.86 ;
        RECT 66.07 70.93 66.43 71.29 ;
        RECT 66.07 62.83 66.43 63.19 ;
        RECT 66.07 61.26 66.43 61.62 ;
        RECT 66.07 59.69 66.43 60.05 ;
        RECT 66.07 51.59 66.43 51.95 ;
        RECT 66.07 50.02 66.43 50.38 ;
        RECT 66.07 48.45 66.43 48.81 ;
        RECT 66.07 40.35 66.43 40.71 ;
        RECT 66.07 38.78 66.43 39.14 ;
        RECT 66.07 37.21 66.43 37.57 ;
        RECT 66.07 29.11 66.43 29.47 ;
        RECT 66.07 27.54 66.43 27.9 ;
        RECT 66.07 25.97 66.43 26.33 ;
        RECT 66.07 17.87 66.43 18.23 ;
        RECT 66.07 16.3 66.43 16.66 ;
        RECT 66.07 14.73 66.43 15.09 ;
        RECT 66.82 90.92 67.18 91.28 ;
        RECT 66.82 90.11 67.18 90.47 ;
        RECT 66.82 89.3 67.18 89.66 ;
        RECT 66.82 88.49 67.18 88.85 ;
        RECT 66.82 87.68 67.18 88.04 ;
        RECT 66.82 79.68 67.18 80.04 ;
        RECT 66.82 78.87 67.18 79.23 ;
        RECT 66.82 78.06 67.18 78.42 ;
        RECT 66.82 77.25 67.18 77.61 ;
        RECT 66.82 76.44 67.18 76.8 ;
        RECT 66.82 68.44 67.18 68.8 ;
        RECT 66.82 67.63 67.18 67.99 ;
        RECT 66.82 66.82 67.18 67.18 ;
        RECT 66.82 66.01 67.18 66.37 ;
        RECT 66.82 65.2 67.18 65.56 ;
        RECT 66.82 57.2 67.18 57.56 ;
        RECT 66.82 56.39 67.18 56.75 ;
        RECT 66.82 55.58 67.18 55.94 ;
        RECT 66.82 54.77 67.18 55.13 ;
        RECT 66.82 53.96 67.18 54.32 ;
        RECT 66.82 45.96 67.18 46.32 ;
        RECT 66.82 45.15 67.18 45.51 ;
        RECT 66.82 44.34 67.18 44.7 ;
        RECT 66.82 43.53 67.18 43.89 ;
        RECT 66.82 42.72 67.18 43.08 ;
        RECT 66.82 34.72 67.18 35.08 ;
        RECT 66.82 33.91 67.18 34.27 ;
        RECT 66.82 33.1 67.18 33.46 ;
        RECT 66.82 32.29 67.18 32.65 ;
        RECT 66.82 31.48 67.18 31.84 ;
        RECT 66.82 23.48 67.18 23.84 ;
        RECT 66.82 22.67 67.18 23.03 ;
        RECT 66.82 21.86 67.18 22.22 ;
        RECT 66.82 21.05 67.18 21.41 ;
        RECT 66.82 20.24 67.18 20.6 ;
        RECT 66.82 12.24 67.18 12.6 ;
        RECT 66.82 11.43 67.18 11.79 ;
        RECT 66.82 10.62 67.18 10.98 ;
        RECT 66.82 9.81 67.18 10.17 ;
        RECT 66.82 9 67.18 9.36 ;
        RECT 66.88 85.31 67.24 85.67 ;
        RECT 66.88 83.74 67.24 84.1 ;
        RECT 66.88 82.17 67.24 82.53 ;
        RECT 66.88 74.07 67.24 74.43 ;
        RECT 66.88 72.5 67.24 72.86 ;
        RECT 66.88 70.93 67.24 71.29 ;
        RECT 66.88 62.83 67.24 63.19 ;
        RECT 66.88 61.26 67.24 61.62 ;
        RECT 66.88 59.69 67.24 60.05 ;
        RECT 66.88 51.59 67.24 51.95 ;
        RECT 66.88 50.02 67.24 50.38 ;
        RECT 66.88 48.45 67.24 48.81 ;
        RECT 66.88 40.35 67.24 40.71 ;
        RECT 66.88 38.78 67.24 39.14 ;
        RECT 66.88 37.21 67.24 37.57 ;
        RECT 66.88 29.11 67.24 29.47 ;
        RECT 66.88 27.54 67.24 27.9 ;
        RECT 66.88 25.97 67.24 26.33 ;
        RECT 66.88 17.87 67.24 18.23 ;
        RECT 66.88 16.3 67.24 16.66 ;
        RECT 66.88 14.73 67.24 15.09 ;
        RECT 67.69 85.31 68.05 85.67 ;
        RECT 67.69 83.74 68.05 84.1 ;
        RECT 67.69 82.17 68.05 82.53 ;
        RECT 67.69 74.07 68.05 74.43 ;
        RECT 67.69 72.5 68.05 72.86 ;
        RECT 67.69 70.93 68.05 71.29 ;
        RECT 67.69 62.83 68.05 63.19 ;
        RECT 67.69 61.26 68.05 61.62 ;
        RECT 67.69 59.69 68.05 60.05 ;
        RECT 67.69 51.59 68.05 51.95 ;
        RECT 67.69 50.02 68.05 50.38 ;
        RECT 67.69 48.45 68.05 48.81 ;
        RECT 67.69 40.35 68.05 40.71 ;
        RECT 67.69 38.78 68.05 39.14 ;
        RECT 67.69 37.21 68.05 37.57 ;
        RECT 67.69 29.11 68.05 29.47 ;
        RECT 67.69 27.54 68.05 27.9 ;
        RECT 67.69 25.97 68.05 26.33 ;
        RECT 67.69 17.87 68.05 18.23 ;
        RECT 67.69 16.3 68.05 16.66 ;
        RECT 67.69 14.73 68.05 15.09 ;
        RECT 68.39 90.92 68.75 91.28 ;
        RECT 68.39 90.11 68.75 90.47 ;
        RECT 68.39 89.3 68.75 89.66 ;
        RECT 68.39 88.49 68.75 88.85 ;
        RECT 68.39 87.68 68.75 88.04 ;
        RECT 68.39 79.68 68.75 80.04 ;
        RECT 68.39 78.87 68.75 79.23 ;
        RECT 68.39 78.06 68.75 78.42 ;
        RECT 68.39 77.25 68.75 77.61 ;
        RECT 68.39 76.44 68.75 76.8 ;
        RECT 68.39 68.44 68.75 68.8 ;
        RECT 68.39 67.63 68.75 67.99 ;
        RECT 68.39 66.82 68.75 67.18 ;
        RECT 68.39 66.01 68.75 66.37 ;
        RECT 68.39 65.2 68.75 65.56 ;
        RECT 68.39 57.2 68.75 57.56 ;
        RECT 68.39 56.39 68.75 56.75 ;
        RECT 68.39 55.58 68.75 55.94 ;
        RECT 68.39 54.77 68.75 55.13 ;
        RECT 68.39 53.96 68.75 54.32 ;
        RECT 68.39 45.96 68.75 46.32 ;
        RECT 68.39 45.15 68.75 45.51 ;
        RECT 68.39 44.34 68.75 44.7 ;
        RECT 68.39 43.53 68.75 43.89 ;
        RECT 68.39 42.72 68.75 43.08 ;
        RECT 68.39 34.72 68.75 35.08 ;
        RECT 68.39 33.91 68.75 34.27 ;
        RECT 68.39 33.1 68.75 33.46 ;
        RECT 68.39 32.29 68.75 32.65 ;
        RECT 68.39 31.48 68.75 31.84 ;
        RECT 68.39 23.48 68.75 23.84 ;
        RECT 68.39 22.67 68.75 23.03 ;
        RECT 68.39 21.86 68.75 22.22 ;
        RECT 68.39 21.05 68.75 21.41 ;
        RECT 68.39 20.24 68.75 20.6 ;
        RECT 68.39 12.24 68.75 12.6 ;
        RECT 68.39 11.43 68.75 11.79 ;
        RECT 68.39 10.62 68.75 10.98 ;
        RECT 68.39 9.81 68.75 10.17 ;
        RECT 68.39 9 68.75 9.36 ;
        RECT 68.5 85.31 68.86 85.67 ;
        RECT 68.5 83.74 68.86 84.1 ;
        RECT 68.5 82.17 68.86 82.53 ;
        RECT 68.5 74.07 68.86 74.43 ;
        RECT 68.5 72.5 68.86 72.86 ;
        RECT 68.5 70.93 68.86 71.29 ;
        RECT 68.5 62.83 68.86 63.19 ;
        RECT 68.5 61.26 68.86 61.62 ;
        RECT 68.5 59.69 68.86 60.05 ;
        RECT 68.5 51.59 68.86 51.95 ;
        RECT 68.5 50.02 68.86 50.38 ;
        RECT 68.5 48.45 68.86 48.81 ;
        RECT 68.5 40.35 68.86 40.71 ;
        RECT 68.5 38.78 68.86 39.14 ;
        RECT 68.5 37.21 68.86 37.57 ;
        RECT 68.5 29.11 68.86 29.47 ;
        RECT 68.5 27.54 68.86 27.9 ;
        RECT 68.5 25.97 68.86 26.33 ;
        RECT 68.5 17.87 68.86 18.23 ;
        RECT 68.5 16.3 68.86 16.66 ;
        RECT 68.5 14.73 68.86 15.09 ;
        RECT 70.82 90.93 71.18 91.29 ;
        RECT 70.82 89.36 71.18 89.72 ;
        RECT 70.82 87.79 71.18 88.15 ;
        RECT 70.82 79.69 71.18 80.05 ;
        RECT 70.82 78.12 71.18 78.48 ;
        RECT 70.82 76.55 71.18 76.91 ;
        RECT 70.82 68.45 71.18 68.81 ;
        RECT 70.82 66.88 71.18 67.24 ;
        RECT 70.82 65.31 71.18 65.67 ;
        RECT 70.82 57.21 71.18 57.57 ;
        RECT 70.82 55.64 71.18 56 ;
        RECT 70.82 54.07 71.18 54.43 ;
        RECT 70.82 45.97 71.18 46.33 ;
        RECT 70.82 44.4 71.18 44.76 ;
        RECT 70.82 42.83 71.18 43.19 ;
        RECT 70.82 34.73 71.18 35.09 ;
        RECT 70.82 33.16 71.18 33.52 ;
        RECT 70.82 31.59 71.18 31.95 ;
        RECT 70.82 23.49 71.18 23.85 ;
        RECT 70.82 21.92 71.18 22.28 ;
        RECT 70.82 20.35 71.18 20.71 ;
        RECT 70.82 12.25 71.18 12.61 ;
        RECT 70.82 10.68 71.18 11.04 ;
        RECT 70.82 9.11 71.18 9.47 ;
        RECT 70.93 85.3 71.29 85.66 ;
        RECT 70.93 84.49 71.29 84.85 ;
        RECT 70.93 83.68 71.29 84.04 ;
        RECT 70.93 82.87 71.29 83.23 ;
        RECT 70.93 82.06 71.29 82.42 ;
        RECT 70.93 74.06 71.29 74.42 ;
        RECT 70.93 73.25 71.29 73.61 ;
        RECT 70.93 72.44 71.29 72.8 ;
        RECT 70.93 71.63 71.29 71.99 ;
        RECT 70.93 70.82 71.29 71.18 ;
        RECT 70.93 62.82 71.29 63.18 ;
        RECT 70.93 62.01 71.29 62.37 ;
        RECT 70.93 61.2 71.29 61.56 ;
        RECT 70.93 60.39 71.29 60.75 ;
        RECT 70.93 59.58 71.29 59.94 ;
        RECT 70.93 51.58 71.29 51.94 ;
        RECT 70.93 50.77 71.29 51.13 ;
        RECT 70.93 49.96 71.29 50.32 ;
        RECT 70.93 49.15 71.29 49.51 ;
        RECT 70.93 48.34 71.29 48.7 ;
        RECT 70.93 40.34 71.29 40.7 ;
        RECT 70.93 39.53 71.29 39.89 ;
        RECT 70.93 38.72 71.29 39.08 ;
        RECT 70.93 37.91 71.29 38.27 ;
        RECT 70.93 37.1 71.29 37.46 ;
        RECT 70.93 29.1 71.29 29.46 ;
        RECT 70.93 28.29 71.29 28.65 ;
        RECT 70.93 27.48 71.29 27.84 ;
        RECT 70.93 26.67 71.29 27.03 ;
        RECT 70.93 25.86 71.29 26.22 ;
        RECT 70.93 17.86 71.29 18.22 ;
        RECT 70.93 17.05 71.29 17.41 ;
        RECT 70.93 16.24 71.29 16.6 ;
        RECT 70.93 15.43 71.29 15.79 ;
        RECT 70.93 14.62 71.29 14.98 ;
        RECT 71.63 90.93 71.99 91.29 ;
        RECT 71.63 89.36 71.99 89.72 ;
        RECT 71.63 87.79 71.99 88.15 ;
        RECT 71.63 79.69 71.99 80.05 ;
        RECT 71.63 78.12 71.99 78.48 ;
        RECT 71.63 76.55 71.99 76.91 ;
        RECT 71.63 68.45 71.99 68.81 ;
        RECT 71.63 66.88 71.99 67.24 ;
        RECT 71.63 65.31 71.99 65.67 ;
        RECT 71.63 57.21 71.99 57.57 ;
        RECT 71.63 55.64 71.99 56 ;
        RECT 71.63 54.07 71.99 54.43 ;
        RECT 71.63 45.97 71.99 46.33 ;
        RECT 71.63 44.4 71.99 44.76 ;
        RECT 71.63 42.83 71.99 43.19 ;
        RECT 71.63 34.73 71.99 35.09 ;
        RECT 71.63 33.16 71.99 33.52 ;
        RECT 71.63 31.59 71.99 31.95 ;
        RECT 71.63 23.49 71.99 23.85 ;
        RECT 71.63 21.92 71.99 22.28 ;
        RECT 71.63 20.35 71.99 20.71 ;
        RECT 71.63 12.25 71.99 12.61 ;
        RECT 71.63 10.68 71.99 11.04 ;
        RECT 71.63 9.11 71.99 9.47 ;
        RECT 72.44 90.93 72.8 91.29 ;
        RECT 72.44 89.36 72.8 89.72 ;
        RECT 72.44 87.79 72.8 88.15 ;
        RECT 72.44 79.69 72.8 80.05 ;
        RECT 72.44 78.12 72.8 78.48 ;
        RECT 72.44 76.55 72.8 76.91 ;
        RECT 72.44 68.45 72.8 68.81 ;
        RECT 72.44 66.88 72.8 67.24 ;
        RECT 72.44 65.31 72.8 65.67 ;
        RECT 72.44 57.21 72.8 57.57 ;
        RECT 72.44 55.64 72.8 56 ;
        RECT 72.44 54.07 72.8 54.43 ;
        RECT 72.44 45.97 72.8 46.33 ;
        RECT 72.44 44.4 72.8 44.76 ;
        RECT 72.44 42.83 72.8 43.19 ;
        RECT 72.44 34.73 72.8 35.09 ;
        RECT 72.44 33.16 72.8 33.52 ;
        RECT 72.44 31.59 72.8 31.95 ;
        RECT 72.44 23.49 72.8 23.85 ;
        RECT 72.44 21.92 72.8 22.28 ;
        RECT 72.44 20.35 72.8 20.71 ;
        RECT 72.44 12.25 72.8 12.61 ;
        RECT 72.44 10.68 72.8 11.04 ;
        RECT 72.44 9.11 72.8 9.47 ;
        RECT 72.5 85.3 72.86 85.66 ;
        RECT 72.5 84.49 72.86 84.85 ;
        RECT 72.5 83.68 72.86 84.04 ;
        RECT 72.5 82.87 72.86 83.23 ;
        RECT 72.5 82.06 72.86 82.42 ;
        RECT 72.5 74.06 72.86 74.42 ;
        RECT 72.5 73.25 72.86 73.61 ;
        RECT 72.5 72.44 72.86 72.8 ;
        RECT 72.5 71.63 72.86 71.99 ;
        RECT 72.5 70.82 72.86 71.18 ;
        RECT 72.5 62.82 72.86 63.18 ;
        RECT 72.5 62.01 72.86 62.37 ;
        RECT 72.5 61.2 72.86 61.56 ;
        RECT 72.5 60.39 72.86 60.75 ;
        RECT 72.5 59.58 72.86 59.94 ;
        RECT 72.5 51.58 72.86 51.94 ;
        RECT 72.5 50.77 72.86 51.13 ;
        RECT 72.5 49.96 72.86 50.32 ;
        RECT 72.5 49.15 72.86 49.51 ;
        RECT 72.5 48.34 72.86 48.7 ;
        RECT 72.5 40.34 72.86 40.7 ;
        RECT 72.5 39.53 72.86 39.89 ;
        RECT 72.5 38.72 72.86 39.08 ;
        RECT 72.5 37.91 72.86 38.27 ;
        RECT 72.5 37.1 72.86 37.46 ;
        RECT 72.5 29.1 72.86 29.46 ;
        RECT 72.5 28.29 72.86 28.65 ;
        RECT 72.5 27.48 72.86 27.84 ;
        RECT 72.5 26.67 72.86 27.03 ;
        RECT 72.5 25.86 72.86 26.22 ;
        RECT 72.5 17.86 72.86 18.22 ;
        RECT 72.5 17.05 72.86 17.41 ;
        RECT 72.5 16.24 72.86 16.6 ;
        RECT 72.5 15.43 72.86 15.79 ;
        RECT 72.5 14.62 72.86 14.98 ;
        RECT 73.25 90.93 73.61 91.29 ;
        RECT 73.25 89.36 73.61 89.72 ;
        RECT 73.25 87.79 73.61 88.15 ;
        RECT 73.25 79.69 73.61 80.05 ;
        RECT 73.25 78.12 73.61 78.48 ;
        RECT 73.25 76.55 73.61 76.91 ;
        RECT 73.25 68.45 73.61 68.81 ;
        RECT 73.25 66.88 73.61 67.24 ;
        RECT 73.25 65.31 73.61 65.67 ;
        RECT 73.25 57.21 73.61 57.57 ;
        RECT 73.25 55.64 73.61 56 ;
        RECT 73.25 54.07 73.61 54.43 ;
        RECT 73.25 45.97 73.61 46.33 ;
        RECT 73.25 44.4 73.61 44.76 ;
        RECT 73.25 42.83 73.61 43.19 ;
        RECT 73.25 34.73 73.61 35.09 ;
        RECT 73.25 33.16 73.61 33.52 ;
        RECT 73.25 31.59 73.61 31.95 ;
        RECT 73.25 23.49 73.61 23.85 ;
        RECT 73.25 21.92 73.61 22.28 ;
        RECT 73.25 20.35 73.61 20.71 ;
        RECT 73.25 12.25 73.61 12.61 ;
        RECT 73.25 10.68 73.61 11.04 ;
        RECT 73.25 9.11 73.61 9.47 ;
        RECT 74.06 90.93 74.42 91.29 ;
        RECT 74.06 89.36 74.42 89.72 ;
        RECT 74.06 87.79 74.42 88.15 ;
        RECT 74.06 79.69 74.42 80.05 ;
        RECT 74.06 78.12 74.42 78.48 ;
        RECT 74.06 76.55 74.42 76.91 ;
        RECT 74.06 68.45 74.42 68.81 ;
        RECT 74.06 66.88 74.42 67.24 ;
        RECT 74.06 65.31 74.42 65.67 ;
        RECT 74.06 57.21 74.42 57.57 ;
        RECT 74.06 55.64 74.42 56 ;
        RECT 74.06 54.07 74.42 54.43 ;
        RECT 74.06 45.97 74.42 46.33 ;
        RECT 74.06 44.4 74.42 44.76 ;
        RECT 74.06 42.83 74.42 43.19 ;
        RECT 74.06 34.73 74.42 35.09 ;
        RECT 74.06 33.16 74.42 33.52 ;
        RECT 74.06 31.59 74.42 31.95 ;
        RECT 74.06 23.49 74.42 23.85 ;
        RECT 74.06 21.92 74.42 22.28 ;
        RECT 74.06 20.35 74.42 20.71 ;
        RECT 74.06 12.25 74.42 12.61 ;
        RECT 74.06 10.68 74.42 11.04 ;
        RECT 74.06 9.11 74.42 9.47 ;
        RECT 74.07 85.3 74.43 85.66 ;
        RECT 74.07 84.49 74.43 84.85 ;
        RECT 74.07 83.68 74.43 84.04 ;
        RECT 74.07 82.87 74.43 83.23 ;
        RECT 74.07 82.06 74.43 82.42 ;
        RECT 74.07 74.06 74.43 74.42 ;
        RECT 74.07 73.25 74.43 73.61 ;
        RECT 74.07 72.44 74.43 72.8 ;
        RECT 74.07 71.63 74.43 71.99 ;
        RECT 74.07 70.82 74.43 71.18 ;
        RECT 74.07 62.82 74.43 63.18 ;
        RECT 74.07 62.01 74.43 62.37 ;
        RECT 74.07 61.2 74.43 61.56 ;
        RECT 74.07 60.39 74.43 60.75 ;
        RECT 74.07 59.58 74.43 59.94 ;
        RECT 74.07 51.58 74.43 51.94 ;
        RECT 74.07 50.77 74.43 51.13 ;
        RECT 74.07 49.96 74.43 50.32 ;
        RECT 74.07 49.15 74.43 49.51 ;
        RECT 74.07 48.34 74.43 48.7 ;
        RECT 74.07 40.34 74.43 40.7 ;
        RECT 74.07 39.53 74.43 39.89 ;
        RECT 74.07 38.72 74.43 39.08 ;
        RECT 74.07 37.91 74.43 38.27 ;
        RECT 74.07 37.1 74.43 37.46 ;
        RECT 74.07 29.1 74.43 29.46 ;
        RECT 74.07 28.29 74.43 28.65 ;
        RECT 74.07 27.48 74.43 27.84 ;
        RECT 74.07 26.67 74.43 27.03 ;
        RECT 74.07 25.86 74.43 26.22 ;
        RECT 74.07 17.86 74.43 18.22 ;
        RECT 74.07 17.05 74.43 17.41 ;
        RECT 74.07 16.24 74.43 16.6 ;
        RECT 74.07 15.43 74.43 15.79 ;
        RECT 74.07 14.62 74.43 14.98 ;
        RECT 76.49 90.92 76.85 91.28 ;
        RECT 76.49 90.11 76.85 90.47 ;
        RECT 76.49 89.3 76.85 89.66 ;
        RECT 76.49 88.49 76.85 88.85 ;
        RECT 76.49 87.68 76.85 88.04 ;
        RECT 76.49 79.68 76.85 80.04 ;
        RECT 76.49 78.87 76.85 79.23 ;
        RECT 76.49 78.06 76.85 78.42 ;
        RECT 76.49 77.25 76.85 77.61 ;
        RECT 76.49 76.44 76.85 76.8 ;
        RECT 76.49 68.44 76.85 68.8 ;
        RECT 76.49 67.63 76.85 67.99 ;
        RECT 76.49 66.82 76.85 67.18 ;
        RECT 76.49 66.01 76.85 66.37 ;
        RECT 76.49 65.2 76.85 65.56 ;
        RECT 76.49 57.2 76.85 57.56 ;
        RECT 76.49 56.39 76.85 56.75 ;
        RECT 76.49 55.58 76.85 55.94 ;
        RECT 76.49 54.77 76.85 55.13 ;
        RECT 76.49 53.96 76.85 54.32 ;
        RECT 76.49 45.96 76.85 46.32 ;
        RECT 76.49 45.15 76.85 45.51 ;
        RECT 76.49 44.34 76.85 44.7 ;
        RECT 76.49 43.53 76.85 43.89 ;
        RECT 76.49 42.72 76.85 43.08 ;
        RECT 76.49 34.72 76.85 35.08 ;
        RECT 76.49 33.91 76.85 34.27 ;
        RECT 76.49 33.1 76.85 33.46 ;
        RECT 76.49 32.29 76.85 32.65 ;
        RECT 76.49 31.48 76.85 31.84 ;
        RECT 76.49 23.48 76.85 23.84 ;
        RECT 76.49 22.67 76.85 23.03 ;
        RECT 76.49 21.86 76.85 22.22 ;
        RECT 76.49 21.05 76.85 21.41 ;
        RECT 76.49 20.24 76.85 20.6 ;
        RECT 76.49 12.24 76.85 12.6 ;
        RECT 76.49 11.43 76.85 11.79 ;
        RECT 76.49 10.62 76.85 10.98 ;
        RECT 76.49 9.81 76.85 10.17 ;
        RECT 76.49 9 76.85 9.36 ;
        RECT 76.5 85.31 76.86 85.67 ;
        RECT 76.5 83.74 76.86 84.1 ;
        RECT 76.5 82.17 76.86 82.53 ;
        RECT 76.5 74.07 76.86 74.43 ;
        RECT 76.5 72.5 76.86 72.86 ;
        RECT 76.5 70.93 76.86 71.29 ;
        RECT 76.5 62.83 76.86 63.19 ;
        RECT 76.5 61.26 76.86 61.62 ;
        RECT 76.5 59.69 76.86 60.05 ;
        RECT 76.5 51.59 76.86 51.95 ;
        RECT 76.5 50.02 76.86 50.38 ;
        RECT 76.5 48.45 76.86 48.81 ;
        RECT 76.5 40.35 76.86 40.71 ;
        RECT 76.5 38.78 76.86 39.14 ;
        RECT 76.5 37.21 76.86 37.57 ;
        RECT 76.5 29.11 76.86 29.47 ;
        RECT 76.5 27.54 76.86 27.9 ;
        RECT 76.5 25.97 76.86 26.33 ;
        RECT 76.5 17.87 76.86 18.23 ;
        RECT 76.5 16.3 76.86 16.66 ;
        RECT 76.5 14.73 76.86 15.09 ;
        RECT 77.31 85.31 77.67 85.67 ;
        RECT 77.31 83.74 77.67 84.1 ;
        RECT 77.31 82.17 77.67 82.53 ;
        RECT 77.31 74.07 77.67 74.43 ;
        RECT 77.31 72.5 77.67 72.86 ;
        RECT 77.31 70.93 77.67 71.29 ;
        RECT 77.31 62.83 77.67 63.19 ;
        RECT 77.31 61.26 77.67 61.62 ;
        RECT 77.31 59.69 77.67 60.05 ;
        RECT 77.31 51.59 77.67 51.95 ;
        RECT 77.31 50.02 77.67 50.38 ;
        RECT 77.31 48.45 77.67 48.81 ;
        RECT 77.31 40.35 77.67 40.71 ;
        RECT 77.31 38.78 77.67 39.14 ;
        RECT 77.31 37.21 77.67 37.57 ;
        RECT 77.31 29.11 77.67 29.47 ;
        RECT 77.31 27.54 77.67 27.9 ;
        RECT 77.31 25.97 77.67 26.33 ;
        RECT 77.31 17.87 77.67 18.23 ;
        RECT 77.31 16.3 77.67 16.66 ;
        RECT 77.31 14.73 77.67 15.09 ;
        RECT 78.06 90.92 78.42 91.28 ;
        RECT 78.06 90.11 78.42 90.47 ;
        RECT 78.06 89.3 78.42 89.66 ;
        RECT 78.06 88.49 78.42 88.85 ;
        RECT 78.06 87.68 78.42 88.04 ;
        RECT 78.06 79.68 78.42 80.04 ;
        RECT 78.06 78.87 78.42 79.23 ;
        RECT 78.06 78.06 78.42 78.42 ;
        RECT 78.06 77.25 78.42 77.61 ;
        RECT 78.06 76.44 78.42 76.8 ;
        RECT 78.06 68.44 78.42 68.8 ;
        RECT 78.06 67.63 78.42 67.99 ;
        RECT 78.06 66.82 78.42 67.18 ;
        RECT 78.06 66.01 78.42 66.37 ;
        RECT 78.06 65.2 78.42 65.56 ;
        RECT 78.06 57.2 78.42 57.56 ;
        RECT 78.06 56.39 78.42 56.75 ;
        RECT 78.06 55.58 78.42 55.94 ;
        RECT 78.06 54.77 78.42 55.13 ;
        RECT 78.06 53.96 78.42 54.32 ;
        RECT 78.06 45.96 78.42 46.32 ;
        RECT 78.06 45.15 78.42 45.51 ;
        RECT 78.06 44.34 78.42 44.7 ;
        RECT 78.06 43.53 78.42 43.89 ;
        RECT 78.06 42.72 78.42 43.08 ;
        RECT 78.06 34.72 78.42 35.08 ;
        RECT 78.06 33.91 78.42 34.27 ;
        RECT 78.06 33.1 78.42 33.46 ;
        RECT 78.06 32.29 78.42 32.65 ;
        RECT 78.06 31.48 78.42 31.84 ;
        RECT 78.06 23.48 78.42 23.84 ;
        RECT 78.06 22.67 78.42 23.03 ;
        RECT 78.06 21.86 78.42 22.22 ;
        RECT 78.06 21.05 78.42 21.41 ;
        RECT 78.06 20.24 78.42 20.6 ;
        RECT 78.06 12.24 78.42 12.6 ;
        RECT 78.06 11.43 78.42 11.79 ;
        RECT 78.06 10.62 78.42 10.98 ;
        RECT 78.06 9.81 78.42 10.17 ;
        RECT 78.06 9 78.42 9.36 ;
        RECT 78.12 85.31 78.48 85.67 ;
        RECT 78.12 83.74 78.48 84.1 ;
        RECT 78.12 82.17 78.48 82.53 ;
        RECT 78.12 74.07 78.48 74.43 ;
        RECT 78.12 72.5 78.48 72.86 ;
        RECT 78.12 70.93 78.48 71.29 ;
        RECT 78.12 62.83 78.48 63.19 ;
        RECT 78.12 61.26 78.48 61.62 ;
        RECT 78.12 59.69 78.48 60.05 ;
        RECT 78.12 51.59 78.48 51.95 ;
        RECT 78.12 50.02 78.48 50.38 ;
        RECT 78.12 48.45 78.48 48.81 ;
        RECT 78.12 40.35 78.48 40.71 ;
        RECT 78.12 38.78 78.48 39.14 ;
        RECT 78.12 37.21 78.48 37.57 ;
        RECT 78.12 29.11 78.48 29.47 ;
        RECT 78.12 27.54 78.48 27.9 ;
        RECT 78.12 25.97 78.48 26.33 ;
        RECT 78.12 17.87 78.48 18.23 ;
        RECT 78.12 16.3 78.48 16.66 ;
        RECT 78.12 14.73 78.48 15.09 ;
        RECT 78.93 85.31 79.29 85.67 ;
        RECT 78.93 83.74 79.29 84.1 ;
        RECT 78.93 82.17 79.29 82.53 ;
        RECT 78.93 74.07 79.29 74.43 ;
        RECT 78.93 72.5 79.29 72.86 ;
        RECT 78.93 70.93 79.29 71.29 ;
        RECT 78.93 62.83 79.29 63.19 ;
        RECT 78.93 61.26 79.29 61.62 ;
        RECT 78.93 59.69 79.29 60.05 ;
        RECT 78.93 51.59 79.29 51.95 ;
        RECT 78.93 50.02 79.29 50.38 ;
        RECT 78.93 48.45 79.29 48.81 ;
        RECT 78.93 40.35 79.29 40.71 ;
        RECT 78.93 38.78 79.29 39.14 ;
        RECT 78.93 37.21 79.29 37.57 ;
        RECT 78.93 29.11 79.29 29.47 ;
        RECT 78.93 27.54 79.29 27.9 ;
        RECT 78.93 25.97 79.29 26.33 ;
        RECT 78.93 17.87 79.29 18.23 ;
        RECT 78.93 16.3 79.29 16.66 ;
        RECT 78.93 14.73 79.29 15.09 ;
        RECT 79.63 90.92 79.99 91.28 ;
        RECT 79.63 90.11 79.99 90.47 ;
        RECT 79.63 89.3 79.99 89.66 ;
        RECT 79.63 88.49 79.99 88.85 ;
        RECT 79.63 87.68 79.99 88.04 ;
        RECT 79.63 79.68 79.99 80.04 ;
        RECT 79.63 78.87 79.99 79.23 ;
        RECT 79.63 78.06 79.99 78.42 ;
        RECT 79.63 77.25 79.99 77.61 ;
        RECT 79.63 76.44 79.99 76.8 ;
        RECT 79.63 68.44 79.99 68.8 ;
        RECT 79.63 67.63 79.99 67.99 ;
        RECT 79.63 66.82 79.99 67.18 ;
        RECT 79.63 66.01 79.99 66.37 ;
        RECT 79.63 65.2 79.99 65.56 ;
        RECT 79.63 57.2 79.99 57.56 ;
        RECT 79.63 56.39 79.99 56.75 ;
        RECT 79.63 55.58 79.99 55.94 ;
        RECT 79.63 54.77 79.99 55.13 ;
        RECT 79.63 53.96 79.99 54.32 ;
        RECT 79.63 45.96 79.99 46.32 ;
        RECT 79.63 45.15 79.99 45.51 ;
        RECT 79.63 44.34 79.99 44.7 ;
        RECT 79.63 43.53 79.99 43.89 ;
        RECT 79.63 42.72 79.99 43.08 ;
        RECT 79.63 34.72 79.99 35.08 ;
        RECT 79.63 33.91 79.99 34.27 ;
        RECT 79.63 33.1 79.99 33.46 ;
        RECT 79.63 32.29 79.99 32.65 ;
        RECT 79.63 31.48 79.99 31.84 ;
        RECT 79.63 23.48 79.99 23.84 ;
        RECT 79.63 22.67 79.99 23.03 ;
        RECT 79.63 21.86 79.99 22.22 ;
        RECT 79.63 21.05 79.99 21.41 ;
        RECT 79.63 20.24 79.99 20.6 ;
        RECT 79.63 12.24 79.99 12.6 ;
        RECT 79.63 11.43 79.99 11.79 ;
        RECT 79.63 10.62 79.99 10.98 ;
        RECT 79.63 9.81 79.99 10.17 ;
        RECT 79.63 9 79.99 9.36 ;
        RECT 79.74 85.31 80.1 85.67 ;
        RECT 79.74 83.74 80.1 84.1 ;
        RECT 79.74 82.17 80.1 82.53 ;
        RECT 79.74 74.07 80.1 74.43 ;
        RECT 79.74 72.5 80.1 72.86 ;
        RECT 79.74 70.93 80.1 71.29 ;
        RECT 79.74 62.83 80.1 63.19 ;
        RECT 79.74 61.26 80.1 61.62 ;
        RECT 79.74 59.69 80.1 60.05 ;
        RECT 79.74 51.59 80.1 51.95 ;
        RECT 79.74 50.02 80.1 50.38 ;
        RECT 79.74 48.45 80.1 48.81 ;
        RECT 79.74 40.35 80.1 40.71 ;
        RECT 79.74 38.78 80.1 39.14 ;
        RECT 79.74 37.21 80.1 37.57 ;
        RECT 79.74 29.11 80.1 29.47 ;
        RECT 79.74 27.54 80.1 27.9 ;
        RECT 79.74 25.97 80.1 26.33 ;
        RECT 79.74 17.87 80.1 18.23 ;
        RECT 79.74 16.3 80.1 16.66 ;
        RECT 79.74 14.73 80.1 15.09 ;
        RECT 82.06 90.93 82.42 91.29 ;
        RECT 82.06 89.36 82.42 89.72 ;
        RECT 82.06 87.79 82.42 88.15 ;
        RECT 82.06 79.69 82.42 80.05 ;
        RECT 82.06 78.12 82.42 78.48 ;
        RECT 82.06 76.55 82.42 76.91 ;
        RECT 82.06 68.45 82.42 68.81 ;
        RECT 82.06 66.88 82.42 67.24 ;
        RECT 82.06 65.31 82.42 65.67 ;
        RECT 82.06 57.21 82.42 57.57 ;
        RECT 82.06 55.64 82.42 56 ;
        RECT 82.06 54.07 82.42 54.43 ;
        RECT 82.06 45.97 82.42 46.33 ;
        RECT 82.06 44.4 82.42 44.76 ;
        RECT 82.06 42.83 82.42 43.19 ;
        RECT 82.06 34.73 82.42 35.09 ;
        RECT 82.06 33.16 82.42 33.52 ;
        RECT 82.06 31.59 82.42 31.95 ;
        RECT 82.06 23.49 82.42 23.85 ;
        RECT 82.06 21.92 82.42 22.28 ;
        RECT 82.06 20.35 82.42 20.71 ;
        RECT 82.06 12.25 82.42 12.61 ;
        RECT 82.06 10.68 82.42 11.04 ;
        RECT 82.06 9.11 82.42 9.47 ;
        RECT 82.17 85.3 82.53 85.66 ;
        RECT 82.17 84.49 82.53 84.85 ;
        RECT 82.17 83.68 82.53 84.04 ;
        RECT 82.17 82.87 82.53 83.23 ;
        RECT 82.17 82.06 82.53 82.42 ;
        RECT 82.17 74.06 82.53 74.42 ;
        RECT 82.17 73.25 82.53 73.61 ;
        RECT 82.17 72.44 82.53 72.8 ;
        RECT 82.17 71.63 82.53 71.99 ;
        RECT 82.17 70.82 82.53 71.18 ;
        RECT 82.17 62.82 82.53 63.18 ;
        RECT 82.17 62.01 82.53 62.37 ;
        RECT 82.17 61.2 82.53 61.56 ;
        RECT 82.17 60.39 82.53 60.75 ;
        RECT 82.17 59.58 82.53 59.94 ;
        RECT 82.17 51.58 82.53 51.94 ;
        RECT 82.17 50.77 82.53 51.13 ;
        RECT 82.17 49.96 82.53 50.32 ;
        RECT 82.17 49.15 82.53 49.51 ;
        RECT 82.17 48.34 82.53 48.7 ;
        RECT 82.17 40.34 82.53 40.7 ;
        RECT 82.17 39.53 82.53 39.89 ;
        RECT 82.17 38.72 82.53 39.08 ;
        RECT 82.17 37.91 82.53 38.27 ;
        RECT 82.17 37.1 82.53 37.46 ;
        RECT 82.17 29.1 82.53 29.46 ;
        RECT 82.17 28.29 82.53 28.65 ;
        RECT 82.17 27.48 82.53 27.84 ;
        RECT 82.17 26.67 82.53 27.03 ;
        RECT 82.17 25.86 82.53 26.22 ;
        RECT 82.17 17.86 82.53 18.22 ;
        RECT 82.17 17.05 82.53 17.41 ;
        RECT 82.17 16.24 82.53 16.6 ;
        RECT 82.17 15.43 82.53 15.79 ;
        RECT 82.17 14.62 82.53 14.98 ;
        RECT 82.87 90.93 83.23 91.29 ;
        RECT 82.87 89.36 83.23 89.72 ;
        RECT 82.87 87.79 83.23 88.15 ;
        RECT 82.87 79.69 83.23 80.05 ;
        RECT 82.87 78.12 83.23 78.48 ;
        RECT 82.87 76.55 83.23 76.91 ;
        RECT 82.87 68.45 83.23 68.81 ;
        RECT 82.87 66.88 83.23 67.24 ;
        RECT 82.87 65.31 83.23 65.67 ;
        RECT 82.87 57.21 83.23 57.57 ;
        RECT 82.87 55.64 83.23 56 ;
        RECT 82.87 54.07 83.23 54.43 ;
        RECT 82.87 45.97 83.23 46.33 ;
        RECT 82.87 44.4 83.23 44.76 ;
        RECT 82.87 42.83 83.23 43.19 ;
        RECT 82.87 34.73 83.23 35.09 ;
        RECT 33.1 54.77 33.46 55.13 ;
        RECT 33.1 53.96 33.46 54.32 ;
        RECT 33.1 45.96 33.46 46.32 ;
        RECT 33.1 45.15 33.46 45.51 ;
        RECT 33.1 44.34 33.46 44.7 ;
        RECT 33.1 43.53 33.46 43.89 ;
        RECT 33.1 42.72 33.46 43.08 ;
        RECT 33.1 34.72 33.46 35.08 ;
        RECT 33.1 33.91 33.46 34.27 ;
        RECT 33.1 33.1 33.46 33.46 ;
        RECT 33.1 32.29 33.46 32.65 ;
        RECT 33.1 31.48 33.46 31.84 ;
        RECT 33.1 23.48 33.46 23.84 ;
        RECT 33.1 22.67 33.46 23.03 ;
        RECT 33.1 21.86 33.46 22.22 ;
        RECT 33.1 21.05 33.46 21.41 ;
        RECT 33.1 20.24 33.46 20.6 ;
        RECT 33.1 12.24 33.46 12.6 ;
        RECT 33.1 11.43 33.46 11.79 ;
        RECT 33.1 10.62 33.46 10.98 ;
        RECT 33.1 9.81 33.46 10.17 ;
        RECT 33.1 9 33.46 9.36 ;
        RECT 33.16 85.31 33.52 85.67 ;
        RECT 33.16 83.74 33.52 84.1 ;
        RECT 33.16 82.17 33.52 82.53 ;
        RECT 33.16 74.07 33.52 74.43 ;
        RECT 33.16 72.5 33.52 72.86 ;
        RECT 33.16 70.93 33.52 71.29 ;
        RECT 33.16 62.83 33.52 63.19 ;
        RECT 33.16 61.26 33.52 61.62 ;
        RECT 33.16 59.69 33.52 60.05 ;
        RECT 33.16 51.59 33.52 51.95 ;
        RECT 33.16 50.02 33.52 50.38 ;
        RECT 33.16 48.45 33.52 48.81 ;
        RECT 33.16 40.35 33.52 40.71 ;
        RECT 33.16 38.78 33.52 39.14 ;
        RECT 33.16 37.21 33.52 37.57 ;
        RECT 33.16 29.11 33.52 29.47 ;
        RECT 33.16 27.54 33.52 27.9 ;
        RECT 33.16 25.97 33.52 26.33 ;
        RECT 33.16 17.87 33.52 18.23 ;
        RECT 33.16 16.3 33.52 16.66 ;
        RECT 33.16 14.73 33.52 15.09 ;
        RECT 33.97 85.31 34.33 85.67 ;
        RECT 33.97 83.74 34.33 84.1 ;
        RECT 33.97 82.17 34.33 82.53 ;
        RECT 33.97 74.07 34.33 74.43 ;
        RECT 33.97 72.5 34.33 72.86 ;
        RECT 33.97 70.93 34.33 71.29 ;
        RECT 33.97 62.83 34.33 63.19 ;
        RECT 33.97 61.26 34.33 61.62 ;
        RECT 33.97 59.69 34.33 60.05 ;
        RECT 33.97 51.59 34.33 51.95 ;
        RECT 33.97 50.02 34.33 50.38 ;
        RECT 33.97 48.45 34.33 48.81 ;
        RECT 33.97 40.35 34.33 40.71 ;
        RECT 33.97 38.78 34.33 39.14 ;
        RECT 33.97 37.21 34.33 37.57 ;
        RECT 33.97 29.11 34.33 29.47 ;
        RECT 33.97 27.54 34.33 27.9 ;
        RECT 33.97 25.97 34.33 26.33 ;
        RECT 33.97 17.87 34.33 18.23 ;
        RECT 33.97 16.3 34.33 16.66 ;
        RECT 33.97 14.73 34.33 15.09 ;
        RECT 34.67 90.92 35.03 91.28 ;
        RECT 34.67 90.11 35.03 90.47 ;
        RECT 34.67 89.3 35.03 89.66 ;
        RECT 34.67 88.49 35.03 88.85 ;
        RECT 34.67 87.68 35.03 88.04 ;
        RECT 34.67 79.68 35.03 80.04 ;
        RECT 34.67 78.87 35.03 79.23 ;
        RECT 34.67 78.06 35.03 78.42 ;
        RECT 34.67 77.25 35.03 77.61 ;
        RECT 34.67 76.44 35.03 76.8 ;
        RECT 34.67 68.44 35.03 68.8 ;
        RECT 34.67 67.63 35.03 67.99 ;
        RECT 34.67 66.82 35.03 67.18 ;
        RECT 34.67 66.01 35.03 66.37 ;
        RECT 34.67 65.2 35.03 65.56 ;
        RECT 34.67 57.2 35.03 57.56 ;
        RECT 34.67 56.39 35.03 56.75 ;
        RECT 34.67 55.58 35.03 55.94 ;
        RECT 34.67 54.77 35.03 55.13 ;
        RECT 34.67 53.96 35.03 54.32 ;
        RECT 34.67 45.96 35.03 46.32 ;
        RECT 34.67 45.15 35.03 45.51 ;
        RECT 34.67 44.34 35.03 44.7 ;
        RECT 34.67 43.53 35.03 43.89 ;
        RECT 34.67 42.72 35.03 43.08 ;
        RECT 34.67 34.72 35.03 35.08 ;
        RECT 34.67 33.91 35.03 34.27 ;
        RECT 34.67 33.1 35.03 33.46 ;
        RECT 34.67 32.29 35.03 32.65 ;
        RECT 34.67 31.48 35.03 31.84 ;
        RECT 34.67 23.48 35.03 23.84 ;
        RECT 34.67 22.67 35.03 23.03 ;
        RECT 34.67 21.86 35.03 22.22 ;
        RECT 34.67 21.05 35.03 21.41 ;
        RECT 34.67 20.24 35.03 20.6 ;
        RECT 34.67 12.24 35.03 12.6 ;
        RECT 34.67 11.43 35.03 11.79 ;
        RECT 34.67 10.62 35.03 10.98 ;
        RECT 34.67 9.81 35.03 10.17 ;
        RECT 34.67 9 35.03 9.36 ;
        RECT 34.78 85.31 35.14 85.67 ;
        RECT 34.78 83.74 35.14 84.1 ;
        RECT 34.78 82.17 35.14 82.53 ;
        RECT 34.78 74.07 35.14 74.43 ;
        RECT 34.78 72.5 35.14 72.86 ;
        RECT 34.78 70.93 35.14 71.29 ;
        RECT 34.78 62.83 35.14 63.19 ;
        RECT 34.78 61.26 35.14 61.62 ;
        RECT 34.78 59.69 35.14 60.05 ;
        RECT 34.78 51.59 35.14 51.95 ;
        RECT 34.78 50.02 35.14 50.38 ;
        RECT 34.78 48.45 35.14 48.81 ;
        RECT 34.78 40.35 35.14 40.71 ;
        RECT 34.78 38.78 35.14 39.14 ;
        RECT 34.78 37.21 35.14 37.57 ;
        RECT 34.78 29.11 35.14 29.47 ;
        RECT 34.78 27.54 35.14 27.9 ;
        RECT 34.78 25.97 35.14 26.33 ;
        RECT 34.78 17.87 35.14 18.23 ;
        RECT 34.78 16.3 35.14 16.66 ;
        RECT 34.78 14.73 35.14 15.09 ;
        RECT 37.1 90.93 37.46 91.29 ;
        RECT 37.1 89.36 37.46 89.72 ;
        RECT 37.1 87.79 37.46 88.15 ;
        RECT 37.1 79.69 37.46 80.05 ;
        RECT 37.1 78.12 37.46 78.48 ;
        RECT 37.1 76.55 37.46 76.91 ;
        RECT 37.1 68.45 37.46 68.81 ;
        RECT 37.1 66.88 37.46 67.24 ;
        RECT 37.1 65.31 37.46 65.67 ;
        RECT 37.1 57.21 37.46 57.57 ;
        RECT 37.1 55.64 37.46 56 ;
        RECT 37.1 54.07 37.46 54.43 ;
        RECT 37.1 45.97 37.46 46.33 ;
        RECT 37.1 44.4 37.46 44.76 ;
        RECT 37.1 42.83 37.46 43.19 ;
        RECT 37.1 34.73 37.46 35.09 ;
        RECT 37.1 33.16 37.46 33.52 ;
        RECT 37.1 31.59 37.46 31.95 ;
        RECT 37.1 23.49 37.46 23.85 ;
        RECT 37.1 21.92 37.46 22.28 ;
        RECT 37.1 20.35 37.46 20.71 ;
        RECT 37.1 12.25 37.46 12.61 ;
        RECT 37.1 10.68 37.46 11.04 ;
        RECT 37.1 9.11 37.46 9.47 ;
        RECT 37.21 85.3 37.57 85.66 ;
        RECT 37.21 84.49 37.57 84.85 ;
        RECT 37.21 83.68 37.57 84.04 ;
        RECT 37.21 82.87 37.57 83.23 ;
        RECT 37.21 82.06 37.57 82.42 ;
        RECT 37.21 74.06 37.57 74.42 ;
        RECT 37.21 73.25 37.57 73.61 ;
        RECT 37.21 72.44 37.57 72.8 ;
        RECT 37.21 71.63 37.57 71.99 ;
        RECT 37.21 70.82 37.57 71.18 ;
        RECT 37.21 62.82 37.57 63.18 ;
        RECT 37.21 62.01 37.57 62.37 ;
        RECT 37.21 61.2 37.57 61.56 ;
        RECT 37.21 60.39 37.57 60.75 ;
        RECT 37.21 59.58 37.57 59.94 ;
        RECT 37.21 51.58 37.57 51.94 ;
        RECT 37.21 50.77 37.57 51.13 ;
        RECT 37.21 49.96 37.57 50.32 ;
        RECT 37.21 49.15 37.57 49.51 ;
        RECT 37.21 48.34 37.57 48.7 ;
        RECT 37.21 40.34 37.57 40.7 ;
        RECT 37.21 39.53 37.57 39.89 ;
        RECT 37.21 38.72 37.57 39.08 ;
        RECT 37.21 37.91 37.57 38.27 ;
        RECT 37.21 37.1 37.57 37.46 ;
        RECT 37.21 29.1 37.57 29.46 ;
        RECT 37.21 28.29 37.57 28.65 ;
        RECT 37.21 27.48 37.57 27.84 ;
        RECT 37.21 26.67 37.57 27.03 ;
        RECT 37.21 25.86 37.57 26.22 ;
        RECT 37.21 17.86 37.57 18.22 ;
        RECT 37.21 17.05 37.57 17.41 ;
        RECT 37.21 16.24 37.57 16.6 ;
        RECT 37.21 15.43 37.57 15.79 ;
        RECT 37.21 14.62 37.57 14.98 ;
        RECT 37.91 90.93 38.27 91.29 ;
        RECT 37.91 89.36 38.27 89.72 ;
        RECT 37.91 87.79 38.27 88.15 ;
        RECT 37.91 79.69 38.27 80.05 ;
        RECT 37.91 78.12 38.27 78.48 ;
        RECT 37.91 76.55 38.27 76.91 ;
        RECT 37.91 68.45 38.27 68.81 ;
        RECT 37.91 66.88 38.27 67.24 ;
        RECT 37.91 65.31 38.27 65.67 ;
        RECT 37.91 57.21 38.27 57.57 ;
        RECT 37.91 55.64 38.27 56 ;
        RECT 37.91 54.07 38.27 54.43 ;
        RECT 37.91 45.97 38.27 46.33 ;
        RECT 37.91 44.4 38.27 44.76 ;
        RECT 37.91 42.83 38.27 43.19 ;
        RECT 37.91 34.73 38.27 35.09 ;
        RECT 37.91 33.16 38.27 33.52 ;
        RECT 37.91 31.59 38.27 31.95 ;
        RECT 37.91 23.49 38.27 23.85 ;
        RECT 37.91 21.92 38.27 22.28 ;
        RECT 37.91 20.35 38.27 20.71 ;
        RECT 37.91 12.25 38.27 12.61 ;
        RECT 37.91 10.68 38.27 11.04 ;
        RECT 37.91 9.11 38.27 9.47 ;
        RECT 38.72 90.93 39.08 91.29 ;
        RECT 38.72 89.36 39.08 89.72 ;
        RECT 38.72 87.79 39.08 88.15 ;
        RECT 38.72 79.69 39.08 80.05 ;
        RECT 38.72 78.12 39.08 78.48 ;
        RECT 38.72 76.55 39.08 76.91 ;
        RECT 38.72 68.45 39.08 68.81 ;
        RECT 38.72 66.88 39.08 67.24 ;
        RECT 38.72 65.31 39.08 65.67 ;
        RECT 38.72 57.21 39.08 57.57 ;
        RECT 38.72 55.64 39.08 56 ;
        RECT 38.72 54.07 39.08 54.43 ;
        RECT 38.72 45.97 39.08 46.33 ;
        RECT 38.72 44.4 39.08 44.76 ;
        RECT 38.72 42.83 39.08 43.19 ;
        RECT 38.72 34.73 39.08 35.09 ;
        RECT 38.72 33.16 39.08 33.52 ;
        RECT 38.72 31.59 39.08 31.95 ;
        RECT 38.72 23.49 39.08 23.85 ;
        RECT 38.72 21.92 39.08 22.28 ;
        RECT 38.72 20.35 39.08 20.71 ;
        RECT 38.72 12.25 39.08 12.61 ;
        RECT 38.72 10.68 39.08 11.04 ;
        RECT 38.72 9.11 39.08 9.47 ;
        RECT 38.78 85.3 39.14 85.66 ;
        RECT 38.78 84.49 39.14 84.85 ;
        RECT 38.78 83.68 39.14 84.04 ;
        RECT 38.78 82.87 39.14 83.23 ;
        RECT 38.78 82.06 39.14 82.42 ;
        RECT 38.78 74.06 39.14 74.42 ;
        RECT 38.78 73.25 39.14 73.61 ;
        RECT 38.78 72.44 39.14 72.8 ;
        RECT 38.78 71.63 39.14 71.99 ;
        RECT 38.78 70.82 39.14 71.18 ;
        RECT 38.78 62.82 39.14 63.18 ;
        RECT 38.78 62.01 39.14 62.37 ;
        RECT 38.78 61.2 39.14 61.56 ;
        RECT 38.78 60.39 39.14 60.75 ;
        RECT 38.78 59.58 39.14 59.94 ;
        RECT 38.78 51.58 39.14 51.94 ;
        RECT 38.78 50.77 39.14 51.13 ;
        RECT 38.78 49.96 39.14 50.32 ;
        RECT 38.78 49.15 39.14 49.51 ;
        RECT 38.78 48.34 39.14 48.7 ;
        RECT 38.78 40.34 39.14 40.7 ;
        RECT 38.78 39.53 39.14 39.89 ;
        RECT 38.78 38.72 39.14 39.08 ;
        RECT 38.78 37.91 39.14 38.27 ;
        RECT 38.78 37.1 39.14 37.46 ;
        RECT 38.78 29.1 39.14 29.46 ;
        RECT 38.78 28.29 39.14 28.65 ;
        RECT 38.78 27.48 39.14 27.84 ;
        RECT 38.78 26.67 39.14 27.03 ;
        RECT 38.78 25.86 39.14 26.22 ;
        RECT 38.78 17.86 39.14 18.22 ;
        RECT 38.78 17.05 39.14 17.41 ;
        RECT 38.78 16.24 39.14 16.6 ;
        RECT 38.78 15.43 39.14 15.79 ;
        RECT 38.78 14.62 39.14 14.98 ;
        RECT 39.53 90.93 39.89 91.29 ;
        RECT 39.53 89.36 39.89 89.72 ;
        RECT 39.53 87.79 39.89 88.15 ;
        RECT 39.53 79.69 39.89 80.05 ;
        RECT 39.53 78.12 39.89 78.48 ;
        RECT 39.53 76.55 39.89 76.91 ;
        RECT 39.53 68.45 39.89 68.81 ;
        RECT 39.53 66.88 39.89 67.24 ;
        RECT 39.53 65.31 39.89 65.67 ;
        RECT 39.53 57.21 39.89 57.57 ;
        RECT 39.53 55.64 39.89 56 ;
        RECT 39.53 54.07 39.89 54.43 ;
        RECT 39.53 45.97 39.89 46.33 ;
        RECT 39.53 44.4 39.89 44.76 ;
        RECT 39.53 42.83 39.89 43.19 ;
        RECT 39.53 34.73 39.89 35.09 ;
        RECT 39.53 33.16 39.89 33.52 ;
        RECT 39.53 31.59 39.89 31.95 ;
        RECT 39.53 23.49 39.89 23.85 ;
        RECT 39.53 21.92 39.89 22.28 ;
        RECT 39.53 20.35 39.89 20.71 ;
        RECT 39.53 12.25 39.89 12.61 ;
        RECT 39.53 10.68 39.89 11.04 ;
        RECT 39.53 9.11 39.89 9.47 ;
        RECT 40.34 90.93 40.7 91.29 ;
        RECT 40.34 89.36 40.7 89.72 ;
        RECT 40.34 87.79 40.7 88.15 ;
        RECT 40.34 79.69 40.7 80.05 ;
        RECT 40.34 78.12 40.7 78.48 ;
        RECT 40.34 76.55 40.7 76.91 ;
        RECT 40.34 68.45 40.7 68.81 ;
        RECT 40.34 66.88 40.7 67.24 ;
        RECT 40.34 65.31 40.7 65.67 ;
        RECT 40.34 57.21 40.7 57.57 ;
        RECT 40.34 55.64 40.7 56 ;
        RECT 40.34 54.07 40.7 54.43 ;
        RECT 40.34 45.97 40.7 46.33 ;
        RECT 40.34 44.4 40.7 44.76 ;
        RECT 40.34 42.83 40.7 43.19 ;
        RECT 40.34 34.73 40.7 35.09 ;
        RECT 40.34 33.16 40.7 33.52 ;
        RECT 40.34 31.59 40.7 31.95 ;
        RECT 40.34 23.49 40.7 23.85 ;
        RECT 40.34 21.92 40.7 22.28 ;
        RECT 40.34 20.35 40.7 20.71 ;
        RECT 40.34 12.25 40.7 12.61 ;
        RECT 40.34 10.68 40.7 11.04 ;
        RECT 40.34 9.11 40.7 9.47 ;
        RECT 40.35 85.3 40.71 85.66 ;
        RECT 40.35 84.49 40.71 84.85 ;
        RECT 40.35 83.68 40.71 84.04 ;
        RECT 40.35 82.87 40.71 83.23 ;
        RECT 40.35 82.06 40.71 82.42 ;
        RECT 40.35 74.06 40.71 74.42 ;
        RECT 40.35 73.25 40.71 73.61 ;
        RECT 40.35 72.44 40.71 72.8 ;
        RECT 40.35 71.63 40.71 71.99 ;
        RECT 40.35 70.82 40.71 71.18 ;
        RECT 40.35 62.82 40.71 63.18 ;
        RECT 40.35 62.01 40.71 62.37 ;
        RECT 40.35 61.2 40.71 61.56 ;
        RECT 40.35 60.39 40.71 60.75 ;
        RECT 40.35 59.58 40.71 59.94 ;
        RECT 40.35 51.58 40.71 51.94 ;
        RECT 40.35 50.77 40.71 51.13 ;
        RECT 40.35 49.96 40.71 50.32 ;
        RECT 40.35 49.15 40.71 49.51 ;
        RECT 40.35 48.34 40.71 48.7 ;
        RECT 40.35 40.34 40.71 40.7 ;
        RECT 40.35 39.53 40.71 39.89 ;
        RECT 40.35 38.72 40.71 39.08 ;
        RECT 40.35 37.91 40.71 38.27 ;
        RECT 40.35 37.1 40.71 37.46 ;
        RECT 40.35 29.1 40.71 29.46 ;
        RECT 40.35 28.29 40.71 28.65 ;
        RECT 40.35 27.48 40.71 27.84 ;
        RECT 40.35 26.67 40.71 27.03 ;
        RECT 40.35 25.86 40.71 26.22 ;
        RECT 40.35 17.86 40.71 18.22 ;
        RECT 40.35 17.05 40.71 17.41 ;
        RECT 40.35 16.24 40.71 16.6 ;
        RECT 40.35 15.43 40.71 15.79 ;
        RECT 40.35 14.62 40.71 14.98 ;
        RECT 42.77 90.92 43.13 91.28 ;
        RECT 42.77 90.11 43.13 90.47 ;
        RECT 42.77 89.3 43.13 89.66 ;
        RECT 42.77 88.49 43.13 88.85 ;
        RECT 42.77 87.68 43.13 88.04 ;
        RECT 42.77 79.68 43.13 80.04 ;
        RECT 42.77 78.87 43.13 79.23 ;
        RECT 42.77 78.06 43.13 78.42 ;
        RECT 42.77 77.25 43.13 77.61 ;
        RECT 42.77 76.44 43.13 76.8 ;
        RECT 42.77 68.44 43.13 68.8 ;
        RECT 42.77 67.63 43.13 67.99 ;
        RECT 42.77 66.82 43.13 67.18 ;
        RECT 42.77 66.01 43.13 66.37 ;
        RECT 42.77 65.2 43.13 65.56 ;
        RECT 42.77 57.2 43.13 57.56 ;
        RECT 42.77 56.39 43.13 56.75 ;
        RECT 42.77 55.58 43.13 55.94 ;
        RECT 42.77 54.77 43.13 55.13 ;
        RECT 42.77 53.96 43.13 54.32 ;
        RECT 42.77 45.96 43.13 46.32 ;
        RECT 42.77 45.15 43.13 45.51 ;
        RECT 42.77 44.34 43.13 44.7 ;
        RECT 42.77 43.53 43.13 43.89 ;
        RECT 42.77 42.72 43.13 43.08 ;
        RECT 42.77 34.72 43.13 35.08 ;
        RECT 42.77 33.91 43.13 34.27 ;
        RECT 42.77 33.1 43.13 33.46 ;
        RECT 42.77 32.29 43.13 32.65 ;
        RECT 42.77 31.48 43.13 31.84 ;
        RECT 42.77 23.48 43.13 23.84 ;
        RECT 42.77 22.67 43.13 23.03 ;
        RECT 42.77 21.86 43.13 22.22 ;
        RECT 42.77 21.05 43.13 21.41 ;
        RECT 42.77 20.24 43.13 20.6 ;
        RECT 42.77 12.24 43.13 12.6 ;
        RECT 42.77 11.43 43.13 11.79 ;
        RECT 42.77 10.62 43.13 10.98 ;
        RECT 42.77 9.81 43.13 10.17 ;
        RECT 42.77 9 43.13 9.36 ;
        RECT 42.78 85.31 43.14 85.67 ;
        RECT 42.78 83.74 43.14 84.1 ;
        RECT 42.78 82.17 43.14 82.53 ;
        RECT 42.78 74.07 43.14 74.43 ;
        RECT 42.78 72.5 43.14 72.86 ;
        RECT 42.78 70.93 43.14 71.29 ;
        RECT 42.78 62.83 43.14 63.19 ;
        RECT 42.78 61.26 43.14 61.62 ;
        RECT 42.78 59.69 43.14 60.05 ;
        RECT 42.78 51.59 43.14 51.95 ;
        RECT 42.78 50.02 43.14 50.38 ;
        RECT 42.78 48.45 43.14 48.81 ;
        RECT 42.78 40.35 43.14 40.71 ;
        RECT 42.78 38.78 43.14 39.14 ;
        RECT 42.78 37.21 43.14 37.57 ;
        RECT 42.78 29.11 43.14 29.47 ;
        RECT 42.78 27.54 43.14 27.9 ;
        RECT 42.78 25.97 43.14 26.33 ;
        RECT 42.78 17.87 43.14 18.23 ;
        RECT 42.78 16.3 43.14 16.66 ;
        RECT 42.78 14.73 43.14 15.09 ;
        RECT 43.59 85.31 43.95 85.67 ;
        RECT 43.59 83.74 43.95 84.1 ;
        RECT 43.59 82.17 43.95 82.53 ;
        RECT 43.59 74.07 43.95 74.43 ;
        RECT 43.59 72.5 43.95 72.86 ;
        RECT 43.59 70.93 43.95 71.29 ;
        RECT 43.59 62.83 43.95 63.19 ;
        RECT 43.59 61.26 43.95 61.62 ;
        RECT 43.59 59.69 43.95 60.05 ;
        RECT 43.59 51.59 43.95 51.95 ;
        RECT 43.59 50.02 43.95 50.38 ;
        RECT 43.59 48.45 43.95 48.81 ;
        RECT 43.59 40.35 43.95 40.71 ;
        RECT 43.59 38.78 43.95 39.14 ;
        RECT 43.59 37.21 43.95 37.57 ;
        RECT 43.59 29.11 43.95 29.47 ;
        RECT 43.59 27.54 43.95 27.9 ;
        RECT 43.59 25.97 43.95 26.33 ;
        RECT 43.59 17.87 43.95 18.23 ;
        RECT 43.59 16.3 43.95 16.66 ;
        RECT 43.59 14.73 43.95 15.09 ;
        RECT 44.34 90.92 44.7 91.28 ;
        RECT 44.34 90.11 44.7 90.47 ;
        RECT 44.34 89.3 44.7 89.66 ;
        RECT 44.34 88.49 44.7 88.85 ;
        RECT 44.34 87.68 44.7 88.04 ;
        RECT 44.34 79.68 44.7 80.04 ;
        RECT 44.34 78.87 44.7 79.23 ;
        RECT 44.34 78.06 44.7 78.42 ;
        RECT 44.34 77.25 44.7 77.61 ;
        RECT 44.34 76.44 44.7 76.8 ;
        RECT 44.34 68.44 44.7 68.8 ;
        RECT 44.34 67.63 44.7 67.99 ;
        RECT 44.34 66.82 44.7 67.18 ;
        RECT 44.34 66.01 44.7 66.37 ;
        RECT 44.34 65.2 44.7 65.56 ;
        RECT 44.34 57.2 44.7 57.56 ;
        RECT 44.34 56.39 44.7 56.75 ;
        RECT 44.34 55.58 44.7 55.94 ;
        RECT 44.34 54.77 44.7 55.13 ;
        RECT 44.34 53.96 44.7 54.32 ;
        RECT 44.34 45.96 44.7 46.32 ;
        RECT 44.34 45.15 44.7 45.51 ;
        RECT 44.34 44.34 44.7 44.7 ;
        RECT 44.34 43.53 44.7 43.89 ;
        RECT 44.34 42.72 44.7 43.08 ;
        RECT 44.34 34.72 44.7 35.08 ;
        RECT 44.34 33.91 44.7 34.27 ;
        RECT 44.34 33.1 44.7 33.46 ;
        RECT 44.34 32.29 44.7 32.65 ;
        RECT 44.34 31.48 44.7 31.84 ;
        RECT 44.34 23.48 44.7 23.84 ;
        RECT 44.34 22.67 44.7 23.03 ;
        RECT 44.34 21.86 44.7 22.22 ;
        RECT 44.34 21.05 44.7 21.41 ;
        RECT 44.34 20.24 44.7 20.6 ;
        RECT 44.34 12.24 44.7 12.6 ;
        RECT 44.34 11.43 44.7 11.79 ;
        RECT 44.34 10.62 44.7 10.98 ;
        RECT 44.34 9.81 44.7 10.17 ;
        RECT 44.34 9 44.7 9.36 ;
        RECT 44.4 85.31 44.76 85.67 ;
        RECT 44.4 83.74 44.76 84.1 ;
        RECT 44.4 82.17 44.76 82.53 ;
        RECT 44.4 74.07 44.76 74.43 ;
        RECT 44.4 72.5 44.76 72.86 ;
        RECT 44.4 70.93 44.76 71.29 ;
        RECT 44.4 62.83 44.76 63.19 ;
        RECT 44.4 61.26 44.76 61.62 ;
        RECT 44.4 59.69 44.76 60.05 ;
        RECT 44.4 51.59 44.76 51.95 ;
        RECT 44.4 50.02 44.76 50.38 ;
        RECT 44.4 48.45 44.76 48.81 ;
        RECT 44.4 40.35 44.76 40.71 ;
        RECT 44.4 38.78 44.76 39.14 ;
        RECT 44.4 37.21 44.76 37.57 ;
        RECT 44.4 29.11 44.76 29.47 ;
        RECT 44.4 27.54 44.76 27.9 ;
        RECT 44.4 25.97 44.76 26.33 ;
        RECT 44.4 17.87 44.76 18.23 ;
        RECT 44.4 16.3 44.76 16.66 ;
        RECT 44.4 14.73 44.76 15.09 ;
        RECT 45.21 85.31 45.57 85.67 ;
        RECT 45.21 83.74 45.57 84.1 ;
        RECT 45.21 82.17 45.57 82.53 ;
        RECT 45.21 74.07 45.57 74.43 ;
        RECT 45.21 72.5 45.57 72.86 ;
        RECT 45.21 70.93 45.57 71.29 ;
        RECT 45.21 62.83 45.57 63.19 ;
        RECT 45.21 61.26 45.57 61.62 ;
        RECT 45.21 59.69 45.57 60.05 ;
        RECT 45.21 51.59 45.57 51.95 ;
        RECT 45.21 50.02 45.57 50.38 ;
        RECT 45.21 48.45 45.57 48.81 ;
        RECT 45.21 40.35 45.57 40.71 ;
        RECT 45.21 38.78 45.57 39.14 ;
        RECT 45.21 37.21 45.57 37.57 ;
        RECT 45.21 29.11 45.57 29.47 ;
        RECT 45.21 27.54 45.57 27.9 ;
        RECT 45.21 25.97 45.57 26.33 ;
        RECT 45.21 17.87 45.57 18.23 ;
        RECT 45.21 16.3 45.57 16.66 ;
        RECT 45.21 14.73 45.57 15.09 ;
        RECT 45.91 90.92 46.27 91.28 ;
        RECT 45.91 90.11 46.27 90.47 ;
        RECT 45.91 89.3 46.27 89.66 ;
        RECT 45.91 88.49 46.27 88.85 ;
        RECT 45.91 87.68 46.27 88.04 ;
        RECT 45.91 79.68 46.27 80.04 ;
        RECT 45.91 78.87 46.27 79.23 ;
        RECT 45.91 78.06 46.27 78.42 ;
        RECT 45.91 77.25 46.27 77.61 ;
        RECT 45.91 76.44 46.27 76.8 ;
        RECT 45.91 68.44 46.27 68.8 ;
        RECT 45.91 67.63 46.27 67.99 ;
        RECT 45.91 66.82 46.27 67.18 ;
        RECT 45.91 66.01 46.27 66.37 ;
        RECT 45.91 65.2 46.27 65.56 ;
        RECT 45.91 57.2 46.27 57.56 ;
        RECT 45.91 56.39 46.27 56.75 ;
        RECT 45.91 55.58 46.27 55.94 ;
        RECT 45.91 54.77 46.27 55.13 ;
        RECT 45.91 53.96 46.27 54.32 ;
        RECT 45.91 45.96 46.27 46.32 ;
        RECT 45.91 45.15 46.27 45.51 ;
        RECT 45.91 44.34 46.27 44.7 ;
        RECT 45.91 43.53 46.27 43.89 ;
        RECT 45.91 42.72 46.27 43.08 ;
        RECT 45.91 34.72 46.27 35.08 ;
        RECT 45.91 33.91 46.27 34.27 ;
        RECT 45.91 33.1 46.27 33.46 ;
        RECT 45.91 32.29 46.27 32.65 ;
        RECT 45.91 31.48 46.27 31.84 ;
        RECT 45.91 23.48 46.27 23.84 ;
        RECT 45.91 22.67 46.27 23.03 ;
        RECT 45.91 21.86 46.27 22.22 ;
        RECT 45.91 21.05 46.27 21.41 ;
        RECT 45.91 20.24 46.27 20.6 ;
        RECT 45.91 12.24 46.27 12.6 ;
        RECT 45.91 11.43 46.27 11.79 ;
        RECT 45.91 10.62 46.27 10.98 ;
        RECT 45.91 9.81 46.27 10.17 ;
        RECT 45.91 9 46.27 9.36 ;
        RECT 46.02 85.31 46.38 85.67 ;
        RECT 46.02 83.74 46.38 84.1 ;
        RECT 46.02 82.17 46.38 82.53 ;
        RECT 46.02 74.07 46.38 74.43 ;
        RECT 46.02 72.5 46.38 72.86 ;
        RECT 46.02 70.93 46.38 71.29 ;
        RECT 46.02 62.83 46.38 63.19 ;
        RECT 46.02 61.26 46.38 61.62 ;
        RECT 46.02 59.69 46.38 60.05 ;
        RECT 46.02 51.59 46.38 51.95 ;
        RECT 46.02 50.02 46.38 50.38 ;
        RECT 46.02 48.45 46.38 48.81 ;
        RECT 46.02 40.35 46.38 40.71 ;
        RECT 46.02 38.78 46.38 39.14 ;
        RECT 46.02 37.21 46.38 37.57 ;
        RECT 46.02 29.11 46.38 29.47 ;
        RECT 46.02 27.54 46.38 27.9 ;
        RECT 46.02 25.97 46.38 26.33 ;
        RECT 46.02 17.87 46.38 18.23 ;
        RECT 46.02 16.3 46.38 16.66 ;
        RECT 46.02 14.73 46.38 15.09 ;
        RECT 48.34 90.93 48.7 91.29 ;
        RECT 48.34 89.36 48.7 89.72 ;
        RECT 48.34 87.79 48.7 88.15 ;
        RECT 48.34 79.69 48.7 80.05 ;
        RECT 48.34 78.12 48.7 78.48 ;
        RECT 48.34 76.55 48.7 76.91 ;
        RECT 48.34 68.45 48.7 68.81 ;
        RECT 48.34 66.88 48.7 67.24 ;
        RECT 48.34 65.31 48.7 65.67 ;
        RECT 48.34 57.21 48.7 57.57 ;
        RECT 48.34 55.64 48.7 56 ;
        RECT 48.34 54.07 48.7 54.43 ;
        RECT 48.34 45.97 48.7 46.33 ;
        RECT 48.34 44.4 48.7 44.76 ;
        RECT 48.34 42.83 48.7 43.19 ;
        RECT 48.34 34.73 48.7 35.09 ;
        RECT 48.34 33.16 48.7 33.52 ;
        RECT 48.34 31.59 48.7 31.95 ;
        RECT 48.34 23.49 48.7 23.85 ;
        RECT 48.34 21.92 48.7 22.28 ;
        RECT 48.34 20.35 48.7 20.71 ;
        RECT 48.34 12.25 48.7 12.61 ;
        RECT 48.34 10.68 48.7 11.04 ;
        RECT 48.34 9.11 48.7 9.47 ;
        RECT 48.45 85.3 48.81 85.66 ;
        RECT 48.45 84.49 48.81 84.85 ;
        RECT 48.45 83.68 48.81 84.04 ;
        RECT 48.45 82.87 48.81 83.23 ;
        RECT 48.45 82.06 48.81 82.42 ;
        RECT 48.45 74.06 48.81 74.42 ;
        RECT 48.45 73.25 48.81 73.61 ;
        RECT 48.45 72.44 48.81 72.8 ;
        RECT 48.45 71.63 48.81 71.99 ;
        RECT 48.45 70.82 48.81 71.18 ;
        RECT 48.45 62.82 48.81 63.18 ;
        RECT 48.45 62.01 48.81 62.37 ;
        RECT 48.45 61.2 48.81 61.56 ;
        RECT 48.45 60.39 48.81 60.75 ;
        RECT 48.45 59.58 48.81 59.94 ;
        RECT 48.45 51.58 48.81 51.94 ;
        RECT 48.45 50.77 48.81 51.13 ;
        RECT 48.45 49.96 48.81 50.32 ;
        RECT 48.45 49.15 48.81 49.51 ;
        RECT 48.45 48.34 48.81 48.7 ;
        RECT 48.45 40.34 48.81 40.7 ;
        RECT 48.45 39.53 48.81 39.89 ;
        RECT 48.45 38.72 48.81 39.08 ;
        RECT 48.45 37.91 48.81 38.27 ;
        RECT 48.45 37.1 48.81 37.46 ;
        RECT 48.45 29.1 48.81 29.46 ;
        RECT 48.45 28.29 48.81 28.65 ;
        RECT 48.45 27.48 48.81 27.84 ;
        RECT 48.45 26.67 48.81 27.03 ;
        RECT 48.45 25.86 48.81 26.22 ;
        RECT 48.45 17.86 48.81 18.22 ;
        RECT 48.45 17.05 48.81 17.41 ;
        RECT 48.45 16.24 48.81 16.6 ;
        RECT 48.45 15.43 48.81 15.79 ;
        RECT 48.45 14.62 48.81 14.98 ;
        RECT 49.15 90.93 49.51 91.29 ;
        RECT 49.15 89.36 49.51 89.72 ;
        RECT 49.15 87.79 49.51 88.15 ;
        RECT 49.15 79.69 49.51 80.05 ;
        RECT 49.15 78.12 49.51 78.48 ;
        RECT 49.15 76.55 49.51 76.91 ;
        RECT 49.15 68.45 49.51 68.81 ;
        RECT 49.15 66.88 49.51 67.24 ;
        RECT 49.15 65.31 49.51 65.67 ;
        RECT 49.15 57.21 49.51 57.57 ;
        RECT 49.15 55.64 49.51 56 ;
        RECT 49.15 54.07 49.51 54.43 ;
        RECT 49.15 45.97 49.51 46.33 ;
        RECT 49.15 44.4 49.51 44.76 ;
        RECT 49.15 42.83 49.51 43.19 ;
        RECT 49.15 34.73 49.51 35.09 ;
        RECT 49.15 33.16 49.51 33.52 ;
        RECT 49.15 31.59 49.51 31.95 ;
        RECT 49.15 23.49 49.51 23.85 ;
        RECT 49.15 21.92 49.51 22.28 ;
        RECT 49.15 20.35 49.51 20.71 ;
        RECT 49.15 12.25 49.51 12.61 ;
        RECT 49.15 10.68 49.51 11.04 ;
        RECT 49.15 9.11 49.51 9.47 ;
        RECT 49.96 90.93 50.32 91.29 ;
        RECT 49.96 89.36 50.32 89.72 ;
        RECT 49.96 87.79 50.32 88.15 ;
        RECT 49.96 79.69 50.32 80.05 ;
        RECT 49.96 78.12 50.32 78.48 ;
        RECT 49.96 76.55 50.32 76.91 ;
        RECT 49.96 68.45 50.32 68.81 ;
        RECT 49.96 66.88 50.32 67.24 ;
        RECT 49.96 65.31 50.32 65.67 ;
        RECT 49.96 57.21 50.32 57.57 ;
        RECT 49.96 55.64 50.32 56 ;
        RECT 49.96 54.07 50.32 54.43 ;
        RECT 49.96 45.97 50.32 46.33 ;
        RECT 49.96 44.4 50.32 44.76 ;
        RECT 49.96 42.83 50.32 43.19 ;
        RECT 49.96 34.73 50.32 35.09 ;
        RECT 49.96 33.16 50.32 33.52 ;
        RECT 49.96 31.59 50.32 31.95 ;
        RECT 49.96 23.49 50.32 23.85 ;
        RECT 49.96 21.92 50.32 22.28 ;
        RECT 49.96 20.35 50.32 20.71 ;
        RECT 49.96 12.25 50.32 12.61 ;
        RECT 49.96 10.68 50.32 11.04 ;
        RECT 49.96 9.11 50.32 9.47 ;
        RECT 50.02 85.3 50.38 85.66 ;
        RECT 50.02 84.49 50.38 84.85 ;
        RECT 50.02 83.68 50.38 84.04 ;
        RECT 50.02 82.87 50.38 83.23 ;
        RECT 50.02 82.06 50.38 82.42 ;
        RECT 50.02 74.06 50.38 74.42 ;
        RECT 50.02 73.25 50.38 73.61 ;
        RECT 50.02 72.44 50.38 72.8 ;
        RECT 50.02 71.63 50.38 71.99 ;
        RECT 50.02 70.82 50.38 71.18 ;
        RECT 50.02 62.82 50.38 63.18 ;
        RECT 50.02 62.01 50.38 62.37 ;
        RECT 50.02 61.2 50.38 61.56 ;
        RECT 50.02 60.39 50.38 60.75 ;
        RECT 50.02 59.58 50.38 59.94 ;
        RECT 50.02 51.58 50.38 51.94 ;
        RECT 50.02 50.77 50.38 51.13 ;
        RECT 50.02 49.96 50.38 50.32 ;
        RECT 50.02 49.15 50.38 49.51 ;
        RECT 50.02 48.34 50.38 48.7 ;
        RECT 50.02 40.34 50.38 40.7 ;
        RECT 50.02 39.53 50.38 39.89 ;
        RECT 50.02 38.72 50.38 39.08 ;
        RECT 50.02 37.91 50.38 38.27 ;
        RECT 50.02 37.1 50.38 37.46 ;
        RECT 50.02 29.1 50.38 29.46 ;
        RECT 50.02 28.29 50.38 28.65 ;
        RECT 50.02 27.48 50.38 27.84 ;
        RECT 50.02 26.67 50.38 27.03 ;
        RECT 50.02 25.86 50.38 26.22 ;
        RECT 50.02 17.86 50.38 18.22 ;
        RECT 50.02 17.05 50.38 17.41 ;
        RECT 50.02 16.24 50.38 16.6 ;
        RECT 50.02 15.43 50.38 15.79 ;
        RECT 50.02 14.62 50.38 14.98 ;
        RECT 50.77 90.93 51.13 91.29 ;
        RECT 50.77 89.36 51.13 89.72 ;
        RECT 50.77 87.79 51.13 88.15 ;
        RECT 50.77 79.69 51.13 80.05 ;
        RECT 50.77 78.12 51.13 78.48 ;
        RECT 50.77 76.55 51.13 76.91 ;
        RECT 50.77 68.45 51.13 68.81 ;
        RECT 50.77 66.88 51.13 67.24 ;
        RECT 50.77 65.31 51.13 65.67 ;
        RECT 50.77 57.21 51.13 57.57 ;
        RECT 50.77 55.64 51.13 56 ;
        RECT 50.77 54.07 51.13 54.43 ;
        RECT 50.77 45.97 51.13 46.33 ;
        RECT 50.77 44.4 51.13 44.76 ;
        RECT 50.77 42.83 51.13 43.19 ;
        RECT 50.77 34.73 51.13 35.09 ;
        RECT 50.77 33.16 51.13 33.52 ;
        RECT 50.77 31.59 51.13 31.95 ;
        RECT 50.77 23.49 51.13 23.85 ;
        RECT 50.77 21.92 51.13 22.28 ;
        RECT 50.77 20.35 51.13 20.71 ;
        RECT 50.77 12.25 51.13 12.61 ;
        RECT 50.77 10.68 51.13 11.04 ;
        RECT 50.77 9.11 51.13 9.47 ;
        RECT 51.58 90.93 51.94 91.29 ;
        RECT 51.58 89.36 51.94 89.72 ;
        RECT 51.58 87.79 51.94 88.15 ;
        RECT 51.58 79.69 51.94 80.05 ;
        RECT 51.58 78.12 51.94 78.48 ;
        RECT 51.58 76.55 51.94 76.91 ;
        RECT 51.58 68.45 51.94 68.81 ;
        RECT 51.58 66.88 51.94 67.24 ;
        RECT 51.58 65.31 51.94 65.67 ;
        RECT 51.58 57.21 51.94 57.57 ;
        RECT 51.58 55.64 51.94 56 ;
        RECT 51.58 54.07 51.94 54.43 ;
        RECT 51.58 45.97 51.94 46.33 ;
        RECT 51.58 44.4 51.94 44.76 ;
        RECT 51.58 42.83 51.94 43.19 ;
        RECT 51.58 34.73 51.94 35.09 ;
        RECT 51.58 33.16 51.94 33.52 ;
        RECT 51.58 31.59 51.94 31.95 ;
        RECT 51.58 23.49 51.94 23.85 ;
        RECT 51.58 21.92 51.94 22.28 ;
        RECT 51.58 20.35 51.94 20.71 ;
        RECT 51.58 12.25 51.94 12.61 ;
        RECT 51.58 10.68 51.94 11.04 ;
        RECT 51.58 9.11 51.94 9.47 ;
        RECT 51.59 85.3 51.95 85.66 ;
        RECT 51.59 84.49 51.95 84.85 ;
        RECT 51.59 83.68 51.95 84.04 ;
        RECT 51.59 82.87 51.95 83.23 ;
        RECT 51.59 82.06 51.95 82.42 ;
        RECT 51.59 74.06 51.95 74.42 ;
        RECT 51.59 73.25 51.95 73.61 ;
        RECT 51.59 72.44 51.95 72.8 ;
        RECT 51.59 71.63 51.95 71.99 ;
        RECT 51.59 70.82 51.95 71.18 ;
        RECT 51.59 62.82 51.95 63.18 ;
        RECT 51.59 62.01 51.95 62.37 ;
        RECT 51.59 61.2 51.95 61.56 ;
        RECT 51.59 60.39 51.95 60.75 ;
        RECT 51.59 59.58 51.95 59.94 ;
        RECT 51.59 51.58 51.95 51.94 ;
        RECT 51.59 50.77 51.95 51.13 ;
        RECT 51.59 49.96 51.95 50.32 ;
        RECT 51.59 49.15 51.95 49.51 ;
        RECT 51.59 48.34 51.95 48.7 ;
        RECT 51.59 40.34 51.95 40.7 ;
        RECT 51.59 39.53 51.95 39.89 ;
        RECT 51.59 38.72 51.95 39.08 ;
        RECT 51.59 37.91 51.95 38.27 ;
        RECT 51.59 37.1 51.95 37.46 ;
        RECT 51.59 29.1 51.95 29.46 ;
        RECT 51.59 28.29 51.95 28.65 ;
        RECT 51.59 27.48 51.95 27.84 ;
        RECT 51.59 26.67 51.95 27.03 ;
        RECT 51.59 25.86 51.95 26.22 ;
        RECT 51.59 17.86 51.95 18.22 ;
        RECT 51.59 17.05 51.95 17.41 ;
        RECT 51.59 16.24 51.95 16.6 ;
        RECT 51.59 15.43 51.95 15.79 ;
        RECT 51.59 14.62 51.95 14.98 ;
        RECT 54.01 90.92 54.37 91.28 ;
        RECT 54.01 90.11 54.37 90.47 ;
        RECT 54.01 89.3 54.37 89.66 ;
        RECT 54.01 88.49 54.37 88.85 ;
        RECT 54.01 87.68 54.37 88.04 ;
        RECT 54.01 79.68 54.37 80.04 ;
        RECT 54.01 78.87 54.37 79.23 ;
        RECT 54.01 78.06 54.37 78.42 ;
        RECT 54.01 77.25 54.37 77.61 ;
        RECT 54.01 76.44 54.37 76.8 ;
        RECT 54.01 68.44 54.37 68.8 ;
        RECT 54.01 67.63 54.37 67.99 ;
        RECT 54.01 66.82 54.37 67.18 ;
        RECT 54.01 66.01 54.37 66.37 ;
        RECT 54.01 65.2 54.37 65.56 ;
        RECT 54.01 57.2 54.37 57.56 ;
        RECT 54.01 56.39 54.37 56.75 ;
        RECT 54.01 55.58 54.37 55.94 ;
        RECT 54.01 54.77 54.37 55.13 ;
        RECT 54.01 53.96 54.37 54.32 ;
        RECT 54.01 45.96 54.37 46.32 ;
        RECT 54.01 45.15 54.37 45.51 ;
        RECT 54.01 44.34 54.37 44.7 ;
        RECT 54.01 43.53 54.37 43.89 ;
        RECT 54.01 42.72 54.37 43.08 ;
        RECT 54.01 34.72 54.37 35.08 ;
        RECT 54.01 33.91 54.37 34.27 ;
        RECT 54.01 33.1 54.37 33.46 ;
        RECT 54.01 32.29 54.37 32.65 ;
        RECT 54.01 31.48 54.37 31.84 ;
        RECT 54.01 23.48 54.37 23.84 ;
        RECT 54.01 22.67 54.37 23.03 ;
        RECT 54.01 21.86 54.37 22.22 ;
        RECT 54.01 21.05 54.37 21.41 ;
        RECT 54.01 20.24 54.37 20.6 ;
        RECT 54.01 12.24 54.37 12.6 ;
        RECT 54.01 11.43 54.37 11.79 ;
        RECT 54.01 10.62 54.37 10.98 ;
        RECT 54.01 9.81 54.37 10.17 ;
        RECT 54.01 9 54.37 9.36 ;
        RECT 54.02 85.31 54.38 85.67 ;
        RECT 54.02 83.74 54.38 84.1 ;
        RECT 54.02 82.17 54.38 82.53 ;
        RECT 54.02 74.07 54.38 74.43 ;
        RECT 54.02 72.5 54.38 72.86 ;
        RECT 54.02 70.93 54.38 71.29 ;
        RECT 54.02 62.83 54.38 63.19 ;
        RECT 54.02 61.26 54.38 61.62 ;
        RECT 54.02 59.69 54.38 60.05 ;
        RECT 54.02 51.59 54.38 51.95 ;
        RECT 54.02 50.02 54.38 50.38 ;
        RECT 54.02 48.45 54.38 48.81 ;
        RECT 54.02 40.35 54.38 40.71 ;
        RECT 54.02 38.78 54.38 39.14 ;
        RECT 54.02 37.21 54.38 37.57 ;
        RECT 54.02 29.11 54.38 29.47 ;
        RECT 54.02 27.54 54.38 27.9 ;
        RECT 54.02 25.97 54.38 26.33 ;
        RECT 54.02 17.87 54.38 18.23 ;
        RECT 54.02 16.3 54.38 16.66 ;
        RECT 54.02 14.73 54.38 15.09 ;
        RECT 54.83 85.31 55.19 85.67 ;
        RECT 54.83 83.74 55.19 84.1 ;
        RECT 54.83 82.17 55.19 82.53 ;
        RECT 54.83 74.07 55.19 74.43 ;
        RECT 54.83 72.5 55.19 72.86 ;
        RECT 54.83 70.93 55.19 71.29 ;
        RECT 54.83 62.83 55.19 63.19 ;
        RECT 54.83 61.26 55.19 61.62 ;
        RECT 54.83 59.69 55.19 60.05 ;
        RECT 54.83 51.59 55.19 51.95 ;
        RECT 54.83 50.02 55.19 50.38 ;
        RECT 54.83 48.45 55.19 48.81 ;
        RECT 54.83 40.35 55.19 40.71 ;
        RECT 54.83 38.78 55.19 39.14 ;
        RECT 54.83 37.21 55.19 37.57 ;
        RECT 54.83 29.11 55.19 29.47 ;
        RECT 54.83 27.54 55.19 27.9 ;
        RECT 54.83 25.97 55.19 26.33 ;
        RECT 54.83 17.87 55.19 18.23 ;
        RECT 54.83 16.3 55.19 16.66 ;
        RECT 54.83 14.73 55.19 15.09 ;
        RECT 55.58 90.92 55.94 91.28 ;
        RECT 55.58 90.11 55.94 90.47 ;
        RECT 55.58 89.3 55.94 89.66 ;
        RECT 55.58 88.49 55.94 88.85 ;
        RECT 55.58 87.68 55.94 88.04 ;
        RECT 55.58 79.68 55.94 80.04 ;
        RECT 55.58 78.87 55.94 79.23 ;
        RECT 55.58 78.06 55.94 78.42 ;
        RECT 55.58 77.25 55.94 77.61 ;
        RECT 55.58 76.44 55.94 76.8 ;
        RECT 55.58 68.44 55.94 68.8 ;
        RECT 55.58 67.63 55.94 67.99 ;
        RECT 55.58 66.82 55.94 67.18 ;
        RECT 55.58 66.01 55.94 66.37 ;
        RECT 55.58 65.2 55.94 65.56 ;
        RECT 55.58 57.2 55.94 57.56 ;
        RECT 55.58 56.39 55.94 56.75 ;
        RECT 55.58 55.58 55.94 55.94 ;
        RECT 55.58 54.77 55.94 55.13 ;
        RECT 55.58 53.96 55.94 54.32 ;
        RECT 55.58 45.96 55.94 46.32 ;
        RECT 55.58 45.15 55.94 45.51 ;
        RECT 55.58 44.34 55.94 44.7 ;
        RECT 55.58 43.53 55.94 43.89 ;
        RECT 55.58 42.72 55.94 43.08 ;
        RECT 55.58 34.72 55.94 35.08 ;
        RECT 55.58 33.91 55.94 34.27 ;
        RECT 55.58 33.1 55.94 33.46 ;
        RECT 55.58 32.29 55.94 32.65 ;
        RECT 55.58 31.48 55.94 31.84 ;
        RECT 55.58 23.48 55.94 23.84 ;
        RECT 55.58 22.67 55.94 23.03 ;
        RECT 55.58 21.86 55.94 22.22 ;
        RECT 55.58 21.05 55.94 21.41 ;
        RECT 55.58 20.24 55.94 20.6 ;
        RECT 55.58 12.24 55.94 12.6 ;
        RECT 55.58 11.43 55.94 11.79 ;
        RECT 55.58 10.62 55.94 10.98 ;
        RECT 55.58 9.81 55.94 10.17 ;
        RECT 55.58 9 55.94 9.36 ;
        RECT 55.64 85.31 56 85.67 ;
        RECT 55.64 83.74 56 84.1 ;
        RECT 55.64 82.17 56 82.53 ;
        RECT 55.64 74.07 56 74.43 ;
        RECT 55.64 72.5 56 72.86 ;
        RECT 55.64 70.93 56 71.29 ;
        RECT 55.64 62.83 56 63.19 ;
        RECT 55.64 61.26 56 61.62 ;
        RECT 55.64 59.69 56 60.05 ;
        RECT 55.64 51.59 56 51.95 ;
        RECT 55.64 50.02 56 50.38 ;
        RECT 55.64 48.45 56 48.81 ;
        RECT 55.64 40.35 56 40.71 ;
        RECT 55.64 38.78 56 39.14 ;
        RECT 55.64 37.21 56 37.57 ;
        RECT 55.64 29.11 56 29.47 ;
        RECT 55.64 27.54 56 27.9 ;
        RECT 55.64 25.97 56 26.33 ;
        RECT 55.64 17.87 56 18.23 ;
        RECT 55.64 16.3 56 16.66 ;
        RECT 55.64 14.73 56 15.09 ;
        RECT 56.45 85.31 56.81 85.67 ;
        RECT 56.45 83.74 56.81 84.1 ;
        RECT 56.45 82.17 56.81 82.53 ;
        RECT 56.45 74.07 56.81 74.43 ;
        RECT 56.45 72.5 56.81 72.86 ;
        RECT 56.45 70.93 56.81 71.29 ;
        RECT 56.45 62.83 56.81 63.19 ;
        RECT 56.45 61.26 56.81 61.62 ;
        RECT 56.45 59.69 56.81 60.05 ;
        RECT 56.45 51.59 56.81 51.95 ;
        RECT 56.45 50.02 56.81 50.38 ;
        RECT 56.45 48.45 56.81 48.81 ;
        RECT 56.45 40.35 56.81 40.71 ;
        RECT 56.45 38.78 56.81 39.14 ;
        RECT 56.45 37.21 56.81 37.57 ;
        RECT 56.45 29.11 56.81 29.47 ;
        RECT 56.45 27.54 56.81 27.9 ;
        RECT 56.45 25.97 56.81 26.33 ;
        RECT 56.45 17.87 56.81 18.23 ;
        RECT 56.45 16.3 56.81 16.66 ;
        RECT 56.45 14.73 56.81 15.09 ;
        RECT 57.15 90.92 57.51 91.28 ;
        RECT 57.15 90.11 57.51 90.47 ;
        RECT 57.15 89.3 57.51 89.66 ;
        RECT 57.15 88.49 57.51 88.85 ;
        RECT 57.15 87.68 57.51 88.04 ;
        RECT 57.15 79.68 57.51 80.04 ;
        RECT 57.15 78.87 57.51 79.23 ;
        RECT 57.15 78.06 57.51 78.42 ;
        RECT 57.15 77.25 57.51 77.61 ;
        RECT 57.15 76.44 57.51 76.8 ;
        RECT 57.15 68.44 57.51 68.8 ;
        RECT 57.15 67.63 57.51 67.99 ;
        RECT 57.15 66.82 57.51 67.18 ;
        RECT 57.15 66.01 57.51 66.37 ;
        RECT 57.15 65.2 57.51 65.56 ;
        RECT 57.15 57.2 57.51 57.56 ;
        RECT 57.15 56.39 57.51 56.75 ;
        RECT 57.15 55.58 57.51 55.94 ;
        RECT 57.15 54.77 57.51 55.13 ;
        RECT 57.15 53.96 57.51 54.32 ;
        RECT 57.15 45.96 57.51 46.32 ;
        RECT 57.15 45.15 57.51 45.51 ;
        RECT 57.15 44.34 57.51 44.7 ;
        RECT 57.15 43.53 57.51 43.89 ;
        RECT 57.15 42.72 57.51 43.08 ;
        RECT 57.15 34.72 57.51 35.08 ;
        RECT 57.15 33.91 57.51 34.27 ;
        RECT 57.15 33.1 57.51 33.46 ;
        RECT 57.15 32.29 57.51 32.65 ;
        RECT 57.15 31.48 57.51 31.84 ;
        RECT 57.15 23.48 57.51 23.84 ;
        RECT 57.15 22.67 57.51 23.03 ;
        RECT 57.15 21.86 57.51 22.22 ;
        RECT 57.15 21.05 57.51 21.41 ;
        RECT 57.15 20.24 57.51 20.6 ;
        RECT 57.15 12.24 57.51 12.6 ;
        RECT 9.05 90.92 9.41 91.28 ;
        RECT 9.05 90.11 9.41 90.47 ;
        RECT 9.05 89.3 9.41 89.66 ;
        RECT 9.05 88.49 9.41 88.85 ;
        RECT 9.05 87.68 9.41 88.04 ;
        RECT 9.05 79.68 9.41 80.04 ;
        RECT 9.05 78.87 9.41 79.23 ;
        RECT 9.05 78.06 9.41 78.42 ;
        RECT 9.05 77.25 9.41 77.61 ;
        RECT 9.05 76.44 9.41 76.8 ;
        RECT 9.05 68.44 9.41 68.8 ;
        RECT 9.05 67.63 9.41 67.99 ;
        RECT 9.05 66.82 9.41 67.18 ;
        RECT 9.05 66.01 9.41 66.37 ;
        RECT 9.05 65.2 9.41 65.56 ;
        RECT 9.05 57.2 9.41 57.56 ;
        RECT 9.05 56.39 9.41 56.75 ;
        RECT 9.05 55.58 9.41 55.94 ;
        RECT 9.05 54.77 9.41 55.13 ;
        RECT 9.05 53.96 9.41 54.32 ;
        RECT 9.05 45.96 9.41 46.32 ;
        RECT 9.05 45.15 9.41 45.51 ;
        RECT 9.05 44.34 9.41 44.7 ;
        RECT 9.05 43.53 9.41 43.89 ;
        RECT 9.05 42.72 9.41 43.08 ;
        RECT 9.05 34.72 9.41 35.08 ;
        RECT 9.05 33.91 9.41 34.27 ;
        RECT 9.05 33.1 9.41 33.46 ;
        RECT 9.05 32.29 9.41 32.65 ;
        RECT 9.05 31.48 9.41 31.84 ;
        RECT 9.05 23.48 9.41 23.84 ;
        RECT 9.05 22.67 9.41 23.03 ;
        RECT 9.05 21.86 9.41 22.22 ;
        RECT 9.05 21.05 9.41 21.41 ;
        RECT 9.05 20.24 9.41 20.6 ;
        RECT 9.05 12.24 9.41 12.6 ;
        RECT 9.05 11.43 9.41 11.79 ;
        RECT 9.05 10.62 9.41 10.98 ;
        RECT 9.05 9.81 9.41 10.17 ;
        RECT 9.05 9 9.41 9.36 ;
        RECT 9.06 85.31 9.42 85.67 ;
        RECT 9.06 83.74 9.42 84.1 ;
        RECT 9.06 82.17 9.42 82.53 ;
        RECT 9.06 74.07 9.42 74.43 ;
        RECT 9.06 72.5 9.42 72.86 ;
        RECT 9.06 70.93 9.42 71.29 ;
        RECT 9.06 62.83 9.42 63.19 ;
        RECT 9.06 61.26 9.42 61.62 ;
        RECT 9.06 59.69 9.42 60.05 ;
        RECT 9.06 51.59 9.42 51.95 ;
        RECT 9.06 50.02 9.42 50.38 ;
        RECT 9.06 48.45 9.42 48.81 ;
        RECT 9.06 40.35 9.42 40.71 ;
        RECT 9.06 38.78 9.42 39.14 ;
        RECT 9.06 37.21 9.42 37.57 ;
        RECT 9.06 29.11 9.42 29.47 ;
        RECT 9.06 27.54 9.42 27.9 ;
        RECT 9.06 25.97 9.42 26.33 ;
        RECT 9.06 17.87 9.42 18.23 ;
        RECT 9.06 16.3 9.42 16.66 ;
        RECT 9.06 14.73 9.42 15.09 ;
        RECT 9.87 85.31 10.23 85.67 ;
        RECT 9.87 83.74 10.23 84.1 ;
        RECT 9.87 82.17 10.23 82.53 ;
        RECT 9.87 74.07 10.23 74.43 ;
        RECT 9.87 72.5 10.23 72.86 ;
        RECT 9.87 70.93 10.23 71.29 ;
        RECT 9.87 62.83 10.23 63.19 ;
        RECT 9.87 61.26 10.23 61.62 ;
        RECT 9.87 59.69 10.23 60.05 ;
        RECT 9.87 51.59 10.23 51.95 ;
        RECT 9.87 50.02 10.23 50.38 ;
        RECT 9.87 48.45 10.23 48.81 ;
        RECT 9.87 40.35 10.23 40.71 ;
        RECT 9.87 38.78 10.23 39.14 ;
        RECT 9.87 37.21 10.23 37.57 ;
        RECT 9.87 29.11 10.23 29.47 ;
        RECT 9.87 27.54 10.23 27.9 ;
        RECT 9.87 25.97 10.23 26.33 ;
        RECT 9.87 17.87 10.23 18.23 ;
        RECT 9.87 16.3 10.23 16.66 ;
        RECT 9.87 14.73 10.23 15.09 ;
        RECT 10.62 90.92 10.98 91.28 ;
        RECT 10.62 90.11 10.98 90.47 ;
        RECT 10.62 89.3 10.98 89.66 ;
        RECT 10.62 88.49 10.98 88.85 ;
        RECT 10.62 87.68 10.98 88.04 ;
        RECT 10.62 79.68 10.98 80.04 ;
        RECT 10.62 78.87 10.98 79.23 ;
        RECT 10.62 78.06 10.98 78.42 ;
        RECT 10.62 77.25 10.98 77.61 ;
        RECT 10.62 76.44 10.98 76.8 ;
        RECT 10.62 68.44 10.98 68.8 ;
        RECT 10.62 67.63 10.98 67.99 ;
        RECT 10.62 66.82 10.98 67.18 ;
        RECT 10.62 66.01 10.98 66.37 ;
        RECT 10.62 65.2 10.98 65.56 ;
        RECT 10.62 57.2 10.98 57.56 ;
        RECT 10.62 56.39 10.98 56.75 ;
        RECT 10.62 55.58 10.98 55.94 ;
        RECT 10.62 54.77 10.98 55.13 ;
        RECT 10.62 53.96 10.98 54.32 ;
        RECT 10.62 45.96 10.98 46.32 ;
        RECT 10.62 45.15 10.98 45.51 ;
        RECT 10.62 44.34 10.98 44.7 ;
        RECT 10.62 43.53 10.98 43.89 ;
        RECT 10.62 42.72 10.98 43.08 ;
        RECT 10.62 34.72 10.98 35.08 ;
        RECT 10.62 33.91 10.98 34.27 ;
        RECT 10.62 33.1 10.98 33.46 ;
        RECT 10.62 32.29 10.98 32.65 ;
        RECT 10.62 31.48 10.98 31.84 ;
        RECT 10.62 23.48 10.98 23.84 ;
        RECT 10.62 22.67 10.98 23.03 ;
        RECT 10.62 21.86 10.98 22.22 ;
        RECT 10.62 21.05 10.98 21.41 ;
        RECT 10.62 20.24 10.98 20.6 ;
        RECT 10.62 12.24 10.98 12.6 ;
        RECT 10.62 11.43 10.98 11.79 ;
        RECT 10.62 10.62 10.98 10.98 ;
        RECT 10.62 9.81 10.98 10.17 ;
        RECT 10.62 9 10.98 9.36 ;
        RECT 10.68 85.31 11.04 85.67 ;
        RECT 10.68 83.74 11.04 84.1 ;
        RECT 10.68 82.17 11.04 82.53 ;
        RECT 10.68 74.07 11.04 74.43 ;
        RECT 10.68 72.5 11.04 72.86 ;
        RECT 10.68 70.93 11.04 71.29 ;
        RECT 10.68 62.83 11.04 63.19 ;
        RECT 10.68 61.26 11.04 61.62 ;
        RECT 10.68 59.69 11.04 60.05 ;
        RECT 10.68 51.59 11.04 51.95 ;
        RECT 10.68 50.02 11.04 50.38 ;
        RECT 10.68 48.45 11.04 48.81 ;
        RECT 10.68 40.35 11.04 40.71 ;
        RECT 10.68 38.78 11.04 39.14 ;
        RECT 10.68 37.21 11.04 37.57 ;
        RECT 10.68 29.11 11.04 29.47 ;
        RECT 10.68 27.54 11.04 27.9 ;
        RECT 10.68 25.97 11.04 26.33 ;
        RECT 10.68 17.87 11.04 18.23 ;
        RECT 10.68 16.3 11.04 16.66 ;
        RECT 10.68 14.73 11.04 15.09 ;
        RECT 11.49 85.31 11.85 85.67 ;
        RECT 11.49 83.74 11.85 84.1 ;
        RECT 11.49 82.17 11.85 82.53 ;
        RECT 11.49 74.07 11.85 74.43 ;
        RECT 11.49 72.5 11.85 72.86 ;
        RECT 11.49 70.93 11.85 71.29 ;
        RECT 11.49 62.83 11.85 63.19 ;
        RECT 11.49 61.26 11.85 61.62 ;
        RECT 11.49 59.69 11.85 60.05 ;
        RECT 11.49 51.59 11.85 51.95 ;
        RECT 11.49 50.02 11.85 50.38 ;
        RECT 11.49 48.45 11.85 48.81 ;
        RECT 11.49 40.35 11.85 40.71 ;
        RECT 11.49 38.78 11.85 39.14 ;
        RECT 11.49 37.21 11.85 37.57 ;
        RECT 11.49 29.11 11.85 29.47 ;
        RECT 11.49 27.54 11.85 27.9 ;
        RECT 11.49 25.97 11.85 26.33 ;
        RECT 11.49 17.87 11.85 18.23 ;
        RECT 11.49 16.3 11.85 16.66 ;
        RECT 11.49 14.73 11.85 15.09 ;
        RECT 12.19 90.92 12.55 91.28 ;
        RECT 12.19 90.11 12.55 90.47 ;
        RECT 12.19 89.3 12.55 89.66 ;
        RECT 12.19 88.49 12.55 88.85 ;
        RECT 12.19 87.68 12.55 88.04 ;
        RECT 12.19 79.68 12.55 80.04 ;
        RECT 12.19 78.87 12.55 79.23 ;
        RECT 12.19 78.06 12.55 78.42 ;
        RECT 12.19 77.25 12.55 77.61 ;
        RECT 12.19 76.44 12.55 76.8 ;
        RECT 12.19 68.44 12.55 68.8 ;
        RECT 12.19 67.63 12.55 67.99 ;
        RECT 12.19 66.82 12.55 67.18 ;
        RECT 12.19 66.01 12.55 66.37 ;
        RECT 12.19 65.2 12.55 65.56 ;
        RECT 12.19 57.2 12.55 57.56 ;
        RECT 12.19 56.39 12.55 56.75 ;
        RECT 12.19 55.58 12.55 55.94 ;
        RECT 12.19 54.77 12.55 55.13 ;
        RECT 12.19 53.96 12.55 54.32 ;
        RECT 12.19 45.96 12.55 46.32 ;
        RECT 12.19 45.15 12.55 45.51 ;
        RECT 12.19 44.34 12.55 44.7 ;
        RECT 12.19 43.53 12.55 43.89 ;
        RECT 12.19 42.72 12.55 43.08 ;
        RECT 12.19 34.72 12.55 35.08 ;
        RECT 12.19 33.91 12.55 34.27 ;
        RECT 12.19 33.1 12.55 33.46 ;
        RECT 12.19 32.29 12.55 32.65 ;
        RECT 12.19 31.48 12.55 31.84 ;
        RECT 12.19 23.48 12.55 23.84 ;
        RECT 12.19 22.67 12.55 23.03 ;
        RECT 12.19 21.86 12.55 22.22 ;
        RECT 12.19 21.05 12.55 21.41 ;
        RECT 12.19 20.24 12.55 20.6 ;
        RECT 12.19 12.24 12.55 12.6 ;
        RECT 12.19 11.43 12.55 11.79 ;
        RECT 12.19 10.62 12.55 10.98 ;
        RECT 12.19 9.81 12.55 10.17 ;
        RECT 12.19 9 12.55 9.36 ;
        RECT 12.3 85.31 12.66 85.67 ;
        RECT 12.3 83.74 12.66 84.1 ;
        RECT 12.3 82.17 12.66 82.53 ;
        RECT 12.3 74.07 12.66 74.43 ;
        RECT 12.3 72.5 12.66 72.86 ;
        RECT 12.3 70.93 12.66 71.29 ;
        RECT 12.3 62.83 12.66 63.19 ;
        RECT 12.3 61.26 12.66 61.62 ;
        RECT 12.3 59.69 12.66 60.05 ;
        RECT 12.3 51.59 12.66 51.95 ;
        RECT 12.3 50.02 12.66 50.38 ;
        RECT 12.3 48.45 12.66 48.81 ;
        RECT 12.3 40.35 12.66 40.71 ;
        RECT 12.3 38.78 12.66 39.14 ;
        RECT 12.3 37.21 12.66 37.57 ;
        RECT 12.3 29.11 12.66 29.47 ;
        RECT 12.3 27.54 12.66 27.9 ;
        RECT 12.3 25.97 12.66 26.33 ;
        RECT 12.3 17.87 12.66 18.23 ;
        RECT 12.3 16.3 12.66 16.66 ;
        RECT 12.3 14.73 12.66 15.09 ;
        RECT 14.62 90.93 14.98 91.29 ;
        RECT 14.62 89.36 14.98 89.72 ;
        RECT 14.62 87.79 14.98 88.15 ;
        RECT 14.62 79.69 14.98 80.05 ;
        RECT 14.62 78.12 14.98 78.48 ;
        RECT 14.62 76.55 14.98 76.91 ;
        RECT 14.62 68.45 14.98 68.81 ;
        RECT 14.62 66.88 14.98 67.24 ;
        RECT 14.62 65.31 14.98 65.67 ;
        RECT 14.62 57.21 14.98 57.57 ;
        RECT 14.62 55.64 14.98 56 ;
        RECT 14.62 54.07 14.98 54.43 ;
        RECT 14.62 45.97 14.98 46.33 ;
        RECT 14.62 44.4 14.98 44.76 ;
        RECT 14.62 42.83 14.98 43.19 ;
        RECT 14.62 34.73 14.98 35.09 ;
        RECT 14.62 33.16 14.98 33.52 ;
        RECT 14.62 31.59 14.98 31.95 ;
        RECT 14.62 23.49 14.98 23.85 ;
        RECT 14.62 21.92 14.98 22.28 ;
        RECT 14.62 20.35 14.98 20.71 ;
        RECT 14.62 12.25 14.98 12.61 ;
        RECT 14.62 10.68 14.98 11.04 ;
        RECT 14.62 9.11 14.98 9.47 ;
        RECT 14.73 85.3 15.09 85.66 ;
        RECT 14.73 84.49 15.09 84.85 ;
        RECT 14.73 83.68 15.09 84.04 ;
        RECT 14.73 82.87 15.09 83.23 ;
        RECT 14.73 82.06 15.09 82.42 ;
        RECT 14.73 74.06 15.09 74.42 ;
        RECT 14.73 73.25 15.09 73.61 ;
        RECT 14.73 72.44 15.09 72.8 ;
        RECT 14.73 71.63 15.09 71.99 ;
        RECT 14.73 70.82 15.09 71.18 ;
        RECT 14.73 62.82 15.09 63.18 ;
        RECT 14.73 62.01 15.09 62.37 ;
        RECT 14.73 61.2 15.09 61.56 ;
        RECT 14.73 60.39 15.09 60.75 ;
        RECT 14.73 59.58 15.09 59.94 ;
        RECT 14.73 51.58 15.09 51.94 ;
        RECT 14.73 50.77 15.09 51.13 ;
        RECT 14.73 49.96 15.09 50.32 ;
        RECT 14.73 49.15 15.09 49.51 ;
        RECT 14.73 48.34 15.09 48.7 ;
        RECT 14.73 40.34 15.09 40.7 ;
        RECT 14.73 39.53 15.09 39.89 ;
        RECT 14.73 38.72 15.09 39.08 ;
        RECT 14.73 37.91 15.09 38.27 ;
        RECT 14.73 37.1 15.09 37.46 ;
        RECT 14.73 29.1 15.09 29.46 ;
        RECT 14.73 28.29 15.09 28.65 ;
        RECT 14.73 27.48 15.09 27.84 ;
        RECT 14.73 26.67 15.09 27.03 ;
        RECT 14.73 25.86 15.09 26.22 ;
        RECT 14.73 17.86 15.09 18.22 ;
        RECT 14.73 17.05 15.09 17.41 ;
        RECT 14.73 16.24 15.09 16.6 ;
        RECT 14.73 15.43 15.09 15.79 ;
        RECT 14.73 14.62 15.09 14.98 ;
        RECT 15.43 90.93 15.79 91.29 ;
        RECT 15.43 89.36 15.79 89.72 ;
        RECT 15.43 87.79 15.79 88.15 ;
        RECT 15.43 79.69 15.79 80.05 ;
        RECT 15.43 78.12 15.79 78.48 ;
        RECT 15.43 76.55 15.79 76.91 ;
        RECT 15.43 68.45 15.79 68.81 ;
        RECT 15.43 66.88 15.79 67.24 ;
        RECT 15.43 65.31 15.79 65.67 ;
        RECT 15.43 57.21 15.79 57.57 ;
        RECT 15.43 55.64 15.79 56 ;
        RECT 15.43 54.07 15.79 54.43 ;
        RECT 15.43 45.97 15.79 46.33 ;
        RECT 15.43 44.4 15.79 44.76 ;
        RECT 15.43 42.83 15.79 43.19 ;
        RECT 15.43 34.73 15.79 35.09 ;
        RECT 15.43 33.16 15.79 33.52 ;
        RECT 15.43 31.59 15.79 31.95 ;
        RECT 15.43 23.49 15.79 23.85 ;
        RECT 15.43 21.92 15.79 22.28 ;
        RECT 15.43 20.35 15.79 20.71 ;
        RECT 15.43 12.25 15.79 12.61 ;
        RECT 15.43 10.68 15.79 11.04 ;
        RECT 15.43 9.11 15.79 9.47 ;
        RECT 16.24 90.93 16.6 91.29 ;
        RECT 16.24 89.36 16.6 89.72 ;
        RECT 16.24 87.79 16.6 88.15 ;
        RECT 16.24 79.69 16.6 80.05 ;
        RECT 16.24 78.12 16.6 78.48 ;
        RECT 16.24 76.55 16.6 76.91 ;
        RECT 16.24 68.45 16.6 68.81 ;
        RECT 16.24 66.88 16.6 67.24 ;
        RECT 16.24 65.31 16.6 65.67 ;
        RECT 16.24 57.21 16.6 57.57 ;
        RECT 16.24 55.64 16.6 56 ;
        RECT 16.24 54.07 16.6 54.43 ;
        RECT 16.24 45.97 16.6 46.33 ;
        RECT 16.24 44.4 16.6 44.76 ;
        RECT 16.24 42.83 16.6 43.19 ;
        RECT 16.24 34.73 16.6 35.09 ;
        RECT 16.24 33.16 16.6 33.52 ;
        RECT 16.24 31.59 16.6 31.95 ;
        RECT 16.24 23.49 16.6 23.85 ;
        RECT 16.24 21.92 16.6 22.28 ;
        RECT 16.24 20.35 16.6 20.71 ;
        RECT 16.24 12.25 16.6 12.61 ;
        RECT 16.24 10.68 16.6 11.04 ;
        RECT 16.24 9.11 16.6 9.47 ;
        RECT 16.3 85.3 16.66 85.66 ;
        RECT 16.3 84.49 16.66 84.85 ;
        RECT 16.3 83.68 16.66 84.04 ;
        RECT 16.3 82.87 16.66 83.23 ;
        RECT 16.3 82.06 16.66 82.42 ;
        RECT 16.3 74.06 16.66 74.42 ;
        RECT 16.3 73.25 16.66 73.61 ;
        RECT 16.3 72.44 16.66 72.8 ;
        RECT 16.3 71.63 16.66 71.99 ;
        RECT 16.3 70.82 16.66 71.18 ;
        RECT 16.3 62.82 16.66 63.18 ;
        RECT 16.3 62.01 16.66 62.37 ;
        RECT 16.3 61.2 16.66 61.56 ;
        RECT 16.3 60.39 16.66 60.75 ;
        RECT 16.3 59.58 16.66 59.94 ;
        RECT 16.3 51.58 16.66 51.94 ;
        RECT 16.3 50.77 16.66 51.13 ;
        RECT 16.3 49.96 16.66 50.32 ;
        RECT 16.3 49.15 16.66 49.51 ;
        RECT 16.3 48.34 16.66 48.7 ;
        RECT 16.3 40.34 16.66 40.7 ;
        RECT 16.3 39.53 16.66 39.89 ;
        RECT 16.3 38.72 16.66 39.08 ;
        RECT 16.3 37.91 16.66 38.27 ;
        RECT 16.3 37.1 16.66 37.46 ;
        RECT 16.3 29.1 16.66 29.46 ;
        RECT 16.3 28.29 16.66 28.65 ;
        RECT 16.3 27.48 16.66 27.84 ;
        RECT 16.3 26.67 16.66 27.03 ;
        RECT 16.3 25.86 16.66 26.22 ;
        RECT 16.3 17.86 16.66 18.22 ;
        RECT 16.3 17.05 16.66 17.41 ;
        RECT 16.3 16.24 16.66 16.6 ;
        RECT 16.3 15.43 16.66 15.79 ;
        RECT 16.3 14.62 16.66 14.98 ;
        RECT 17.05 90.93 17.41 91.29 ;
        RECT 17.05 89.36 17.41 89.72 ;
        RECT 17.05 87.79 17.41 88.15 ;
        RECT 17.05 79.69 17.41 80.05 ;
        RECT 17.05 78.12 17.41 78.48 ;
        RECT 17.05 76.55 17.41 76.91 ;
        RECT 17.05 68.45 17.41 68.81 ;
        RECT 17.05 66.88 17.41 67.24 ;
        RECT 17.05 65.31 17.41 65.67 ;
        RECT 17.05 57.21 17.41 57.57 ;
        RECT 17.05 55.64 17.41 56 ;
        RECT 17.05 54.07 17.41 54.43 ;
        RECT 17.05 45.97 17.41 46.33 ;
        RECT 17.05 44.4 17.41 44.76 ;
        RECT 17.05 42.83 17.41 43.19 ;
        RECT 17.05 34.73 17.41 35.09 ;
        RECT 17.05 33.16 17.41 33.52 ;
        RECT 17.05 31.59 17.41 31.95 ;
        RECT 17.05 23.49 17.41 23.85 ;
        RECT 17.05 21.92 17.41 22.28 ;
        RECT 17.05 20.35 17.41 20.71 ;
        RECT 17.05 12.25 17.41 12.61 ;
        RECT 17.05 10.68 17.41 11.04 ;
        RECT 17.05 9.11 17.41 9.47 ;
        RECT 17.86 90.93 18.22 91.29 ;
        RECT 17.86 89.36 18.22 89.72 ;
        RECT 17.86 87.79 18.22 88.15 ;
        RECT 17.86 79.69 18.22 80.05 ;
        RECT 17.86 78.12 18.22 78.48 ;
        RECT 17.86 76.55 18.22 76.91 ;
        RECT 17.86 68.45 18.22 68.81 ;
        RECT 17.86 66.88 18.22 67.24 ;
        RECT 17.86 65.31 18.22 65.67 ;
        RECT 17.86 57.21 18.22 57.57 ;
        RECT 17.86 55.64 18.22 56 ;
        RECT 17.86 54.07 18.22 54.43 ;
        RECT 17.86 45.97 18.22 46.33 ;
        RECT 17.86 44.4 18.22 44.76 ;
        RECT 17.86 42.83 18.22 43.19 ;
        RECT 17.86 34.73 18.22 35.09 ;
        RECT 17.86 33.16 18.22 33.52 ;
        RECT 17.86 31.59 18.22 31.95 ;
        RECT 17.86 23.49 18.22 23.85 ;
        RECT 17.86 21.92 18.22 22.28 ;
        RECT 17.86 20.35 18.22 20.71 ;
        RECT 17.86 12.25 18.22 12.61 ;
        RECT 17.86 10.68 18.22 11.04 ;
        RECT 17.86 9.11 18.22 9.47 ;
        RECT 17.87 85.3 18.23 85.66 ;
        RECT 17.87 84.49 18.23 84.85 ;
        RECT 17.87 83.68 18.23 84.04 ;
        RECT 17.87 82.87 18.23 83.23 ;
        RECT 17.87 82.06 18.23 82.42 ;
        RECT 17.87 74.06 18.23 74.42 ;
        RECT 17.87 73.25 18.23 73.61 ;
        RECT 17.87 72.44 18.23 72.8 ;
        RECT 17.87 71.63 18.23 71.99 ;
        RECT 17.87 70.82 18.23 71.18 ;
        RECT 17.87 62.82 18.23 63.18 ;
        RECT 17.87 62.01 18.23 62.37 ;
        RECT 17.87 61.2 18.23 61.56 ;
        RECT 17.87 60.39 18.23 60.75 ;
        RECT 17.87 59.58 18.23 59.94 ;
        RECT 17.87 51.58 18.23 51.94 ;
        RECT 17.87 50.77 18.23 51.13 ;
        RECT 17.87 49.96 18.23 50.32 ;
        RECT 17.87 49.15 18.23 49.51 ;
        RECT 17.87 48.34 18.23 48.7 ;
        RECT 17.87 40.34 18.23 40.7 ;
        RECT 17.87 39.53 18.23 39.89 ;
        RECT 17.87 38.72 18.23 39.08 ;
        RECT 17.87 37.91 18.23 38.27 ;
        RECT 17.87 37.1 18.23 37.46 ;
        RECT 17.87 29.1 18.23 29.46 ;
        RECT 17.87 28.29 18.23 28.65 ;
        RECT 17.87 27.48 18.23 27.84 ;
        RECT 17.87 26.67 18.23 27.03 ;
        RECT 17.87 25.86 18.23 26.22 ;
        RECT 17.87 17.86 18.23 18.22 ;
        RECT 17.87 17.05 18.23 17.41 ;
        RECT 17.87 16.24 18.23 16.6 ;
        RECT 17.87 15.43 18.23 15.79 ;
        RECT 17.87 14.62 18.23 14.98 ;
        RECT 20.29 90.92 20.65 91.28 ;
        RECT 20.29 90.11 20.65 90.47 ;
        RECT 20.29 89.3 20.65 89.66 ;
        RECT 20.29 88.49 20.65 88.85 ;
        RECT 20.29 87.68 20.65 88.04 ;
        RECT 20.29 79.68 20.65 80.04 ;
        RECT 20.29 78.87 20.65 79.23 ;
        RECT 20.29 78.06 20.65 78.42 ;
        RECT 20.29 77.25 20.65 77.61 ;
        RECT 20.29 76.44 20.65 76.8 ;
        RECT 20.29 68.44 20.65 68.8 ;
        RECT 20.29 67.63 20.65 67.99 ;
        RECT 20.29 66.82 20.65 67.18 ;
        RECT 20.29 66.01 20.65 66.37 ;
        RECT 20.29 65.2 20.65 65.56 ;
        RECT 20.29 57.2 20.65 57.56 ;
        RECT 20.29 56.39 20.65 56.75 ;
        RECT 20.29 55.58 20.65 55.94 ;
        RECT 20.29 54.77 20.65 55.13 ;
        RECT 20.29 53.96 20.65 54.32 ;
        RECT 20.29 45.96 20.65 46.32 ;
        RECT 20.29 45.15 20.65 45.51 ;
        RECT 20.29 44.34 20.65 44.7 ;
        RECT 20.29 43.53 20.65 43.89 ;
        RECT 20.29 42.72 20.65 43.08 ;
        RECT 20.29 34.72 20.65 35.08 ;
        RECT 20.29 33.91 20.65 34.27 ;
        RECT 20.29 33.1 20.65 33.46 ;
        RECT 20.29 32.29 20.65 32.65 ;
        RECT 20.29 31.48 20.65 31.84 ;
        RECT 20.29 23.48 20.65 23.84 ;
        RECT 20.29 22.67 20.65 23.03 ;
        RECT 20.29 21.86 20.65 22.22 ;
        RECT 20.29 21.05 20.65 21.41 ;
        RECT 20.29 20.24 20.65 20.6 ;
        RECT 20.29 12.24 20.65 12.6 ;
        RECT 20.29 11.43 20.65 11.79 ;
        RECT 20.29 10.62 20.65 10.98 ;
        RECT 20.29 9.81 20.65 10.17 ;
        RECT 20.29 9 20.65 9.36 ;
        RECT 20.3 85.31 20.66 85.67 ;
        RECT 20.3 83.74 20.66 84.1 ;
        RECT 20.3 82.17 20.66 82.53 ;
        RECT 20.3 74.07 20.66 74.43 ;
        RECT 20.3 72.5 20.66 72.86 ;
        RECT 20.3 70.93 20.66 71.29 ;
        RECT 20.3 62.83 20.66 63.19 ;
        RECT 20.3 61.26 20.66 61.62 ;
        RECT 20.3 59.69 20.66 60.05 ;
        RECT 20.3 51.59 20.66 51.95 ;
        RECT 20.3 50.02 20.66 50.38 ;
        RECT 20.3 48.45 20.66 48.81 ;
        RECT 20.3 40.35 20.66 40.71 ;
        RECT 20.3 38.78 20.66 39.14 ;
        RECT 20.3 37.21 20.66 37.57 ;
        RECT 20.3 29.11 20.66 29.47 ;
        RECT 20.3 27.54 20.66 27.9 ;
        RECT 20.3 25.97 20.66 26.33 ;
        RECT 20.3 17.87 20.66 18.23 ;
        RECT 20.3 16.3 20.66 16.66 ;
        RECT 20.3 14.73 20.66 15.09 ;
        RECT 21.11 85.31 21.47 85.67 ;
        RECT 21.11 83.74 21.47 84.1 ;
        RECT 21.11 82.17 21.47 82.53 ;
        RECT 21.11 74.07 21.47 74.43 ;
        RECT 21.11 72.5 21.47 72.86 ;
        RECT 21.11 70.93 21.47 71.29 ;
        RECT 21.11 62.83 21.47 63.19 ;
        RECT 21.11 61.26 21.47 61.62 ;
        RECT 21.11 59.69 21.47 60.05 ;
        RECT 21.11 51.59 21.47 51.95 ;
        RECT 21.11 50.02 21.47 50.38 ;
        RECT 21.11 48.45 21.47 48.81 ;
        RECT 21.11 40.35 21.47 40.71 ;
        RECT 21.11 38.78 21.47 39.14 ;
        RECT 21.11 37.21 21.47 37.57 ;
        RECT 21.11 29.11 21.47 29.47 ;
        RECT 21.11 27.54 21.47 27.9 ;
        RECT 21.11 25.97 21.47 26.33 ;
        RECT 21.11 17.87 21.47 18.23 ;
        RECT 21.11 16.3 21.47 16.66 ;
        RECT 21.11 14.73 21.47 15.09 ;
        RECT 21.86 90.92 22.22 91.28 ;
        RECT 21.86 90.11 22.22 90.47 ;
        RECT 21.86 89.3 22.22 89.66 ;
        RECT 21.86 88.49 22.22 88.85 ;
        RECT 21.86 87.68 22.22 88.04 ;
        RECT 21.86 79.68 22.22 80.04 ;
        RECT 21.86 78.87 22.22 79.23 ;
        RECT 21.86 78.06 22.22 78.42 ;
        RECT 21.86 77.25 22.22 77.61 ;
        RECT 21.86 76.44 22.22 76.8 ;
        RECT 21.86 68.44 22.22 68.8 ;
        RECT 21.86 67.63 22.22 67.99 ;
        RECT 21.86 66.82 22.22 67.18 ;
        RECT 21.86 66.01 22.22 66.37 ;
        RECT 21.86 65.2 22.22 65.56 ;
        RECT 21.86 57.2 22.22 57.56 ;
        RECT 21.86 56.39 22.22 56.75 ;
        RECT 21.86 55.58 22.22 55.94 ;
        RECT 21.86 54.77 22.22 55.13 ;
        RECT 21.86 53.96 22.22 54.32 ;
        RECT 21.86 45.96 22.22 46.32 ;
        RECT 21.86 45.15 22.22 45.51 ;
        RECT 21.86 44.34 22.22 44.7 ;
        RECT 21.86 43.53 22.22 43.89 ;
        RECT 21.86 42.72 22.22 43.08 ;
        RECT 21.86 34.72 22.22 35.08 ;
        RECT 21.86 33.91 22.22 34.27 ;
        RECT 21.86 33.1 22.22 33.46 ;
        RECT 21.86 32.29 22.22 32.65 ;
        RECT 21.86 31.48 22.22 31.84 ;
        RECT 21.86 23.48 22.22 23.84 ;
        RECT 21.86 22.67 22.22 23.03 ;
        RECT 21.86 21.86 22.22 22.22 ;
        RECT 21.86 21.05 22.22 21.41 ;
        RECT 21.86 20.24 22.22 20.6 ;
        RECT 21.86 12.24 22.22 12.6 ;
        RECT 21.86 11.43 22.22 11.79 ;
        RECT 21.86 10.62 22.22 10.98 ;
        RECT 21.86 9.81 22.22 10.17 ;
        RECT 21.86 9 22.22 9.36 ;
        RECT 21.92 85.31 22.28 85.67 ;
        RECT 21.92 83.74 22.28 84.1 ;
        RECT 21.92 82.17 22.28 82.53 ;
        RECT 21.92 74.07 22.28 74.43 ;
        RECT 21.92 72.5 22.28 72.86 ;
        RECT 21.92 70.93 22.28 71.29 ;
        RECT 21.92 62.83 22.28 63.19 ;
        RECT 21.92 61.26 22.28 61.62 ;
        RECT 21.92 59.69 22.28 60.05 ;
        RECT 21.92 51.59 22.28 51.95 ;
        RECT 21.92 50.02 22.28 50.38 ;
        RECT 21.92 48.45 22.28 48.81 ;
        RECT 21.92 40.35 22.28 40.71 ;
        RECT 21.92 38.78 22.28 39.14 ;
        RECT 21.92 37.21 22.28 37.57 ;
        RECT 21.92 29.11 22.28 29.47 ;
        RECT 21.92 27.54 22.28 27.9 ;
        RECT 21.92 25.97 22.28 26.33 ;
        RECT 21.92 17.87 22.28 18.23 ;
        RECT 21.92 16.3 22.28 16.66 ;
        RECT 21.92 14.73 22.28 15.09 ;
        RECT 22.73 85.31 23.09 85.67 ;
        RECT 22.73 83.74 23.09 84.1 ;
        RECT 22.73 82.17 23.09 82.53 ;
        RECT 22.73 74.07 23.09 74.43 ;
        RECT 22.73 72.5 23.09 72.86 ;
        RECT 22.73 70.93 23.09 71.29 ;
        RECT 22.73 62.83 23.09 63.19 ;
        RECT 22.73 61.26 23.09 61.62 ;
        RECT 22.73 59.69 23.09 60.05 ;
        RECT 22.73 51.59 23.09 51.95 ;
        RECT 22.73 50.02 23.09 50.38 ;
        RECT 22.73 48.45 23.09 48.81 ;
        RECT 22.73 40.35 23.09 40.71 ;
        RECT 22.73 38.78 23.09 39.14 ;
        RECT 22.73 37.21 23.09 37.57 ;
        RECT 22.73 29.11 23.09 29.47 ;
        RECT 22.73 27.54 23.09 27.9 ;
        RECT 22.73 25.97 23.09 26.33 ;
        RECT 22.73 17.87 23.09 18.23 ;
        RECT 22.73 16.3 23.09 16.66 ;
        RECT 22.73 14.73 23.09 15.09 ;
        RECT 23.43 90.92 23.79 91.28 ;
        RECT 23.43 90.11 23.79 90.47 ;
        RECT 23.43 89.3 23.79 89.66 ;
        RECT 23.43 88.49 23.79 88.85 ;
        RECT 23.43 87.68 23.79 88.04 ;
        RECT 23.43 79.68 23.79 80.04 ;
        RECT 23.43 78.87 23.79 79.23 ;
        RECT 23.43 78.06 23.79 78.42 ;
        RECT 23.43 77.25 23.79 77.61 ;
        RECT 23.43 76.44 23.79 76.8 ;
        RECT 23.43 68.44 23.79 68.8 ;
        RECT 23.43 67.63 23.79 67.99 ;
        RECT 23.43 66.82 23.79 67.18 ;
        RECT 23.43 66.01 23.79 66.37 ;
        RECT 23.43 65.2 23.79 65.56 ;
        RECT 23.43 57.2 23.79 57.56 ;
        RECT 23.43 56.39 23.79 56.75 ;
        RECT 23.43 55.58 23.79 55.94 ;
        RECT 23.43 54.77 23.79 55.13 ;
        RECT 23.43 53.96 23.79 54.32 ;
        RECT 23.43 45.96 23.79 46.32 ;
        RECT 23.43 45.15 23.79 45.51 ;
        RECT 23.43 44.34 23.79 44.7 ;
        RECT 23.43 43.53 23.79 43.89 ;
        RECT 23.43 42.72 23.79 43.08 ;
        RECT 23.43 34.72 23.79 35.08 ;
        RECT 23.43 33.91 23.79 34.27 ;
        RECT 23.43 33.1 23.79 33.46 ;
        RECT 23.43 32.29 23.79 32.65 ;
        RECT 23.43 31.48 23.79 31.84 ;
        RECT 23.43 23.48 23.79 23.84 ;
        RECT 23.43 22.67 23.79 23.03 ;
        RECT 23.43 21.86 23.79 22.22 ;
        RECT 23.43 21.05 23.79 21.41 ;
        RECT 23.43 20.24 23.79 20.6 ;
        RECT 23.43 12.24 23.79 12.6 ;
        RECT 23.43 11.43 23.79 11.79 ;
        RECT 23.43 10.62 23.79 10.98 ;
        RECT 23.43 9.81 23.79 10.17 ;
        RECT 23.43 9 23.79 9.36 ;
        RECT 23.54 85.31 23.9 85.67 ;
        RECT 23.54 83.74 23.9 84.1 ;
        RECT 23.54 82.17 23.9 82.53 ;
        RECT 23.54 74.07 23.9 74.43 ;
        RECT 23.54 72.5 23.9 72.86 ;
        RECT 23.54 70.93 23.9 71.29 ;
        RECT 23.54 62.83 23.9 63.19 ;
        RECT 23.54 61.26 23.9 61.62 ;
        RECT 23.54 59.69 23.9 60.05 ;
        RECT 23.54 51.59 23.9 51.95 ;
        RECT 23.54 50.02 23.9 50.38 ;
        RECT 23.54 48.45 23.9 48.81 ;
        RECT 23.54 40.35 23.9 40.71 ;
        RECT 23.54 38.78 23.9 39.14 ;
        RECT 23.54 37.21 23.9 37.57 ;
        RECT 23.54 29.11 23.9 29.47 ;
        RECT 23.54 27.54 23.9 27.9 ;
        RECT 23.54 25.97 23.9 26.33 ;
        RECT 23.54 17.87 23.9 18.23 ;
        RECT 23.54 16.3 23.9 16.66 ;
        RECT 23.54 14.73 23.9 15.09 ;
        RECT 25.86 90.93 26.22 91.29 ;
        RECT 25.86 89.36 26.22 89.72 ;
        RECT 25.86 87.79 26.22 88.15 ;
        RECT 25.86 79.69 26.22 80.05 ;
        RECT 25.86 78.12 26.22 78.48 ;
        RECT 25.86 76.55 26.22 76.91 ;
        RECT 25.86 68.45 26.22 68.81 ;
        RECT 25.86 66.88 26.22 67.24 ;
        RECT 25.86 65.31 26.22 65.67 ;
        RECT 25.86 57.21 26.22 57.57 ;
        RECT 25.86 55.64 26.22 56 ;
        RECT 25.86 54.07 26.22 54.43 ;
        RECT 25.86 45.97 26.22 46.33 ;
        RECT 25.86 44.4 26.22 44.76 ;
        RECT 25.86 42.83 26.22 43.19 ;
        RECT 25.86 34.73 26.22 35.09 ;
        RECT 25.86 33.16 26.22 33.52 ;
        RECT 25.86 31.59 26.22 31.95 ;
        RECT 25.86 23.49 26.22 23.85 ;
        RECT 25.86 21.92 26.22 22.28 ;
        RECT 25.86 20.35 26.22 20.71 ;
        RECT 25.86 12.25 26.22 12.61 ;
        RECT 25.86 10.68 26.22 11.04 ;
        RECT 25.86 9.11 26.22 9.47 ;
        RECT 25.97 85.3 26.33 85.66 ;
        RECT 25.97 84.49 26.33 84.85 ;
        RECT 25.97 83.68 26.33 84.04 ;
        RECT 25.97 82.87 26.33 83.23 ;
        RECT 25.97 82.06 26.33 82.42 ;
        RECT 25.97 74.06 26.33 74.42 ;
        RECT 25.97 73.25 26.33 73.61 ;
        RECT 25.97 72.44 26.33 72.8 ;
        RECT 25.97 71.63 26.33 71.99 ;
        RECT 25.97 70.82 26.33 71.18 ;
        RECT 25.97 62.82 26.33 63.18 ;
        RECT 25.97 62.01 26.33 62.37 ;
        RECT 25.97 61.2 26.33 61.56 ;
        RECT 25.97 60.39 26.33 60.75 ;
        RECT 25.97 59.58 26.33 59.94 ;
        RECT 25.97 51.58 26.33 51.94 ;
        RECT 25.97 50.77 26.33 51.13 ;
        RECT 25.97 49.96 26.33 50.32 ;
        RECT 25.97 49.15 26.33 49.51 ;
        RECT 25.97 48.34 26.33 48.7 ;
        RECT 25.97 40.34 26.33 40.7 ;
        RECT 25.97 39.53 26.33 39.89 ;
        RECT 25.97 38.72 26.33 39.08 ;
        RECT 25.97 37.91 26.33 38.27 ;
        RECT 25.97 37.1 26.33 37.46 ;
        RECT 25.97 29.1 26.33 29.46 ;
        RECT 25.97 28.29 26.33 28.65 ;
        RECT 25.97 27.48 26.33 27.84 ;
        RECT 25.97 26.67 26.33 27.03 ;
        RECT 25.97 25.86 26.33 26.22 ;
        RECT 25.97 17.86 26.33 18.22 ;
        RECT 25.97 17.05 26.33 17.41 ;
        RECT 25.97 16.24 26.33 16.6 ;
        RECT 25.97 15.43 26.33 15.79 ;
        RECT 25.97 14.62 26.33 14.98 ;
        RECT 26.67 90.93 27.03 91.29 ;
        RECT 26.67 89.36 27.03 89.72 ;
        RECT 26.67 87.79 27.03 88.15 ;
        RECT 26.67 79.69 27.03 80.05 ;
        RECT 26.67 78.12 27.03 78.48 ;
        RECT 26.67 76.55 27.03 76.91 ;
        RECT 26.67 68.45 27.03 68.81 ;
        RECT 26.67 66.88 27.03 67.24 ;
        RECT 26.67 65.31 27.03 65.67 ;
        RECT 26.67 57.21 27.03 57.57 ;
        RECT 26.67 55.64 27.03 56 ;
        RECT 26.67 54.07 27.03 54.43 ;
        RECT 26.67 45.97 27.03 46.33 ;
        RECT 26.67 44.4 27.03 44.76 ;
        RECT 26.67 42.83 27.03 43.19 ;
        RECT 26.67 34.73 27.03 35.09 ;
        RECT 26.67 33.16 27.03 33.52 ;
        RECT 26.67 31.59 27.03 31.95 ;
        RECT 26.67 23.49 27.03 23.85 ;
        RECT 26.67 21.92 27.03 22.28 ;
        RECT 26.67 20.35 27.03 20.71 ;
        RECT 26.67 12.25 27.03 12.61 ;
        RECT 26.67 10.68 27.03 11.04 ;
        RECT 26.67 9.11 27.03 9.47 ;
        RECT 27.48 90.93 27.84 91.29 ;
        RECT 27.48 89.36 27.84 89.72 ;
        RECT 27.48 87.79 27.84 88.15 ;
        RECT 27.48 79.69 27.84 80.05 ;
        RECT 27.48 78.12 27.84 78.48 ;
        RECT 27.48 76.55 27.84 76.91 ;
        RECT 27.48 68.45 27.84 68.81 ;
        RECT 27.48 66.88 27.84 67.24 ;
        RECT 27.48 65.31 27.84 65.67 ;
        RECT 27.48 57.21 27.84 57.57 ;
        RECT 27.48 55.64 27.84 56 ;
        RECT 27.48 54.07 27.84 54.43 ;
        RECT 27.48 45.97 27.84 46.33 ;
        RECT 27.48 44.4 27.84 44.76 ;
        RECT 27.48 42.83 27.84 43.19 ;
        RECT 27.48 34.73 27.84 35.09 ;
        RECT 27.48 33.16 27.84 33.52 ;
        RECT 27.48 31.59 27.84 31.95 ;
        RECT 27.48 23.49 27.84 23.85 ;
        RECT 27.48 21.92 27.84 22.28 ;
        RECT 27.48 20.35 27.84 20.71 ;
        RECT 27.48 12.25 27.84 12.61 ;
        RECT 27.48 10.68 27.84 11.04 ;
        RECT 27.48 9.11 27.84 9.47 ;
        RECT 27.54 85.3 27.9 85.66 ;
        RECT 27.54 84.49 27.9 84.85 ;
        RECT 27.54 83.68 27.9 84.04 ;
        RECT 27.54 82.87 27.9 83.23 ;
        RECT 27.54 82.06 27.9 82.42 ;
        RECT 27.54 74.06 27.9 74.42 ;
        RECT 27.54 73.25 27.9 73.61 ;
        RECT 27.54 72.44 27.9 72.8 ;
        RECT 27.54 71.63 27.9 71.99 ;
        RECT 27.54 70.82 27.9 71.18 ;
        RECT 27.54 62.82 27.9 63.18 ;
        RECT 27.54 62.01 27.9 62.37 ;
        RECT 27.54 61.2 27.9 61.56 ;
        RECT 27.54 60.39 27.9 60.75 ;
        RECT 27.54 59.58 27.9 59.94 ;
        RECT 27.54 51.58 27.9 51.94 ;
        RECT 27.54 50.77 27.9 51.13 ;
        RECT 27.54 49.96 27.9 50.32 ;
        RECT 27.54 49.15 27.9 49.51 ;
        RECT 27.54 48.34 27.9 48.7 ;
        RECT 27.54 40.34 27.9 40.7 ;
        RECT 27.54 39.53 27.9 39.89 ;
        RECT 27.54 38.72 27.9 39.08 ;
        RECT 27.54 37.91 27.9 38.27 ;
        RECT 27.54 37.1 27.9 37.46 ;
        RECT 27.54 29.1 27.9 29.46 ;
        RECT 27.54 28.29 27.9 28.65 ;
        RECT 27.54 27.48 27.9 27.84 ;
        RECT 27.54 26.67 27.9 27.03 ;
        RECT 27.54 25.86 27.9 26.22 ;
        RECT 27.54 17.86 27.9 18.22 ;
        RECT 27.54 17.05 27.9 17.41 ;
        RECT 27.54 16.24 27.9 16.6 ;
        RECT 27.54 15.43 27.9 15.79 ;
        RECT 27.54 14.62 27.9 14.98 ;
        RECT 28.29 90.93 28.65 91.29 ;
        RECT 28.29 89.36 28.65 89.72 ;
        RECT 28.29 87.79 28.65 88.15 ;
        RECT 28.29 79.69 28.65 80.05 ;
        RECT 28.29 78.12 28.65 78.48 ;
        RECT 28.29 76.55 28.65 76.91 ;
        RECT 28.29 68.45 28.65 68.81 ;
        RECT 28.29 66.88 28.65 67.24 ;
        RECT 28.29 65.31 28.65 65.67 ;
        RECT 28.29 57.21 28.65 57.57 ;
        RECT 28.29 55.64 28.65 56 ;
        RECT 28.29 54.07 28.65 54.43 ;
        RECT 28.29 45.97 28.65 46.33 ;
        RECT 28.29 44.4 28.65 44.76 ;
        RECT 28.29 42.83 28.65 43.19 ;
        RECT 28.29 34.73 28.65 35.09 ;
        RECT 28.29 33.16 28.65 33.52 ;
        RECT 28.29 31.59 28.65 31.95 ;
        RECT 28.29 23.49 28.65 23.85 ;
        RECT 28.29 21.92 28.65 22.28 ;
        RECT 28.29 20.35 28.65 20.71 ;
        RECT 28.29 12.25 28.65 12.61 ;
        RECT 28.29 10.68 28.65 11.04 ;
        RECT 28.29 9.11 28.65 9.47 ;
        RECT 29.1 90.93 29.46 91.29 ;
        RECT 29.1 89.36 29.46 89.72 ;
        RECT 29.1 87.79 29.46 88.15 ;
        RECT 29.1 79.69 29.46 80.05 ;
        RECT 29.1 78.12 29.46 78.48 ;
        RECT 29.1 76.55 29.46 76.91 ;
        RECT 29.1 68.45 29.46 68.81 ;
        RECT 29.1 66.88 29.46 67.24 ;
        RECT 29.1 65.31 29.46 65.67 ;
        RECT 29.1 57.21 29.46 57.57 ;
        RECT 29.1 55.64 29.46 56 ;
        RECT 29.1 54.07 29.46 54.43 ;
        RECT 29.1 45.97 29.46 46.33 ;
        RECT 29.1 44.4 29.46 44.76 ;
        RECT 29.1 42.83 29.46 43.19 ;
        RECT 29.1 34.73 29.46 35.09 ;
        RECT 29.1 33.16 29.46 33.52 ;
        RECT 29.1 31.59 29.46 31.95 ;
        RECT 29.1 23.49 29.46 23.85 ;
        RECT 29.1 21.92 29.46 22.28 ;
        RECT 29.1 20.35 29.46 20.71 ;
        RECT 29.1 12.25 29.46 12.61 ;
        RECT 29.1 10.68 29.46 11.04 ;
        RECT 29.1 9.11 29.46 9.47 ;
        RECT 29.11 85.3 29.47 85.66 ;
        RECT 29.11 84.49 29.47 84.85 ;
        RECT 29.11 83.68 29.47 84.04 ;
        RECT 29.11 82.87 29.47 83.23 ;
        RECT 29.11 82.06 29.47 82.42 ;
        RECT 29.11 74.06 29.47 74.42 ;
        RECT 29.11 73.25 29.47 73.61 ;
        RECT 29.11 72.44 29.47 72.8 ;
        RECT 29.11 71.63 29.47 71.99 ;
        RECT 29.11 70.82 29.47 71.18 ;
        RECT 29.11 62.82 29.47 63.18 ;
        RECT 29.11 62.01 29.47 62.37 ;
        RECT 29.11 61.2 29.47 61.56 ;
        RECT 29.11 60.39 29.47 60.75 ;
        RECT 29.11 59.58 29.47 59.94 ;
        RECT 29.11 51.58 29.47 51.94 ;
        RECT 29.11 50.77 29.47 51.13 ;
        RECT 29.11 49.96 29.47 50.32 ;
        RECT 29.11 49.15 29.47 49.51 ;
        RECT 29.11 48.34 29.47 48.7 ;
        RECT 29.11 40.34 29.47 40.7 ;
        RECT 29.11 39.53 29.47 39.89 ;
        RECT 29.11 38.72 29.47 39.08 ;
        RECT 29.11 37.91 29.47 38.27 ;
        RECT 29.11 37.1 29.47 37.46 ;
        RECT 29.11 29.1 29.47 29.46 ;
        RECT 29.11 28.29 29.47 28.65 ;
        RECT 29.11 27.48 29.47 27.84 ;
        RECT 29.11 26.67 29.47 27.03 ;
        RECT 29.11 25.86 29.47 26.22 ;
        RECT 29.11 17.86 29.47 18.22 ;
        RECT 29.11 17.05 29.47 17.41 ;
        RECT 29.11 16.24 29.47 16.6 ;
        RECT 29.11 15.43 29.47 15.79 ;
        RECT 29.11 14.62 29.47 14.98 ;
        RECT 31.53 90.92 31.89 91.28 ;
        RECT 31.53 90.11 31.89 90.47 ;
        RECT 31.53 89.3 31.89 89.66 ;
        RECT 31.53 88.49 31.89 88.85 ;
        RECT 31.53 87.68 31.89 88.04 ;
        RECT 31.53 79.68 31.89 80.04 ;
        RECT 31.53 78.87 31.89 79.23 ;
        RECT 31.53 78.06 31.89 78.42 ;
        RECT 31.53 77.25 31.89 77.61 ;
        RECT 31.53 76.44 31.89 76.8 ;
        RECT 31.53 68.44 31.89 68.8 ;
        RECT 31.53 67.63 31.89 67.99 ;
        RECT 31.53 66.82 31.89 67.18 ;
        RECT 31.53 66.01 31.89 66.37 ;
        RECT 31.53 65.2 31.89 65.56 ;
        RECT 31.53 57.2 31.89 57.56 ;
        RECT 31.53 56.39 31.89 56.75 ;
        RECT 31.53 55.58 31.89 55.94 ;
        RECT 31.53 54.77 31.89 55.13 ;
        RECT 31.53 53.96 31.89 54.32 ;
        RECT 31.53 45.96 31.89 46.32 ;
        RECT 31.53 45.15 31.89 45.51 ;
        RECT 31.53 44.34 31.89 44.7 ;
        RECT 31.53 43.53 31.89 43.89 ;
        RECT 31.53 42.72 31.89 43.08 ;
        RECT 31.53 34.72 31.89 35.08 ;
        RECT 31.53 33.91 31.89 34.27 ;
        RECT 31.53 33.1 31.89 33.46 ;
        RECT 31.53 32.29 31.89 32.65 ;
        RECT 31.53 31.48 31.89 31.84 ;
        RECT 31.53 23.48 31.89 23.84 ;
        RECT 31.53 22.67 31.89 23.03 ;
        RECT 31.53 21.86 31.89 22.22 ;
        RECT 31.53 21.05 31.89 21.41 ;
        RECT 31.53 20.24 31.89 20.6 ;
        RECT 31.53 12.24 31.89 12.6 ;
        RECT 31.53 11.43 31.89 11.79 ;
        RECT 31.53 10.62 31.89 10.98 ;
        RECT 31.53 9.81 31.89 10.17 ;
        RECT 31.53 9 31.89 9.36 ;
        RECT 31.54 85.31 31.9 85.67 ;
        RECT 31.54 83.74 31.9 84.1 ;
        RECT 31.54 82.17 31.9 82.53 ;
        RECT 31.54 74.07 31.9 74.43 ;
        RECT 31.54 72.5 31.9 72.86 ;
        RECT 31.54 70.93 31.9 71.29 ;
        RECT 31.54 62.83 31.9 63.19 ;
        RECT 31.54 61.26 31.9 61.62 ;
        RECT 31.54 59.69 31.9 60.05 ;
        RECT 31.54 51.59 31.9 51.95 ;
        RECT 31.54 50.02 31.9 50.38 ;
        RECT 31.54 48.45 31.9 48.81 ;
        RECT 31.54 40.35 31.9 40.71 ;
        RECT 31.54 38.78 31.9 39.14 ;
        RECT 31.54 37.21 31.9 37.57 ;
        RECT 31.54 29.11 31.9 29.47 ;
        RECT 31.54 27.54 31.9 27.9 ;
        RECT 31.54 25.97 31.9 26.33 ;
        RECT 31.54 17.87 31.9 18.23 ;
        RECT 31.54 16.3 31.9 16.66 ;
        RECT 31.54 14.73 31.9 15.09 ;
        RECT 32.35 85.31 32.71 85.67 ;
        RECT 32.35 83.74 32.71 84.1 ;
        RECT 32.35 82.17 32.71 82.53 ;
        RECT 32.35 74.07 32.71 74.43 ;
        RECT 32.35 72.5 32.71 72.86 ;
        RECT 32.35 70.93 32.71 71.29 ;
        RECT 32.35 62.83 32.71 63.19 ;
        RECT 32.35 61.26 32.71 61.62 ;
        RECT 32.35 59.69 32.71 60.05 ;
        RECT 32.35 51.59 32.71 51.95 ;
        RECT 32.35 50.02 32.71 50.38 ;
        RECT 32.35 48.45 32.71 48.81 ;
        RECT 32.35 40.35 32.71 40.71 ;
        RECT 32.35 38.78 32.71 39.14 ;
        RECT 32.35 37.21 32.71 37.57 ;
        RECT 32.35 29.11 32.71 29.47 ;
        RECT 32.35 27.54 32.71 27.9 ;
        RECT 32.35 25.97 32.71 26.33 ;
        RECT 32.35 17.87 32.71 18.23 ;
        RECT 32.35 16.3 32.71 16.66 ;
        RECT 32.35 14.73 32.71 15.09 ;
        RECT 33.1 90.92 33.46 91.28 ;
        RECT 33.1 90.11 33.46 90.47 ;
        RECT 33.1 89.3 33.46 89.66 ;
        RECT 33.1 88.49 33.46 88.85 ;
        RECT 33.1 87.68 33.46 88.04 ;
        RECT 33.1 79.68 33.46 80.04 ;
        RECT 33.1 78.87 33.46 79.23 ;
        RECT 33.1 78.06 33.46 78.42 ;
        RECT 33.1 77.25 33.46 77.61 ;
        RECT 33.1 76.44 33.46 76.8 ;
        RECT 33.1 68.44 33.46 68.8 ;
        RECT 33.1 67.63 33.46 67.99 ;
        RECT 33.1 66.82 33.46 67.18 ;
        RECT 33.1 66.01 33.46 66.37 ;
        RECT 33.1 65.2 33.46 65.56 ;
        RECT 33.1 57.2 33.46 57.56 ;
        RECT 33.1 56.39 33.46 56.75 ;
        RECT 33.1 55.58 33.46 55.94 ;
      LAYER V4 ;
        RECT 80.65 58.725 80.91 58.985 ;
        RECT 80.65 57.965 80.91 58.225 ;
        RECT 80.65 57.205 80.91 57.465 ;
        RECT 80.65 56.445 80.91 56.705 ;
        RECT 80.65 55.685 80.91 55.945 ;
        RECT 80.65 54.925 80.91 55.185 ;
        RECT 80.65 54.165 80.91 54.425 ;
        RECT 80.65 53.405 80.91 53.665 ;
        RECT 80.65 52.645 80.91 52.905 ;
        RECT 80.65 51.885 80.91 52.145 ;
        RECT 80.65 51.125 80.91 51.385 ;
        RECT 80.65 50.365 80.91 50.625 ;
        RECT 80.65 49.605 80.91 49.865 ;
        RECT 80.65 48.845 80.91 49.105 ;
        RECT 80.65 48.085 80.91 48.345 ;
        RECT 80.65 47.325 80.91 47.585 ;
        RECT 80.65 46.565 80.91 46.825 ;
        RECT 80.65 45.805 80.91 46.065 ;
        RECT 80.65 45.045 80.91 45.305 ;
        RECT 80.65 44.285 80.91 44.545 ;
        RECT 80.65 43.525 80.91 43.785 ;
        RECT 80.65 42.765 80.91 43.025 ;
        RECT 80.65 42.005 80.91 42.265 ;
        RECT 80.65 41.245 80.91 41.505 ;
        RECT 80.65 40.485 80.91 40.745 ;
        RECT 80.65 39.725 80.91 39.985 ;
        RECT 80.65 38.965 80.91 39.225 ;
        RECT 80.65 38.205 80.91 38.465 ;
        RECT 80.65 37.445 80.91 37.705 ;
        RECT 80.65 36.685 80.91 36.945 ;
        RECT 81.41 58.725 81.67 58.985 ;
        RECT 81.41 57.965 81.67 58.225 ;
        RECT 81.41 57.205 81.67 57.465 ;
        RECT 81.41 56.445 81.67 56.705 ;
        RECT 81.41 55.685 81.67 55.945 ;
        RECT 81.41 54.925 81.67 55.185 ;
        RECT 81.41 54.165 81.67 54.425 ;
        RECT 81.41 53.405 81.67 53.665 ;
        RECT 81.41 52.645 81.67 52.905 ;
        RECT 81.41 51.885 81.67 52.145 ;
        RECT 81.41 51.125 81.67 51.385 ;
        RECT 81.41 50.365 81.67 50.625 ;
        RECT 81.41 49.605 81.67 49.865 ;
        RECT 81.41 48.845 81.67 49.105 ;
        RECT 81.41 48.085 81.67 48.345 ;
        RECT 81.41 47.325 81.67 47.585 ;
        RECT 81.41 46.565 81.67 46.825 ;
        RECT 81.41 45.805 81.67 46.065 ;
        RECT 81.41 45.045 81.67 45.305 ;
        RECT 81.41 44.285 81.67 44.545 ;
        RECT 81.41 43.525 81.67 43.785 ;
        RECT 81.41 42.765 81.67 43.025 ;
        RECT 81.41 42.005 81.67 42.265 ;
        RECT 81.41 41.245 81.67 41.505 ;
        RECT 81.41 40.485 81.67 40.745 ;
        RECT 81.41 39.725 81.67 39.985 ;
        RECT 81.41 38.965 81.67 39.225 ;
        RECT 81.41 38.205 81.67 38.465 ;
        RECT 81.41 37.445 81.67 37.705 ;
        RECT 81.41 36.685 81.67 36.945 ;
        RECT 82.17 58.725 82.43 58.985 ;
        RECT 82.17 57.965 82.43 58.225 ;
        RECT 82.17 57.205 82.43 57.465 ;
        RECT 82.17 56.445 82.43 56.705 ;
        RECT 82.17 55.685 82.43 55.945 ;
        RECT 82.17 54.925 82.43 55.185 ;
        RECT 82.17 54.165 82.43 54.425 ;
        RECT 82.17 53.405 82.43 53.665 ;
        RECT 82.17 52.645 82.43 52.905 ;
        RECT 82.17 51.885 82.43 52.145 ;
        RECT 82.17 51.125 82.43 51.385 ;
        RECT 82.17 50.365 82.43 50.625 ;
        RECT 82.17 49.605 82.43 49.865 ;
        RECT 82.17 48.845 82.43 49.105 ;
        RECT 82.17 48.085 82.43 48.345 ;
        RECT 82.17 47.325 82.43 47.585 ;
        RECT 82.17 46.565 82.43 46.825 ;
        RECT 82.17 45.805 82.43 46.065 ;
        RECT 82.17 45.045 82.43 45.305 ;
        RECT 82.17 44.285 82.43 44.545 ;
        RECT 82.17 43.525 82.43 43.785 ;
        RECT 82.17 42.765 82.43 43.025 ;
        RECT 82.17 42.005 82.43 42.265 ;
        RECT 82.17 41.245 82.43 41.505 ;
        RECT 82.17 40.485 82.43 40.745 ;
        RECT 82.17 39.725 82.43 39.985 ;
        RECT 82.17 38.965 82.43 39.225 ;
        RECT 82.17 38.205 82.43 38.465 ;
        RECT 82.17 37.445 82.43 37.705 ;
        RECT 82.17 36.685 82.43 36.945 ;
        RECT 82.93 58.725 83.19 58.985 ;
        RECT 82.93 57.965 83.19 58.225 ;
        RECT 82.93 57.205 83.19 57.465 ;
        RECT 82.93 56.445 83.19 56.705 ;
        RECT 82.93 55.685 83.19 55.945 ;
        RECT 82.93 54.925 83.19 55.185 ;
        RECT 82.93 54.165 83.19 54.425 ;
        RECT 82.93 53.405 83.19 53.665 ;
        RECT 82.93 52.645 83.19 52.905 ;
        RECT 82.93 51.885 83.19 52.145 ;
        RECT 82.93 51.125 83.19 51.385 ;
        RECT 82.93 50.365 83.19 50.625 ;
        RECT 82.93 49.605 83.19 49.865 ;
        RECT 82.93 48.845 83.19 49.105 ;
        RECT 82.93 48.085 83.19 48.345 ;
        RECT 82.93 47.325 83.19 47.585 ;
        RECT 82.93 46.565 83.19 46.825 ;
        RECT 82.93 45.805 83.19 46.065 ;
        RECT 82.93 45.045 83.19 45.305 ;
        RECT 82.93 44.285 83.19 44.545 ;
        RECT 82.93 43.525 83.19 43.785 ;
        RECT 82.93 42.765 83.19 43.025 ;
        RECT 82.93 42.005 83.19 42.265 ;
        RECT 82.93 41.245 83.19 41.505 ;
        RECT 82.93 40.485 83.19 40.745 ;
        RECT 82.93 39.725 83.19 39.985 ;
        RECT 82.93 38.965 83.19 39.225 ;
        RECT 82.93 38.205 83.19 38.465 ;
        RECT 82.93 37.445 83.19 37.705 ;
        RECT 82.93 36.685 83.19 36.945 ;
        RECT 83.69 58.725 83.95 58.985 ;
        RECT 83.69 57.965 83.95 58.225 ;
        RECT 83.69 57.205 83.95 57.465 ;
        RECT 83.69 56.445 83.95 56.705 ;
        RECT 83.69 55.685 83.95 55.945 ;
        RECT 83.69 54.925 83.95 55.185 ;
        RECT 83.69 54.165 83.95 54.425 ;
        RECT 83.69 53.405 83.95 53.665 ;
        RECT 83.69 52.645 83.95 52.905 ;
        RECT 83.69 51.885 83.95 52.145 ;
        RECT 83.69 51.125 83.95 51.385 ;
        RECT 83.69 50.365 83.95 50.625 ;
        RECT 83.69 49.605 83.95 49.865 ;
        RECT 83.69 48.845 83.95 49.105 ;
        RECT 83.69 48.085 83.95 48.345 ;
        RECT 83.69 47.325 83.95 47.585 ;
        RECT 83.69 46.565 83.95 46.825 ;
        RECT 83.69 45.805 83.95 46.065 ;
        RECT 83.69 45.045 83.95 45.305 ;
        RECT 83.69 44.285 83.95 44.545 ;
        RECT 83.69 43.525 83.95 43.785 ;
        RECT 83.69 42.765 83.95 43.025 ;
        RECT 83.69 42.005 83.95 42.265 ;
        RECT 83.69 41.245 83.95 41.505 ;
        RECT 83.69 40.485 83.95 40.745 ;
        RECT 83.69 39.725 83.95 39.985 ;
        RECT 83.69 38.965 83.95 39.225 ;
        RECT 83.69 38.205 83.95 38.465 ;
        RECT 83.69 37.445 83.95 37.705 ;
        RECT 83.69 36.685 83.95 36.945 ;
        RECT 84.45 58.725 84.71 58.985 ;
        RECT 84.45 57.965 84.71 58.225 ;
        RECT 84.45 57.205 84.71 57.465 ;
        RECT 84.45 56.445 84.71 56.705 ;
        RECT 84.45 55.685 84.71 55.945 ;
        RECT 84.45 54.925 84.71 55.185 ;
        RECT 84.45 54.165 84.71 54.425 ;
        RECT 84.45 53.405 84.71 53.665 ;
        RECT 84.45 52.645 84.71 52.905 ;
        RECT 84.45 51.885 84.71 52.145 ;
        RECT 84.45 51.125 84.71 51.385 ;
        RECT 84.45 50.365 84.71 50.625 ;
        RECT 84.45 49.605 84.71 49.865 ;
        RECT 84.45 48.845 84.71 49.105 ;
        RECT 84.45 48.085 84.71 48.345 ;
        RECT 84.45 47.325 84.71 47.585 ;
        RECT 84.45 46.565 84.71 46.825 ;
        RECT 84.45 45.805 84.71 46.065 ;
        RECT 84.45 45.045 84.71 45.305 ;
        RECT 84.45 44.285 84.71 44.545 ;
        RECT 84.45 43.525 84.71 43.785 ;
        RECT 84.45 42.765 84.71 43.025 ;
        RECT 84.45 42.005 84.71 42.265 ;
        RECT 84.45 41.245 84.71 41.505 ;
        RECT 84.45 40.485 84.71 40.745 ;
        RECT 84.45 39.725 84.71 39.985 ;
        RECT 84.45 38.965 84.71 39.225 ;
        RECT 84.45 38.205 84.71 38.465 ;
        RECT 84.45 37.445 84.71 37.705 ;
        RECT 84.45 36.685 84.71 36.945 ;
        RECT 85.21 58.725 85.47 58.985 ;
        RECT 85.21 57.965 85.47 58.225 ;
        RECT 85.21 57.205 85.47 57.465 ;
        RECT 85.21 56.445 85.47 56.705 ;
        RECT 85.21 55.685 85.47 55.945 ;
        RECT 85.21 54.925 85.47 55.185 ;
        RECT 85.21 54.165 85.47 54.425 ;
        RECT 85.21 53.405 85.47 53.665 ;
        RECT 85.21 52.645 85.47 52.905 ;
        RECT 85.21 51.885 85.47 52.145 ;
        RECT 85.21 51.125 85.47 51.385 ;
        RECT 85.21 50.365 85.47 50.625 ;
        RECT 85.21 49.605 85.47 49.865 ;
        RECT 85.21 48.845 85.47 49.105 ;
        RECT 85.21 48.085 85.47 48.345 ;
        RECT 85.21 47.325 85.47 47.585 ;
        RECT 85.21 46.565 85.47 46.825 ;
        RECT 85.21 45.805 85.47 46.065 ;
        RECT 85.21 45.045 85.47 45.305 ;
        RECT 85.21 44.285 85.47 44.545 ;
        RECT 85.21 43.525 85.47 43.785 ;
        RECT 85.21 42.765 85.47 43.025 ;
        RECT 85.21 42.005 85.47 42.265 ;
        RECT 85.21 41.245 85.47 41.505 ;
        RECT 85.21 40.485 85.47 40.745 ;
        RECT 85.21 39.725 85.47 39.985 ;
        RECT 85.21 38.965 85.47 39.225 ;
        RECT 85.21 38.205 85.47 38.465 ;
        RECT 85.21 37.445 85.47 37.705 ;
        RECT 85.21 36.685 85.47 36.945 ;
        RECT 85.97 58.725 86.23 58.985 ;
        RECT 85.97 57.965 86.23 58.225 ;
        RECT 85.97 57.205 86.23 57.465 ;
        RECT 85.97 56.445 86.23 56.705 ;
        RECT 85.97 55.685 86.23 55.945 ;
        RECT 85.97 54.925 86.23 55.185 ;
        RECT 85.97 54.165 86.23 54.425 ;
        RECT 85.97 53.405 86.23 53.665 ;
        RECT 85.97 52.645 86.23 52.905 ;
        RECT 85.97 51.885 86.23 52.145 ;
        RECT 85.97 51.125 86.23 51.385 ;
        RECT 85.97 50.365 86.23 50.625 ;
        RECT 85.97 49.605 86.23 49.865 ;
        RECT 85.97 48.845 86.23 49.105 ;
        RECT 85.97 48.085 86.23 48.345 ;
        RECT 85.97 47.325 86.23 47.585 ;
        RECT 85.97 46.565 86.23 46.825 ;
        RECT 85.97 45.805 86.23 46.065 ;
        RECT 85.97 45.045 86.23 45.305 ;
        RECT 85.97 44.285 86.23 44.545 ;
        RECT 85.97 43.525 86.23 43.785 ;
        RECT 85.97 42.765 86.23 43.025 ;
        RECT 85.97 42.005 86.23 42.265 ;
        RECT 85.97 41.245 86.23 41.505 ;
        RECT 85.97 40.485 86.23 40.745 ;
        RECT 85.97 39.725 86.23 39.985 ;
        RECT 85.97 38.965 86.23 39.225 ;
        RECT 85.97 38.205 86.23 38.465 ;
        RECT 85.97 37.445 86.23 37.705 ;
        RECT 85.97 36.685 86.23 36.945 ;
        RECT 86.73 58.725 86.99 58.985 ;
        RECT 86.73 57.965 86.99 58.225 ;
        RECT 86.73 57.205 86.99 57.465 ;
        RECT 86.73 56.445 86.99 56.705 ;
        RECT 86.73 55.685 86.99 55.945 ;
        RECT 86.73 54.925 86.99 55.185 ;
        RECT 86.73 54.165 86.99 54.425 ;
        RECT 86.73 53.405 86.99 53.665 ;
        RECT 86.73 52.645 86.99 52.905 ;
        RECT 86.73 51.885 86.99 52.145 ;
        RECT 86.73 51.125 86.99 51.385 ;
        RECT 86.73 50.365 86.99 50.625 ;
        RECT 86.73 49.605 86.99 49.865 ;
        RECT 86.73 48.845 86.99 49.105 ;
        RECT 86.73 48.085 86.99 48.345 ;
        RECT 86.73 47.325 86.99 47.585 ;
        RECT 86.73 46.565 86.99 46.825 ;
        RECT 86.73 45.805 86.99 46.065 ;
        RECT 86.73 45.045 86.99 45.305 ;
        RECT 86.73 44.285 86.99 44.545 ;
        RECT 86.73 43.525 86.99 43.785 ;
        RECT 86.73 42.765 86.99 43.025 ;
        RECT 86.73 42.005 86.99 42.265 ;
        RECT 86.73 41.245 86.99 41.505 ;
        RECT 86.73 40.485 86.99 40.745 ;
        RECT 86.73 39.725 86.99 39.985 ;
        RECT 86.73 38.965 86.99 39.225 ;
        RECT 86.73 38.205 86.99 38.465 ;
        RECT 86.73 37.445 86.99 37.705 ;
        RECT 86.73 36.685 86.99 36.945 ;
        RECT 87.49 58.725 87.75 58.985 ;
        RECT 87.49 57.965 87.75 58.225 ;
        RECT 87.49 57.205 87.75 57.465 ;
        RECT 87.49 56.445 87.75 56.705 ;
        RECT 87.49 55.685 87.75 55.945 ;
        RECT 87.49 54.925 87.75 55.185 ;
        RECT 87.49 54.165 87.75 54.425 ;
        RECT 87.49 53.405 87.75 53.665 ;
        RECT 87.49 52.645 87.75 52.905 ;
        RECT 87.49 51.885 87.75 52.145 ;
        RECT 87.49 51.125 87.75 51.385 ;
        RECT 87.49 50.365 87.75 50.625 ;
        RECT 87.49 49.605 87.75 49.865 ;
        RECT 87.49 48.845 87.75 49.105 ;
        RECT 87.49 48.085 87.75 48.345 ;
        RECT 87.49 47.325 87.75 47.585 ;
        RECT 87.49 46.565 87.75 46.825 ;
        RECT 87.49 45.805 87.75 46.065 ;
        RECT 87.49 45.045 87.75 45.305 ;
        RECT 87.49 44.285 87.75 44.545 ;
        RECT 87.49 43.525 87.75 43.785 ;
        RECT 87.49 42.765 87.75 43.025 ;
        RECT 87.49 42.005 87.75 42.265 ;
        RECT 87.49 41.245 87.75 41.505 ;
        RECT 87.49 40.485 87.75 40.745 ;
        RECT 87.49 39.725 87.75 39.985 ;
        RECT 87.49 38.965 87.75 39.225 ;
        RECT 87.49 38.205 87.75 38.465 ;
        RECT 87.49 37.445 87.75 37.705 ;
        RECT 87.49 36.685 87.75 36.945 ;
        RECT 88.25 58.725 88.51 58.985 ;
        RECT 88.25 57.965 88.51 58.225 ;
        RECT 88.25 57.205 88.51 57.465 ;
        RECT 88.25 56.445 88.51 56.705 ;
        RECT 88.25 55.685 88.51 55.945 ;
        RECT 88.25 54.925 88.51 55.185 ;
        RECT 88.25 54.165 88.51 54.425 ;
        RECT 88.25 53.405 88.51 53.665 ;
        RECT 88.25 52.645 88.51 52.905 ;
        RECT 88.25 51.885 88.51 52.145 ;
        RECT 88.25 51.125 88.51 51.385 ;
        RECT 88.25 50.365 88.51 50.625 ;
        RECT 88.25 49.605 88.51 49.865 ;
        RECT 88.25 48.845 88.51 49.105 ;
        RECT 88.25 48.085 88.51 48.345 ;
        RECT 88.25 47.325 88.51 47.585 ;
        RECT 88.25 46.565 88.51 46.825 ;
        RECT 88.25 45.805 88.51 46.065 ;
        RECT 88.25 45.045 88.51 45.305 ;
        RECT 88.25 44.285 88.51 44.545 ;
        RECT 88.25 43.525 88.51 43.785 ;
        RECT 88.25 42.765 88.51 43.025 ;
        RECT 88.25 42.005 88.51 42.265 ;
        RECT 88.25 41.245 88.51 41.505 ;
        RECT 88.25 40.485 88.51 40.745 ;
        RECT 88.25 39.725 88.51 39.985 ;
        RECT 88.25 38.965 88.51 39.225 ;
        RECT 88.25 38.205 88.51 38.465 ;
        RECT 88.25 37.445 88.51 37.705 ;
        RECT 88.25 36.685 88.51 36.945 ;
        RECT 89.01 58.725 89.27 58.985 ;
        RECT 89.01 57.965 89.27 58.225 ;
        RECT 89.01 57.205 89.27 57.465 ;
        RECT 89.01 56.445 89.27 56.705 ;
        RECT 89.01 55.685 89.27 55.945 ;
        RECT 89.01 54.925 89.27 55.185 ;
        RECT 89.01 54.165 89.27 54.425 ;
        RECT 89.01 53.405 89.27 53.665 ;
        RECT 89.01 52.645 89.27 52.905 ;
        RECT 89.01 51.885 89.27 52.145 ;
        RECT 89.01 51.125 89.27 51.385 ;
        RECT 89.01 50.365 89.27 50.625 ;
        RECT 89.01 49.605 89.27 49.865 ;
        RECT 89.01 48.845 89.27 49.105 ;
        RECT 89.01 48.085 89.27 48.345 ;
        RECT 89.01 47.325 89.27 47.585 ;
        RECT 89.01 46.565 89.27 46.825 ;
        RECT 89.01 45.805 89.27 46.065 ;
        RECT 89.01 45.045 89.27 45.305 ;
        RECT 89.01 44.285 89.27 44.545 ;
        RECT 89.01 43.525 89.27 43.785 ;
        RECT 89.01 42.765 89.27 43.025 ;
        RECT 89.01 42.005 89.27 42.265 ;
        RECT 89.01 41.245 89.27 41.505 ;
        RECT 89.01 40.485 89.27 40.745 ;
        RECT 89.01 39.725 89.27 39.985 ;
        RECT 89.01 38.965 89.27 39.225 ;
        RECT 89.01 38.205 89.27 38.465 ;
        RECT 89.01 37.445 89.27 37.705 ;
        RECT 89.01 36.685 89.27 36.945 ;
        RECT 89.77 58.725 90.03 58.985 ;
        RECT 89.77 57.965 90.03 58.225 ;
        RECT 89.77 57.205 90.03 57.465 ;
        RECT 89.77 56.445 90.03 56.705 ;
        RECT 89.77 55.685 90.03 55.945 ;
        RECT 89.77 54.925 90.03 55.185 ;
        RECT 89.77 54.165 90.03 54.425 ;
        RECT 89.77 53.405 90.03 53.665 ;
        RECT 89.77 52.645 90.03 52.905 ;
        RECT 89.77 51.885 90.03 52.145 ;
        RECT 89.77 51.125 90.03 51.385 ;
        RECT 89.77 50.365 90.03 50.625 ;
        RECT 89.77 49.605 90.03 49.865 ;
        RECT 89.77 48.845 90.03 49.105 ;
        RECT 89.77 48.085 90.03 48.345 ;
        RECT 89.77 47.325 90.03 47.585 ;
        RECT 89.77 46.565 90.03 46.825 ;
        RECT 89.77 45.805 90.03 46.065 ;
        RECT 89.77 45.045 90.03 45.305 ;
        RECT 89.77 44.285 90.03 44.545 ;
        RECT 89.77 43.525 90.03 43.785 ;
        RECT 89.77 42.765 90.03 43.025 ;
        RECT 89.77 42.005 90.03 42.265 ;
        RECT 89.77 41.245 90.03 41.505 ;
        RECT 89.77 40.485 90.03 40.745 ;
        RECT 89.77 39.725 90.03 39.985 ;
        RECT 89.77 38.965 90.03 39.225 ;
        RECT 89.77 38.205 90.03 38.465 ;
        RECT 89.77 37.445 90.03 37.705 ;
        RECT 89.77 36.685 90.03 36.945 ;
        RECT 90.53 58.725 90.79 58.985 ;
        RECT 90.53 57.965 90.79 58.225 ;
        RECT 90.53 57.205 90.79 57.465 ;
        RECT 90.53 56.445 90.79 56.705 ;
        RECT 90.53 55.685 90.79 55.945 ;
        RECT 90.53 54.925 90.79 55.185 ;
        RECT 90.53 54.165 90.79 54.425 ;
        RECT 90.53 53.405 90.79 53.665 ;
        RECT 90.53 52.645 90.79 52.905 ;
        RECT 90.53 51.885 90.79 52.145 ;
        RECT 90.53 51.125 90.79 51.385 ;
        RECT 90.53 50.365 90.79 50.625 ;
        RECT 90.53 49.605 90.79 49.865 ;
        RECT 90.53 48.845 90.79 49.105 ;
        RECT 90.53 48.085 90.79 48.345 ;
        RECT 90.53 47.325 90.79 47.585 ;
        RECT 90.53 46.565 90.79 46.825 ;
        RECT 90.53 45.805 90.79 46.065 ;
        RECT 90.53 45.045 90.79 45.305 ;
        RECT 90.53 44.285 90.79 44.545 ;
        RECT 90.53 43.525 90.79 43.785 ;
        RECT 90.53 42.765 90.79 43.025 ;
        RECT 90.53 42.005 90.79 42.265 ;
        RECT 90.53 41.245 90.79 41.505 ;
        RECT 90.53 40.485 90.79 40.745 ;
        RECT 90.53 39.725 90.79 39.985 ;
        RECT 90.53 38.965 90.79 39.225 ;
        RECT 90.53 38.205 90.79 38.465 ;
        RECT 90.53 37.445 90.79 37.705 ;
        RECT 90.53 36.685 90.79 36.945 ;
        RECT 91.29 58.725 91.55 58.985 ;
        RECT 91.29 57.965 91.55 58.225 ;
        RECT 91.29 57.205 91.55 57.465 ;
        RECT 91.29 56.445 91.55 56.705 ;
        RECT 91.29 55.685 91.55 55.945 ;
        RECT 91.29 54.925 91.55 55.185 ;
        RECT 91.29 54.165 91.55 54.425 ;
        RECT 91.29 53.405 91.55 53.665 ;
        RECT 91.29 52.645 91.55 52.905 ;
        RECT 91.29 51.885 91.55 52.145 ;
        RECT 91.29 51.125 91.55 51.385 ;
        RECT 91.29 50.365 91.55 50.625 ;
        RECT 91.29 49.605 91.55 49.865 ;
        RECT 91.29 48.845 91.55 49.105 ;
        RECT 91.29 48.085 91.55 48.345 ;
        RECT 91.29 47.325 91.55 47.585 ;
        RECT 91.29 46.565 91.55 46.825 ;
        RECT 91.29 45.805 91.55 46.065 ;
        RECT 91.29 45.045 91.55 45.305 ;
        RECT 91.29 44.285 91.55 44.545 ;
        RECT 91.29 43.525 91.55 43.785 ;
        RECT 91.29 42.765 91.55 43.025 ;
        RECT 91.29 42.005 91.55 42.265 ;
        RECT 91.29 41.245 91.55 41.505 ;
        RECT 91.29 40.485 91.55 40.745 ;
        RECT 91.29 39.725 91.55 39.985 ;
        RECT 91.29 38.965 91.55 39.225 ;
        RECT 91.29 38.205 91.55 38.465 ;
        RECT 91.29 37.445 91.55 37.705 ;
        RECT 91.29 36.685 91.55 36.945 ;
        RECT 92.05 58.725 92.31 58.985 ;
        RECT 92.05 57.965 92.31 58.225 ;
        RECT 92.05 57.205 92.31 57.465 ;
        RECT 92.05 56.445 92.31 56.705 ;
        RECT 92.05 55.685 92.31 55.945 ;
        RECT 92.05 54.925 92.31 55.185 ;
        RECT 92.05 54.165 92.31 54.425 ;
        RECT 92.05 53.405 92.31 53.665 ;
        RECT 92.05 52.645 92.31 52.905 ;
        RECT 92.05 51.885 92.31 52.145 ;
        RECT 92.05 51.125 92.31 51.385 ;
        RECT 92.05 50.365 92.31 50.625 ;
        RECT 92.05 49.605 92.31 49.865 ;
        RECT 92.05 48.845 92.31 49.105 ;
        RECT 92.05 48.085 92.31 48.345 ;
        RECT 92.05 47.325 92.31 47.585 ;
        RECT 92.05 46.565 92.31 46.825 ;
        RECT 92.05 45.805 92.31 46.065 ;
        RECT 92.05 45.045 92.31 45.305 ;
        RECT 92.05 44.285 92.31 44.545 ;
        RECT 92.05 43.525 92.31 43.785 ;
        RECT 92.05 42.765 92.31 43.025 ;
        RECT 92.05 42.005 92.31 42.265 ;
        RECT 92.05 41.245 92.31 41.505 ;
        RECT 92.05 40.485 92.31 40.745 ;
        RECT 92.05 39.725 92.31 39.985 ;
        RECT 92.05 38.965 92.31 39.225 ;
        RECT 92.05 38.205 92.31 38.465 ;
        RECT 92.05 37.445 92.31 37.705 ;
        RECT 92.05 36.685 92.31 36.945 ;
        RECT 92.81 58.725 93.07 58.985 ;
        RECT 92.81 57.965 93.07 58.225 ;
        RECT 92.81 57.205 93.07 57.465 ;
        RECT 92.81 56.445 93.07 56.705 ;
        RECT 92.81 55.685 93.07 55.945 ;
        RECT 92.81 54.925 93.07 55.185 ;
        RECT 92.81 54.165 93.07 54.425 ;
        RECT 92.81 53.405 93.07 53.665 ;
        RECT 92.81 52.645 93.07 52.905 ;
        RECT 92.81 51.885 93.07 52.145 ;
        RECT 92.81 51.125 93.07 51.385 ;
        RECT 92.81 50.365 93.07 50.625 ;
        RECT 92.81 49.605 93.07 49.865 ;
        RECT 92.81 48.845 93.07 49.105 ;
        RECT 92.81 48.085 93.07 48.345 ;
        RECT 92.81 47.325 93.07 47.585 ;
        RECT 92.81 46.565 93.07 46.825 ;
        RECT 92.81 45.805 93.07 46.065 ;
        RECT 92.81 45.045 93.07 45.305 ;
        RECT 92.81 44.285 93.07 44.545 ;
        RECT 92.81 43.525 93.07 43.785 ;
        RECT 92.81 42.765 93.07 43.025 ;
        RECT 92.81 42.005 93.07 42.265 ;
        RECT 92.81 41.245 93.07 41.505 ;
        RECT 92.81 40.485 93.07 40.745 ;
        RECT 92.81 39.725 93.07 39.985 ;
        RECT 92.81 38.965 93.07 39.225 ;
        RECT 92.81 38.205 93.07 38.465 ;
        RECT 92.81 37.445 93.07 37.705 ;
        RECT 92.81 36.685 93.07 36.945 ;
        RECT 93.57 58.725 93.83 58.985 ;
        RECT 93.57 57.965 93.83 58.225 ;
        RECT 93.57 57.205 93.83 57.465 ;
        RECT 93.57 56.445 93.83 56.705 ;
        RECT 93.57 55.685 93.83 55.945 ;
        RECT 93.57 54.925 93.83 55.185 ;
        RECT 93.57 54.165 93.83 54.425 ;
        RECT 93.57 53.405 93.83 53.665 ;
        RECT 93.57 52.645 93.83 52.905 ;
        RECT 93.57 51.885 93.83 52.145 ;
        RECT 93.57 51.125 93.83 51.385 ;
        RECT 93.57 50.365 93.83 50.625 ;
        RECT 93.57 49.605 93.83 49.865 ;
        RECT 93.57 48.845 93.83 49.105 ;
        RECT 93.57 48.085 93.83 48.345 ;
        RECT 93.57 47.325 93.83 47.585 ;
        RECT 93.57 46.565 93.83 46.825 ;
        RECT 93.57 45.805 93.83 46.065 ;
        RECT 93.57 45.045 93.83 45.305 ;
        RECT 93.57 44.285 93.83 44.545 ;
        RECT 93.57 43.525 93.83 43.785 ;
        RECT 93.57 42.765 93.83 43.025 ;
        RECT 93.57 42.005 93.83 42.265 ;
        RECT 93.57 41.245 93.83 41.505 ;
        RECT 93.57 40.485 93.83 40.745 ;
        RECT 93.57 39.725 93.83 39.985 ;
        RECT 93.57 38.965 93.83 39.225 ;
        RECT 93.57 38.205 93.83 38.465 ;
        RECT 93.57 37.445 93.83 37.705 ;
        RECT 93.57 36.685 93.83 36.945 ;
        RECT 94.33 58.725 94.59 58.985 ;
        RECT 94.33 57.965 94.59 58.225 ;
        RECT 94.33 57.205 94.59 57.465 ;
        RECT 94.33 56.445 94.59 56.705 ;
        RECT 94.33 55.685 94.59 55.945 ;
        RECT 94.33 54.925 94.59 55.185 ;
        RECT 94.33 54.165 94.59 54.425 ;
        RECT 94.33 53.405 94.59 53.665 ;
        RECT 94.33 52.645 94.59 52.905 ;
        RECT 94.33 51.885 94.59 52.145 ;
        RECT 94.33 51.125 94.59 51.385 ;
        RECT 94.33 50.365 94.59 50.625 ;
        RECT 94.33 49.605 94.59 49.865 ;
        RECT 94.33 48.845 94.59 49.105 ;
        RECT 94.33 48.085 94.59 48.345 ;
        RECT 94.33 47.325 94.59 47.585 ;
        RECT 94.33 46.565 94.59 46.825 ;
        RECT 94.33 45.805 94.59 46.065 ;
        RECT 94.33 45.045 94.59 45.305 ;
        RECT 94.33 44.285 94.59 44.545 ;
        RECT 94.33 43.525 94.59 43.785 ;
        RECT 94.33 42.765 94.59 43.025 ;
        RECT 94.33 42.005 94.59 42.265 ;
        RECT 94.33 41.245 94.59 41.505 ;
        RECT 94.33 40.485 94.59 40.745 ;
        RECT 94.33 39.725 94.59 39.985 ;
        RECT 94.33 38.965 94.59 39.225 ;
        RECT 94.33 38.205 94.59 38.465 ;
        RECT 94.33 37.445 94.59 37.705 ;
        RECT 94.33 36.685 94.59 36.945 ;
        RECT 95.09 58.725 95.35 58.985 ;
        RECT 95.09 57.965 95.35 58.225 ;
        RECT 95.09 57.205 95.35 57.465 ;
        RECT 95.09 56.445 95.35 56.705 ;
        RECT 95.09 55.685 95.35 55.945 ;
        RECT 95.09 54.925 95.35 55.185 ;
        RECT 95.09 54.165 95.35 54.425 ;
        RECT 95.09 53.405 95.35 53.665 ;
        RECT 95.09 52.645 95.35 52.905 ;
        RECT 95.09 51.885 95.35 52.145 ;
        RECT 95.09 51.125 95.35 51.385 ;
        RECT 95.09 50.365 95.35 50.625 ;
        RECT 95.09 49.605 95.35 49.865 ;
        RECT 95.09 48.845 95.35 49.105 ;
        RECT 95.09 48.085 95.35 48.345 ;
        RECT 95.09 47.325 95.35 47.585 ;
        RECT 95.09 46.565 95.35 46.825 ;
        RECT 95.09 45.805 95.35 46.065 ;
        RECT 95.09 45.045 95.35 45.305 ;
        RECT 95.09 44.285 95.35 44.545 ;
        RECT 95.09 43.525 95.35 43.785 ;
        RECT 95.09 42.765 95.35 43.025 ;
        RECT 95.09 42.005 95.35 42.265 ;
        RECT 95.09 41.245 95.35 41.505 ;
        RECT 95.09 40.485 95.35 40.745 ;
        RECT 95.09 39.725 95.35 39.985 ;
        RECT 95.09 38.965 95.35 39.225 ;
        RECT 95.09 38.205 95.35 38.465 ;
        RECT 95.09 37.445 95.35 37.705 ;
        RECT 95.09 36.685 95.35 36.945 ;
        RECT 54.81 43.525 55.07 43.785 ;
        RECT 54.81 42.765 55.07 43.025 ;
        RECT 54.81 42.005 55.07 42.265 ;
        RECT 54.81 41.245 55.07 41.505 ;
        RECT 54.81 40.485 55.07 40.745 ;
        RECT 54.81 39.725 55.07 39.985 ;
        RECT 54.81 38.965 55.07 39.225 ;
        RECT 54.81 38.205 55.07 38.465 ;
        RECT 54.81 37.445 55.07 37.705 ;
        RECT 54.81 36.685 55.07 36.945 ;
        RECT 55.57 58.725 55.83 58.985 ;
        RECT 55.57 57.965 55.83 58.225 ;
        RECT 55.57 57.205 55.83 57.465 ;
        RECT 55.57 56.445 55.83 56.705 ;
        RECT 55.57 55.685 55.83 55.945 ;
        RECT 55.57 54.925 55.83 55.185 ;
        RECT 55.57 54.165 55.83 54.425 ;
        RECT 55.57 53.405 55.83 53.665 ;
        RECT 55.57 52.645 55.83 52.905 ;
        RECT 55.57 51.885 55.83 52.145 ;
        RECT 55.57 51.125 55.83 51.385 ;
        RECT 55.57 50.365 55.83 50.625 ;
        RECT 55.57 49.605 55.83 49.865 ;
        RECT 55.57 48.845 55.83 49.105 ;
        RECT 55.57 48.085 55.83 48.345 ;
        RECT 55.57 47.325 55.83 47.585 ;
        RECT 55.57 46.565 55.83 46.825 ;
        RECT 55.57 45.805 55.83 46.065 ;
        RECT 55.57 45.045 55.83 45.305 ;
        RECT 55.57 44.285 55.83 44.545 ;
        RECT 55.57 43.525 55.83 43.785 ;
        RECT 55.57 42.765 55.83 43.025 ;
        RECT 55.57 42.005 55.83 42.265 ;
        RECT 55.57 41.245 55.83 41.505 ;
        RECT 55.57 40.485 55.83 40.745 ;
        RECT 55.57 39.725 55.83 39.985 ;
        RECT 55.57 38.965 55.83 39.225 ;
        RECT 55.57 38.205 55.83 38.465 ;
        RECT 55.57 37.445 55.83 37.705 ;
        RECT 55.57 36.685 55.83 36.945 ;
        RECT 56.33 58.725 56.59 58.985 ;
        RECT 56.33 57.965 56.59 58.225 ;
        RECT 56.33 57.205 56.59 57.465 ;
        RECT 56.33 56.445 56.59 56.705 ;
        RECT 56.33 55.685 56.59 55.945 ;
        RECT 56.33 54.925 56.59 55.185 ;
        RECT 56.33 54.165 56.59 54.425 ;
        RECT 56.33 53.405 56.59 53.665 ;
        RECT 56.33 52.645 56.59 52.905 ;
        RECT 56.33 51.885 56.59 52.145 ;
        RECT 56.33 51.125 56.59 51.385 ;
        RECT 56.33 50.365 56.59 50.625 ;
        RECT 56.33 49.605 56.59 49.865 ;
        RECT 56.33 48.845 56.59 49.105 ;
        RECT 56.33 48.085 56.59 48.345 ;
        RECT 56.33 47.325 56.59 47.585 ;
        RECT 56.33 46.565 56.59 46.825 ;
        RECT 56.33 45.805 56.59 46.065 ;
        RECT 56.33 45.045 56.59 45.305 ;
        RECT 56.33 44.285 56.59 44.545 ;
        RECT 56.33 43.525 56.59 43.785 ;
        RECT 56.33 42.765 56.59 43.025 ;
        RECT 56.33 42.005 56.59 42.265 ;
        RECT 56.33 41.245 56.59 41.505 ;
        RECT 56.33 40.485 56.59 40.745 ;
        RECT 56.33 39.725 56.59 39.985 ;
        RECT 56.33 38.965 56.59 39.225 ;
        RECT 56.33 38.205 56.59 38.465 ;
        RECT 56.33 37.445 56.59 37.705 ;
        RECT 56.33 36.685 56.59 36.945 ;
        RECT 57.09 58.725 57.35 58.985 ;
        RECT 57.09 57.965 57.35 58.225 ;
        RECT 57.09 57.205 57.35 57.465 ;
        RECT 57.09 56.445 57.35 56.705 ;
        RECT 57.09 55.685 57.35 55.945 ;
        RECT 57.09 54.925 57.35 55.185 ;
        RECT 57.09 54.165 57.35 54.425 ;
        RECT 57.09 53.405 57.35 53.665 ;
        RECT 57.09 52.645 57.35 52.905 ;
        RECT 57.09 51.885 57.35 52.145 ;
        RECT 57.09 51.125 57.35 51.385 ;
        RECT 57.09 50.365 57.35 50.625 ;
        RECT 57.09 49.605 57.35 49.865 ;
        RECT 57.09 48.845 57.35 49.105 ;
        RECT 57.09 48.085 57.35 48.345 ;
        RECT 57.09 47.325 57.35 47.585 ;
        RECT 57.09 46.565 57.35 46.825 ;
        RECT 57.09 45.805 57.35 46.065 ;
        RECT 57.09 45.045 57.35 45.305 ;
        RECT 57.09 44.285 57.35 44.545 ;
        RECT 57.09 43.525 57.35 43.785 ;
        RECT 57.09 42.765 57.35 43.025 ;
        RECT 57.09 42.005 57.35 42.265 ;
        RECT 57.09 41.245 57.35 41.505 ;
        RECT 57.09 40.485 57.35 40.745 ;
        RECT 57.09 39.725 57.35 39.985 ;
        RECT 57.09 38.965 57.35 39.225 ;
        RECT 57.09 38.205 57.35 38.465 ;
        RECT 57.09 37.445 57.35 37.705 ;
        RECT 57.09 36.685 57.35 36.945 ;
        RECT 57.85 58.725 58.11 58.985 ;
        RECT 57.85 57.965 58.11 58.225 ;
        RECT 57.85 57.205 58.11 57.465 ;
        RECT 57.85 56.445 58.11 56.705 ;
        RECT 57.85 55.685 58.11 55.945 ;
        RECT 57.85 54.925 58.11 55.185 ;
        RECT 57.85 54.165 58.11 54.425 ;
        RECT 57.85 53.405 58.11 53.665 ;
        RECT 57.85 52.645 58.11 52.905 ;
        RECT 57.85 51.885 58.11 52.145 ;
        RECT 57.85 51.125 58.11 51.385 ;
        RECT 57.85 50.365 58.11 50.625 ;
        RECT 57.85 49.605 58.11 49.865 ;
        RECT 57.85 48.845 58.11 49.105 ;
        RECT 57.85 48.085 58.11 48.345 ;
        RECT 57.85 47.325 58.11 47.585 ;
        RECT 57.85 46.565 58.11 46.825 ;
        RECT 57.85 45.805 58.11 46.065 ;
        RECT 57.85 45.045 58.11 45.305 ;
        RECT 57.85 44.285 58.11 44.545 ;
        RECT 57.85 43.525 58.11 43.785 ;
        RECT 57.85 42.765 58.11 43.025 ;
        RECT 57.85 42.005 58.11 42.265 ;
        RECT 57.85 41.245 58.11 41.505 ;
        RECT 57.85 40.485 58.11 40.745 ;
        RECT 57.85 39.725 58.11 39.985 ;
        RECT 57.85 38.965 58.11 39.225 ;
        RECT 57.85 38.205 58.11 38.465 ;
        RECT 57.85 37.445 58.11 37.705 ;
        RECT 57.85 36.685 58.11 36.945 ;
        RECT 58.61 58.725 58.87 58.985 ;
        RECT 58.61 57.965 58.87 58.225 ;
        RECT 58.61 57.205 58.87 57.465 ;
        RECT 58.61 56.445 58.87 56.705 ;
        RECT 58.61 55.685 58.87 55.945 ;
        RECT 58.61 54.925 58.87 55.185 ;
        RECT 58.61 54.165 58.87 54.425 ;
        RECT 58.61 53.405 58.87 53.665 ;
        RECT 58.61 52.645 58.87 52.905 ;
        RECT 58.61 51.885 58.87 52.145 ;
        RECT 58.61 51.125 58.87 51.385 ;
        RECT 58.61 50.365 58.87 50.625 ;
        RECT 58.61 49.605 58.87 49.865 ;
        RECT 58.61 48.845 58.87 49.105 ;
        RECT 58.61 48.085 58.87 48.345 ;
        RECT 58.61 47.325 58.87 47.585 ;
        RECT 58.61 46.565 58.87 46.825 ;
        RECT 58.61 45.805 58.87 46.065 ;
        RECT 58.61 45.045 58.87 45.305 ;
        RECT 58.61 44.285 58.87 44.545 ;
        RECT 58.61 43.525 58.87 43.785 ;
        RECT 58.61 42.765 58.87 43.025 ;
        RECT 58.61 42.005 58.87 42.265 ;
        RECT 58.61 41.245 58.87 41.505 ;
        RECT 58.61 40.485 58.87 40.745 ;
        RECT 58.61 39.725 58.87 39.985 ;
        RECT 58.61 38.965 58.87 39.225 ;
        RECT 58.61 38.205 58.87 38.465 ;
        RECT 58.61 37.445 58.87 37.705 ;
        RECT 58.61 36.685 58.87 36.945 ;
        RECT 59.37 58.725 59.63 58.985 ;
        RECT 59.37 57.965 59.63 58.225 ;
        RECT 59.37 57.205 59.63 57.465 ;
        RECT 59.37 56.445 59.63 56.705 ;
        RECT 59.37 55.685 59.63 55.945 ;
        RECT 59.37 54.925 59.63 55.185 ;
        RECT 59.37 54.165 59.63 54.425 ;
        RECT 59.37 53.405 59.63 53.665 ;
        RECT 59.37 52.645 59.63 52.905 ;
        RECT 59.37 51.885 59.63 52.145 ;
        RECT 59.37 51.125 59.63 51.385 ;
        RECT 59.37 50.365 59.63 50.625 ;
        RECT 59.37 49.605 59.63 49.865 ;
        RECT 59.37 48.845 59.63 49.105 ;
        RECT 59.37 48.085 59.63 48.345 ;
        RECT 59.37 47.325 59.63 47.585 ;
        RECT 59.37 46.565 59.63 46.825 ;
        RECT 59.37 45.805 59.63 46.065 ;
        RECT 59.37 45.045 59.63 45.305 ;
        RECT 59.37 44.285 59.63 44.545 ;
        RECT 59.37 43.525 59.63 43.785 ;
        RECT 59.37 42.765 59.63 43.025 ;
        RECT 59.37 42.005 59.63 42.265 ;
        RECT 59.37 41.245 59.63 41.505 ;
        RECT 59.37 40.485 59.63 40.745 ;
        RECT 59.37 39.725 59.63 39.985 ;
        RECT 59.37 38.965 59.63 39.225 ;
        RECT 59.37 38.205 59.63 38.465 ;
        RECT 59.37 37.445 59.63 37.705 ;
        RECT 59.37 36.685 59.63 36.945 ;
        RECT 60.13 58.725 60.39 58.985 ;
        RECT 60.13 57.965 60.39 58.225 ;
        RECT 60.13 57.205 60.39 57.465 ;
        RECT 60.13 56.445 60.39 56.705 ;
        RECT 60.13 55.685 60.39 55.945 ;
        RECT 60.13 54.925 60.39 55.185 ;
        RECT 60.13 54.165 60.39 54.425 ;
        RECT 60.13 53.405 60.39 53.665 ;
        RECT 60.13 52.645 60.39 52.905 ;
        RECT 60.13 51.885 60.39 52.145 ;
        RECT 60.13 51.125 60.39 51.385 ;
        RECT 60.13 50.365 60.39 50.625 ;
        RECT 60.13 49.605 60.39 49.865 ;
        RECT 60.13 48.845 60.39 49.105 ;
        RECT 60.13 48.085 60.39 48.345 ;
        RECT 60.13 47.325 60.39 47.585 ;
        RECT 60.13 46.565 60.39 46.825 ;
        RECT 60.13 45.805 60.39 46.065 ;
        RECT 60.13 45.045 60.39 45.305 ;
        RECT 60.13 44.285 60.39 44.545 ;
        RECT 60.13 43.525 60.39 43.785 ;
        RECT 60.13 42.765 60.39 43.025 ;
        RECT 60.13 42.005 60.39 42.265 ;
        RECT 60.13 41.245 60.39 41.505 ;
        RECT 60.13 40.485 60.39 40.745 ;
        RECT 60.13 39.725 60.39 39.985 ;
        RECT 60.13 38.965 60.39 39.225 ;
        RECT 60.13 38.205 60.39 38.465 ;
        RECT 60.13 37.445 60.39 37.705 ;
        RECT 60.13 36.685 60.39 36.945 ;
        RECT 60.89 58.725 61.15 58.985 ;
        RECT 60.89 57.965 61.15 58.225 ;
        RECT 60.89 57.205 61.15 57.465 ;
        RECT 60.89 56.445 61.15 56.705 ;
        RECT 60.89 55.685 61.15 55.945 ;
        RECT 60.89 54.925 61.15 55.185 ;
        RECT 60.89 54.165 61.15 54.425 ;
        RECT 60.89 53.405 61.15 53.665 ;
        RECT 60.89 52.645 61.15 52.905 ;
        RECT 60.89 51.885 61.15 52.145 ;
        RECT 60.89 51.125 61.15 51.385 ;
        RECT 60.89 50.365 61.15 50.625 ;
        RECT 60.89 49.605 61.15 49.865 ;
        RECT 60.89 48.845 61.15 49.105 ;
        RECT 60.89 48.085 61.15 48.345 ;
        RECT 60.89 47.325 61.15 47.585 ;
        RECT 60.89 46.565 61.15 46.825 ;
        RECT 60.89 45.805 61.15 46.065 ;
        RECT 60.89 45.045 61.15 45.305 ;
        RECT 60.89 44.285 61.15 44.545 ;
        RECT 60.89 43.525 61.15 43.785 ;
        RECT 60.89 42.765 61.15 43.025 ;
        RECT 60.89 42.005 61.15 42.265 ;
        RECT 60.89 41.245 61.15 41.505 ;
        RECT 60.89 40.485 61.15 40.745 ;
        RECT 60.89 39.725 61.15 39.985 ;
        RECT 60.89 38.965 61.15 39.225 ;
        RECT 60.89 38.205 61.15 38.465 ;
        RECT 60.89 37.445 61.15 37.705 ;
        RECT 60.89 36.685 61.15 36.945 ;
        RECT 61.65 58.725 61.91 58.985 ;
        RECT 61.65 57.965 61.91 58.225 ;
        RECT 61.65 57.205 61.91 57.465 ;
        RECT 61.65 56.445 61.91 56.705 ;
        RECT 61.65 55.685 61.91 55.945 ;
        RECT 61.65 54.925 61.91 55.185 ;
        RECT 61.65 54.165 61.91 54.425 ;
        RECT 61.65 53.405 61.91 53.665 ;
        RECT 61.65 52.645 61.91 52.905 ;
        RECT 61.65 51.885 61.91 52.145 ;
        RECT 61.65 51.125 61.91 51.385 ;
        RECT 61.65 50.365 61.91 50.625 ;
        RECT 61.65 49.605 61.91 49.865 ;
        RECT 61.65 48.845 61.91 49.105 ;
        RECT 61.65 48.085 61.91 48.345 ;
        RECT 61.65 47.325 61.91 47.585 ;
        RECT 61.65 46.565 61.91 46.825 ;
        RECT 61.65 45.805 61.91 46.065 ;
        RECT 61.65 45.045 61.91 45.305 ;
        RECT 61.65 44.285 61.91 44.545 ;
        RECT 61.65 43.525 61.91 43.785 ;
        RECT 61.65 42.765 61.91 43.025 ;
        RECT 61.65 42.005 61.91 42.265 ;
        RECT 61.65 41.245 61.91 41.505 ;
        RECT 61.65 40.485 61.91 40.745 ;
        RECT 61.65 39.725 61.91 39.985 ;
        RECT 61.65 38.965 61.91 39.225 ;
        RECT 61.65 38.205 61.91 38.465 ;
        RECT 61.65 37.445 61.91 37.705 ;
        RECT 61.65 36.685 61.91 36.945 ;
        RECT 62.41 58.725 62.67 58.985 ;
        RECT 62.41 57.965 62.67 58.225 ;
        RECT 62.41 57.205 62.67 57.465 ;
        RECT 62.41 56.445 62.67 56.705 ;
        RECT 62.41 55.685 62.67 55.945 ;
        RECT 62.41 54.925 62.67 55.185 ;
        RECT 62.41 54.165 62.67 54.425 ;
        RECT 62.41 53.405 62.67 53.665 ;
        RECT 62.41 52.645 62.67 52.905 ;
        RECT 62.41 51.885 62.67 52.145 ;
        RECT 62.41 51.125 62.67 51.385 ;
        RECT 62.41 50.365 62.67 50.625 ;
        RECT 62.41 49.605 62.67 49.865 ;
        RECT 62.41 48.845 62.67 49.105 ;
        RECT 62.41 48.085 62.67 48.345 ;
        RECT 62.41 47.325 62.67 47.585 ;
        RECT 62.41 46.565 62.67 46.825 ;
        RECT 62.41 45.805 62.67 46.065 ;
        RECT 62.41 45.045 62.67 45.305 ;
        RECT 62.41 44.285 62.67 44.545 ;
        RECT 62.41 43.525 62.67 43.785 ;
        RECT 62.41 42.765 62.67 43.025 ;
        RECT 62.41 42.005 62.67 42.265 ;
        RECT 62.41 41.245 62.67 41.505 ;
        RECT 62.41 40.485 62.67 40.745 ;
        RECT 62.41 39.725 62.67 39.985 ;
        RECT 62.41 38.965 62.67 39.225 ;
        RECT 62.41 38.205 62.67 38.465 ;
        RECT 62.41 37.445 62.67 37.705 ;
        RECT 62.41 36.685 62.67 36.945 ;
        RECT 63.17 58.725 63.43 58.985 ;
        RECT 63.17 57.965 63.43 58.225 ;
        RECT 63.17 57.205 63.43 57.465 ;
        RECT 63.17 56.445 63.43 56.705 ;
        RECT 63.17 55.685 63.43 55.945 ;
        RECT 63.17 54.925 63.43 55.185 ;
        RECT 63.17 54.165 63.43 54.425 ;
        RECT 63.17 53.405 63.43 53.665 ;
        RECT 63.17 52.645 63.43 52.905 ;
        RECT 63.17 51.885 63.43 52.145 ;
        RECT 63.17 51.125 63.43 51.385 ;
        RECT 63.17 50.365 63.43 50.625 ;
        RECT 63.17 49.605 63.43 49.865 ;
        RECT 63.17 48.845 63.43 49.105 ;
        RECT 63.17 48.085 63.43 48.345 ;
        RECT 63.17 47.325 63.43 47.585 ;
        RECT 63.17 46.565 63.43 46.825 ;
        RECT 63.17 45.805 63.43 46.065 ;
        RECT 63.17 45.045 63.43 45.305 ;
        RECT 63.17 44.285 63.43 44.545 ;
        RECT 63.17 43.525 63.43 43.785 ;
        RECT 63.17 42.765 63.43 43.025 ;
        RECT 63.17 42.005 63.43 42.265 ;
        RECT 63.17 41.245 63.43 41.505 ;
        RECT 63.17 40.485 63.43 40.745 ;
        RECT 63.17 39.725 63.43 39.985 ;
        RECT 63.17 38.965 63.43 39.225 ;
        RECT 63.17 38.205 63.43 38.465 ;
        RECT 63.17 37.445 63.43 37.705 ;
        RECT 63.17 36.685 63.43 36.945 ;
        RECT 63.93 58.725 64.19 58.985 ;
        RECT 63.93 57.965 64.19 58.225 ;
        RECT 63.93 57.205 64.19 57.465 ;
        RECT 63.93 56.445 64.19 56.705 ;
        RECT 63.93 55.685 64.19 55.945 ;
        RECT 63.93 54.925 64.19 55.185 ;
        RECT 63.93 54.165 64.19 54.425 ;
        RECT 63.93 53.405 64.19 53.665 ;
        RECT 63.93 52.645 64.19 52.905 ;
        RECT 63.93 51.885 64.19 52.145 ;
        RECT 63.93 51.125 64.19 51.385 ;
        RECT 63.93 50.365 64.19 50.625 ;
        RECT 63.93 49.605 64.19 49.865 ;
        RECT 63.93 48.845 64.19 49.105 ;
        RECT 63.93 48.085 64.19 48.345 ;
        RECT 63.93 47.325 64.19 47.585 ;
        RECT 63.93 46.565 64.19 46.825 ;
        RECT 63.93 45.805 64.19 46.065 ;
        RECT 63.93 45.045 64.19 45.305 ;
        RECT 63.93 44.285 64.19 44.545 ;
        RECT 63.93 43.525 64.19 43.785 ;
        RECT 63.93 42.765 64.19 43.025 ;
        RECT 63.93 42.005 64.19 42.265 ;
        RECT 63.93 41.245 64.19 41.505 ;
        RECT 63.93 40.485 64.19 40.745 ;
        RECT 63.93 39.725 64.19 39.985 ;
        RECT 63.93 38.965 64.19 39.225 ;
        RECT 63.93 38.205 64.19 38.465 ;
        RECT 63.93 37.445 64.19 37.705 ;
        RECT 63.93 36.685 64.19 36.945 ;
        RECT 64.69 58.725 64.95 58.985 ;
        RECT 64.69 57.965 64.95 58.225 ;
        RECT 64.69 57.205 64.95 57.465 ;
        RECT 64.69 56.445 64.95 56.705 ;
        RECT 64.69 55.685 64.95 55.945 ;
        RECT 64.69 54.925 64.95 55.185 ;
        RECT 64.69 54.165 64.95 54.425 ;
        RECT 64.69 53.405 64.95 53.665 ;
        RECT 64.69 52.645 64.95 52.905 ;
        RECT 64.69 51.885 64.95 52.145 ;
        RECT 64.69 51.125 64.95 51.385 ;
        RECT 64.69 50.365 64.95 50.625 ;
        RECT 64.69 49.605 64.95 49.865 ;
        RECT 64.69 48.845 64.95 49.105 ;
        RECT 64.69 48.085 64.95 48.345 ;
        RECT 64.69 47.325 64.95 47.585 ;
        RECT 64.69 46.565 64.95 46.825 ;
        RECT 64.69 45.805 64.95 46.065 ;
        RECT 64.69 45.045 64.95 45.305 ;
        RECT 64.69 44.285 64.95 44.545 ;
        RECT 64.69 43.525 64.95 43.785 ;
        RECT 64.69 42.765 64.95 43.025 ;
        RECT 64.69 42.005 64.95 42.265 ;
        RECT 64.69 41.245 64.95 41.505 ;
        RECT 64.69 40.485 64.95 40.745 ;
        RECT 64.69 39.725 64.95 39.985 ;
        RECT 64.69 38.965 64.95 39.225 ;
        RECT 64.69 38.205 64.95 38.465 ;
        RECT 64.69 37.445 64.95 37.705 ;
        RECT 64.69 36.685 64.95 36.945 ;
        RECT 65.45 58.725 65.71 58.985 ;
        RECT 65.45 57.965 65.71 58.225 ;
        RECT 65.45 57.205 65.71 57.465 ;
        RECT 65.45 56.445 65.71 56.705 ;
        RECT 65.45 55.685 65.71 55.945 ;
        RECT 65.45 54.925 65.71 55.185 ;
        RECT 65.45 54.165 65.71 54.425 ;
        RECT 65.45 53.405 65.71 53.665 ;
        RECT 65.45 52.645 65.71 52.905 ;
        RECT 65.45 51.885 65.71 52.145 ;
        RECT 65.45 51.125 65.71 51.385 ;
        RECT 65.45 50.365 65.71 50.625 ;
        RECT 65.45 49.605 65.71 49.865 ;
        RECT 65.45 48.845 65.71 49.105 ;
        RECT 65.45 48.085 65.71 48.345 ;
        RECT 65.45 47.325 65.71 47.585 ;
        RECT 65.45 46.565 65.71 46.825 ;
        RECT 65.45 45.805 65.71 46.065 ;
        RECT 65.45 45.045 65.71 45.305 ;
        RECT 65.45 44.285 65.71 44.545 ;
        RECT 65.45 43.525 65.71 43.785 ;
        RECT 65.45 42.765 65.71 43.025 ;
        RECT 65.45 42.005 65.71 42.265 ;
        RECT 65.45 41.245 65.71 41.505 ;
        RECT 65.45 40.485 65.71 40.745 ;
        RECT 65.45 39.725 65.71 39.985 ;
        RECT 65.45 38.965 65.71 39.225 ;
        RECT 65.45 38.205 65.71 38.465 ;
        RECT 65.45 37.445 65.71 37.705 ;
        RECT 65.45 36.685 65.71 36.945 ;
        RECT 66.21 58.725 66.47 58.985 ;
        RECT 66.21 57.965 66.47 58.225 ;
        RECT 66.21 57.205 66.47 57.465 ;
        RECT 66.21 56.445 66.47 56.705 ;
        RECT 66.21 55.685 66.47 55.945 ;
        RECT 66.21 54.925 66.47 55.185 ;
        RECT 66.21 54.165 66.47 54.425 ;
        RECT 66.21 53.405 66.47 53.665 ;
        RECT 66.21 52.645 66.47 52.905 ;
        RECT 66.21 51.885 66.47 52.145 ;
        RECT 66.21 51.125 66.47 51.385 ;
        RECT 66.21 50.365 66.47 50.625 ;
        RECT 66.21 49.605 66.47 49.865 ;
        RECT 66.21 48.845 66.47 49.105 ;
        RECT 66.21 48.085 66.47 48.345 ;
        RECT 66.21 47.325 66.47 47.585 ;
        RECT 66.21 46.565 66.47 46.825 ;
        RECT 66.21 45.805 66.47 46.065 ;
        RECT 66.21 45.045 66.47 45.305 ;
        RECT 66.21 44.285 66.47 44.545 ;
        RECT 66.21 43.525 66.47 43.785 ;
        RECT 66.21 42.765 66.47 43.025 ;
        RECT 66.21 42.005 66.47 42.265 ;
        RECT 66.21 41.245 66.47 41.505 ;
        RECT 66.21 40.485 66.47 40.745 ;
        RECT 66.21 39.725 66.47 39.985 ;
        RECT 66.21 38.965 66.47 39.225 ;
        RECT 66.21 38.205 66.47 38.465 ;
        RECT 66.21 37.445 66.47 37.705 ;
        RECT 66.21 36.685 66.47 36.945 ;
        RECT 66.97 58.725 67.23 58.985 ;
        RECT 66.97 57.965 67.23 58.225 ;
        RECT 66.97 57.205 67.23 57.465 ;
        RECT 66.97 56.445 67.23 56.705 ;
        RECT 66.97 55.685 67.23 55.945 ;
        RECT 66.97 54.925 67.23 55.185 ;
        RECT 66.97 54.165 67.23 54.425 ;
        RECT 66.97 53.405 67.23 53.665 ;
        RECT 66.97 52.645 67.23 52.905 ;
        RECT 66.97 51.885 67.23 52.145 ;
        RECT 66.97 51.125 67.23 51.385 ;
        RECT 66.97 50.365 67.23 50.625 ;
        RECT 66.97 49.605 67.23 49.865 ;
        RECT 66.97 48.845 67.23 49.105 ;
        RECT 66.97 48.085 67.23 48.345 ;
        RECT 66.97 47.325 67.23 47.585 ;
        RECT 66.97 46.565 67.23 46.825 ;
        RECT 66.97 45.805 67.23 46.065 ;
        RECT 66.97 45.045 67.23 45.305 ;
        RECT 66.97 44.285 67.23 44.545 ;
        RECT 66.97 43.525 67.23 43.785 ;
        RECT 66.97 42.765 67.23 43.025 ;
        RECT 66.97 42.005 67.23 42.265 ;
        RECT 66.97 41.245 67.23 41.505 ;
        RECT 66.97 40.485 67.23 40.745 ;
        RECT 66.97 39.725 67.23 39.985 ;
        RECT 66.97 38.965 67.23 39.225 ;
        RECT 66.97 38.205 67.23 38.465 ;
        RECT 66.97 37.445 67.23 37.705 ;
        RECT 66.97 36.685 67.23 36.945 ;
        RECT 67.73 58.725 67.99 58.985 ;
        RECT 67.73 57.965 67.99 58.225 ;
        RECT 67.73 57.205 67.99 57.465 ;
        RECT 67.73 56.445 67.99 56.705 ;
        RECT 67.73 55.685 67.99 55.945 ;
        RECT 67.73 54.925 67.99 55.185 ;
        RECT 67.73 54.165 67.99 54.425 ;
        RECT 67.73 53.405 67.99 53.665 ;
        RECT 67.73 52.645 67.99 52.905 ;
        RECT 67.73 51.885 67.99 52.145 ;
        RECT 67.73 51.125 67.99 51.385 ;
        RECT 67.73 50.365 67.99 50.625 ;
        RECT 67.73 49.605 67.99 49.865 ;
        RECT 67.73 48.845 67.99 49.105 ;
        RECT 67.73 48.085 67.99 48.345 ;
        RECT 67.73 47.325 67.99 47.585 ;
        RECT 67.73 46.565 67.99 46.825 ;
        RECT 67.73 45.805 67.99 46.065 ;
        RECT 67.73 45.045 67.99 45.305 ;
        RECT 67.73 44.285 67.99 44.545 ;
        RECT 67.73 43.525 67.99 43.785 ;
        RECT 67.73 42.765 67.99 43.025 ;
        RECT 67.73 42.005 67.99 42.265 ;
        RECT 67.73 41.245 67.99 41.505 ;
        RECT 67.73 40.485 67.99 40.745 ;
        RECT 67.73 39.725 67.99 39.985 ;
        RECT 67.73 38.965 67.99 39.225 ;
        RECT 67.73 38.205 67.99 38.465 ;
        RECT 67.73 37.445 67.99 37.705 ;
        RECT 67.73 36.685 67.99 36.945 ;
        RECT 68.49 58.725 68.75 58.985 ;
        RECT 68.49 57.965 68.75 58.225 ;
        RECT 68.49 57.205 68.75 57.465 ;
        RECT 68.49 56.445 68.75 56.705 ;
        RECT 68.49 55.685 68.75 55.945 ;
        RECT 68.49 54.925 68.75 55.185 ;
        RECT 68.49 54.165 68.75 54.425 ;
        RECT 68.49 53.405 68.75 53.665 ;
        RECT 68.49 52.645 68.75 52.905 ;
        RECT 68.49 51.885 68.75 52.145 ;
        RECT 68.49 51.125 68.75 51.385 ;
        RECT 68.49 50.365 68.75 50.625 ;
        RECT 68.49 49.605 68.75 49.865 ;
        RECT 68.49 48.845 68.75 49.105 ;
        RECT 68.49 48.085 68.75 48.345 ;
        RECT 68.49 47.325 68.75 47.585 ;
        RECT 68.49 46.565 68.75 46.825 ;
        RECT 68.49 45.805 68.75 46.065 ;
        RECT 68.49 45.045 68.75 45.305 ;
        RECT 68.49 44.285 68.75 44.545 ;
        RECT 68.49 43.525 68.75 43.785 ;
        RECT 68.49 42.765 68.75 43.025 ;
        RECT 68.49 42.005 68.75 42.265 ;
        RECT 68.49 41.245 68.75 41.505 ;
        RECT 68.49 40.485 68.75 40.745 ;
        RECT 68.49 39.725 68.75 39.985 ;
        RECT 68.49 38.965 68.75 39.225 ;
        RECT 68.49 38.205 68.75 38.465 ;
        RECT 68.49 37.445 68.75 37.705 ;
        RECT 68.49 36.685 68.75 36.945 ;
        RECT 69.25 58.725 69.51 58.985 ;
        RECT 69.25 57.965 69.51 58.225 ;
        RECT 69.25 57.205 69.51 57.465 ;
        RECT 69.25 56.445 69.51 56.705 ;
        RECT 69.25 55.685 69.51 55.945 ;
        RECT 69.25 54.925 69.51 55.185 ;
        RECT 69.25 54.165 69.51 54.425 ;
        RECT 69.25 53.405 69.51 53.665 ;
        RECT 69.25 52.645 69.51 52.905 ;
        RECT 69.25 51.885 69.51 52.145 ;
        RECT 69.25 51.125 69.51 51.385 ;
        RECT 69.25 50.365 69.51 50.625 ;
        RECT 69.25 49.605 69.51 49.865 ;
        RECT 69.25 48.845 69.51 49.105 ;
        RECT 69.25 48.085 69.51 48.345 ;
        RECT 69.25 47.325 69.51 47.585 ;
        RECT 69.25 46.565 69.51 46.825 ;
        RECT 69.25 45.805 69.51 46.065 ;
        RECT 69.25 45.045 69.51 45.305 ;
        RECT 69.25 44.285 69.51 44.545 ;
        RECT 69.25 43.525 69.51 43.785 ;
        RECT 69.25 42.765 69.51 43.025 ;
        RECT 69.25 42.005 69.51 42.265 ;
        RECT 69.25 41.245 69.51 41.505 ;
        RECT 69.25 40.485 69.51 40.745 ;
        RECT 69.25 39.725 69.51 39.985 ;
        RECT 69.25 38.965 69.51 39.225 ;
        RECT 69.25 38.205 69.51 38.465 ;
        RECT 69.25 37.445 69.51 37.705 ;
        RECT 69.25 36.685 69.51 36.945 ;
        RECT 70.01 58.725 70.27 58.985 ;
        RECT 70.01 57.965 70.27 58.225 ;
        RECT 70.01 57.205 70.27 57.465 ;
        RECT 70.01 56.445 70.27 56.705 ;
        RECT 70.01 55.685 70.27 55.945 ;
        RECT 70.01 54.925 70.27 55.185 ;
        RECT 70.01 54.165 70.27 54.425 ;
        RECT 70.01 53.405 70.27 53.665 ;
        RECT 70.01 52.645 70.27 52.905 ;
        RECT 70.01 51.885 70.27 52.145 ;
        RECT 70.01 51.125 70.27 51.385 ;
        RECT 70.01 50.365 70.27 50.625 ;
        RECT 70.01 49.605 70.27 49.865 ;
        RECT 70.01 48.845 70.27 49.105 ;
        RECT 70.01 48.085 70.27 48.345 ;
        RECT 70.01 47.325 70.27 47.585 ;
        RECT 70.01 46.565 70.27 46.825 ;
        RECT 70.01 45.805 70.27 46.065 ;
        RECT 70.01 45.045 70.27 45.305 ;
        RECT 70.01 44.285 70.27 44.545 ;
        RECT 70.01 43.525 70.27 43.785 ;
        RECT 70.01 42.765 70.27 43.025 ;
        RECT 70.01 42.005 70.27 42.265 ;
        RECT 70.01 41.245 70.27 41.505 ;
        RECT 70.01 40.485 70.27 40.745 ;
        RECT 70.01 39.725 70.27 39.985 ;
        RECT 70.01 38.965 70.27 39.225 ;
        RECT 70.01 38.205 70.27 38.465 ;
        RECT 70.01 37.445 70.27 37.705 ;
        RECT 70.01 36.685 70.27 36.945 ;
        RECT 70.77 58.725 71.03 58.985 ;
        RECT 70.77 57.965 71.03 58.225 ;
        RECT 70.77 57.205 71.03 57.465 ;
        RECT 70.77 56.445 71.03 56.705 ;
        RECT 70.77 55.685 71.03 55.945 ;
        RECT 70.77 54.925 71.03 55.185 ;
        RECT 70.77 54.165 71.03 54.425 ;
        RECT 70.77 53.405 71.03 53.665 ;
        RECT 70.77 52.645 71.03 52.905 ;
        RECT 70.77 51.885 71.03 52.145 ;
        RECT 70.77 51.125 71.03 51.385 ;
        RECT 70.77 50.365 71.03 50.625 ;
        RECT 70.77 49.605 71.03 49.865 ;
        RECT 70.77 48.845 71.03 49.105 ;
        RECT 70.77 48.085 71.03 48.345 ;
        RECT 70.77 47.325 71.03 47.585 ;
        RECT 70.77 46.565 71.03 46.825 ;
        RECT 70.77 45.805 71.03 46.065 ;
        RECT 70.77 45.045 71.03 45.305 ;
        RECT 70.77 44.285 71.03 44.545 ;
        RECT 70.77 43.525 71.03 43.785 ;
        RECT 70.77 42.765 71.03 43.025 ;
        RECT 70.77 42.005 71.03 42.265 ;
        RECT 70.77 41.245 71.03 41.505 ;
        RECT 70.77 40.485 71.03 40.745 ;
        RECT 70.77 39.725 71.03 39.985 ;
        RECT 70.77 38.965 71.03 39.225 ;
        RECT 70.77 38.205 71.03 38.465 ;
        RECT 70.77 37.445 71.03 37.705 ;
        RECT 70.77 36.685 71.03 36.945 ;
        RECT 71.53 58.725 71.79 58.985 ;
        RECT 71.53 57.965 71.79 58.225 ;
        RECT 71.53 57.205 71.79 57.465 ;
        RECT 71.53 56.445 71.79 56.705 ;
        RECT 71.53 55.685 71.79 55.945 ;
        RECT 71.53 54.925 71.79 55.185 ;
        RECT 71.53 54.165 71.79 54.425 ;
        RECT 71.53 53.405 71.79 53.665 ;
        RECT 71.53 52.645 71.79 52.905 ;
        RECT 71.53 51.885 71.79 52.145 ;
        RECT 71.53 51.125 71.79 51.385 ;
        RECT 71.53 50.365 71.79 50.625 ;
        RECT 71.53 49.605 71.79 49.865 ;
        RECT 71.53 48.845 71.79 49.105 ;
        RECT 71.53 48.085 71.79 48.345 ;
        RECT 71.53 47.325 71.79 47.585 ;
        RECT 71.53 46.565 71.79 46.825 ;
        RECT 71.53 45.805 71.79 46.065 ;
        RECT 71.53 45.045 71.79 45.305 ;
        RECT 71.53 44.285 71.79 44.545 ;
        RECT 71.53 43.525 71.79 43.785 ;
        RECT 71.53 42.765 71.79 43.025 ;
        RECT 71.53 42.005 71.79 42.265 ;
        RECT 71.53 41.245 71.79 41.505 ;
        RECT 71.53 40.485 71.79 40.745 ;
        RECT 71.53 39.725 71.79 39.985 ;
        RECT 71.53 38.965 71.79 39.225 ;
        RECT 71.53 38.205 71.79 38.465 ;
        RECT 71.53 37.445 71.79 37.705 ;
        RECT 71.53 36.685 71.79 36.945 ;
        RECT 72.29 58.725 72.55 58.985 ;
        RECT 72.29 57.965 72.55 58.225 ;
        RECT 72.29 57.205 72.55 57.465 ;
        RECT 72.29 56.445 72.55 56.705 ;
        RECT 72.29 55.685 72.55 55.945 ;
        RECT 72.29 54.925 72.55 55.185 ;
        RECT 72.29 54.165 72.55 54.425 ;
        RECT 72.29 53.405 72.55 53.665 ;
        RECT 72.29 52.645 72.55 52.905 ;
        RECT 72.29 51.885 72.55 52.145 ;
        RECT 72.29 51.125 72.55 51.385 ;
        RECT 72.29 50.365 72.55 50.625 ;
        RECT 72.29 49.605 72.55 49.865 ;
        RECT 72.29 48.845 72.55 49.105 ;
        RECT 72.29 48.085 72.55 48.345 ;
        RECT 72.29 47.325 72.55 47.585 ;
        RECT 72.29 46.565 72.55 46.825 ;
        RECT 72.29 45.805 72.55 46.065 ;
        RECT 72.29 45.045 72.55 45.305 ;
        RECT 72.29 44.285 72.55 44.545 ;
        RECT 72.29 43.525 72.55 43.785 ;
        RECT 72.29 42.765 72.55 43.025 ;
        RECT 72.29 42.005 72.55 42.265 ;
        RECT 72.29 41.245 72.55 41.505 ;
        RECT 72.29 40.485 72.55 40.745 ;
        RECT 72.29 39.725 72.55 39.985 ;
        RECT 72.29 38.965 72.55 39.225 ;
        RECT 72.29 38.205 72.55 38.465 ;
        RECT 72.29 37.445 72.55 37.705 ;
        RECT 72.29 36.685 72.55 36.945 ;
        RECT 73.05 58.725 73.31 58.985 ;
        RECT 73.05 57.965 73.31 58.225 ;
        RECT 73.05 57.205 73.31 57.465 ;
        RECT 73.05 56.445 73.31 56.705 ;
        RECT 73.05 55.685 73.31 55.945 ;
        RECT 73.05 54.925 73.31 55.185 ;
        RECT 73.05 54.165 73.31 54.425 ;
        RECT 73.05 53.405 73.31 53.665 ;
        RECT 73.05 52.645 73.31 52.905 ;
        RECT 73.05 51.885 73.31 52.145 ;
        RECT 73.05 51.125 73.31 51.385 ;
        RECT 73.05 50.365 73.31 50.625 ;
        RECT 73.05 49.605 73.31 49.865 ;
        RECT 73.05 48.845 73.31 49.105 ;
        RECT 73.05 48.085 73.31 48.345 ;
        RECT 73.05 47.325 73.31 47.585 ;
        RECT 73.05 46.565 73.31 46.825 ;
        RECT 73.05 45.805 73.31 46.065 ;
        RECT 73.05 45.045 73.31 45.305 ;
        RECT 73.05 44.285 73.31 44.545 ;
        RECT 73.05 43.525 73.31 43.785 ;
        RECT 73.05 42.765 73.31 43.025 ;
        RECT 73.05 42.005 73.31 42.265 ;
        RECT 73.05 41.245 73.31 41.505 ;
        RECT 73.05 40.485 73.31 40.745 ;
        RECT 73.05 39.725 73.31 39.985 ;
        RECT 73.05 38.965 73.31 39.225 ;
        RECT 73.05 38.205 73.31 38.465 ;
        RECT 73.05 37.445 73.31 37.705 ;
        RECT 73.05 36.685 73.31 36.945 ;
        RECT 73.81 58.725 74.07 58.985 ;
        RECT 73.81 57.965 74.07 58.225 ;
        RECT 73.81 57.205 74.07 57.465 ;
        RECT 73.81 56.445 74.07 56.705 ;
        RECT 73.81 55.685 74.07 55.945 ;
        RECT 73.81 54.925 74.07 55.185 ;
        RECT 73.81 54.165 74.07 54.425 ;
        RECT 73.81 53.405 74.07 53.665 ;
        RECT 73.81 52.645 74.07 52.905 ;
        RECT 73.81 51.885 74.07 52.145 ;
        RECT 73.81 51.125 74.07 51.385 ;
        RECT 73.81 50.365 74.07 50.625 ;
        RECT 73.81 49.605 74.07 49.865 ;
        RECT 73.81 48.845 74.07 49.105 ;
        RECT 73.81 48.085 74.07 48.345 ;
        RECT 73.81 47.325 74.07 47.585 ;
        RECT 73.81 46.565 74.07 46.825 ;
        RECT 73.81 45.805 74.07 46.065 ;
        RECT 73.81 45.045 74.07 45.305 ;
        RECT 73.81 44.285 74.07 44.545 ;
        RECT 73.81 43.525 74.07 43.785 ;
        RECT 73.81 42.765 74.07 43.025 ;
        RECT 73.81 42.005 74.07 42.265 ;
        RECT 73.81 41.245 74.07 41.505 ;
        RECT 73.81 40.485 74.07 40.745 ;
        RECT 73.81 39.725 74.07 39.985 ;
        RECT 73.81 38.965 74.07 39.225 ;
        RECT 73.81 38.205 74.07 38.465 ;
        RECT 73.81 37.445 74.07 37.705 ;
        RECT 73.81 36.685 74.07 36.945 ;
        RECT 74.57 58.725 74.83 58.985 ;
        RECT 74.57 57.965 74.83 58.225 ;
        RECT 74.57 57.205 74.83 57.465 ;
        RECT 74.57 56.445 74.83 56.705 ;
        RECT 74.57 55.685 74.83 55.945 ;
        RECT 74.57 54.925 74.83 55.185 ;
        RECT 74.57 54.165 74.83 54.425 ;
        RECT 74.57 53.405 74.83 53.665 ;
        RECT 74.57 52.645 74.83 52.905 ;
        RECT 74.57 51.885 74.83 52.145 ;
        RECT 74.57 51.125 74.83 51.385 ;
        RECT 74.57 50.365 74.83 50.625 ;
        RECT 74.57 49.605 74.83 49.865 ;
        RECT 74.57 48.845 74.83 49.105 ;
        RECT 74.57 48.085 74.83 48.345 ;
        RECT 74.57 47.325 74.83 47.585 ;
        RECT 74.57 46.565 74.83 46.825 ;
        RECT 74.57 45.805 74.83 46.065 ;
        RECT 74.57 45.045 74.83 45.305 ;
        RECT 74.57 44.285 74.83 44.545 ;
        RECT 74.57 43.525 74.83 43.785 ;
        RECT 74.57 42.765 74.83 43.025 ;
        RECT 74.57 42.005 74.83 42.265 ;
        RECT 74.57 41.245 74.83 41.505 ;
        RECT 74.57 40.485 74.83 40.745 ;
        RECT 74.57 39.725 74.83 39.985 ;
        RECT 74.57 38.965 74.83 39.225 ;
        RECT 74.57 38.205 74.83 38.465 ;
        RECT 74.57 37.445 74.83 37.705 ;
        RECT 74.57 36.685 74.83 36.945 ;
        RECT 75.33 58.725 75.59 58.985 ;
        RECT 75.33 57.965 75.59 58.225 ;
        RECT 75.33 57.205 75.59 57.465 ;
        RECT 75.33 56.445 75.59 56.705 ;
        RECT 75.33 55.685 75.59 55.945 ;
        RECT 75.33 54.925 75.59 55.185 ;
        RECT 75.33 54.165 75.59 54.425 ;
        RECT 75.33 53.405 75.59 53.665 ;
        RECT 75.33 52.645 75.59 52.905 ;
        RECT 75.33 51.885 75.59 52.145 ;
        RECT 75.33 51.125 75.59 51.385 ;
        RECT 75.33 50.365 75.59 50.625 ;
        RECT 75.33 49.605 75.59 49.865 ;
        RECT 75.33 48.845 75.59 49.105 ;
        RECT 75.33 48.085 75.59 48.345 ;
        RECT 75.33 47.325 75.59 47.585 ;
        RECT 75.33 46.565 75.59 46.825 ;
        RECT 75.33 45.805 75.59 46.065 ;
        RECT 75.33 45.045 75.59 45.305 ;
        RECT 75.33 44.285 75.59 44.545 ;
        RECT 75.33 43.525 75.59 43.785 ;
        RECT 75.33 42.765 75.59 43.025 ;
        RECT 75.33 42.005 75.59 42.265 ;
        RECT 75.33 41.245 75.59 41.505 ;
        RECT 75.33 40.485 75.59 40.745 ;
        RECT 75.33 39.725 75.59 39.985 ;
        RECT 75.33 38.965 75.59 39.225 ;
        RECT 75.33 38.205 75.59 38.465 ;
        RECT 75.33 37.445 75.59 37.705 ;
        RECT 75.33 36.685 75.59 36.945 ;
        RECT 76.09 58.725 76.35 58.985 ;
        RECT 76.09 57.965 76.35 58.225 ;
        RECT 76.09 57.205 76.35 57.465 ;
        RECT 76.09 56.445 76.35 56.705 ;
        RECT 76.09 55.685 76.35 55.945 ;
        RECT 76.09 54.925 76.35 55.185 ;
        RECT 76.09 54.165 76.35 54.425 ;
        RECT 76.09 53.405 76.35 53.665 ;
        RECT 76.09 52.645 76.35 52.905 ;
        RECT 76.09 51.885 76.35 52.145 ;
        RECT 76.09 51.125 76.35 51.385 ;
        RECT 76.09 50.365 76.35 50.625 ;
        RECT 76.09 49.605 76.35 49.865 ;
        RECT 76.09 48.845 76.35 49.105 ;
        RECT 76.09 48.085 76.35 48.345 ;
        RECT 76.09 47.325 76.35 47.585 ;
        RECT 76.09 46.565 76.35 46.825 ;
        RECT 76.09 45.805 76.35 46.065 ;
        RECT 76.09 45.045 76.35 45.305 ;
        RECT 76.09 44.285 76.35 44.545 ;
        RECT 76.09 43.525 76.35 43.785 ;
        RECT 76.09 42.765 76.35 43.025 ;
        RECT 76.09 42.005 76.35 42.265 ;
        RECT 76.09 41.245 76.35 41.505 ;
        RECT 76.09 40.485 76.35 40.745 ;
        RECT 76.09 39.725 76.35 39.985 ;
        RECT 76.09 38.965 76.35 39.225 ;
        RECT 76.09 38.205 76.35 38.465 ;
        RECT 76.09 37.445 76.35 37.705 ;
        RECT 76.09 36.685 76.35 36.945 ;
        RECT 76.85 58.725 77.11 58.985 ;
        RECT 76.85 57.965 77.11 58.225 ;
        RECT 76.85 57.205 77.11 57.465 ;
        RECT 76.85 56.445 77.11 56.705 ;
        RECT 76.85 55.685 77.11 55.945 ;
        RECT 76.85 54.925 77.11 55.185 ;
        RECT 76.85 54.165 77.11 54.425 ;
        RECT 76.85 53.405 77.11 53.665 ;
        RECT 76.85 52.645 77.11 52.905 ;
        RECT 76.85 51.885 77.11 52.145 ;
        RECT 76.85 51.125 77.11 51.385 ;
        RECT 76.85 50.365 77.11 50.625 ;
        RECT 76.85 49.605 77.11 49.865 ;
        RECT 76.85 48.845 77.11 49.105 ;
        RECT 76.85 48.085 77.11 48.345 ;
        RECT 76.85 47.325 77.11 47.585 ;
        RECT 76.85 46.565 77.11 46.825 ;
        RECT 76.85 45.805 77.11 46.065 ;
        RECT 76.85 45.045 77.11 45.305 ;
        RECT 76.85 44.285 77.11 44.545 ;
        RECT 76.85 43.525 77.11 43.785 ;
        RECT 76.85 42.765 77.11 43.025 ;
        RECT 76.85 42.005 77.11 42.265 ;
        RECT 76.85 41.245 77.11 41.505 ;
        RECT 76.85 40.485 77.11 40.745 ;
        RECT 76.85 39.725 77.11 39.985 ;
        RECT 76.85 38.965 77.11 39.225 ;
        RECT 76.85 38.205 77.11 38.465 ;
        RECT 76.85 37.445 77.11 37.705 ;
        RECT 76.85 36.685 77.11 36.945 ;
        RECT 77.61 58.725 77.87 58.985 ;
        RECT 77.61 57.965 77.87 58.225 ;
        RECT 77.61 57.205 77.87 57.465 ;
        RECT 77.61 56.445 77.87 56.705 ;
        RECT 77.61 55.685 77.87 55.945 ;
        RECT 77.61 54.925 77.87 55.185 ;
        RECT 77.61 54.165 77.87 54.425 ;
        RECT 77.61 53.405 77.87 53.665 ;
        RECT 77.61 52.645 77.87 52.905 ;
        RECT 77.61 51.885 77.87 52.145 ;
        RECT 77.61 51.125 77.87 51.385 ;
        RECT 77.61 50.365 77.87 50.625 ;
        RECT 77.61 49.605 77.87 49.865 ;
        RECT 77.61 48.845 77.87 49.105 ;
        RECT 77.61 48.085 77.87 48.345 ;
        RECT 77.61 47.325 77.87 47.585 ;
        RECT 77.61 46.565 77.87 46.825 ;
        RECT 77.61 45.805 77.87 46.065 ;
        RECT 77.61 45.045 77.87 45.305 ;
        RECT 77.61 44.285 77.87 44.545 ;
        RECT 77.61 43.525 77.87 43.785 ;
        RECT 77.61 42.765 77.87 43.025 ;
        RECT 77.61 42.005 77.87 42.265 ;
        RECT 77.61 41.245 77.87 41.505 ;
        RECT 77.61 40.485 77.87 40.745 ;
        RECT 77.61 39.725 77.87 39.985 ;
        RECT 77.61 38.965 77.87 39.225 ;
        RECT 77.61 38.205 77.87 38.465 ;
        RECT 77.61 37.445 77.87 37.705 ;
        RECT 77.61 36.685 77.87 36.945 ;
        RECT 78.37 58.725 78.63 58.985 ;
        RECT 78.37 57.965 78.63 58.225 ;
        RECT 78.37 57.205 78.63 57.465 ;
        RECT 78.37 56.445 78.63 56.705 ;
        RECT 78.37 55.685 78.63 55.945 ;
        RECT 78.37 54.925 78.63 55.185 ;
        RECT 78.37 54.165 78.63 54.425 ;
        RECT 78.37 53.405 78.63 53.665 ;
        RECT 78.37 52.645 78.63 52.905 ;
        RECT 78.37 51.885 78.63 52.145 ;
        RECT 78.37 51.125 78.63 51.385 ;
        RECT 78.37 50.365 78.63 50.625 ;
        RECT 78.37 49.605 78.63 49.865 ;
        RECT 78.37 48.845 78.63 49.105 ;
        RECT 78.37 48.085 78.63 48.345 ;
        RECT 78.37 47.325 78.63 47.585 ;
        RECT 78.37 46.565 78.63 46.825 ;
        RECT 78.37 45.805 78.63 46.065 ;
        RECT 78.37 45.045 78.63 45.305 ;
        RECT 78.37 44.285 78.63 44.545 ;
        RECT 78.37 43.525 78.63 43.785 ;
        RECT 78.37 42.765 78.63 43.025 ;
        RECT 78.37 42.005 78.63 42.265 ;
        RECT 78.37 41.245 78.63 41.505 ;
        RECT 78.37 40.485 78.63 40.745 ;
        RECT 78.37 39.725 78.63 39.985 ;
        RECT 78.37 38.965 78.63 39.225 ;
        RECT 78.37 38.205 78.63 38.465 ;
        RECT 78.37 37.445 78.63 37.705 ;
        RECT 78.37 36.685 78.63 36.945 ;
        RECT 79.13 58.725 79.39 58.985 ;
        RECT 79.13 57.965 79.39 58.225 ;
        RECT 79.13 57.205 79.39 57.465 ;
        RECT 79.13 56.445 79.39 56.705 ;
        RECT 79.13 55.685 79.39 55.945 ;
        RECT 79.13 54.925 79.39 55.185 ;
        RECT 79.13 54.165 79.39 54.425 ;
        RECT 79.13 53.405 79.39 53.665 ;
        RECT 79.13 52.645 79.39 52.905 ;
        RECT 79.13 51.885 79.39 52.145 ;
        RECT 79.13 51.125 79.39 51.385 ;
        RECT 79.13 50.365 79.39 50.625 ;
        RECT 79.13 49.605 79.39 49.865 ;
        RECT 79.13 48.845 79.39 49.105 ;
        RECT 79.13 48.085 79.39 48.345 ;
        RECT 79.13 47.325 79.39 47.585 ;
        RECT 79.13 46.565 79.39 46.825 ;
        RECT 79.13 45.805 79.39 46.065 ;
        RECT 79.13 45.045 79.39 45.305 ;
        RECT 79.13 44.285 79.39 44.545 ;
        RECT 79.13 43.525 79.39 43.785 ;
        RECT 79.13 42.765 79.39 43.025 ;
        RECT 79.13 42.005 79.39 42.265 ;
        RECT 79.13 41.245 79.39 41.505 ;
        RECT 79.13 40.485 79.39 40.745 ;
        RECT 79.13 39.725 79.39 39.985 ;
        RECT 79.13 38.965 79.39 39.225 ;
        RECT 79.13 38.205 79.39 38.465 ;
        RECT 79.13 37.445 79.39 37.705 ;
        RECT 79.13 36.685 79.39 36.945 ;
        RECT 79.89 58.725 80.15 58.985 ;
        RECT 79.89 57.965 80.15 58.225 ;
        RECT 79.89 57.205 80.15 57.465 ;
        RECT 79.89 56.445 80.15 56.705 ;
        RECT 79.89 55.685 80.15 55.945 ;
        RECT 79.89 54.925 80.15 55.185 ;
        RECT 79.89 54.165 80.15 54.425 ;
        RECT 79.89 53.405 80.15 53.665 ;
        RECT 79.89 52.645 80.15 52.905 ;
        RECT 79.89 51.885 80.15 52.145 ;
        RECT 79.89 51.125 80.15 51.385 ;
        RECT 79.89 50.365 80.15 50.625 ;
        RECT 79.89 49.605 80.15 49.865 ;
        RECT 79.89 48.845 80.15 49.105 ;
        RECT 79.89 48.085 80.15 48.345 ;
        RECT 79.89 47.325 80.15 47.585 ;
        RECT 79.89 46.565 80.15 46.825 ;
        RECT 79.89 45.805 80.15 46.065 ;
        RECT 79.89 45.045 80.15 45.305 ;
        RECT 79.89 44.285 80.15 44.545 ;
        RECT 79.89 43.525 80.15 43.785 ;
        RECT 79.89 42.765 80.15 43.025 ;
        RECT 79.89 42.005 80.15 42.265 ;
        RECT 79.89 41.245 80.15 41.505 ;
        RECT 79.89 40.485 80.15 40.745 ;
        RECT 79.89 39.725 80.15 39.985 ;
        RECT 79.89 38.965 80.15 39.225 ;
        RECT 79.89 38.205 80.15 38.465 ;
        RECT 79.89 37.445 80.15 37.705 ;
        RECT 79.89 36.685 80.15 36.945 ;
        RECT 29.73 51.125 29.99 51.385 ;
        RECT 29.73 50.365 29.99 50.625 ;
        RECT 29.73 49.605 29.99 49.865 ;
        RECT 29.73 48.845 29.99 49.105 ;
        RECT 29.73 48.085 29.99 48.345 ;
        RECT 29.73 47.325 29.99 47.585 ;
        RECT 29.73 46.565 29.99 46.825 ;
        RECT 29.73 45.805 29.99 46.065 ;
        RECT 29.73 45.045 29.99 45.305 ;
        RECT 29.73 44.285 29.99 44.545 ;
        RECT 29.73 43.525 29.99 43.785 ;
        RECT 29.73 42.765 29.99 43.025 ;
        RECT 29.73 42.005 29.99 42.265 ;
        RECT 29.73 41.245 29.99 41.505 ;
        RECT 29.73 40.485 29.99 40.745 ;
        RECT 29.73 39.725 29.99 39.985 ;
        RECT 29.73 38.965 29.99 39.225 ;
        RECT 29.73 38.205 29.99 38.465 ;
        RECT 29.73 37.445 29.99 37.705 ;
        RECT 29.73 36.685 29.99 36.945 ;
        RECT 30.49 58.725 30.75 58.985 ;
        RECT 30.49 57.965 30.75 58.225 ;
        RECT 30.49 57.205 30.75 57.465 ;
        RECT 30.49 56.445 30.75 56.705 ;
        RECT 30.49 55.685 30.75 55.945 ;
        RECT 30.49 54.925 30.75 55.185 ;
        RECT 30.49 54.165 30.75 54.425 ;
        RECT 30.49 53.405 30.75 53.665 ;
        RECT 30.49 52.645 30.75 52.905 ;
        RECT 30.49 51.885 30.75 52.145 ;
        RECT 30.49 51.125 30.75 51.385 ;
        RECT 30.49 50.365 30.75 50.625 ;
        RECT 30.49 49.605 30.75 49.865 ;
        RECT 30.49 48.845 30.75 49.105 ;
        RECT 30.49 48.085 30.75 48.345 ;
        RECT 30.49 47.325 30.75 47.585 ;
        RECT 30.49 46.565 30.75 46.825 ;
        RECT 30.49 45.805 30.75 46.065 ;
        RECT 30.49 45.045 30.75 45.305 ;
        RECT 30.49 44.285 30.75 44.545 ;
        RECT 30.49 43.525 30.75 43.785 ;
        RECT 30.49 42.765 30.75 43.025 ;
        RECT 30.49 42.005 30.75 42.265 ;
        RECT 30.49 41.245 30.75 41.505 ;
        RECT 30.49 40.485 30.75 40.745 ;
        RECT 30.49 39.725 30.75 39.985 ;
        RECT 30.49 38.965 30.75 39.225 ;
        RECT 30.49 38.205 30.75 38.465 ;
        RECT 30.49 37.445 30.75 37.705 ;
        RECT 30.49 36.685 30.75 36.945 ;
        RECT 31.25 58.725 31.51 58.985 ;
        RECT 31.25 57.965 31.51 58.225 ;
        RECT 31.25 57.205 31.51 57.465 ;
        RECT 31.25 56.445 31.51 56.705 ;
        RECT 31.25 55.685 31.51 55.945 ;
        RECT 31.25 54.925 31.51 55.185 ;
        RECT 31.25 54.165 31.51 54.425 ;
        RECT 31.25 53.405 31.51 53.665 ;
        RECT 31.25 52.645 31.51 52.905 ;
        RECT 31.25 51.885 31.51 52.145 ;
        RECT 31.25 51.125 31.51 51.385 ;
        RECT 31.25 50.365 31.51 50.625 ;
        RECT 31.25 49.605 31.51 49.865 ;
        RECT 31.25 48.845 31.51 49.105 ;
        RECT 31.25 48.085 31.51 48.345 ;
        RECT 31.25 47.325 31.51 47.585 ;
        RECT 31.25 46.565 31.51 46.825 ;
        RECT 31.25 45.805 31.51 46.065 ;
        RECT 31.25 45.045 31.51 45.305 ;
        RECT 31.25 44.285 31.51 44.545 ;
        RECT 31.25 43.525 31.51 43.785 ;
        RECT 31.25 42.765 31.51 43.025 ;
        RECT 31.25 42.005 31.51 42.265 ;
        RECT 31.25 41.245 31.51 41.505 ;
        RECT 31.25 40.485 31.51 40.745 ;
        RECT 31.25 39.725 31.51 39.985 ;
        RECT 31.25 38.965 31.51 39.225 ;
        RECT 31.25 38.205 31.51 38.465 ;
        RECT 31.25 37.445 31.51 37.705 ;
        RECT 31.25 36.685 31.51 36.945 ;
        RECT 32.01 58.725 32.27 58.985 ;
        RECT 32.01 57.965 32.27 58.225 ;
        RECT 32.01 57.205 32.27 57.465 ;
        RECT 32.01 56.445 32.27 56.705 ;
        RECT 32.01 55.685 32.27 55.945 ;
        RECT 32.01 54.925 32.27 55.185 ;
        RECT 32.01 54.165 32.27 54.425 ;
        RECT 32.01 53.405 32.27 53.665 ;
        RECT 32.01 52.645 32.27 52.905 ;
        RECT 32.01 51.885 32.27 52.145 ;
        RECT 32.01 51.125 32.27 51.385 ;
        RECT 32.01 50.365 32.27 50.625 ;
        RECT 32.01 49.605 32.27 49.865 ;
        RECT 32.01 48.845 32.27 49.105 ;
        RECT 32.01 48.085 32.27 48.345 ;
        RECT 32.01 47.325 32.27 47.585 ;
        RECT 32.01 46.565 32.27 46.825 ;
        RECT 32.01 45.805 32.27 46.065 ;
        RECT 32.01 45.045 32.27 45.305 ;
        RECT 32.01 44.285 32.27 44.545 ;
        RECT 32.01 43.525 32.27 43.785 ;
        RECT 32.01 42.765 32.27 43.025 ;
        RECT 32.01 42.005 32.27 42.265 ;
        RECT 32.01 41.245 32.27 41.505 ;
        RECT 32.01 40.485 32.27 40.745 ;
        RECT 32.01 39.725 32.27 39.985 ;
        RECT 32.01 38.965 32.27 39.225 ;
        RECT 32.01 38.205 32.27 38.465 ;
        RECT 32.01 37.445 32.27 37.705 ;
        RECT 32.01 36.685 32.27 36.945 ;
        RECT 32.77 58.725 33.03 58.985 ;
        RECT 32.77 57.965 33.03 58.225 ;
        RECT 32.77 57.205 33.03 57.465 ;
        RECT 32.77 56.445 33.03 56.705 ;
        RECT 32.77 55.685 33.03 55.945 ;
        RECT 32.77 54.925 33.03 55.185 ;
        RECT 32.77 54.165 33.03 54.425 ;
        RECT 32.77 53.405 33.03 53.665 ;
        RECT 32.77 52.645 33.03 52.905 ;
        RECT 32.77 51.885 33.03 52.145 ;
        RECT 32.77 51.125 33.03 51.385 ;
        RECT 32.77 50.365 33.03 50.625 ;
        RECT 32.77 49.605 33.03 49.865 ;
        RECT 32.77 48.845 33.03 49.105 ;
        RECT 32.77 48.085 33.03 48.345 ;
        RECT 32.77 47.325 33.03 47.585 ;
        RECT 32.77 46.565 33.03 46.825 ;
        RECT 32.77 45.805 33.03 46.065 ;
        RECT 32.77 45.045 33.03 45.305 ;
        RECT 32.77 44.285 33.03 44.545 ;
        RECT 32.77 43.525 33.03 43.785 ;
        RECT 32.77 42.765 33.03 43.025 ;
        RECT 32.77 42.005 33.03 42.265 ;
        RECT 32.77 41.245 33.03 41.505 ;
        RECT 32.77 40.485 33.03 40.745 ;
        RECT 32.77 39.725 33.03 39.985 ;
        RECT 32.77 38.965 33.03 39.225 ;
        RECT 32.77 38.205 33.03 38.465 ;
        RECT 32.77 37.445 33.03 37.705 ;
        RECT 32.77 36.685 33.03 36.945 ;
        RECT 33.53 58.725 33.79 58.985 ;
        RECT 33.53 57.965 33.79 58.225 ;
        RECT 33.53 57.205 33.79 57.465 ;
        RECT 33.53 56.445 33.79 56.705 ;
        RECT 33.53 55.685 33.79 55.945 ;
        RECT 33.53 54.925 33.79 55.185 ;
        RECT 33.53 54.165 33.79 54.425 ;
        RECT 33.53 53.405 33.79 53.665 ;
        RECT 33.53 52.645 33.79 52.905 ;
        RECT 33.53 51.885 33.79 52.145 ;
        RECT 33.53 51.125 33.79 51.385 ;
        RECT 33.53 50.365 33.79 50.625 ;
        RECT 33.53 49.605 33.79 49.865 ;
        RECT 33.53 48.845 33.79 49.105 ;
        RECT 33.53 48.085 33.79 48.345 ;
        RECT 33.53 47.325 33.79 47.585 ;
        RECT 33.53 46.565 33.79 46.825 ;
        RECT 33.53 45.805 33.79 46.065 ;
        RECT 33.53 45.045 33.79 45.305 ;
        RECT 33.53 44.285 33.79 44.545 ;
        RECT 33.53 43.525 33.79 43.785 ;
        RECT 33.53 42.765 33.79 43.025 ;
        RECT 33.53 42.005 33.79 42.265 ;
        RECT 33.53 41.245 33.79 41.505 ;
        RECT 33.53 40.485 33.79 40.745 ;
        RECT 33.53 39.725 33.79 39.985 ;
        RECT 33.53 38.965 33.79 39.225 ;
        RECT 33.53 38.205 33.79 38.465 ;
        RECT 33.53 37.445 33.79 37.705 ;
        RECT 33.53 36.685 33.79 36.945 ;
        RECT 34.29 58.725 34.55 58.985 ;
        RECT 34.29 57.965 34.55 58.225 ;
        RECT 34.29 57.205 34.55 57.465 ;
        RECT 34.29 56.445 34.55 56.705 ;
        RECT 34.29 55.685 34.55 55.945 ;
        RECT 34.29 54.925 34.55 55.185 ;
        RECT 34.29 54.165 34.55 54.425 ;
        RECT 34.29 53.405 34.55 53.665 ;
        RECT 34.29 52.645 34.55 52.905 ;
        RECT 34.29 51.885 34.55 52.145 ;
        RECT 34.29 51.125 34.55 51.385 ;
        RECT 34.29 50.365 34.55 50.625 ;
        RECT 34.29 49.605 34.55 49.865 ;
        RECT 34.29 48.845 34.55 49.105 ;
        RECT 34.29 48.085 34.55 48.345 ;
        RECT 34.29 47.325 34.55 47.585 ;
        RECT 34.29 46.565 34.55 46.825 ;
        RECT 34.29 45.805 34.55 46.065 ;
        RECT 34.29 45.045 34.55 45.305 ;
        RECT 34.29 44.285 34.55 44.545 ;
        RECT 34.29 43.525 34.55 43.785 ;
        RECT 34.29 42.765 34.55 43.025 ;
        RECT 34.29 42.005 34.55 42.265 ;
        RECT 34.29 41.245 34.55 41.505 ;
        RECT 34.29 40.485 34.55 40.745 ;
        RECT 34.29 39.725 34.55 39.985 ;
        RECT 34.29 38.965 34.55 39.225 ;
        RECT 34.29 38.205 34.55 38.465 ;
        RECT 34.29 37.445 34.55 37.705 ;
        RECT 34.29 36.685 34.55 36.945 ;
        RECT 35.05 58.725 35.31 58.985 ;
        RECT 35.05 57.965 35.31 58.225 ;
        RECT 35.05 57.205 35.31 57.465 ;
        RECT 35.05 56.445 35.31 56.705 ;
        RECT 35.05 55.685 35.31 55.945 ;
        RECT 35.05 54.925 35.31 55.185 ;
        RECT 35.05 54.165 35.31 54.425 ;
        RECT 35.05 53.405 35.31 53.665 ;
        RECT 35.05 52.645 35.31 52.905 ;
        RECT 35.05 51.885 35.31 52.145 ;
        RECT 35.05 51.125 35.31 51.385 ;
        RECT 35.05 50.365 35.31 50.625 ;
        RECT 35.05 49.605 35.31 49.865 ;
        RECT 35.05 48.845 35.31 49.105 ;
        RECT 35.05 48.085 35.31 48.345 ;
        RECT 35.05 47.325 35.31 47.585 ;
        RECT 35.05 46.565 35.31 46.825 ;
        RECT 35.05 45.805 35.31 46.065 ;
        RECT 35.05 45.045 35.31 45.305 ;
        RECT 35.05 44.285 35.31 44.545 ;
        RECT 35.05 43.525 35.31 43.785 ;
        RECT 35.05 42.765 35.31 43.025 ;
        RECT 35.05 42.005 35.31 42.265 ;
        RECT 35.05 41.245 35.31 41.505 ;
        RECT 35.05 40.485 35.31 40.745 ;
        RECT 35.05 39.725 35.31 39.985 ;
        RECT 35.05 38.965 35.31 39.225 ;
        RECT 35.05 38.205 35.31 38.465 ;
        RECT 35.05 37.445 35.31 37.705 ;
        RECT 35.05 36.685 35.31 36.945 ;
        RECT 35.81 58.725 36.07 58.985 ;
        RECT 35.81 57.965 36.07 58.225 ;
        RECT 35.81 57.205 36.07 57.465 ;
        RECT 35.81 56.445 36.07 56.705 ;
        RECT 35.81 55.685 36.07 55.945 ;
        RECT 35.81 54.925 36.07 55.185 ;
        RECT 35.81 54.165 36.07 54.425 ;
        RECT 35.81 53.405 36.07 53.665 ;
        RECT 35.81 52.645 36.07 52.905 ;
        RECT 35.81 51.885 36.07 52.145 ;
        RECT 35.81 51.125 36.07 51.385 ;
        RECT 35.81 50.365 36.07 50.625 ;
        RECT 35.81 49.605 36.07 49.865 ;
        RECT 35.81 48.845 36.07 49.105 ;
        RECT 35.81 48.085 36.07 48.345 ;
        RECT 35.81 47.325 36.07 47.585 ;
        RECT 35.81 46.565 36.07 46.825 ;
        RECT 35.81 45.805 36.07 46.065 ;
        RECT 35.81 45.045 36.07 45.305 ;
        RECT 35.81 44.285 36.07 44.545 ;
        RECT 35.81 43.525 36.07 43.785 ;
        RECT 35.81 42.765 36.07 43.025 ;
        RECT 35.81 42.005 36.07 42.265 ;
        RECT 35.81 41.245 36.07 41.505 ;
        RECT 35.81 40.485 36.07 40.745 ;
        RECT 35.81 39.725 36.07 39.985 ;
        RECT 35.81 38.965 36.07 39.225 ;
        RECT 35.81 38.205 36.07 38.465 ;
        RECT 35.81 37.445 36.07 37.705 ;
        RECT 35.81 36.685 36.07 36.945 ;
        RECT 36.57 58.725 36.83 58.985 ;
        RECT 36.57 57.965 36.83 58.225 ;
        RECT 36.57 57.205 36.83 57.465 ;
        RECT 36.57 56.445 36.83 56.705 ;
        RECT 36.57 55.685 36.83 55.945 ;
        RECT 36.57 54.925 36.83 55.185 ;
        RECT 36.57 54.165 36.83 54.425 ;
        RECT 36.57 53.405 36.83 53.665 ;
        RECT 36.57 52.645 36.83 52.905 ;
        RECT 36.57 51.885 36.83 52.145 ;
        RECT 36.57 51.125 36.83 51.385 ;
        RECT 36.57 50.365 36.83 50.625 ;
        RECT 36.57 49.605 36.83 49.865 ;
        RECT 36.57 48.845 36.83 49.105 ;
        RECT 36.57 48.085 36.83 48.345 ;
        RECT 36.57 47.325 36.83 47.585 ;
        RECT 36.57 46.565 36.83 46.825 ;
        RECT 36.57 45.805 36.83 46.065 ;
        RECT 36.57 45.045 36.83 45.305 ;
        RECT 36.57 44.285 36.83 44.545 ;
        RECT 36.57 43.525 36.83 43.785 ;
        RECT 36.57 42.765 36.83 43.025 ;
        RECT 36.57 42.005 36.83 42.265 ;
        RECT 36.57 41.245 36.83 41.505 ;
        RECT 36.57 40.485 36.83 40.745 ;
        RECT 36.57 39.725 36.83 39.985 ;
        RECT 36.57 38.965 36.83 39.225 ;
        RECT 36.57 38.205 36.83 38.465 ;
        RECT 36.57 37.445 36.83 37.705 ;
        RECT 36.57 36.685 36.83 36.945 ;
        RECT 37.33 58.725 37.59 58.985 ;
        RECT 37.33 57.965 37.59 58.225 ;
        RECT 37.33 57.205 37.59 57.465 ;
        RECT 37.33 56.445 37.59 56.705 ;
        RECT 37.33 55.685 37.59 55.945 ;
        RECT 37.33 54.925 37.59 55.185 ;
        RECT 37.33 54.165 37.59 54.425 ;
        RECT 37.33 53.405 37.59 53.665 ;
        RECT 37.33 52.645 37.59 52.905 ;
        RECT 37.33 51.885 37.59 52.145 ;
        RECT 37.33 51.125 37.59 51.385 ;
        RECT 37.33 50.365 37.59 50.625 ;
        RECT 37.33 49.605 37.59 49.865 ;
        RECT 37.33 48.845 37.59 49.105 ;
        RECT 37.33 48.085 37.59 48.345 ;
        RECT 37.33 47.325 37.59 47.585 ;
        RECT 37.33 46.565 37.59 46.825 ;
        RECT 37.33 45.805 37.59 46.065 ;
        RECT 37.33 45.045 37.59 45.305 ;
        RECT 37.33 44.285 37.59 44.545 ;
        RECT 37.33 43.525 37.59 43.785 ;
        RECT 37.33 42.765 37.59 43.025 ;
        RECT 37.33 42.005 37.59 42.265 ;
        RECT 37.33 41.245 37.59 41.505 ;
        RECT 37.33 40.485 37.59 40.745 ;
        RECT 37.33 39.725 37.59 39.985 ;
        RECT 37.33 38.965 37.59 39.225 ;
        RECT 37.33 38.205 37.59 38.465 ;
        RECT 37.33 37.445 37.59 37.705 ;
        RECT 37.33 36.685 37.59 36.945 ;
        RECT 38.09 58.725 38.35 58.985 ;
        RECT 38.09 57.965 38.35 58.225 ;
        RECT 38.09 57.205 38.35 57.465 ;
        RECT 38.09 56.445 38.35 56.705 ;
        RECT 38.09 55.685 38.35 55.945 ;
        RECT 38.09 54.925 38.35 55.185 ;
        RECT 38.09 54.165 38.35 54.425 ;
        RECT 38.09 53.405 38.35 53.665 ;
        RECT 38.09 52.645 38.35 52.905 ;
        RECT 38.09 51.885 38.35 52.145 ;
        RECT 38.09 51.125 38.35 51.385 ;
        RECT 38.09 50.365 38.35 50.625 ;
        RECT 38.09 49.605 38.35 49.865 ;
        RECT 38.09 48.845 38.35 49.105 ;
        RECT 38.09 48.085 38.35 48.345 ;
        RECT 38.09 47.325 38.35 47.585 ;
        RECT 38.09 46.565 38.35 46.825 ;
        RECT 38.09 45.805 38.35 46.065 ;
        RECT 38.09 45.045 38.35 45.305 ;
        RECT 38.09 44.285 38.35 44.545 ;
        RECT 38.09 43.525 38.35 43.785 ;
        RECT 38.09 42.765 38.35 43.025 ;
        RECT 38.09 42.005 38.35 42.265 ;
        RECT 38.09 41.245 38.35 41.505 ;
        RECT 38.09 40.485 38.35 40.745 ;
        RECT 38.09 39.725 38.35 39.985 ;
        RECT 38.09 38.965 38.35 39.225 ;
        RECT 38.09 38.205 38.35 38.465 ;
        RECT 38.09 37.445 38.35 37.705 ;
        RECT 38.09 36.685 38.35 36.945 ;
        RECT 38.85 58.725 39.11 58.985 ;
        RECT 38.85 57.965 39.11 58.225 ;
        RECT 38.85 57.205 39.11 57.465 ;
        RECT 38.85 56.445 39.11 56.705 ;
        RECT 38.85 55.685 39.11 55.945 ;
        RECT 38.85 54.925 39.11 55.185 ;
        RECT 38.85 54.165 39.11 54.425 ;
        RECT 38.85 53.405 39.11 53.665 ;
        RECT 38.85 52.645 39.11 52.905 ;
        RECT 38.85 51.885 39.11 52.145 ;
        RECT 38.85 51.125 39.11 51.385 ;
        RECT 38.85 50.365 39.11 50.625 ;
        RECT 38.85 49.605 39.11 49.865 ;
        RECT 38.85 48.845 39.11 49.105 ;
        RECT 38.85 48.085 39.11 48.345 ;
        RECT 38.85 47.325 39.11 47.585 ;
        RECT 38.85 46.565 39.11 46.825 ;
        RECT 38.85 45.805 39.11 46.065 ;
        RECT 38.85 45.045 39.11 45.305 ;
        RECT 38.85 44.285 39.11 44.545 ;
        RECT 38.85 43.525 39.11 43.785 ;
        RECT 38.85 42.765 39.11 43.025 ;
        RECT 38.85 42.005 39.11 42.265 ;
        RECT 38.85 41.245 39.11 41.505 ;
        RECT 38.85 40.485 39.11 40.745 ;
        RECT 38.85 39.725 39.11 39.985 ;
        RECT 38.85 38.965 39.11 39.225 ;
        RECT 38.85 38.205 39.11 38.465 ;
        RECT 38.85 37.445 39.11 37.705 ;
        RECT 38.85 36.685 39.11 36.945 ;
        RECT 39.61 58.725 39.87 58.985 ;
        RECT 39.61 57.965 39.87 58.225 ;
        RECT 39.61 57.205 39.87 57.465 ;
        RECT 39.61 56.445 39.87 56.705 ;
        RECT 39.61 55.685 39.87 55.945 ;
        RECT 39.61 54.925 39.87 55.185 ;
        RECT 39.61 54.165 39.87 54.425 ;
        RECT 39.61 53.405 39.87 53.665 ;
        RECT 39.61 52.645 39.87 52.905 ;
        RECT 39.61 51.885 39.87 52.145 ;
        RECT 39.61 51.125 39.87 51.385 ;
        RECT 39.61 50.365 39.87 50.625 ;
        RECT 39.61 49.605 39.87 49.865 ;
        RECT 39.61 48.845 39.87 49.105 ;
        RECT 39.61 48.085 39.87 48.345 ;
        RECT 39.61 47.325 39.87 47.585 ;
        RECT 39.61 46.565 39.87 46.825 ;
        RECT 39.61 45.805 39.87 46.065 ;
        RECT 39.61 45.045 39.87 45.305 ;
        RECT 39.61 44.285 39.87 44.545 ;
        RECT 39.61 43.525 39.87 43.785 ;
        RECT 39.61 42.765 39.87 43.025 ;
        RECT 39.61 42.005 39.87 42.265 ;
        RECT 39.61 41.245 39.87 41.505 ;
        RECT 39.61 40.485 39.87 40.745 ;
        RECT 39.61 39.725 39.87 39.985 ;
        RECT 39.61 38.965 39.87 39.225 ;
        RECT 39.61 38.205 39.87 38.465 ;
        RECT 39.61 37.445 39.87 37.705 ;
        RECT 39.61 36.685 39.87 36.945 ;
        RECT 40.37 58.725 40.63 58.985 ;
        RECT 40.37 57.965 40.63 58.225 ;
        RECT 40.37 57.205 40.63 57.465 ;
        RECT 40.37 56.445 40.63 56.705 ;
        RECT 40.37 55.685 40.63 55.945 ;
        RECT 40.37 54.925 40.63 55.185 ;
        RECT 40.37 54.165 40.63 54.425 ;
        RECT 40.37 53.405 40.63 53.665 ;
        RECT 40.37 52.645 40.63 52.905 ;
        RECT 40.37 51.885 40.63 52.145 ;
        RECT 40.37 51.125 40.63 51.385 ;
        RECT 40.37 50.365 40.63 50.625 ;
        RECT 40.37 49.605 40.63 49.865 ;
        RECT 40.37 48.845 40.63 49.105 ;
        RECT 40.37 48.085 40.63 48.345 ;
        RECT 40.37 47.325 40.63 47.585 ;
        RECT 40.37 46.565 40.63 46.825 ;
        RECT 40.37 45.805 40.63 46.065 ;
        RECT 40.37 45.045 40.63 45.305 ;
        RECT 40.37 44.285 40.63 44.545 ;
        RECT 40.37 43.525 40.63 43.785 ;
        RECT 40.37 42.765 40.63 43.025 ;
        RECT 40.37 42.005 40.63 42.265 ;
        RECT 40.37 41.245 40.63 41.505 ;
        RECT 40.37 40.485 40.63 40.745 ;
        RECT 40.37 39.725 40.63 39.985 ;
        RECT 40.37 38.965 40.63 39.225 ;
        RECT 40.37 38.205 40.63 38.465 ;
        RECT 40.37 37.445 40.63 37.705 ;
        RECT 40.37 36.685 40.63 36.945 ;
        RECT 41.13 58.725 41.39 58.985 ;
        RECT 41.13 57.965 41.39 58.225 ;
        RECT 41.13 57.205 41.39 57.465 ;
        RECT 41.13 56.445 41.39 56.705 ;
        RECT 41.13 55.685 41.39 55.945 ;
        RECT 41.13 54.925 41.39 55.185 ;
        RECT 41.13 54.165 41.39 54.425 ;
        RECT 41.13 53.405 41.39 53.665 ;
        RECT 41.13 52.645 41.39 52.905 ;
        RECT 41.13 51.885 41.39 52.145 ;
        RECT 41.13 51.125 41.39 51.385 ;
        RECT 41.13 50.365 41.39 50.625 ;
        RECT 41.13 49.605 41.39 49.865 ;
        RECT 41.13 48.845 41.39 49.105 ;
        RECT 41.13 48.085 41.39 48.345 ;
        RECT 41.13 47.325 41.39 47.585 ;
        RECT 41.13 46.565 41.39 46.825 ;
        RECT 41.13 45.805 41.39 46.065 ;
        RECT 41.13 45.045 41.39 45.305 ;
        RECT 41.13 44.285 41.39 44.545 ;
        RECT 41.13 43.525 41.39 43.785 ;
        RECT 41.13 42.765 41.39 43.025 ;
        RECT 41.13 42.005 41.39 42.265 ;
        RECT 41.13 41.245 41.39 41.505 ;
        RECT 41.13 40.485 41.39 40.745 ;
        RECT 41.13 39.725 41.39 39.985 ;
        RECT 41.13 38.965 41.39 39.225 ;
        RECT 41.13 38.205 41.39 38.465 ;
        RECT 41.13 37.445 41.39 37.705 ;
        RECT 41.13 36.685 41.39 36.945 ;
        RECT 41.89 58.725 42.15 58.985 ;
        RECT 41.89 57.965 42.15 58.225 ;
        RECT 41.89 57.205 42.15 57.465 ;
        RECT 41.89 56.445 42.15 56.705 ;
        RECT 41.89 55.685 42.15 55.945 ;
        RECT 41.89 54.925 42.15 55.185 ;
        RECT 41.89 54.165 42.15 54.425 ;
        RECT 41.89 53.405 42.15 53.665 ;
        RECT 41.89 52.645 42.15 52.905 ;
        RECT 41.89 51.885 42.15 52.145 ;
        RECT 41.89 51.125 42.15 51.385 ;
        RECT 41.89 50.365 42.15 50.625 ;
        RECT 41.89 49.605 42.15 49.865 ;
        RECT 41.89 48.845 42.15 49.105 ;
        RECT 41.89 48.085 42.15 48.345 ;
        RECT 41.89 47.325 42.15 47.585 ;
        RECT 41.89 46.565 42.15 46.825 ;
        RECT 41.89 45.805 42.15 46.065 ;
        RECT 41.89 45.045 42.15 45.305 ;
        RECT 41.89 44.285 42.15 44.545 ;
        RECT 41.89 43.525 42.15 43.785 ;
        RECT 41.89 42.765 42.15 43.025 ;
        RECT 41.89 42.005 42.15 42.265 ;
        RECT 41.89 41.245 42.15 41.505 ;
        RECT 41.89 40.485 42.15 40.745 ;
        RECT 41.89 39.725 42.15 39.985 ;
        RECT 41.89 38.965 42.15 39.225 ;
        RECT 41.89 38.205 42.15 38.465 ;
        RECT 41.89 37.445 42.15 37.705 ;
        RECT 41.89 36.685 42.15 36.945 ;
        RECT 42.65 58.725 42.91 58.985 ;
        RECT 42.65 57.965 42.91 58.225 ;
        RECT 42.65 57.205 42.91 57.465 ;
        RECT 42.65 56.445 42.91 56.705 ;
        RECT 42.65 55.685 42.91 55.945 ;
        RECT 42.65 54.925 42.91 55.185 ;
        RECT 42.65 54.165 42.91 54.425 ;
        RECT 42.65 53.405 42.91 53.665 ;
        RECT 42.65 52.645 42.91 52.905 ;
        RECT 42.65 51.885 42.91 52.145 ;
        RECT 42.65 51.125 42.91 51.385 ;
        RECT 42.65 50.365 42.91 50.625 ;
        RECT 42.65 49.605 42.91 49.865 ;
        RECT 42.65 48.845 42.91 49.105 ;
        RECT 42.65 48.085 42.91 48.345 ;
        RECT 42.65 47.325 42.91 47.585 ;
        RECT 42.65 46.565 42.91 46.825 ;
        RECT 42.65 45.805 42.91 46.065 ;
        RECT 42.65 45.045 42.91 45.305 ;
        RECT 42.65 44.285 42.91 44.545 ;
        RECT 42.65 43.525 42.91 43.785 ;
        RECT 42.65 42.765 42.91 43.025 ;
        RECT 42.65 42.005 42.91 42.265 ;
        RECT 42.65 41.245 42.91 41.505 ;
        RECT 42.65 40.485 42.91 40.745 ;
        RECT 42.65 39.725 42.91 39.985 ;
        RECT 42.65 38.965 42.91 39.225 ;
        RECT 42.65 38.205 42.91 38.465 ;
        RECT 42.65 37.445 42.91 37.705 ;
        RECT 42.65 36.685 42.91 36.945 ;
        RECT 43.41 58.725 43.67 58.985 ;
        RECT 43.41 57.965 43.67 58.225 ;
        RECT 43.41 57.205 43.67 57.465 ;
        RECT 43.41 56.445 43.67 56.705 ;
        RECT 43.41 55.685 43.67 55.945 ;
        RECT 43.41 54.925 43.67 55.185 ;
        RECT 43.41 54.165 43.67 54.425 ;
        RECT 43.41 53.405 43.67 53.665 ;
        RECT 43.41 52.645 43.67 52.905 ;
        RECT 43.41 51.885 43.67 52.145 ;
        RECT 43.41 51.125 43.67 51.385 ;
        RECT 43.41 50.365 43.67 50.625 ;
        RECT 43.41 49.605 43.67 49.865 ;
        RECT 43.41 48.845 43.67 49.105 ;
        RECT 43.41 48.085 43.67 48.345 ;
        RECT 43.41 47.325 43.67 47.585 ;
        RECT 43.41 46.565 43.67 46.825 ;
        RECT 43.41 45.805 43.67 46.065 ;
        RECT 43.41 45.045 43.67 45.305 ;
        RECT 43.41 44.285 43.67 44.545 ;
        RECT 43.41 43.525 43.67 43.785 ;
        RECT 43.41 42.765 43.67 43.025 ;
        RECT 43.41 42.005 43.67 42.265 ;
        RECT 43.41 41.245 43.67 41.505 ;
        RECT 43.41 40.485 43.67 40.745 ;
        RECT 43.41 39.725 43.67 39.985 ;
        RECT 43.41 38.965 43.67 39.225 ;
        RECT 43.41 38.205 43.67 38.465 ;
        RECT 43.41 37.445 43.67 37.705 ;
        RECT 43.41 36.685 43.67 36.945 ;
        RECT 44.17 58.725 44.43 58.985 ;
        RECT 44.17 57.965 44.43 58.225 ;
        RECT 44.17 57.205 44.43 57.465 ;
        RECT 44.17 56.445 44.43 56.705 ;
        RECT 44.17 55.685 44.43 55.945 ;
        RECT 44.17 54.925 44.43 55.185 ;
        RECT 44.17 54.165 44.43 54.425 ;
        RECT 44.17 53.405 44.43 53.665 ;
        RECT 44.17 52.645 44.43 52.905 ;
        RECT 44.17 51.885 44.43 52.145 ;
        RECT 44.17 51.125 44.43 51.385 ;
        RECT 44.17 50.365 44.43 50.625 ;
        RECT 44.17 49.605 44.43 49.865 ;
        RECT 44.17 48.845 44.43 49.105 ;
        RECT 44.17 48.085 44.43 48.345 ;
        RECT 44.17 47.325 44.43 47.585 ;
        RECT 44.17 46.565 44.43 46.825 ;
        RECT 44.17 45.805 44.43 46.065 ;
        RECT 44.17 45.045 44.43 45.305 ;
        RECT 44.17 44.285 44.43 44.545 ;
        RECT 44.17 43.525 44.43 43.785 ;
        RECT 44.17 42.765 44.43 43.025 ;
        RECT 44.17 42.005 44.43 42.265 ;
        RECT 44.17 41.245 44.43 41.505 ;
        RECT 44.17 40.485 44.43 40.745 ;
        RECT 44.17 39.725 44.43 39.985 ;
        RECT 44.17 38.965 44.43 39.225 ;
        RECT 44.17 38.205 44.43 38.465 ;
        RECT 44.17 37.445 44.43 37.705 ;
        RECT 44.17 36.685 44.43 36.945 ;
        RECT 44.93 58.725 45.19 58.985 ;
        RECT 44.93 57.965 45.19 58.225 ;
        RECT 44.93 57.205 45.19 57.465 ;
        RECT 44.93 56.445 45.19 56.705 ;
        RECT 44.93 55.685 45.19 55.945 ;
        RECT 44.93 54.925 45.19 55.185 ;
        RECT 44.93 54.165 45.19 54.425 ;
        RECT 44.93 53.405 45.19 53.665 ;
        RECT 44.93 52.645 45.19 52.905 ;
        RECT 44.93 51.885 45.19 52.145 ;
        RECT 44.93 51.125 45.19 51.385 ;
        RECT 44.93 50.365 45.19 50.625 ;
        RECT 44.93 49.605 45.19 49.865 ;
        RECT 44.93 48.845 45.19 49.105 ;
        RECT 44.93 48.085 45.19 48.345 ;
        RECT 44.93 47.325 45.19 47.585 ;
        RECT 44.93 46.565 45.19 46.825 ;
        RECT 44.93 45.805 45.19 46.065 ;
        RECT 44.93 45.045 45.19 45.305 ;
        RECT 44.93 44.285 45.19 44.545 ;
        RECT 44.93 43.525 45.19 43.785 ;
        RECT 44.93 42.765 45.19 43.025 ;
        RECT 44.93 42.005 45.19 42.265 ;
        RECT 44.93 41.245 45.19 41.505 ;
        RECT 44.93 40.485 45.19 40.745 ;
        RECT 44.93 39.725 45.19 39.985 ;
        RECT 44.93 38.965 45.19 39.225 ;
        RECT 44.93 38.205 45.19 38.465 ;
        RECT 44.93 37.445 45.19 37.705 ;
        RECT 44.93 36.685 45.19 36.945 ;
        RECT 45.69 58.725 45.95 58.985 ;
        RECT 45.69 57.965 45.95 58.225 ;
        RECT 45.69 57.205 45.95 57.465 ;
        RECT 45.69 56.445 45.95 56.705 ;
        RECT 45.69 55.685 45.95 55.945 ;
        RECT 45.69 54.925 45.95 55.185 ;
        RECT 45.69 54.165 45.95 54.425 ;
        RECT 45.69 53.405 45.95 53.665 ;
        RECT 45.69 52.645 45.95 52.905 ;
        RECT 45.69 51.885 45.95 52.145 ;
        RECT 45.69 51.125 45.95 51.385 ;
        RECT 45.69 50.365 45.95 50.625 ;
        RECT 45.69 49.605 45.95 49.865 ;
        RECT 45.69 48.845 45.95 49.105 ;
        RECT 45.69 48.085 45.95 48.345 ;
        RECT 45.69 47.325 45.95 47.585 ;
        RECT 45.69 46.565 45.95 46.825 ;
        RECT 45.69 45.805 45.95 46.065 ;
        RECT 45.69 45.045 45.95 45.305 ;
        RECT 45.69 44.285 45.95 44.545 ;
        RECT 45.69 43.525 45.95 43.785 ;
        RECT 45.69 42.765 45.95 43.025 ;
        RECT 45.69 42.005 45.95 42.265 ;
        RECT 45.69 41.245 45.95 41.505 ;
        RECT 45.69 40.485 45.95 40.745 ;
        RECT 45.69 39.725 45.95 39.985 ;
        RECT 45.69 38.965 45.95 39.225 ;
        RECT 45.69 38.205 45.95 38.465 ;
        RECT 45.69 37.445 45.95 37.705 ;
        RECT 45.69 36.685 45.95 36.945 ;
        RECT 46.45 58.725 46.71 58.985 ;
        RECT 46.45 57.965 46.71 58.225 ;
        RECT 46.45 57.205 46.71 57.465 ;
        RECT 46.45 56.445 46.71 56.705 ;
        RECT 46.45 55.685 46.71 55.945 ;
        RECT 46.45 54.925 46.71 55.185 ;
        RECT 46.45 54.165 46.71 54.425 ;
        RECT 46.45 53.405 46.71 53.665 ;
        RECT 46.45 52.645 46.71 52.905 ;
        RECT 46.45 51.885 46.71 52.145 ;
        RECT 46.45 51.125 46.71 51.385 ;
        RECT 46.45 50.365 46.71 50.625 ;
        RECT 46.45 49.605 46.71 49.865 ;
        RECT 46.45 48.845 46.71 49.105 ;
        RECT 46.45 48.085 46.71 48.345 ;
        RECT 46.45 47.325 46.71 47.585 ;
        RECT 46.45 46.565 46.71 46.825 ;
        RECT 46.45 45.805 46.71 46.065 ;
        RECT 46.45 45.045 46.71 45.305 ;
        RECT 46.45 44.285 46.71 44.545 ;
        RECT 46.45 43.525 46.71 43.785 ;
        RECT 46.45 42.765 46.71 43.025 ;
        RECT 46.45 42.005 46.71 42.265 ;
        RECT 46.45 41.245 46.71 41.505 ;
        RECT 46.45 40.485 46.71 40.745 ;
        RECT 46.45 39.725 46.71 39.985 ;
        RECT 46.45 38.965 46.71 39.225 ;
        RECT 46.45 38.205 46.71 38.465 ;
        RECT 46.45 37.445 46.71 37.705 ;
        RECT 46.45 36.685 46.71 36.945 ;
        RECT 47.21 58.725 47.47 58.985 ;
        RECT 47.21 57.965 47.47 58.225 ;
        RECT 47.21 57.205 47.47 57.465 ;
        RECT 47.21 56.445 47.47 56.705 ;
        RECT 47.21 55.685 47.47 55.945 ;
        RECT 47.21 54.925 47.47 55.185 ;
        RECT 47.21 54.165 47.47 54.425 ;
        RECT 47.21 53.405 47.47 53.665 ;
        RECT 47.21 52.645 47.47 52.905 ;
        RECT 47.21 51.885 47.47 52.145 ;
        RECT 47.21 51.125 47.47 51.385 ;
        RECT 47.21 50.365 47.47 50.625 ;
        RECT 47.21 49.605 47.47 49.865 ;
        RECT 47.21 48.845 47.47 49.105 ;
        RECT 47.21 48.085 47.47 48.345 ;
        RECT 47.21 47.325 47.47 47.585 ;
        RECT 47.21 46.565 47.47 46.825 ;
        RECT 47.21 45.805 47.47 46.065 ;
        RECT 47.21 45.045 47.47 45.305 ;
        RECT 47.21 44.285 47.47 44.545 ;
        RECT 47.21 43.525 47.47 43.785 ;
        RECT 47.21 42.765 47.47 43.025 ;
        RECT 47.21 42.005 47.47 42.265 ;
        RECT 47.21 41.245 47.47 41.505 ;
        RECT 47.21 40.485 47.47 40.745 ;
        RECT 47.21 39.725 47.47 39.985 ;
        RECT 47.21 38.965 47.47 39.225 ;
        RECT 47.21 38.205 47.47 38.465 ;
        RECT 47.21 37.445 47.47 37.705 ;
        RECT 47.21 36.685 47.47 36.945 ;
        RECT 47.97 58.725 48.23 58.985 ;
        RECT 47.97 57.965 48.23 58.225 ;
        RECT 47.97 57.205 48.23 57.465 ;
        RECT 47.97 56.445 48.23 56.705 ;
        RECT 47.97 55.685 48.23 55.945 ;
        RECT 47.97 54.925 48.23 55.185 ;
        RECT 47.97 54.165 48.23 54.425 ;
        RECT 47.97 53.405 48.23 53.665 ;
        RECT 47.97 52.645 48.23 52.905 ;
        RECT 47.97 51.885 48.23 52.145 ;
        RECT 47.97 51.125 48.23 51.385 ;
        RECT 47.97 50.365 48.23 50.625 ;
        RECT 47.97 49.605 48.23 49.865 ;
        RECT 47.97 48.845 48.23 49.105 ;
        RECT 47.97 48.085 48.23 48.345 ;
        RECT 47.97 47.325 48.23 47.585 ;
        RECT 47.97 46.565 48.23 46.825 ;
        RECT 47.97 45.805 48.23 46.065 ;
        RECT 47.97 45.045 48.23 45.305 ;
        RECT 47.97 44.285 48.23 44.545 ;
        RECT 47.97 43.525 48.23 43.785 ;
        RECT 47.97 42.765 48.23 43.025 ;
        RECT 47.97 42.005 48.23 42.265 ;
        RECT 47.97 41.245 48.23 41.505 ;
        RECT 47.97 40.485 48.23 40.745 ;
        RECT 47.97 39.725 48.23 39.985 ;
        RECT 47.97 38.965 48.23 39.225 ;
        RECT 47.97 38.205 48.23 38.465 ;
        RECT 47.97 37.445 48.23 37.705 ;
        RECT 47.97 36.685 48.23 36.945 ;
        RECT 48.73 58.725 48.99 58.985 ;
        RECT 48.73 57.965 48.99 58.225 ;
        RECT 48.73 57.205 48.99 57.465 ;
        RECT 48.73 56.445 48.99 56.705 ;
        RECT 48.73 55.685 48.99 55.945 ;
        RECT 48.73 54.925 48.99 55.185 ;
        RECT 48.73 54.165 48.99 54.425 ;
        RECT 48.73 53.405 48.99 53.665 ;
        RECT 48.73 52.645 48.99 52.905 ;
        RECT 48.73 51.885 48.99 52.145 ;
        RECT 48.73 51.125 48.99 51.385 ;
        RECT 48.73 50.365 48.99 50.625 ;
        RECT 48.73 49.605 48.99 49.865 ;
        RECT 48.73 48.845 48.99 49.105 ;
        RECT 48.73 48.085 48.99 48.345 ;
        RECT 48.73 47.325 48.99 47.585 ;
        RECT 48.73 46.565 48.99 46.825 ;
        RECT 48.73 45.805 48.99 46.065 ;
        RECT 48.73 45.045 48.99 45.305 ;
        RECT 48.73 44.285 48.99 44.545 ;
        RECT 48.73 43.525 48.99 43.785 ;
        RECT 48.73 42.765 48.99 43.025 ;
        RECT 48.73 42.005 48.99 42.265 ;
        RECT 48.73 41.245 48.99 41.505 ;
        RECT 48.73 40.485 48.99 40.745 ;
        RECT 48.73 39.725 48.99 39.985 ;
        RECT 48.73 38.965 48.99 39.225 ;
        RECT 48.73 38.205 48.99 38.465 ;
        RECT 48.73 37.445 48.99 37.705 ;
        RECT 48.73 36.685 48.99 36.945 ;
        RECT 49.49 58.725 49.75 58.985 ;
        RECT 49.49 57.965 49.75 58.225 ;
        RECT 49.49 57.205 49.75 57.465 ;
        RECT 49.49 56.445 49.75 56.705 ;
        RECT 49.49 55.685 49.75 55.945 ;
        RECT 49.49 54.925 49.75 55.185 ;
        RECT 49.49 54.165 49.75 54.425 ;
        RECT 49.49 53.405 49.75 53.665 ;
        RECT 49.49 52.645 49.75 52.905 ;
        RECT 49.49 51.885 49.75 52.145 ;
        RECT 49.49 51.125 49.75 51.385 ;
        RECT 49.49 50.365 49.75 50.625 ;
        RECT 49.49 49.605 49.75 49.865 ;
        RECT 49.49 48.845 49.75 49.105 ;
        RECT 49.49 48.085 49.75 48.345 ;
        RECT 49.49 47.325 49.75 47.585 ;
        RECT 49.49 46.565 49.75 46.825 ;
        RECT 49.49 45.805 49.75 46.065 ;
        RECT 49.49 45.045 49.75 45.305 ;
        RECT 49.49 44.285 49.75 44.545 ;
        RECT 49.49 43.525 49.75 43.785 ;
        RECT 49.49 42.765 49.75 43.025 ;
        RECT 49.49 42.005 49.75 42.265 ;
        RECT 49.49 41.245 49.75 41.505 ;
        RECT 49.49 40.485 49.75 40.745 ;
        RECT 49.49 39.725 49.75 39.985 ;
        RECT 49.49 38.965 49.75 39.225 ;
        RECT 49.49 38.205 49.75 38.465 ;
        RECT 49.49 37.445 49.75 37.705 ;
        RECT 49.49 36.685 49.75 36.945 ;
        RECT 50.25 58.725 50.51 58.985 ;
        RECT 50.25 57.965 50.51 58.225 ;
        RECT 50.25 57.205 50.51 57.465 ;
        RECT 50.25 56.445 50.51 56.705 ;
        RECT 50.25 55.685 50.51 55.945 ;
        RECT 50.25 54.925 50.51 55.185 ;
        RECT 50.25 54.165 50.51 54.425 ;
        RECT 50.25 53.405 50.51 53.665 ;
        RECT 50.25 52.645 50.51 52.905 ;
        RECT 50.25 51.885 50.51 52.145 ;
        RECT 50.25 51.125 50.51 51.385 ;
        RECT 50.25 50.365 50.51 50.625 ;
        RECT 50.25 49.605 50.51 49.865 ;
        RECT 50.25 48.845 50.51 49.105 ;
        RECT 50.25 48.085 50.51 48.345 ;
        RECT 50.25 47.325 50.51 47.585 ;
        RECT 50.25 46.565 50.51 46.825 ;
        RECT 50.25 45.805 50.51 46.065 ;
        RECT 50.25 45.045 50.51 45.305 ;
        RECT 50.25 44.285 50.51 44.545 ;
        RECT 50.25 43.525 50.51 43.785 ;
        RECT 50.25 42.765 50.51 43.025 ;
        RECT 50.25 42.005 50.51 42.265 ;
        RECT 50.25 41.245 50.51 41.505 ;
        RECT 50.25 40.485 50.51 40.745 ;
        RECT 50.25 39.725 50.51 39.985 ;
        RECT 50.25 38.965 50.51 39.225 ;
        RECT 50.25 38.205 50.51 38.465 ;
        RECT 50.25 37.445 50.51 37.705 ;
        RECT 50.25 36.685 50.51 36.945 ;
        RECT 51.01 58.725 51.27 58.985 ;
        RECT 51.01 57.965 51.27 58.225 ;
        RECT 51.01 57.205 51.27 57.465 ;
        RECT 51.01 56.445 51.27 56.705 ;
        RECT 51.01 55.685 51.27 55.945 ;
        RECT 51.01 54.925 51.27 55.185 ;
        RECT 51.01 54.165 51.27 54.425 ;
        RECT 51.01 53.405 51.27 53.665 ;
        RECT 51.01 52.645 51.27 52.905 ;
        RECT 51.01 51.885 51.27 52.145 ;
        RECT 51.01 51.125 51.27 51.385 ;
        RECT 51.01 50.365 51.27 50.625 ;
        RECT 51.01 49.605 51.27 49.865 ;
        RECT 51.01 48.845 51.27 49.105 ;
        RECT 51.01 48.085 51.27 48.345 ;
        RECT 51.01 47.325 51.27 47.585 ;
        RECT 51.01 46.565 51.27 46.825 ;
        RECT 51.01 45.805 51.27 46.065 ;
        RECT 51.01 45.045 51.27 45.305 ;
        RECT 51.01 44.285 51.27 44.545 ;
        RECT 51.01 43.525 51.27 43.785 ;
        RECT 51.01 42.765 51.27 43.025 ;
        RECT 51.01 42.005 51.27 42.265 ;
        RECT 51.01 41.245 51.27 41.505 ;
        RECT 51.01 40.485 51.27 40.745 ;
        RECT 51.01 39.725 51.27 39.985 ;
        RECT 51.01 38.965 51.27 39.225 ;
        RECT 51.01 38.205 51.27 38.465 ;
        RECT 51.01 37.445 51.27 37.705 ;
        RECT 51.01 36.685 51.27 36.945 ;
        RECT 51.77 58.725 52.03 58.985 ;
        RECT 51.77 57.965 52.03 58.225 ;
        RECT 51.77 57.205 52.03 57.465 ;
        RECT 51.77 56.445 52.03 56.705 ;
        RECT 51.77 55.685 52.03 55.945 ;
        RECT 51.77 54.925 52.03 55.185 ;
        RECT 51.77 54.165 52.03 54.425 ;
        RECT 51.77 53.405 52.03 53.665 ;
        RECT 51.77 52.645 52.03 52.905 ;
        RECT 51.77 51.885 52.03 52.145 ;
        RECT 51.77 51.125 52.03 51.385 ;
        RECT 51.77 50.365 52.03 50.625 ;
        RECT 51.77 49.605 52.03 49.865 ;
        RECT 51.77 48.845 52.03 49.105 ;
        RECT 51.77 48.085 52.03 48.345 ;
        RECT 51.77 47.325 52.03 47.585 ;
        RECT 51.77 46.565 52.03 46.825 ;
        RECT 51.77 45.805 52.03 46.065 ;
        RECT 51.77 45.045 52.03 45.305 ;
        RECT 51.77 44.285 52.03 44.545 ;
        RECT 51.77 43.525 52.03 43.785 ;
        RECT 51.77 42.765 52.03 43.025 ;
        RECT 51.77 42.005 52.03 42.265 ;
        RECT 51.77 41.245 52.03 41.505 ;
        RECT 51.77 40.485 52.03 40.745 ;
        RECT 51.77 39.725 52.03 39.985 ;
        RECT 51.77 38.965 52.03 39.225 ;
        RECT 51.77 38.205 52.03 38.465 ;
        RECT 51.77 37.445 52.03 37.705 ;
        RECT 51.77 36.685 52.03 36.945 ;
        RECT 52.53 58.725 52.79 58.985 ;
        RECT 52.53 57.965 52.79 58.225 ;
        RECT 52.53 57.205 52.79 57.465 ;
        RECT 52.53 56.445 52.79 56.705 ;
        RECT 52.53 55.685 52.79 55.945 ;
        RECT 52.53 54.925 52.79 55.185 ;
        RECT 52.53 54.165 52.79 54.425 ;
        RECT 52.53 53.405 52.79 53.665 ;
        RECT 52.53 52.645 52.79 52.905 ;
        RECT 52.53 51.885 52.79 52.145 ;
        RECT 52.53 51.125 52.79 51.385 ;
        RECT 52.53 50.365 52.79 50.625 ;
        RECT 52.53 49.605 52.79 49.865 ;
        RECT 52.53 48.845 52.79 49.105 ;
        RECT 52.53 48.085 52.79 48.345 ;
        RECT 52.53 47.325 52.79 47.585 ;
        RECT 52.53 46.565 52.79 46.825 ;
        RECT 52.53 45.805 52.79 46.065 ;
        RECT 52.53 45.045 52.79 45.305 ;
        RECT 52.53 44.285 52.79 44.545 ;
        RECT 52.53 43.525 52.79 43.785 ;
        RECT 52.53 42.765 52.79 43.025 ;
        RECT 52.53 42.005 52.79 42.265 ;
        RECT 52.53 41.245 52.79 41.505 ;
        RECT 52.53 40.485 52.79 40.745 ;
        RECT 52.53 39.725 52.79 39.985 ;
        RECT 52.53 38.965 52.79 39.225 ;
        RECT 52.53 38.205 52.79 38.465 ;
        RECT 52.53 37.445 52.79 37.705 ;
        RECT 52.53 36.685 52.79 36.945 ;
        RECT 53.29 58.725 53.55 58.985 ;
        RECT 53.29 57.965 53.55 58.225 ;
        RECT 53.29 57.205 53.55 57.465 ;
        RECT 53.29 56.445 53.55 56.705 ;
        RECT 53.29 55.685 53.55 55.945 ;
        RECT 53.29 54.925 53.55 55.185 ;
        RECT 53.29 54.165 53.55 54.425 ;
        RECT 53.29 53.405 53.55 53.665 ;
        RECT 53.29 52.645 53.55 52.905 ;
        RECT 53.29 51.885 53.55 52.145 ;
        RECT 53.29 51.125 53.55 51.385 ;
        RECT 53.29 50.365 53.55 50.625 ;
        RECT 53.29 49.605 53.55 49.865 ;
        RECT 53.29 48.845 53.55 49.105 ;
        RECT 53.29 48.085 53.55 48.345 ;
        RECT 53.29 47.325 53.55 47.585 ;
        RECT 53.29 46.565 53.55 46.825 ;
        RECT 53.29 45.805 53.55 46.065 ;
        RECT 53.29 45.045 53.55 45.305 ;
        RECT 53.29 44.285 53.55 44.545 ;
        RECT 53.29 43.525 53.55 43.785 ;
        RECT 53.29 42.765 53.55 43.025 ;
        RECT 53.29 42.005 53.55 42.265 ;
        RECT 53.29 41.245 53.55 41.505 ;
        RECT 53.29 40.485 53.55 40.745 ;
        RECT 53.29 39.725 53.55 39.985 ;
        RECT 53.29 38.965 53.55 39.225 ;
        RECT 53.29 38.205 53.55 38.465 ;
        RECT 53.29 37.445 53.55 37.705 ;
        RECT 53.29 36.685 53.55 36.945 ;
        RECT 54.05 58.725 54.31 58.985 ;
        RECT 54.05 57.965 54.31 58.225 ;
        RECT 54.05 57.205 54.31 57.465 ;
        RECT 54.05 56.445 54.31 56.705 ;
        RECT 54.05 55.685 54.31 55.945 ;
        RECT 54.05 54.925 54.31 55.185 ;
        RECT 54.05 54.165 54.31 54.425 ;
        RECT 54.05 53.405 54.31 53.665 ;
        RECT 54.05 52.645 54.31 52.905 ;
        RECT 54.05 51.885 54.31 52.145 ;
        RECT 54.05 51.125 54.31 51.385 ;
        RECT 54.05 50.365 54.31 50.625 ;
        RECT 54.05 49.605 54.31 49.865 ;
        RECT 54.05 48.845 54.31 49.105 ;
        RECT 54.05 48.085 54.31 48.345 ;
        RECT 54.05 47.325 54.31 47.585 ;
        RECT 54.05 46.565 54.31 46.825 ;
        RECT 54.05 45.805 54.31 46.065 ;
        RECT 54.05 45.045 54.31 45.305 ;
        RECT 54.05 44.285 54.31 44.545 ;
        RECT 54.05 43.525 54.31 43.785 ;
        RECT 54.05 42.765 54.31 43.025 ;
        RECT 54.05 42.005 54.31 42.265 ;
        RECT 54.05 41.245 54.31 41.505 ;
        RECT 54.05 40.485 54.31 40.745 ;
        RECT 54.05 39.725 54.31 39.985 ;
        RECT 54.05 38.965 54.31 39.225 ;
        RECT 54.05 38.205 54.31 38.465 ;
        RECT 54.05 37.445 54.31 37.705 ;
        RECT 54.05 36.685 54.31 36.945 ;
        RECT 54.81 58.725 55.07 58.985 ;
        RECT 54.81 57.965 55.07 58.225 ;
        RECT 54.81 57.205 55.07 57.465 ;
        RECT 54.81 56.445 55.07 56.705 ;
        RECT 54.81 55.685 55.07 55.945 ;
        RECT 54.81 54.925 55.07 55.185 ;
        RECT 54.81 54.165 55.07 54.425 ;
        RECT 54.81 53.405 55.07 53.665 ;
        RECT 54.81 52.645 55.07 52.905 ;
        RECT 54.81 51.885 55.07 52.145 ;
        RECT 54.81 51.125 55.07 51.385 ;
        RECT 54.81 50.365 55.07 50.625 ;
        RECT 54.81 49.605 55.07 49.865 ;
        RECT 54.81 48.845 55.07 49.105 ;
        RECT 54.81 48.085 55.07 48.345 ;
        RECT 54.81 47.325 55.07 47.585 ;
        RECT 54.81 46.565 55.07 46.825 ;
        RECT 54.81 45.805 55.07 46.065 ;
        RECT 54.81 45.045 55.07 45.305 ;
        RECT 54.81 44.285 55.07 44.545 ;
        RECT 4.65 58.725 4.91 58.985 ;
        RECT 4.65 57.965 4.91 58.225 ;
        RECT 4.65 57.205 4.91 57.465 ;
        RECT 4.65 56.445 4.91 56.705 ;
        RECT 4.65 55.685 4.91 55.945 ;
        RECT 4.65 54.925 4.91 55.185 ;
        RECT 4.65 54.165 4.91 54.425 ;
        RECT 4.65 53.405 4.91 53.665 ;
        RECT 4.65 52.645 4.91 52.905 ;
        RECT 4.65 51.885 4.91 52.145 ;
        RECT 4.65 51.125 4.91 51.385 ;
        RECT 4.65 50.365 4.91 50.625 ;
        RECT 4.65 49.605 4.91 49.865 ;
        RECT 4.65 48.845 4.91 49.105 ;
        RECT 4.65 48.085 4.91 48.345 ;
        RECT 4.65 47.325 4.91 47.585 ;
        RECT 4.65 46.565 4.91 46.825 ;
        RECT 4.65 45.805 4.91 46.065 ;
        RECT 4.65 45.045 4.91 45.305 ;
        RECT 4.65 44.285 4.91 44.545 ;
        RECT 4.65 43.525 4.91 43.785 ;
        RECT 4.65 42.765 4.91 43.025 ;
        RECT 4.65 42.005 4.91 42.265 ;
        RECT 4.65 41.245 4.91 41.505 ;
        RECT 4.65 40.485 4.91 40.745 ;
        RECT 4.65 39.725 4.91 39.985 ;
        RECT 4.65 38.965 4.91 39.225 ;
        RECT 4.65 38.205 4.91 38.465 ;
        RECT 4.65 37.445 4.91 37.705 ;
        RECT 4.65 36.685 4.91 36.945 ;
        RECT 5.41 58.725 5.67 58.985 ;
        RECT 5.41 57.965 5.67 58.225 ;
        RECT 5.41 57.205 5.67 57.465 ;
        RECT 5.41 56.445 5.67 56.705 ;
        RECT 5.41 55.685 5.67 55.945 ;
        RECT 5.41 54.925 5.67 55.185 ;
        RECT 5.41 54.165 5.67 54.425 ;
        RECT 5.41 53.405 5.67 53.665 ;
        RECT 5.41 52.645 5.67 52.905 ;
        RECT 5.41 51.885 5.67 52.145 ;
        RECT 5.41 51.125 5.67 51.385 ;
        RECT 5.41 50.365 5.67 50.625 ;
        RECT 5.41 49.605 5.67 49.865 ;
        RECT 5.41 48.845 5.67 49.105 ;
        RECT 5.41 48.085 5.67 48.345 ;
        RECT 5.41 47.325 5.67 47.585 ;
        RECT 5.41 46.565 5.67 46.825 ;
        RECT 5.41 45.805 5.67 46.065 ;
        RECT 5.41 45.045 5.67 45.305 ;
        RECT 5.41 44.285 5.67 44.545 ;
        RECT 5.41 43.525 5.67 43.785 ;
        RECT 5.41 42.765 5.67 43.025 ;
        RECT 5.41 42.005 5.67 42.265 ;
        RECT 5.41 41.245 5.67 41.505 ;
        RECT 5.41 40.485 5.67 40.745 ;
        RECT 5.41 39.725 5.67 39.985 ;
        RECT 5.41 38.965 5.67 39.225 ;
        RECT 5.41 38.205 5.67 38.465 ;
        RECT 5.41 37.445 5.67 37.705 ;
        RECT 5.41 36.685 5.67 36.945 ;
        RECT 6.17 58.725 6.43 58.985 ;
        RECT 6.17 57.965 6.43 58.225 ;
        RECT 6.17 57.205 6.43 57.465 ;
        RECT 6.17 56.445 6.43 56.705 ;
        RECT 6.17 55.685 6.43 55.945 ;
        RECT 6.17 54.925 6.43 55.185 ;
        RECT 6.17 54.165 6.43 54.425 ;
        RECT 6.17 53.405 6.43 53.665 ;
        RECT 6.17 52.645 6.43 52.905 ;
        RECT 6.17 51.885 6.43 52.145 ;
        RECT 6.17 51.125 6.43 51.385 ;
        RECT 6.17 50.365 6.43 50.625 ;
        RECT 6.17 49.605 6.43 49.865 ;
        RECT 6.17 48.845 6.43 49.105 ;
        RECT 6.17 48.085 6.43 48.345 ;
        RECT 6.17 47.325 6.43 47.585 ;
        RECT 6.17 46.565 6.43 46.825 ;
        RECT 6.17 45.805 6.43 46.065 ;
        RECT 6.17 45.045 6.43 45.305 ;
        RECT 6.17 44.285 6.43 44.545 ;
        RECT 6.17 43.525 6.43 43.785 ;
        RECT 6.17 42.765 6.43 43.025 ;
        RECT 6.17 42.005 6.43 42.265 ;
        RECT 6.17 41.245 6.43 41.505 ;
        RECT 6.17 40.485 6.43 40.745 ;
        RECT 6.17 39.725 6.43 39.985 ;
        RECT 6.17 38.965 6.43 39.225 ;
        RECT 6.17 38.205 6.43 38.465 ;
        RECT 6.17 37.445 6.43 37.705 ;
        RECT 6.17 36.685 6.43 36.945 ;
        RECT 6.93 58.725 7.19 58.985 ;
        RECT 6.93 57.965 7.19 58.225 ;
        RECT 6.93 57.205 7.19 57.465 ;
        RECT 6.93 56.445 7.19 56.705 ;
        RECT 6.93 55.685 7.19 55.945 ;
        RECT 6.93 54.925 7.19 55.185 ;
        RECT 6.93 54.165 7.19 54.425 ;
        RECT 6.93 53.405 7.19 53.665 ;
        RECT 6.93 52.645 7.19 52.905 ;
        RECT 6.93 51.885 7.19 52.145 ;
        RECT 6.93 51.125 7.19 51.385 ;
        RECT 6.93 50.365 7.19 50.625 ;
        RECT 6.93 49.605 7.19 49.865 ;
        RECT 6.93 48.845 7.19 49.105 ;
        RECT 6.93 48.085 7.19 48.345 ;
        RECT 6.93 47.325 7.19 47.585 ;
        RECT 6.93 46.565 7.19 46.825 ;
        RECT 6.93 45.805 7.19 46.065 ;
        RECT 6.93 45.045 7.19 45.305 ;
        RECT 6.93 44.285 7.19 44.545 ;
        RECT 6.93 43.525 7.19 43.785 ;
        RECT 6.93 42.765 7.19 43.025 ;
        RECT 6.93 42.005 7.19 42.265 ;
        RECT 6.93 41.245 7.19 41.505 ;
        RECT 6.93 40.485 7.19 40.745 ;
        RECT 6.93 39.725 7.19 39.985 ;
        RECT 6.93 38.965 7.19 39.225 ;
        RECT 6.93 38.205 7.19 38.465 ;
        RECT 6.93 37.445 7.19 37.705 ;
        RECT 6.93 36.685 7.19 36.945 ;
        RECT 7.69 58.725 7.95 58.985 ;
        RECT 7.69 57.965 7.95 58.225 ;
        RECT 7.69 57.205 7.95 57.465 ;
        RECT 7.69 56.445 7.95 56.705 ;
        RECT 7.69 55.685 7.95 55.945 ;
        RECT 7.69 54.925 7.95 55.185 ;
        RECT 7.69 54.165 7.95 54.425 ;
        RECT 7.69 53.405 7.95 53.665 ;
        RECT 7.69 52.645 7.95 52.905 ;
        RECT 7.69 51.885 7.95 52.145 ;
        RECT 7.69 51.125 7.95 51.385 ;
        RECT 7.69 50.365 7.95 50.625 ;
        RECT 7.69 49.605 7.95 49.865 ;
        RECT 7.69 48.845 7.95 49.105 ;
        RECT 7.69 48.085 7.95 48.345 ;
        RECT 7.69 47.325 7.95 47.585 ;
        RECT 7.69 46.565 7.95 46.825 ;
        RECT 7.69 45.805 7.95 46.065 ;
        RECT 7.69 45.045 7.95 45.305 ;
        RECT 7.69 44.285 7.95 44.545 ;
        RECT 7.69 43.525 7.95 43.785 ;
        RECT 7.69 42.765 7.95 43.025 ;
        RECT 7.69 42.005 7.95 42.265 ;
        RECT 7.69 41.245 7.95 41.505 ;
        RECT 7.69 40.485 7.95 40.745 ;
        RECT 7.69 39.725 7.95 39.985 ;
        RECT 7.69 38.965 7.95 39.225 ;
        RECT 7.69 38.205 7.95 38.465 ;
        RECT 7.69 37.445 7.95 37.705 ;
        RECT 7.69 36.685 7.95 36.945 ;
        RECT 8.45 58.725 8.71 58.985 ;
        RECT 8.45 57.965 8.71 58.225 ;
        RECT 8.45 57.205 8.71 57.465 ;
        RECT 8.45 56.445 8.71 56.705 ;
        RECT 8.45 55.685 8.71 55.945 ;
        RECT 8.45 54.925 8.71 55.185 ;
        RECT 8.45 54.165 8.71 54.425 ;
        RECT 8.45 53.405 8.71 53.665 ;
        RECT 8.45 52.645 8.71 52.905 ;
        RECT 8.45 51.885 8.71 52.145 ;
        RECT 8.45 51.125 8.71 51.385 ;
        RECT 8.45 50.365 8.71 50.625 ;
        RECT 8.45 49.605 8.71 49.865 ;
        RECT 8.45 48.845 8.71 49.105 ;
        RECT 8.45 48.085 8.71 48.345 ;
        RECT 8.45 47.325 8.71 47.585 ;
        RECT 8.45 46.565 8.71 46.825 ;
        RECT 8.45 45.805 8.71 46.065 ;
        RECT 8.45 45.045 8.71 45.305 ;
        RECT 8.45 44.285 8.71 44.545 ;
        RECT 8.45 43.525 8.71 43.785 ;
        RECT 8.45 42.765 8.71 43.025 ;
        RECT 8.45 42.005 8.71 42.265 ;
        RECT 8.45 41.245 8.71 41.505 ;
        RECT 8.45 40.485 8.71 40.745 ;
        RECT 8.45 39.725 8.71 39.985 ;
        RECT 8.45 38.965 8.71 39.225 ;
        RECT 8.45 38.205 8.71 38.465 ;
        RECT 8.45 37.445 8.71 37.705 ;
        RECT 8.45 36.685 8.71 36.945 ;
        RECT 9.21 58.725 9.47 58.985 ;
        RECT 9.21 57.965 9.47 58.225 ;
        RECT 9.21 57.205 9.47 57.465 ;
        RECT 9.21 56.445 9.47 56.705 ;
        RECT 9.21 55.685 9.47 55.945 ;
        RECT 9.21 54.925 9.47 55.185 ;
        RECT 9.21 54.165 9.47 54.425 ;
        RECT 9.21 53.405 9.47 53.665 ;
        RECT 9.21 52.645 9.47 52.905 ;
        RECT 9.21 51.885 9.47 52.145 ;
        RECT 9.21 51.125 9.47 51.385 ;
        RECT 9.21 50.365 9.47 50.625 ;
        RECT 9.21 49.605 9.47 49.865 ;
        RECT 9.21 48.845 9.47 49.105 ;
        RECT 9.21 48.085 9.47 48.345 ;
        RECT 9.21 47.325 9.47 47.585 ;
        RECT 9.21 46.565 9.47 46.825 ;
        RECT 9.21 45.805 9.47 46.065 ;
        RECT 9.21 45.045 9.47 45.305 ;
        RECT 9.21 44.285 9.47 44.545 ;
        RECT 9.21 43.525 9.47 43.785 ;
        RECT 9.21 42.765 9.47 43.025 ;
        RECT 9.21 42.005 9.47 42.265 ;
        RECT 9.21 41.245 9.47 41.505 ;
        RECT 9.21 40.485 9.47 40.745 ;
        RECT 9.21 39.725 9.47 39.985 ;
        RECT 9.21 38.965 9.47 39.225 ;
        RECT 9.21 38.205 9.47 38.465 ;
        RECT 9.21 37.445 9.47 37.705 ;
        RECT 9.21 36.685 9.47 36.945 ;
        RECT 9.97 58.725 10.23 58.985 ;
        RECT 9.97 57.965 10.23 58.225 ;
        RECT 9.97 57.205 10.23 57.465 ;
        RECT 9.97 56.445 10.23 56.705 ;
        RECT 9.97 55.685 10.23 55.945 ;
        RECT 9.97 54.925 10.23 55.185 ;
        RECT 9.97 54.165 10.23 54.425 ;
        RECT 9.97 53.405 10.23 53.665 ;
        RECT 9.97 52.645 10.23 52.905 ;
        RECT 9.97 51.885 10.23 52.145 ;
        RECT 9.97 51.125 10.23 51.385 ;
        RECT 9.97 50.365 10.23 50.625 ;
        RECT 9.97 49.605 10.23 49.865 ;
        RECT 9.97 48.845 10.23 49.105 ;
        RECT 9.97 48.085 10.23 48.345 ;
        RECT 9.97 47.325 10.23 47.585 ;
        RECT 9.97 46.565 10.23 46.825 ;
        RECT 9.97 45.805 10.23 46.065 ;
        RECT 9.97 45.045 10.23 45.305 ;
        RECT 9.97 44.285 10.23 44.545 ;
        RECT 9.97 43.525 10.23 43.785 ;
        RECT 9.97 42.765 10.23 43.025 ;
        RECT 9.97 42.005 10.23 42.265 ;
        RECT 9.97 41.245 10.23 41.505 ;
        RECT 9.97 40.485 10.23 40.745 ;
        RECT 9.97 39.725 10.23 39.985 ;
        RECT 9.97 38.965 10.23 39.225 ;
        RECT 9.97 38.205 10.23 38.465 ;
        RECT 9.97 37.445 10.23 37.705 ;
        RECT 9.97 36.685 10.23 36.945 ;
        RECT 10.73 58.725 10.99 58.985 ;
        RECT 10.73 57.965 10.99 58.225 ;
        RECT 10.73 57.205 10.99 57.465 ;
        RECT 10.73 56.445 10.99 56.705 ;
        RECT 10.73 55.685 10.99 55.945 ;
        RECT 10.73 54.925 10.99 55.185 ;
        RECT 10.73 54.165 10.99 54.425 ;
        RECT 10.73 53.405 10.99 53.665 ;
        RECT 10.73 52.645 10.99 52.905 ;
        RECT 10.73 51.885 10.99 52.145 ;
        RECT 10.73 51.125 10.99 51.385 ;
        RECT 10.73 50.365 10.99 50.625 ;
        RECT 10.73 49.605 10.99 49.865 ;
        RECT 10.73 48.845 10.99 49.105 ;
        RECT 10.73 48.085 10.99 48.345 ;
        RECT 10.73 47.325 10.99 47.585 ;
        RECT 10.73 46.565 10.99 46.825 ;
        RECT 10.73 45.805 10.99 46.065 ;
        RECT 10.73 45.045 10.99 45.305 ;
        RECT 10.73 44.285 10.99 44.545 ;
        RECT 10.73 43.525 10.99 43.785 ;
        RECT 10.73 42.765 10.99 43.025 ;
        RECT 10.73 42.005 10.99 42.265 ;
        RECT 10.73 41.245 10.99 41.505 ;
        RECT 10.73 40.485 10.99 40.745 ;
        RECT 10.73 39.725 10.99 39.985 ;
        RECT 10.73 38.965 10.99 39.225 ;
        RECT 10.73 38.205 10.99 38.465 ;
        RECT 10.73 37.445 10.99 37.705 ;
        RECT 10.73 36.685 10.99 36.945 ;
        RECT 11.49 58.725 11.75 58.985 ;
        RECT 11.49 57.965 11.75 58.225 ;
        RECT 11.49 57.205 11.75 57.465 ;
        RECT 11.49 56.445 11.75 56.705 ;
        RECT 11.49 55.685 11.75 55.945 ;
        RECT 11.49 54.925 11.75 55.185 ;
        RECT 11.49 54.165 11.75 54.425 ;
        RECT 11.49 53.405 11.75 53.665 ;
        RECT 11.49 52.645 11.75 52.905 ;
        RECT 11.49 51.885 11.75 52.145 ;
        RECT 11.49 51.125 11.75 51.385 ;
        RECT 11.49 50.365 11.75 50.625 ;
        RECT 11.49 49.605 11.75 49.865 ;
        RECT 11.49 48.845 11.75 49.105 ;
        RECT 11.49 48.085 11.75 48.345 ;
        RECT 11.49 47.325 11.75 47.585 ;
        RECT 11.49 46.565 11.75 46.825 ;
        RECT 11.49 45.805 11.75 46.065 ;
        RECT 11.49 45.045 11.75 45.305 ;
        RECT 11.49 44.285 11.75 44.545 ;
        RECT 11.49 43.525 11.75 43.785 ;
        RECT 11.49 42.765 11.75 43.025 ;
        RECT 11.49 42.005 11.75 42.265 ;
        RECT 11.49 41.245 11.75 41.505 ;
        RECT 11.49 40.485 11.75 40.745 ;
        RECT 11.49 39.725 11.75 39.985 ;
        RECT 11.49 38.965 11.75 39.225 ;
        RECT 11.49 38.205 11.75 38.465 ;
        RECT 11.49 37.445 11.75 37.705 ;
        RECT 11.49 36.685 11.75 36.945 ;
        RECT 12.25 58.725 12.51 58.985 ;
        RECT 12.25 57.965 12.51 58.225 ;
        RECT 12.25 57.205 12.51 57.465 ;
        RECT 12.25 56.445 12.51 56.705 ;
        RECT 12.25 55.685 12.51 55.945 ;
        RECT 12.25 54.925 12.51 55.185 ;
        RECT 12.25 54.165 12.51 54.425 ;
        RECT 12.25 53.405 12.51 53.665 ;
        RECT 12.25 52.645 12.51 52.905 ;
        RECT 12.25 51.885 12.51 52.145 ;
        RECT 12.25 51.125 12.51 51.385 ;
        RECT 12.25 50.365 12.51 50.625 ;
        RECT 12.25 49.605 12.51 49.865 ;
        RECT 12.25 48.845 12.51 49.105 ;
        RECT 12.25 48.085 12.51 48.345 ;
        RECT 12.25 47.325 12.51 47.585 ;
        RECT 12.25 46.565 12.51 46.825 ;
        RECT 12.25 45.805 12.51 46.065 ;
        RECT 12.25 45.045 12.51 45.305 ;
        RECT 12.25 44.285 12.51 44.545 ;
        RECT 12.25 43.525 12.51 43.785 ;
        RECT 12.25 42.765 12.51 43.025 ;
        RECT 12.25 42.005 12.51 42.265 ;
        RECT 12.25 41.245 12.51 41.505 ;
        RECT 12.25 40.485 12.51 40.745 ;
        RECT 12.25 39.725 12.51 39.985 ;
        RECT 12.25 38.965 12.51 39.225 ;
        RECT 12.25 38.205 12.51 38.465 ;
        RECT 12.25 37.445 12.51 37.705 ;
        RECT 12.25 36.685 12.51 36.945 ;
        RECT 13.01 58.725 13.27 58.985 ;
        RECT 13.01 57.965 13.27 58.225 ;
        RECT 13.01 57.205 13.27 57.465 ;
        RECT 13.01 56.445 13.27 56.705 ;
        RECT 13.01 55.685 13.27 55.945 ;
        RECT 13.01 54.925 13.27 55.185 ;
        RECT 13.01 54.165 13.27 54.425 ;
        RECT 13.01 53.405 13.27 53.665 ;
        RECT 13.01 52.645 13.27 52.905 ;
        RECT 13.01 51.885 13.27 52.145 ;
        RECT 13.01 51.125 13.27 51.385 ;
        RECT 13.01 50.365 13.27 50.625 ;
        RECT 13.01 49.605 13.27 49.865 ;
        RECT 13.01 48.845 13.27 49.105 ;
        RECT 13.01 48.085 13.27 48.345 ;
        RECT 13.01 47.325 13.27 47.585 ;
        RECT 13.01 46.565 13.27 46.825 ;
        RECT 13.01 45.805 13.27 46.065 ;
        RECT 13.01 45.045 13.27 45.305 ;
        RECT 13.01 44.285 13.27 44.545 ;
        RECT 13.01 43.525 13.27 43.785 ;
        RECT 13.01 42.765 13.27 43.025 ;
        RECT 13.01 42.005 13.27 42.265 ;
        RECT 13.01 41.245 13.27 41.505 ;
        RECT 13.01 40.485 13.27 40.745 ;
        RECT 13.01 39.725 13.27 39.985 ;
        RECT 13.01 38.965 13.27 39.225 ;
        RECT 13.01 38.205 13.27 38.465 ;
        RECT 13.01 37.445 13.27 37.705 ;
        RECT 13.01 36.685 13.27 36.945 ;
        RECT 13.77 58.725 14.03 58.985 ;
        RECT 13.77 57.965 14.03 58.225 ;
        RECT 13.77 57.205 14.03 57.465 ;
        RECT 13.77 56.445 14.03 56.705 ;
        RECT 13.77 55.685 14.03 55.945 ;
        RECT 13.77 54.925 14.03 55.185 ;
        RECT 13.77 54.165 14.03 54.425 ;
        RECT 13.77 53.405 14.03 53.665 ;
        RECT 13.77 52.645 14.03 52.905 ;
        RECT 13.77 51.885 14.03 52.145 ;
        RECT 13.77 51.125 14.03 51.385 ;
        RECT 13.77 50.365 14.03 50.625 ;
        RECT 13.77 49.605 14.03 49.865 ;
        RECT 13.77 48.845 14.03 49.105 ;
        RECT 13.77 48.085 14.03 48.345 ;
        RECT 13.77 47.325 14.03 47.585 ;
        RECT 13.77 46.565 14.03 46.825 ;
        RECT 13.77 45.805 14.03 46.065 ;
        RECT 13.77 45.045 14.03 45.305 ;
        RECT 13.77 44.285 14.03 44.545 ;
        RECT 13.77 43.525 14.03 43.785 ;
        RECT 13.77 42.765 14.03 43.025 ;
        RECT 13.77 42.005 14.03 42.265 ;
        RECT 13.77 41.245 14.03 41.505 ;
        RECT 13.77 40.485 14.03 40.745 ;
        RECT 13.77 39.725 14.03 39.985 ;
        RECT 13.77 38.965 14.03 39.225 ;
        RECT 13.77 38.205 14.03 38.465 ;
        RECT 13.77 37.445 14.03 37.705 ;
        RECT 13.77 36.685 14.03 36.945 ;
        RECT 14.53 58.725 14.79 58.985 ;
        RECT 14.53 57.965 14.79 58.225 ;
        RECT 14.53 57.205 14.79 57.465 ;
        RECT 14.53 56.445 14.79 56.705 ;
        RECT 14.53 55.685 14.79 55.945 ;
        RECT 14.53 54.925 14.79 55.185 ;
        RECT 14.53 54.165 14.79 54.425 ;
        RECT 14.53 53.405 14.79 53.665 ;
        RECT 14.53 52.645 14.79 52.905 ;
        RECT 14.53 51.885 14.79 52.145 ;
        RECT 14.53 51.125 14.79 51.385 ;
        RECT 14.53 50.365 14.79 50.625 ;
        RECT 14.53 49.605 14.79 49.865 ;
        RECT 14.53 48.845 14.79 49.105 ;
        RECT 14.53 48.085 14.79 48.345 ;
        RECT 14.53 47.325 14.79 47.585 ;
        RECT 14.53 46.565 14.79 46.825 ;
        RECT 14.53 45.805 14.79 46.065 ;
        RECT 14.53 45.045 14.79 45.305 ;
        RECT 14.53 44.285 14.79 44.545 ;
        RECT 14.53 43.525 14.79 43.785 ;
        RECT 14.53 42.765 14.79 43.025 ;
        RECT 14.53 42.005 14.79 42.265 ;
        RECT 14.53 41.245 14.79 41.505 ;
        RECT 14.53 40.485 14.79 40.745 ;
        RECT 14.53 39.725 14.79 39.985 ;
        RECT 14.53 38.965 14.79 39.225 ;
        RECT 14.53 38.205 14.79 38.465 ;
        RECT 14.53 37.445 14.79 37.705 ;
        RECT 14.53 36.685 14.79 36.945 ;
        RECT 15.29 58.725 15.55 58.985 ;
        RECT 15.29 57.965 15.55 58.225 ;
        RECT 15.29 57.205 15.55 57.465 ;
        RECT 15.29 56.445 15.55 56.705 ;
        RECT 15.29 55.685 15.55 55.945 ;
        RECT 15.29 54.925 15.55 55.185 ;
        RECT 15.29 54.165 15.55 54.425 ;
        RECT 15.29 53.405 15.55 53.665 ;
        RECT 15.29 52.645 15.55 52.905 ;
        RECT 15.29 51.885 15.55 52.145 ;
        RECT 15.29 51.125 15.55 51.385 ;
        RECT 15.29 50.365 15.55 50.625 ;
        RECT 15.29 49.605 15.55 49.865 ;
        RECT 15.29 48.845 15.55 49.105 ;
        RECT 15.29 48.085 15.55 48.345 ;
        RECT 15.29 47.325 15.55 47.585 ;
        RECT 15.29 46.565 15.55 46.825 ;
        RECT 15.29 45.805 15.55 46.065 ;
        RECT 15.29 45.045 15.55 45.305 ;
        RECT 15.29 44.285 15.55 44.545 ;
        RECT 15.29 43.525 15.55 43.785 ;
        RECT 15.29 42.765 15.55 43.025 ;
        RECT 15.29 42.005 15.55 42.265 ;
        RECT 15.29 41.245 15.55 41.505 ;
        RECT 15.29 40.485 15.55 40.745 ;
        RECT 15.29 39.725 15.55 39.985 ;
        RECT 15.29 38.965 15.55 39.225 ;
        RECT 15.29 38.205 15.55 38.465 ;
        RECT 15.29 37.445 15.55 37.705 ;
        RECT 15.29 36.685 15.55 36.945 ;
        RECT 16.05 58.725 16.31 58.985 ;
        RECT 16.05 57.965 16.31 58.225 ;
        RECT 16.05 57.205 16.31 57.465 ;
        RECT 16.05 56.445 16.31 56.705 ;
        RECT 16.05 55.685 16.31 55.945 ;
        RECT 16.05 54.925 16.31 55.185 ;
        RECT 16.05 54.165 16.31 54.425 ;
        RECT 16.05 53.405 16.31 53.665 ;
        RECT 16.05 52.645 16.31 52.905 ;
        RECT 16.05 51.885 16.31 52.145 ;
        RECT 16.05 51.125 16.31 51.385 ;
        RECT 16.05 50.365 16.31 50.625 ;
        RECT 16.05 49.605 16.31 49.865 ;
        RECT 16.05 48.845 16.31 49.105 ;
        RECT 16.05 48.085 16.31 48.345 ;
        RECT 16.05 47.325 16.31 47.585 ;
        RECT 16.05 46.565 16.31 46.825 ;
        RECT 16.05 45.805 16.31 46.065 ;
        RECT 16.05 45.045 16.31 45.305 ;
        RECT 16.05 44.285 16.31 44.545 ;
        RECT 16.05 43.525 16.31 43.785 ;
        RECT 16.05 42.765 16.31 43.025 ;
        RECT 16.05 42.005 16.31 42.265 ;
        RECT 16.05 41.245 16.31 41.505 ;
        RECT 16.05 40.485 16.31 40.745 ;
        RECT 16.05 39.725 16.31 39.985 ;
        RECT 16.05 38.965 16.31 39.225 ;
        RECT 16.05 38.205 16.31 38.465 ;
        RECT 16.05 37.445 16.31 37.705 ;
        RECT 16.05 36.685 16.31 36.945 ;
        RECT 16.81 58.725 17.07 58.985 ;
        RECT 16.81 57.965 17.07 58.225 ;
        RECT 16.81 57.205 17.07 57.465 ;
        RECT 16.81 56.445 17.07 56.705 ;
        RECT 16.81 55.685 17.07 55.945 ;
        RECT 16.81 54.925 17.07 55.185 ;
        RECT 16.81 54.165 17.07 54.425 ;
        RECT 16.81 53.405 17.07 53.665 ;
        RECT 16.81 52.645 17.07 52.905 ;
        RECT 16.81 51.885 17.07 52.145 ;
        RECT 16.81 51.125 17.07 51.385 ;
        RECT 16.81 50.365 17.07 50.625 ;
        RECT 16.81 49.605 17.07 49.865 ;
        RECT 16.81 48.845 17.07 49.105 ;
        RECT 16.81 48.085 17.07 48.345 ;
        RECT 16.81 47.325 17.07 47.585 ;
        RECT 16.81 46.565 17.07 46.825 ;
        RECT 16.81 45.805 17.07 46.065 ;
        RECT 16.81 45.045 17.07 45.305 ;
        RECT 16.81 44.285 17.07 44.545 ;
        RECT 16.81 43.525 17.07 43.785 ;
        RECT 16.81 42.765 17.07 43.025 ;
        RECT 16.81 42.005 17.07 42.265 ;
        RECT 16.81 41.245 17.07 41.505 ;
        RECT 16.81 40.485 17.07 40.745 ;
        RECT 16.81 39.725 17.07 39.985 ;
        RECT 16.81 38.965 17.07 39.225 ;
        RECT 16.81 38.205 17.07 38.465 ;
        RECT 16.81 37.445 17.07 37.705 ;
        RECT 16.81 36.685 17.07 36.945 ;
        RECT 17.57 58.725 17.83 58.985 ;
        RECT 17.57 57.965 17.83 58.225 ;
        RECT 17.57 57.205 17.83 57.465 ;
        RECT 17.57 56.445 17.83 56.705 ;
        RECT 17.57 55.685 17.83 55.945 ;
        RECT 17.57 54.925 17.83 55.185 ;
        RECT 17.57 54.165 17.83 54.425 ;
        RECT 17.57 53.405 17.83 53.665 ;
        RECT 17.57 52.645 17.83 52.905 ;
        RECT 17.57 51.885 17.83 52.145 ;
        RECT 17.57 51.125 17.83 51.385 ;
        RECT 17.57 50.365 17.83 50.625 ;
        RECT 17.57 49.605 17.83 49.865 ;
        RECT 17.57 48.845 17.83 49.105 ;
        RECT 17.57 48.085 17.83 48.345 ;
        RECT 17.57 47.325 17.83 47.585 ;
        RECT 17.57 46.565 17.83 46.825 ;
        RECT 17.57 45.805 17.83 46.065 ;
        RECT 17.57 45.045 17.83 45.305 ;
        RECT 17.57 44.285 17.83 44.545 ;
        RECT 17.57 43.525 17.83 43.785 ;
        RECT 17.57 42.765 17.83 43.025 ;
        RECT 17.57 42.005 17.83 42.265 ;
        RECT 17.57 41.245 17.83 41.505 ;
        RECT 17.57 40.485 17.83 40.745 ;
        RECT 17.57 39.725 17.83 39.985 ;
        RECT 17.57 38.965 17.83 39.225 ;
        RECT 17.57 38.205 17.83 38.465 ;
        RECT 17.57 37.445 17.83 37.705 ;
        RECT 17.57 36.685 17.83 36.945 ;
        RECT 18.33 58.725 18.59 58.985 ;
        RECT 18.33 57.965 18.59 58.225 ;
        RECT 18.33 57.205 18.59 57.465 ;
        RECT 18.33 56.445 18.59 56.705 ;
        RECT 18.33 55.685 18.59 55.945 ;
        RECT 18.33 54.925 18.59 55.185 ;
        RECT 18.33 54.165 18.59 54.425 ;
        RECT 18.33 53.405 18.59 53.665 ;
        RECT 18.33 52.645 18.59 52.905 ;
        RECT 18.33 51.885 18.59 52.145 ;
        RECT 18.33 51.125 18.59 51.385 ;
        RECT 18.33 50.365 18.59 50.625 ;
        RECT 18.33 49.605 18.59 49.865 ;
        RECT 18.33 48.845 18.59 49.105 ;
        RECT 18.33 48.085 18.59 48.345 ;
        RECT 18.33 47.325 18.59 47.585 ;
        RECT 18.33 46.565 18.59 46.825 ;
        RECT 18.33 45.805 18.59 46.065 ;
        RECT 18.33 45.045 18.59 45.305 ;
        RECT 18.33 44.285 18.59 44.545 ;
        RECT 18.33 43.525 18.59 43.785 ;
        RECT 18.33 42.765 18.59 43.025 ;
        RECT 18.33 42.005 18.59 42.265 ;
        RECT 18.33 41.245 18.59 41.505 ;
        RECT 18.33 40.485 18.59 40.745 ;
        RECT 18.33 39.725 18.59 39.985 ;
        RECT 18.33 38.965 18.59 39.225 ;
        RECT 18.33 38.205 18.59 38.465 ;
        RECT 18.33 37.445 18.59 37.705 ;
        RECT 18.33 36.685 18.59 36.945 ;
        RECT 19.09 58.725 19.35 58.985 ;
        RECT 19.09 57.965 19.35 58.225 ;
        RECT 19.09 57.205 19.35 57.465 ;
        RECT 19.09 56.445 19.35 56.705 ;
        RECT 19.09 55.685 19.35 55.945 ;
        RECT 19.09 54.925 19.35 55.185 ;
        RECT 19.09 54.165 19.35 54.425 ;
        RECT 19.09 53.405 19.35 53.665 ;
        RECT 19.09 52.645 19.35 52.905 ;
        RECT 19.09 51.885 19.35 52.145 ;
        RECT 19.09 51.125 19.35 51.385 ;
        RECT 19.09 50.365 19.35 50.625 ;
        RECT 19.09 49.605 19.35 49.865 ;
        RECT 19.09 48.845 19.35 49.105 ;
        RECT 19.09 48.085 19.35 48.345 ;
        RECT 19.09 47.325 19.35 47.585 ;
        RECT 19.09 46.565 19.35 46.825 ;
        RECT 19.09 45.805 19.35 46.065 ;
        RECT 19.09 45.045 19.35 45.305 ;
        RECT 19.09 44.285 19.35 44.545 ;
        RECT 19.09 43.525 19.35 43.785 ;
        RECT 19.09 42.765 19.35 43.025 ;
        RECT 19.09 42.005 19.35 42.265 ;
        RECT 19.09 41.245 19.35 41.505 ;
        RECT 19.09 40.485 19.35 40.745 ;
        RECT 19.09 39.725 19.35 39.985 ;
        RECT 19.09 38.965 19.35 39.225 ;
        RECT 19.09 38.205 19.35 38.465 ;
        RECT 19.09 37.445 19.35 37.705 ;
        RECT 19.09 36.685 19.35 36.945 ;
        RECT 19.85 58.725 20.11 58.985 ;
        RECT 19.85 57.965 20.11 58.225 ;
        RECT 19.85 57.205 20.11 57.465 ;
        RECT 19.85 56.445 20.11 56.705 ;
        RECT 19.85 55.685 20.11 55.945 ;
        RECT 19.85 54.925 20.11 55.185 ;
        RECT 19.85 54.165 20.11 54.425 ;
        RECT 19.85 53.405 20.11 53.665 ;
        RECT 19.85 52.645 20.11 52.905 ;
        RECT 19.85 51.885 20.11 52.145 ;
        RECT 19.85 51.125 20.11 51.385 ;
        RECT 19.85 50.365 20.11 50.625 ;
        RECT 19.85 49.605 20.11 49.865 ;
        RECT 19.85 48.845 20.11 49.105 ;
        RECT 19.85 48.085 20.11 48.345 ;
        RECT 19.85 47.325 20.11 47.585 ;
        RECT 19.85 46.565 20.11 46.825 ;
        RECT 19.85 45.805 20.11 46.065 ;
        RECT 19.85 45.045 20.11 45.305 ;
        RECT 19.85 44.285 20.11 44.545 ;
        RECT 19.85 43.525 20.11 43.785 ;
        RECT 19.85 42.765 20.11 43.025 ;
        RECT 19.85 42.005 20.11 42.265 ;
        RECT 19.85 41.245 20.11 41.505 ;
        RECT 19.85 40.485 20.11 40.745 ;
        RECT 19.85 39.725 20.11 39.985 ;
        RECT 19.85 38.965 20.11 39.225 ;
        RECT 19.85 38.205 20.11 38.465 ;
        RECT 19.85 37.445 20.11 37.705 ;
        RECT 19.85 36.685 20.11 36.945 ;
        RECT 20.61 58.725 20.87 58.985 ;
        RECT 20.61 57.965 20.87 58.225 ;
        RECT 20.61 57.205 20.87 57.465 ;
        RECT 20.61 56.445 20.87 56.705 ;
        RECT 20.61 55.685 20.87 55.945 ;
        RECT 20.61 54.925 20.87 55.185 ;
        RECT 20.61 54.165 20.87 54.425 ;
        RECT 20.61 53.405 20.87 53.665 ;
        RECT 20.61 52.645 20.87 52.905 ;
        RECT 20.61 51.885 20.87 52.145 ;
        RECT 20.61 51.125 20.87 51.385 ;
        RECT 20.61 50.365 20.87 50.625 ;
        RECT 20.61 49.605 20.87 49.865 ;
        RECT 20.61 48.845 20.87 49.105 ;
        RECT 20.61 48.085 20.87 48.345 ;
        RECT 20.61 47.325 20.87 47.585 ;
        RECT 20.61 46.565 20.87 46.825 ;
        RECT 20.61 45.805 20.87 46.065 ;
        RECT 20.61 45.045 20.87 45.305 ;
        RECT 20.61 44.285 20.87 44.545 ;
        RECT 20.61 43.525 20.87 43.785 ;
        RECT 20.61 42.765 20.87 43.025 ;
        RECT 20.61 42.005 20.87 42.265 ;
        RECT 20.61 41.245 20.87 41.505 ;
        RECT 20.61 40.485 20.87 40.745 ;
        RECT 20.61 39.725 20.87 39.985 ;
        RECT 20.61 38.965 20.87 39.225 ;
        RECT 20.61 38.205 20.87 38.465 ;
        RECT 20.61 37.445 20.87 37.705 ;
        RECT 20.61 36.685 20.87 36.945 ;
        RECT 21.37 58.725 21.63 58.985 ;
        RECT 21.37 57.965 21.63 58.225 ;
        RECT 21.37 57.205 21.63 57.465 ;
        RECT 21.37 56.445 21.63 56.705 ;
        RECT 21.37 55.685 21.63 55.945 ;
        RECT 21.37 54.925 21.63 55.185 ;
        RECT 21.37 54.165 21.63 54.425 ;
        RECT 21.37 53.405 21.63 53.665 ;
        RECT 21.37 52.645 21.63 52.905 ;
        RECT 21.37 51.885 21.63 52.145 ;
        RECT 21.37 51.125 21.63 51.385 ;
        RECT 21.37 50.365 21.63 50.625 ;
        RECT 21.37 49.605 21.63 49.865 ;
        RECT 21.37 48.845 21.63 49.105 ;
        RECT 21.37 48.085 21.63 48.345 ;
        RECT 21.37 47.325 21.63 47.585 ;
        RECT 21.37 46.565 21.63 46.825 ;
        RECT 21.37 45.805 21.63 46.065 ;
        RECT 21.37 45.045 21.63 45.305 ;
        RECT 21.37 44.285 21.63 44.545 ;
        RECT 21.37 43.525 21.63 43.785 ;
        RECT 21.37 42.765 21.63 43.025 ;
        RECT 21.37 42.005 21.63 42.265 ;
        RECT 21.37 41.245 21.63 41.505 ;
        RECT 21.37 40.485 21.63 40.745 ;
        RECT 21.37 39.725 21.63 39.985 ;
        RECT 21.37 38.965 21.63 39.225 ;
        RECT 21.37 38.205 21.63 38.465 ;
        RECT 21.37 37.445 21.63 37.705 ;
        RECT 21.37 36.685 21.63 36.945 ;
        RECT 22.13 58.725 22.39 58.985 ;
        RECT 22.13 57.965 22.39 58.225 ;
        RECT 22.13 57.205 22.39 57.465 ;
        RECT 22.13 56.445 22.39 56.705 ;
        RECT 22.13 55.685 22.39 55.945 ;
        RECT 22.13 54.925 22.39 55.185 ;
        RECT 22.13 54.165 22.39 54.425 ;
        RECT 22.13 53.405 22.39 53.665 ;
        RECT 22.13 52.645 22.39 52.905 ;
        RECT 22.13 51.885 22.39 52.145 ;
        RECT 22.13 51.125 22.39 51.385 ;
        RECT 22.13 50.365 22.39 50.625 ;
        RECT 22.13 49.605 22.39 49.865 ;
        RECT 22.13 48.845 22.39 49.105 ;
        RECT 22.13 48.085 22.39 48.345 ;
        RECT 22.13 47.325 22.39 47.585 ;
        RECT 22.13 46.565 22.39 46.825 ;
        RECT 22.13 45.805 22.39 46.065 ;
        RECT 22.13 45.045 22.39 45.305 ;
        RECT 22.13 44.285 22.39 44.545 ;
        RECT 22.13 43.525 22.39 43.785 ;
        RECT 22.13 42.765 22.39 43.025 ;
        RECT 22.13 42.005 22.39 42.265 ;
        RECT 22.13 41.245 22.39 41.505 ;
        RECT 22.13 40.485 22.39 40.745 ;
        RECT 22.13 39.725 22.39 39.985 ;
        RECT 22.13 38.965 22.39 39.225 ;
        RECT 22.13 38.205 22.39 38.465 ;
        RECT 22.13 37.445 22.39 37.705 ;
        RECT 22.13 36.685 22.39 36.945 ;
        RECT 22.89 58.725 23.15 58.985 ;
        RECT 22.89 57.965 23.15 58.225 ;
        RECT 22.89 57.205 23.15 57.465 ;
        RECT 22.89 56.445 23.15 56.705 ;
        RECT 22.89 55.685 23.15 55.945 ;
        RECT 22.89 54.925 23.15 55.185 ;
        RECT 22.89 54.165 23.15 54.425 ;
        RECT 22.89 53.405 23.15 53.665 ;
        RECT 22.89 52.645 23.15 52.905 ;
        RECT 22.89 51.885 23.15 52.145 ;
        RECT 22.89 51.125 23.15 51.385 ;
        RECT 22.89 50.365 23.15 50.625 ;
        RECT 22.89 49.605 23.15 49.865 ;
        RECT 22.89 48.845 23.15 49.105 ;
        RECT 22.89 48.085 23.15 48.345 ;
        RECT 22.89 47.325 23.15 47.585 ;
        RECT 22.89 46.565 23.15 46.825 ;
        RECT 22.89 45.805 23.15 46.065 ;
        RECT 22.89 45.045 23.15 45.305 ;
        RECT 22.89 44.285 23.15 44.545 ;
        RECT 22.89 43.525 23.15 43.785 ;
        RECT 22.89 42.765 23.15 43.025 ;
        RECT 22.89 42.005 23.15 42.265 ;
        RECT 22.89 41.245 23.15 41.505 ;
        RECT 22.89 40.485 23.15 40.745 ;
        RECT 22.89 39.725 23.15 39.985 ;
        RECT 22.89 38.965 23.15 39.225 ;
        RECT 22.89 38.205 23.15 38.465 ;
        RECT 22.89 37.445 23.15 37.705 ;
        RECT 22.89 36.685 23.15 36.945 ;
        RECT 23.65 58.725 23.91 58.985 ;
        RECT 23.65 57.965 23.91 58.225 ;
        RECT 23.65 57.205 23.91 57.465 ;
        RECT 23.65 56.445 23.91 56.705 ;
        RECT 23.65 55.685 23.91 55.945 ;
        RECT 23.65 54.925 23.91 55.185 ;
        RECT 23.65 54.165 23.91 54.425 ;
        RECT 23.65 53.405 23.91 53.665 ;
        RECT 23.65 52.645 23.91 52.905 ;
        RECT 23.65 51.885 23.91 52.145 ;
        RECT 23.65 51.125 23.91 51.385 ;
        RECT 23.65 50.365 23.91 50.625 ;
        RECT 23.65 49.605 23.91 49.865 ;
        RECT 23.65 48.845 23.91 49.105 ;
        RECT 23.65 48.085 23.91 48.345 ;
        RECT 23.65 47.325 23.91 47.585 ;
        RECT 23.65 46.565 23.91 46.825 ;
        RECT 23.65 45.805 23.91 46.065 ;
        RECT 23.65 45.045 23.91 45.305 ;
        RECT 23.65 44.285 23.91 44.545 ;
        RECT 23.65 43.525 23.91 43.785 ;
        RECT 23.65 42.765 23.91 43.025 ;
        RECT 23.65 42.005 23.91 42.265 ;
        RECT 23.65 41.245 23.91 41.505 ;
        RECT 23.65 40.485 23.91 40.745 ;
        RECT 23.65 39.725 23.91 39.985 ;
        RECT 23.65 38.965 23.91 39.225 ;
        RECT 23.65 38.205 23.91 38.465 ;
        RECT 23.65 37.445 23.91 37.705 ;
        RECT 23.65 36.685 23.91 36.945 ;
        RECT 24.41 58.725 24.67 58.985 ;
        RECT 24.41 57.965 24.67 58.225 ;
        RECT 24.41 57.205 24.67 57.465 ;
        RECT 24.41 56.445 24.67 56.705 ;
        RECT 24.41 55.685 24.67 55.945 ;
        RECT 24.41 54.925 24.67 55.185 ;
        RECT 24.41 54.165 24.67 54.425 ;
        RECT 24.41 53.405 24.67 53.665 ;
        RECT 24.41 52.645 24.67 52.905 ;
        RECT 24.41 51.885 24.67 52.145 ;
        RECT 24.41 51.125 24.67 51.385 ;
        RECT 24.41 50.365 24.67 50.625 ;
        RECT 24.41 49.605 24.67 49.865 ;
        RECT 24.41 48.845 24.67 49.105 ;
        RECT 24.41 48.085 24.67 48.345 ;
        RECT 24.41 47.325 24.67 47.585 ;
        RECT 24.41 46.565 24.67 46.825 ;
        RECT 24.41 45.805 24.67 46.065 ;
        RECT 24.41 45.045 24.67 45.305 ;
        RECT 24.41 44.285 24.67 44.545 ;
        RECT 24.41 43.525 24.67 43.785 ;
        RECT 24.41 42.765 24.67 43.025 ;
        RECT 24.41 42.005 24.67 42.265 ;
        RECT 24.41 41.245 24.67 41.505 ;
        RECT 24.41 40.485 24.67 40.745 ;
        RECT 24.41 39.725 24.67 39.985 ;
        RECT 24.41 38.965 24.67 39.225 ;
        RECT 24.41 38.205 24.67 38.465 ;
        RECT 24.41 37.445 24.67 37.705 ;
        RECT 24.41 36.685 24.67 36.945 ;
        RECT 25.17 58.725 25.43 58.985 ;
        RECT 25.17 57.965 25.43 58.225 ;
        RECT 25.17 57.205 25.43 57.465 ;
        RECT 25.17 56.445 25.43 56.705 ;
        RECT 25.17 55.685 25.43 55.945 ;
        RECT 25.17 54.925 25.43 55.185 ;
        RECT 25.17 54.165 25.43 54.425 ;
        RECT 25.17 53.405 25.43 53.665 ;
        RECT 25.17 52.645 25.43 52.905 ;
        RECT 25.17 51.885 25.43 52.145 ;
        RECT 25.17 51.125 25.43 51.385 ;
        RECT 25.17 50.365 25.43 50.625 ;
        RECT 25.17 49.605 25.43 49.865 ;
        RECT 25.17 48.845 25.43 49.105 ;
        RECT 25.17 48.085 25.43 48.345 ;
        RECT 25.17 47.325 25.43 47.585 ;
        RECT 25.17 46.565 25.43 46.825 ;
        RECT 25.17 45.805 25.43 46.065 ;
        RECT 25.17 45.045 25.43 45.305 ;
        RECT 25.17 44.285 25.43 44.545 ;
        RECT 25.17 43.525 25.43 43.785 ;
        RECT 25.17 42.765 25.43 43.025 ;
        RECT 25.17 42.005 25.43 42.265 ;
        RECT 25.17 41.245 25.43 41.505 ;
        RECT 25.17 40.485 25.43 40.745 ;
        RECT 25.17 39.725 25.43 39.985 ;
        RECT 25.17 38.965 25.43 39.225 ;
        RECT 25.17 38.205 25.43 38.465 ;
        RECT 25.17 37.445 25.43 37.705 ;
        RECT 25.17 36.685 25.43 36.945 ;
        RECT 25.93 58.725 26.19 58.985 ;
        RECT 25.93 57.965 26.19 58.225 ;
        RECT 25.93 57.205 26.19 57.465 ;
        RECT 25.93 56.445 26.19 56.705 ;
        RECT 25.93 55.685 26.19 55.945 ;
        RECT 25.93 54.925 26.19 55.185 ;
        RECT 25.93 54.165 26.19 54.425 ;
        RECT 25.93 53.405 26.19 53.665 ;
        RECT 25.93 52.645 26.19 52.905 ;
        RECT 25.93 51.885 26.19 52.145 ;
        RECT 25.93 51.125 26.19 51.385 ;
        RECT 25.93 50.365 26.19 50.625 ;
        RECT 25.93 49.605 26.19 49.865 ;
        RECT 25.93 48.845 26.19 49.105 ;
        RECT 25.93 48.085 26.19 48.345 ;
        RECT 25.93 47.325 26.19 47.585 ;
        RECT 25.93 46.565 26.19 46.825 ;
        RECT 25.93 45.805 26.19 46.065 ;
        RECT 25.93 45.045 26.19 45.305 ;
        RECT 25.93 44.285 26.19 44.545 ;
        RECT 25.93 43.525 26.19 43.785 ;
        RECT 25.93 42.765 26.19 43.025 ;
        RECT 25.93 42.005 26.19 42.265 ;
        RECT 25.93 41.245 26.19 41.505 ;
        RECT 25.93 40.485 26.19 40.745 ;
        RECT 25.93 39.725 26.19 39.985 ;
        RECT 25.93 38.965 26.19 39.225 ;
        RECT 25.93 38.205 26.19 38.465 ;
        RECT 25.93 37.445 26.19 37.705 ;
        RECT 25.93 36.685 26.19 36.945 ;
        RECT 26.69 58.725 26.95 58.985 ;
        RECT 26.69 57.965 26.95 58.225 ;
        RECT 26.69 57.205 26.95 57.465 ;
        RECT 26.69 56.445 26.95 56.705 ;
        RECT 26.69 55.685 26.95 55.945 ;
        RECT 26.69 54.925 26.95 55.185 ;
        RECT 26.69 54.165 26.95 54.425 ;
        RECT 26.69 53.405 26.95 53.665 ;
        RECT 26.69 52.645 26.95 52.905 ;
        RECT 26.69 51.885 26.95 52.145 ;
        RECT 26.69 51.125 26.95 51.385 ;
        RECT 26.69 50.365 26.95 50.625 ;
        RECT 26.69 49.605 26.95 49.865 ;
        RECT 26.69 48.845 26.95 49.105 ;
        RECT 26.69 48.085 26.95 48.345 ;
        RECT 26.69 47.325 26.95 47.585 ;
        RECT 26.69 46.565 26.95 46.825 ;
        RECT 26.69 45.805 26.95 46.065 ;
        RECT 26.69 45.045 26.95 45.305 ;
        RECT 26.69 44.285 26.95 44.545 ;
        RECT 26.69 43.525 26.95 43.785 ;
        RECT 26.69 42.765 26.95 43.025 ;
        RECT 26.69 42.005 26.95 42.265 ;
        RECT 26.69 41.245 26.95 41.505 ;
        RECT 26.69 40.485 26.95 40.745 ;
        RECT 26.69 39.725 26.95 39.985 ;
        RECT 26.69 38.965 26.95 39.225 ;
        RECT 26.69 38.205 26.95 38.465 ;
        RECT 26.69 37.445 26.95 37.705 ;
        RECT 26.69 36.685 26.95 36.945 ;
        RECT 27.45 58.725 27.71 58.985 ;
        RECT 27.45 57.965 27.71 58.225 ;
        RECT 27.45 57.205 27.71 57.465 ;
        RECT 27.45 56.445 27.71 56.705 ;
        RECT 27.45 55.685 27.71 55.945 ;
        RECT 27.45 54.925 27.71 55.185 ;
        RECT 27.45 54.165 27.71 54.425 ;
        RECT 27.45 53.405 27.71 53.665 ;
        RECT 27.45 52.645 27.71 52.905 ;
        RECT 27.45 51.885 27.71 52.145 ;
        RECT 27.45 51.125 27.71 51.385 ;
        RECT 27.45 50.365 27.71 50.625 ;
        RECT 27.45 49.605 27.71 49.865 ;
        RECT 27.45 48.845 27.71 49.105 ;
        RECT 27.45 48.085 27.71 48.345 ;
        RECT 27.45 47.325 27.71 47.585 ;
        RECT 27.45 46.565 27.71 46.825 ;
        RECT 27.45 45.805 27.71 46.065 ;
        RECT 27.45 45.045 27.71 45.305 ;
        RECT 27.45 44.285 27.71 44.545 ;
        RECT 27.45 43.525 27.71 43.785 ;
        RECT 27.45 42.765 27.71 43.025 ;
        RECT 27.45 42.005 27.71 42.265 ;
        RECT 27.45 41.245 27.71 41.505 ;
        RECT 27.45 40.485 27.71 40.745 ;
        RECT 27.45 39.725 27.71 39.985 ;
        RECT 27.45 38.965 27.71 39.225 ;
        RECT 27.45 38.205 27.71 38.465 ;
        RECT 27.45 37.445 27.71 37.705 ;
        RECT 27.45 36.685 27.71 36.945 ;
        RECT 28.21 58.725 28.47 58.985 ;
        RECT 28.21 57.965 28.47 58.225 ;
        RECT 28.21 57.205 28.47 57.465 ;
        RECT 28.21 56.445 28.47 56.705 ;
        RECT 28.21 55.685 28.47 55.945 ;
        RECT 28.21 54.925 28.47 55.185 ;
        RECT 28.21 54.165 28.47 54.425 ;
        RECT 28.21 53.405 28.47 53.665 ;
        RECT 28.21 52.645 28.47 52.905 ;
        RECT 28.21 51.885 28.47 52.145 ;
        RECT 28.21 51.125 28.47 51.385 ;
        RECT 28.21 50.365 28.47 50.625 ;
        RECT 28.21 49.605 28.47 49.865 ;
        RECT 28.21 48.845 28.47 49.105 ;
        RECT 28.21 48.085 28.47 48.345 ;
        RECT 28.21 47.325 28.47 47.585 ;
        RECT 28.21 46.565 28.47 46.825 ;
        RECT 28.21 45.805 28.47 46.065 ;
        RECT 28.21 45.045 28.47 45.305 ;
        RECT 28.21 44.285 28.47 44.545 ;
        RECT 28.21 43.525 28.47 43.785 ;
        RECT 28.21 42.765 28.47 43.025 ;
        RECT 28.21 42.005 28.47 42.265 ;
        RECT 28.21 41.245 28.47 41.505 ;
        RECT 28.21 40.485 28.47 40.745 ;
        RECT 28.21 39.725 28.47 39.985 ;
        RECT 28.21 38.965 28.47 39.225 ;
        RECT 28.21 38.205 28.47 38.465 ;
        RECT 28.21 37.445 28.47 37.705 ;
        RECT 28.21 36.685 28.47 36.945 ;
        RECT 28.97 58.725 29.23 58.985 ;
        RECT 28.97 57.965 29.23 58.225 ;
        RECT 28.97 57.205 29.23 57.465 ;
        RECT 28.97 56.445 29.23 56.705 ;
        RECT 28.97 55.685 29.23 55.945 ;
        RECT 28.97 54.925 29.23 55.185 ;
        RECT 28.97 54.165 29.23 54.425 ;
        RECT 28.97 53.405 29.23 53.665 ;
        RECT 28.97 52.645 29.23 52.905 ;
        RECT 28.97 51.885 29.23 52.145 ;
        RECT 28.97 51.125 29.23 51.385 ;
        RECT 28.97 50.365 29.23 50.625 ;
        RECT 28.97 49.605 29.23 49.865 ;
        RECT 28.97 48.845 29.23 49.105 ;
        RECT 28.97 48.085 29.23 48.345 ;
        RECT 28.97 47.325 29.23 47.585 ;
        RECT 28.97 46.565 29.23 46.825 ;
        RECT 28.97 45.805 29.23 46.065 ;
        RECT 28.97 45.045 29.23 45.305 ;
        RECT 28.97 44.285 29.23 44.545 ;
        RECT 28.97 43.525 29.23 43.785 ;
        RECT 28.97 42.765 29.23 43.025 ;
        RECT 28.97 42.005 29.23 42.265 ;
        RECT 28.97 41.245 29.23 41.505 ;
        RECT 28.97 40.485 29.23 40.745 ;
        RECT 28.97 39.725 29.23 39.985 ;
        RECT 28.97 38.965 29.23 39.225 ;
        RECT 28.97 38.205 29.23 38.465 ;
        RECT 28.97 37.445 29.23 37.705 ;
        RECT 28.97 36.685 29.23 36.945 ;
        RECT 29.73 58.725 29.99 58.985 ;
        RECT 29.73 57.965 29.99 58.225 ;
        RECT 29.73 57.205 29.99 57.465 ;
        RECT 29.73 56.445 29.99 56.705 ;
        RECT 29.73 55.685 29.99 55.945 ;
        RECT 29.73 54.925 29.99 55.185 ;
        RECT 29.73 54.165 29.99 54.425 ;
        RECT 29.73 53.405 29.99 53.665 ;
        RECT 29.73 52.645 29.99 52.905 ;
        RECT 29.73 51.885 29.99 52.145 ;
      LAYER V5 ;
        RECT 80.65 58.775 80.91 59.035 ;
        RECT 80.65 58.015 80.91 58.275 ;
        RECT 80.65 57.255 80.91 57.515 ;
        RECT 80.65 56.495 80.91 56.755 ;
        RECT 80.65 55.735 80.91 55.995 ;
        RECT 80.65 54.975 80.91 55.235 ;
        RECT 80.65 54.215 80.91 54.475 ;
        RECT 80.65 53.455 80.91 53.715 ;
        RECT 80.65 52.695 80.91 52.955 ;
        RECT 80.65 51.935 80.91 52.195 ;
        RECT 80.65 51.175 80.91 51.435 ;
        RECT 80.65 50.415 80.91 50.675 ;
        RECT 80.65 49.655 80.91 49.915 ;
        RECT 80.65 48.895 80.91 49.155 ;
        RECT 80.65 48.135 80.91 48.395 ;
        RECT 80.65 47.375 80.91 47.635 ;
        RECT 80.65 46.615 80.91 46.875 ;
        RECT 80.65 45.855 80.91 46.115 ;
        RECT 80.65 45.095 80.91 45.355 ;
        RECT 80.65 44.335 80.91 44.595 ;
        RECT 80.65 43.575 80.91 43.835 ;
        RECT 80.65 42.815 80.91 43.075 ;
        RECT 80.65 42.055 80.91 42.315 ;
        RECT 80.65 41.295 80.91 41.555 ;
        RECT 80.65 40.535 80.91 40.795 ;
        RECT 80.65 39.775 80.91 40.035 ;
        RECT 80.65 39.015 80.91 39.275 ;
        RECT 80.65 38.255 80.91 38.515 ;
        RECT 80.65 37.495 80.91 37.755 ;
        RECT 80.65 36.735 80.91 36.995 ;
        RECT 81.41 58.775 81.67 59.035 ;
        RECT 81.41 58.015 81.67 58.275 ;
        RECT 81.41 57.255 81.67 57.515 ;
        RECT 81.41 56.495 81.67 56.755 ;
        RECT 81.41 55.735 81.67 55.995 ;
        RECT 81.41 54.975 81.67 55.235 ;
        RECT 81.41 54.215 81.67 54.475 ;
        RECT 81.41 53.455 81.67 53.715 ;
        RECT 81.41 52.695 81.67 52.955 ;
        RECT 81.41 51.935 81.67 52.195 ;
        RECT 81.41 51.175 81.67 51.435 ;
        RECT 81.41 50.415 81.67 50.675 ;
        RECT 81.41 49.655 81.67 49.915 ;
        RECT 81.41 48.895 81.67 49.155 ;
        RECT 81.41 48.135 81.67 48.395 ;
        RECT 81.41 47.375 81.67 47.635 ;
        RECT 81.41 46.615 81.67 46.875 ;
        RECT 81.41 45.855 81.67 46.115 ;
        RECT 81.41 45.095 81.67 45.355 ;
        RECT 81.41 44.335 81.67 44.595 ;
        RECT 81.41 43.575 81.67 43.835 ;
        RECT 81.41 42.815 81.67 43.075 ;
        RECT 81.41 42.055 81.67 42.315 ;
        RECT 81.41 41.295 81.67 41.555 ;
        RECT 81.41 40.535 81.67 40.795 ;
        RECT 81.41 39.775 81.67 40.035 ;
        RECT 81.41 39.015 81.67 39.275 ;
        RECT 81.41 38.255 81.67 38.515 ;
        RECT 81.41 37.495 81.67 37.755 ;
        RECT 81.41 36.735 81.67 36.995 ;
        RECT 82.17 58.775 82.43 59.035 ;
        RECT 82.17 58.015 82.43 58.275 ;
        RECT 82.17 57.255 82.43 57.515 ;
        RECT 82.17 56.495 82.43 56.755 ;
        RECT 82.17 55.735 82.43 55.995 ;
        RECT 82.17 54.975 82.43 55.235 ;
        RECT 82.17 54.215 82.43 54.475 ;
        RECT 82.17 53.455 82.43 53.715 ;
        RECT 82.17 52.695 82.43 52.955 ;
        RECT 82.17 51.935 82.43 52.195 ;
        RECT 82.17 51.175 82.43 51.435 ;
        RECT 82.17 50.415 82.43 50.675 ;
        RECT 82.17 49.655 82.43 49.915 ;
        RECT 82.17 48.895 82.43 49.155 ;
        RECT 82.17 48.135 82.43 48.395 ;
        RECT 82.17 47.375 82.43 47.635 ;
        RECT 82.17 46.615 82.43 46.875 ;
        RECT 82.17 45.855 82.43 46.115 ;
        RECT 82.17 45.095 82.43 45.355 ;
        RECT 82.17 44.335 82.43 44.595 ;
        RECT 82.17 43.575 82.43 43.835 ;
        RECT 82.17 42.815 82.43 43.075 ;
        RECT 82.17 42.055 82.43 42.315 ;
        RECT 82.17 41.295 82.43 41.555 ;
        RECT 82.17 40.535 82.43 40.795 ;
        RECT 82.17 39.775 82.43 40.035 ;
        RECT 82.17 39.015 82.43 39.275 ;
        RECT 82.17 38.255 82.43 38.515 ;
        RECT 82.17 37.495 82.43 37.755 ;
        RECT 82.17 36.735 82.43 36.995 ;
        RECT 82.93 58.775 83.19 59.035 ;
        RECT 82.93 58.015 83.19 58.275 ;
        RECT 82.93 57.255 83.19 57.515 ;
        RECT 82.93 56.495 83.19 56.755 ;
        RECT 82.93 55.735 83.19 55.995 ;
        RECT 82.93 54.975 83.19 55.235 ;
        RECT 82.93 54.215 83.19 54.475 ;
        RECT 82.93 53.455 83.19 53.715 ;
        RECT 82.93 52.695 83.19 52.955 ;
        RECT 82.93 51.935 83.19 52.195 ;
        RECT 82.93 51.175 83.19 51.435 ;
        RECT 82.93 50.415 83.19 50.675 ;
        RECT 82.93 49.655 83.19 49.915 ;
        RECT 82.93 48.895 83.19 49.155 ;
        RECT 82.93 48.135 83.19 48.395 ;
        RECT 82.93 47.375 83.19 47.635 ;
        RECT 82.93 46.615 83.19 46.875 ;
        RECT 82.93 45.855 83.19 46.115 ;
        RECT 82.93 45.095 83.19 45.355 ;
        RECT 82.93 44.335 83.19 44.595 ;
        RECT 82.93 43.575 83.19 43.835 ;
        RECT 82.93 42.815 83.19 43.075 ;
        RECT 82.93 42.055 83.19 42.315 ;
        RECT 82.93 41.295 83.19 41.555 ;
        RECT 82.93 40.535 83.19 40.795 ;
        RECT 82.93 39.775 83.19 40.035 ;
        RECT 82.93 39.015 83.19 39.275 ;
        RECT 82.93 38.255 83.19 38.515 ;
        RECT 82.93 37.495 83.19 37.755 ;
        RECT 82.93 36.735 83.19 36.995 ;
        RECT 83.69 58.775 83.95 59.035 ;
        RECT 83.69 58.015 83.95 58.275 ;
        RECT 83.69 57.255 83.95 57.515 ;
        RECT 83.69 56.495 83.95 56.755 ;
        RECT 83.69 55.735 83.95 55.995 ;
        RECT 83.69 54.975 83.95 55.235 ;
        RECT 83.69 54.215 83.95 54.475 ;
        RECT 83.69 53.455 83.95 53.715 ;
        RECT 83.69 52.695 83.95 52.955 ;
        RECT 83.69 51.935 83.95 52.195 ;
        RECT 83.69 51.175 83.95 51.435 ;
        RECT 83.69 50.415 83.95 50.675 ;
        RECT 83.69 49.655 83.95 49.915 ;
        RECT 83.69 48.895 83.95 49.155 ;
        RECT 83.69 48.135 83.95 48.395 ;
        RECT 83.69 47.375 83.95 47.635 ;
        RECT 83.69 46.615 83.95 46.875 ;
        RECT 83.69 45.855 83.95 46.115 ;
        RECT 83.69 45.095 83.95 45.355 ;
        RECT 83.69 44.335 83.95 44.595 ;
        RECT 83.69 43.575 83.95 43.835 ;
        RECT 83.69 42.815 83.95 43.075 ;
        RECT 83.69 42.055 83.95 42.315 ;
        RECT 83.69 41.295 83.95 41.555 ;
        RECT 83.69 40.535 83.95 40.795 ;
        RECT 83.69 39.775 83.95 40.035 ;
        RECT 83.69 39.015 83.95 39.275 ;
        RECT 83.69 38.255 83.95 38.515 ;
        RECT 83.69 37.495 83.95 37.755 ;
        RECT 83.69 36.735 83.95 36.995 ;
        RECT 84.45 58.775 84.71 59.035 ;
        RECT 84.45 58.015 84.71 58.275 ;
        RECT 84.45 57.255 84.71 57.515 ;
        RECT 84.45 56.495 84.71 56.755 ;
        RECT 84.45 55.735 84.71 55.995 ;
        RECT 84.45 54.975 84.71 55.235 ;
        RECT 84.45 54.215 84.71 54.475 ;
        RECT 84.45 53.455 84.71 53.715 ;
        RECT 84.45 52.695 84.71 52.955 ;
        RECT 84.45 51.935 84.71 52.195 ;
        RECT 84.45 51.175 84.71 51.435 ;
        RECT 84.45 50.415 84.71 50.675 ;
        RECT 84.45 49.655 84.71 49.915 ;
        RECT 84.45 48.895 84.71 49.155 ;
        RECT 84.45 48.135 84.71 48.395 ;
        RECT 84.45 47.375 84.71 47.635 ;
        RECT 84.45 46.615 84.71 46.875 ;
        RECT 84.45 45.855 84.71 46.115 ;
        RECT 84.45 45.095 84.71 45.355 ;
        RECT 84.45 44.335 84.71 44.595 ;
        RECT 84.45 43.575 84.71 43.835 ;
        RECT 84.45 42.815 84.71 43.075 ;
        RECT 84.45 42.055 84.71 42.315 ;
        RECT 84.45 41.295 84.71 41.555 ;
        RECT 84.45 40.535 84.71 40.795 ;
        RECT 84.45 39.775 84.71 40.035 ;
        RECT 84.45 39.015 84.71 39.275 ;
        RECT 84.45 38.255 84.71 38.515 ;
        RECT 84.45 37.495 84.71 37.755 ;
        RECT 84.45 36.735 84.71 36.995 ;
        RECT 85.21 58.775 85.47 59.035 ;
        RECT 85.21 58.015 85.47 58.275 ;
        RECT 85.21 57.255 85.47 57.515 ;
        RECT 85.21 56.495 85.47 56.755 ;
        RECT 85.21 55.735 85.47 55.995 ;
        RECT 85.21 54.975 85.47 55.235 ;
        RECT 85.21 54.215 85.47 54.475 ;
        RECT 85.21 53.455 85.47 53.715 ;
        RECT 85.21 52.695 85.47 52.955 ;
        RECT 85.21 51.935 85.47 52.195 ;
        RECT 85.21 51.175 85.47 51.435 ;
        RECT 85.21 50.415 85.47 50.675 ;
        RECT 85.21 49.655 85.47 49.915 ;
        RECT 85.21 48.895 85.47 49.155 ;
        RECT 85.21 48.135 85.47 48.395 ;
        RECT 85.21 47.375 85.47 47.635 ;
        RECT 85.21 46.615 85.47 46.875 ;
        RECT 85.21 45.855 85.47 46.115 ;
        RECT 85.21 45.095 85.47 45.355 ;
        RECT 85.21 44.335 85.47 44.595 ;
        RECT 85.21 43.575 85.47 43.835 ;
        RECT 85.21 42.815 85.47 43.075 ;
        RECT 85.21 42.055 85.47 42.315 ;
        RECT 85.21 41.295 85.47 41.555 ;
        RECT 85.21 40.535 85.47 40.795 ;
        RECT 85.21 39.775 85.47 40.035 ;
        RECT 85.21 39.015 85.47 39.275 ;
        RECT 85.21 38.255 85.47 38.515 ;
        RECT 85.21 37.495 85.47 37.755 ;
        RECT 85.21 36.735 85.47 36.995 ;
        RECT 85.97 58.775 86.23 59.035 ;
        RECT 85.97 58.015 86.23 58.275 ;
        RECT 85.97 57.255 86.23 57.515 ;
        RECT 85.97 56.495 86.23 56.755 ;
        RECT 85.97 55.735 86.23 55.995 ;
        RECT 85.97 54.975 86.23 55.235 ;
        RECT 85.97 54.215 86.23 54.475 ;
        RECT 85.97 53.455 86.23 53.715 ;
        RECT 85.97 52.695 86.23 52.955 ;
        RECT 85.97 51.935 86.23 52.195 ;
        RECT 85.97 51.175 86.23 51.435 ;
        RECT 85.97 50.415 86.23 50.675 ;
        RECT 85.97 49.655 86.23 49.915 ;
        RECT 85.97 48.895 86.23 49.155 ;
        RECT 85.97 48.135 86.23 48.395 ;
        RECT 85.97 47.375 86.23 47.635 ;
        RECT 85.97 46.615 86.23 46.875 ;
        RECT 85.97 45.855 86.23 46.115 ;
        RECT 85.97 45.095 86.23 45.355 ;
        RECT 85.97 44.335 86.23 44.595 ;
        RECT 85.97 43.575 86.23 43.835 ;
        RECT 85.97 42.815 86.23 43.075 ;
        RECT 85.97 42.055 86.23 42.315 ;
        RECT 85.97 41.295 86.23 41.555 ;
        RECT 85.97 40.535 86.23 40.795 ;
        RECT 85.97 39.775 86.23 40.035 ;
        RECT 85.97 39.015 86.23 39.275 ;
        RECT 85.97 38.255 86.23 38.515 ;
        RECT 85.97 37.495 86.23 37.755 ;
        RECT 85.97 36.735 86.23 36.995 ;
        RECT 86.73 58.775 86.99 59.035 ;
        RECT 86.73 58.015 86.99 58.275 ;
        RECT 86.73 57.255 86.99 57.515 ;
        RECT 86.73 56.495 86.99 56.755 ;
        RECT 86.73 55.735 86.99 55.995 ;
        RECT 86.73 54.975 86.99 55.235 ;
        RECT 86.73 54.215 86.99 54.475 ;
        RECT 86.73 53.455 86.99 53.715 ;
        RECT 86.73 52.695 86.99 52.955 ;
        RECT 86.73 51.935 86.99 52.195 ;
        RECT 86.73 51.175 86.99 51.435 ;
        RECT 86.73 50.415 86.99 50.675 ;
        RECT 86.73 49.655 86.99 49.915 ;
        RECT 86.73 48.895 86.99 49.155 ;
        RECT 86.73 48.135 86.99 48.395 ;
        RECT 86.73 47.375 86.99 47.635 ;
        RECT 86.73 46.615 86.99 46.875 ;
        RECT 86.73 45.855 86.99 46.115 ;
        RECT 86.73 45.095 86.99 45.355 ;
        RECT 86.73 44.335 86.99 44.595 ;
        RECT 86.73 43.575 86.99 43.835 ;
        RECT 86.73 42.815 86.99 43.075 ;
        RECT 86.73 42.055 86.99 42.315 ;
        RECT 86.73 41.295 86.99 41.555 ;
        RECT 86.73 40.535 86.99 40.795 ;
        RECT 86.73 39.775 86.99 40.035 ;
        RECT 86.73 39.015 86.99 39.275 ;
        RECT 86.73 38.255 86.99 38.515 ;
        RECT 86.73 37.495 86.99 37.755 ;
        RECT 86.73 36.735 86.99 36.995 ;
        RECT 87.49 58.775 87.75 59.035 ;
        RECT 87.49 58.015 87.75 58.275 ;
        RECT 87.49 57.255 87.75 57.515 ;
        RECT 87.49 56.495 87.75 56.755 ;
        RECT 87.49 55.735 87.75 55.995 ;
        RECT 87.49 54.975 87.75 55.235 ;
        RECT 87.49 54.215 87.75 54.475 ;
        RECT 87.49 53.455 87.75 53.715 ;
        RECT 87.49 52.695 87.75 52.955 ;
        RECT 87.49 51.935 87.75 52.195 ;
        RECT 87.49 51.175 87.75 51.435 ;
        RECT 87.49 50.415 87.75 50.675 ;
        RECT 87.49 49.655 87.75 49.915 ;
        RECT 87.49 48.895 87.75 49.155 ;
        RECT 87.49 48.135 87.75 48.395 ;
        RECT 87.49 47.375 87.75 47.635 ;
        RECT 87.49 46.615 87.75 46.875 ;
        RECT 87.49 45.855 87.75 46.115 ;
        RECT 87.49 45.095 87.75 45.355 ;
        RECT 87.49 44.335 87.75 44.595 ;
        RECT 87.49 43.575 87.75 43.835 ;
        RECT 87.49 42.815 87.75 43.075 ;
        RECT 87.49 42.055 87.75 42.315 ;
        RECT 87.49 41.295 87.75 41.555 ;
        RECT 87.49 40.535 87.75 40.795 ;
        RECT 87.49 39.775 87.75 40.035 ;
        RECT 87.49 39.015 87.75 39.275 ;
        RECT 87.49 38.255 87.75 38.515 ;
        RECT 87.49 37.495 87.75 37.755 ;
        RECT 87.49 36.735 87.75 36.995 ;
        RECT 88.25 58.775 88.51 59.035 ;
        RECT 88.25 58.015 88.51 58.275 ;
        RECT 88.25 57.255 88.51 57.515 ;
        RECT 88.25 56.495 88.51 56.755 ;
        RECT 88.25 55.735 88.51 55.995 ;
        RECT 88.25 54.975 88.51 55.235 ;
        RECT 88.25 54.215 88.51 54.475 ;
        RECT 88.25 53.455 88.51 53.715 ;
        RECT 88.25 52.695 88.51 52.955 ;
        RECT 88.25 51.935 88.51 52.195 ;
        RECT 88.25 51.175 88.51 51.435 ;
        RECT 88.25 50.415 88.51 50.675 ;
        RECT 88.25 49.655 88.51 49.915 ;
        RECT 88.25 48.895 88.51 49.155 ;
        RECT 88.25 48.135 88.51 48.395 ;
        RECT 88.25 47.375 88.51 47.635 ;
        RECT 88.25 46.615 88.51 46.875 ;
        RECT 88.25 45.855 88.51 46.115 ;
        RECT 88.25 45.095 88.51 45.355 ;
        RECT 88.25 44.335 88.51 44.595 ;
        RECT 88.25 43.575 88.51 43.835 ;
        RECT 88.25 42.815 88.51 43.075 ;
        RECT 88.25 42.055 88.51 42.315 ;
        RECT 88.25 41.295 88.51 41.555 ;
        RECT 88.25 40.535 88.51 40.795 ;
        RECT 88.25 39.775 88.51 40.035 ;
        RECT 88.25 39.015 88.51 39.275 ;
        RECT 88.25 38.255 88.51 38.515 ;
        RECT 88.25 37.495 88.51 37.755 ;
        RECT 88.25 36.735 88.51 36.995 ;
        RECT 89.01 58.775 89.27 59.035 ;
        RECT 89.01 58.015 89.27 58.275 ;
        RECT 89.01 57.255 89.27 57.515 ;
        RECT 89.01 56.495 89.27 56.755 ;
        RECT 89.01 55.735 89.27 55.995 ;
        RECT 89.01 54.975 89.27 55.235 ;
        RECT 89.01 54.215 89.27 54.475 ;
        RECT 89.01 53.455 89.27 53.715 ;
        RECT 89.01 52.695 89.27 52.955 ;
        RECT 89.01 51.935 89.27 52.195 ;
        RECT 89.01 51.175 89.27 51.435 ;
        RECT 89.01 50.415 89.27 50.675 ;
        RECT 89.01 49.655 89.27 49.915 ;
        RECT 89.01 48.895 89.27 49.155 ;
        RECT 89.01 48.135 89.27 48.395 ;
        RECT 89.01 47.375 89.27 47.635 ;
        RECT 89.01 46.615 89.27 46.875 ;
        RECT 89.01 45.855 89.27 46.115 ;
        RECT 89.01 45.095 89.27 45.355 ;
        RECT 89.01 44.335 89.27 44.595 ;
        RECT 89.01 43.575 89.27 43.835 ;
        RECT 89.01 42.815 89.27 43.075 ;
        RECT 89.01 42.055 89.27 42.315 ;
        RECT 89.01 41.295 89.27 41.555 ;
        RECT 89.01 40.535 89.27 40.795 ;
        RECT 89.01 39.775 89.27 40.035 ;
        RECT 89.01 39.015 89.27 39.275 ;
        RECT 89.01 38.255 89.27 38.515 ;
        RECT 89.01 37.495 89.27 37.755 ;
        RECT 89.01 36.735 89.27 36.995 ;
        RECT 89.77 58.775 90.03 59.035 ;
        RECT 89.77 58.015 90.03 58.275 ;
        RECT 89.77 57.255 90.03 57.515 ;
        RECT 89.77 56.495 90.03 56.755 ;
        RECT 89.77 55.735 90.03 55.995 ;
        RECT 89.77 54.975 90.03 55.235 ;
        RECT 89.77 54.215 90.03 54.475 ;
        RECT 89.77 53.455 90.03 53.715 ;
        RECT 89.77 52.695 90.03 52.955 ;
        RECT 89.77 51.935 90.03 52.195 ;
        RECT 89.77 51.175 90.03 51.435 ;
        RECT 89.77 50.415 90.03 50.675 ;
        RECT 89.77 49.655 90.03 49.915 ;
        RECT 89.77 48.895 90.03 49.155 ;
        RECT 89.77 48.135 90.03 48.395 ;
        RECT 89.77 47.375 90.03 47.635 ;
        RECT 89.77 46.615 90.03 46.875 ;
        RECT 89.77 45.855 90.03 46.115 ;
        RECT 89.77 45.095 90.03 45.355 ;
        RECT 89.77 44.335 90.03 44.595 ;
        RECT 89.77 43.575 90.03 43.835 ;
        RECT 89.77 42.815 90.03 43.075 ;
        RECT 89.77 42.055 90.03 42.315 ;
        RECT 89.77 41.295 90.03 41.555 ;
        RECT 89.77 40.535 90.03 40.795 ;
        RECT 89.77 39.775 90.03 40.035 ;
        RECT 89.77 39.015 90.03 39.275 ;
        RECT 89.77 38.255 90.03 38.515 ;
        RECT 89.77 37.495 90.03 37.755 ;
        RECT 89.77 36.735 90.03 36.995 ;
        RECT 90.53 58.775 90.79 59.035 ;
        RECT 90.53 58.015 90.79 58.275 ;
        RECT 90.53 57.255 90.79 57.515 ;
        RECT 90.53 56.495 90.79 56.755 ;
        RECT 90.53 55.735 90.79 55.995 ;
        RECT 90.53 54.975 90.79 55.235 ;
        RECT 90.53 54.215 90.79 54.475 ;
        RECT 90.53 53.455 90.79 53.715 ;
        RECT 90.53 52.695 90.79 52.955 ;
        RECT 90.53 51.935 90.79 52.195 ;
        RECT 90.53 51.175 90.79 51.435 ;
        RECT 90.53 50.415 90.79 50.675 ;
        RECT 90.53 49.655 90.79 49.915 ;
        RECT 90.53 48.895 90.79 49.155 ;
        RECT 90.53 48.135 90.79 48.395 ;
        RECT 90.53 47.375 90.79 47.635 ;
        RECT 90.53 46.615 90.79 46.875 ;
        RECT 90.53 45.855 90.79 46.115 ;
        RECT 90.53 45.095 90.79 45.355 ;
        RECT 90.53 44.335 90.79 44.595 ;
        RECT 90.53 43.575 90.79 43.835 ;
        RECT 90.53 42.815 90.79 43.075 ;
        RECT 90.53 42.055 90.79 42.315 ;
        RECT 90.53 41.295 90.79 41.555 ;
        RECT 90.53 40.535 90.79 40.795 ;
        RECT 90.53 39.775 90.79 40.035 ;
        RECT 90.53 39.015 90.79 39.275 ;
        RECT 90.53 38.255 90.79 38.515 ;
        RECT 90.53 37.495 90.79 37.755 ;
        RECT 90.53 36.735 90.79 36.995 ;
        RECT 91.29 58.775 91.55 59.035 ;
        RECT 91.29 58.015 91.55 58.275 ;
        RECT 91.29 57.255 91.55 57.515 ;
        RECT 91.29 56.495 91.55 56.755 ;
        RECT 91.29 55.735 91.55 55.995 ;
        RECT 91.29 54.975 91.55 55.235 ;
        RECT 91.29 54.215 91.55 54.475 ;
        RECT 91.29 53.455 91.55 53.715 ;
        RECT 91.29 52.695 91.55 52.955 ;
        RECT 91.29 51.935 91.55 52.195 ;
        RECT 91.29 51.175 91.55 51.435 ;
        RECT 91.29 50.415 91.55 50.675 ;
        RECT 91.29 49.655 91.55 49.915 ;
        RECT 91.29 48.895 91.55 49.155 ;
        RECT 91.29 48.135 91.55 48.395 ;
        RECT 91.29 47.375 91.55 47.635 ;
        RECT 91.29 46.615 91.55 46.875 ;
        RECT 91.29 45.855 91.55 46.115 ;
        RECT 91.29 45.095 91.55 45.355 ;
        RECT 91.29 44.335 91.55 44.595 ;
        RECT 91.29 43.575 91.55 43.835 ;
        RECT 91.29 42.815 91.55 43.075 ;
        RECT 91.29 42.055 91.55 42.315 ;
        RECT 91.29 41.295 91.55 41.555 ;
        RECT 91.29 40.535 91.55 40.795 ;
        RECT 91.29 39.775 91.55 40.035 ;
        RECT 91.29 39.015 91.55 39.275 ;
        RECT 91.29 38.255 91.55 38.515 ;
        RECT 91.29 37.495 91.55 37.755 ;
        RECT 91.29 36.735 91.55 36.995 ;
        RECT 92.05 58.775 92.31 59.035 ;
        RECT 92.05 58.015 92.31 58.275 ;
        RECT 92.05 57.255 92.31 57.515 ;
        RECT 92.05 56.495 92.31 56.755 ;
        RECT 92.05 55.735 92.31 55.995 ;
        RECT 92.05 54.975 92.31 55.235 ;
        RECT 92.05 54.215 92.31 54.475 ;
        RECT 92.05 53.455 92.31 53.715 ;
        RECT 92.05 52.695 92.31 52.955 ;
        RECT 92.05 51.935 92.31 52.195 ;
        RECT 92.05 51.175 92.31 51.435 ;
        RECT 92.05 50.415 92.31 50.675 ;
        RECT 92.05 49.655 92.31 49.915 ;
        RECT 92.05 48.895 92.31 49.155 ;
        RECT 92.05 48.135 92.31 48.395 ;
        RECT 92.05 47.375 92.31 47.635 ;
        RECT 92.05 46.615 92.31 46.875 ;
        RECT 92.05 45.855 92.31 46.115 ;
        RECT 92.05 45.095 92.31 45.355 ;
        RECT 92.05 44.335 92.31 44.595 ;
        RECT 92.05 43.575 92.31 43.835 ;
        RECT 92.05 42.815 92.31 43.075 ;
        RECT 92.05 42.055 92.31 42.315 ;
        RECT 92.05 41.295 92.31 41.555 ;
        RECT 92.05 40.535 92.31 40.795 ;
        RECT 92.05 39.775 92.31 40.035 ;
        RECT 92.05 39.015 92.31 39.275 ;
        RECT 92.05 38.255 92.31 38.515 ;
        RECT 92.05 37.495 92.31 37.755 ;
        RECT 92.05 36.735 92.31 36.995 ;
        RECT 92.81 58.775 93.07 59.035 ;
        RECT 92.81 58.015 93.07 58.275 ;
        RECT 92.81 57.255 93.07 57.515 ;
        RECT 92.81 56.495 93.07 56.755 ;
        RECT 92.81 55.735 93.07 55.995 ;
        RECT 92.81 54.975 93.07 55.235 ;
        RECT 92.81 54.215 93.07 54.475 ;
        RECT 92.81 53.455 93.07 53.715 ;
        RECT 92.81 52.695 93.07 52.955 ;
        RECT 92.81 51.935 93.07 52.195 ;
        RECT 92.81 51.175 93.07 51.435 ;
        RECT 92.81 50.415 93.07 50.675 ;
        RECT 92.81 49.655 93.07 49.915 ;
        RECT 92.81 48.895 93.07 49.155 ;
        RECT 92.81 48.135 93.07 48.395 ;
        RECT 92.81 47.375 93.07 47.635 ;
        RECT 92.81 46.615 93.07 46.875 ;
        RECT 92.81 45.855 93.07 46.115 ;
        RECT 92.81 45.095 93.07 45.355 ;
        RECT 92.81 44.335 93.07 44.595 ;
        RECT 92.81 43.575 93.07 43.835 ;
        RECT 92.81 42.815 93.07 43.075 ;
        RECT 92.81 42.055 93.07 42.315 ;
        RECT 92.81 41.295 93.07 41.555 ;
        RECT 92.81 40.535 93.07 40.795 ;
        RECT 92.81 39.775 93.07 40.035 ;
        RECT 92.81 39.015 93.07 39.275 ;
        RECT 92.81 38.255 93.07 38.515 ;
        RECT 92.81 37.495 93.07 37.755 ;
        RECT 92.81 36.735 93.07 36.995 ;
        RECT 93.57 58.775 93.83 59.035 ;
        RECT 93.57 58.015 93.83 58.275 ;
        RECT 93.57 57.255 93.83 57.515 ;
        RECT 93.57 56.495 93.83 56.755 ;
        RECT 93.57 55.735 93.83 55.995 ;
        RECT 93.57 54.975 93.83 55.235 ;
        RECT 93.57 54.215 93.83 54.475 ;
        RECT 93.57 53.455 93.83 53.715 ;
        RECT 93.57 52.695 93.83 52.955 ;
        RECT 93.57 51.935 93.83 52.195 ;
        RECT 93.57 51.175 93.83 51.435 ;
        RECT 93.57 50.415 93.83 50.675 ;
        RECT 93.57 49.655 93.83 49.915 ;
        RECT 93.57 48.895 93.83 49.155 ;
        RECT 93.57 48.135 93.83 48.395 ;
        RECT 93.57 47.375 93.83 47.635 ;
        RECT 93.57 46.615 93.83 46.875 ;
        RECT 93.57 45.855 93.83 46.115 ;
        RECT 93.57 45.095 93.83 45.355 ;
        RECT 93.57 44.335 93.83 44.595 ;
        RECT 93.57 43.575 93.83 43.835 ;
        RECT 93.57 42.815 93.83 43.075 ;
        RECT 93.57 42.055 93.83 42.315 ;
        RECT 93.57 41.295 93.83 41.555 ;
        RECT 93.57 40.535 93.83 40.795 ;
        RECT 93.57 39.775 93.83 40.035 ;
        RECT 93.57 39.015 93.83 39.275 ;
        RECT 93.57 38.255 93.83 38.515 ;
        RECT 93.57 37.495 93.83 37.755 ;
        RECT 93.57 36.735 93.83 36.995 ;
        RECT 94.33 58.775 94.59 59.035 ;
        RECT 94.33 58.015 94.59 58.275 ;
        RECT 94.33 57.255 94.59 57.515 ;
        RECT 94.33 56.495 94.59 56.755 ;
        RECT 94.33 55.735 94.59 55.995 ;
        RECT 94.33 54.975 94.59 55.235 ;
        RECT 94.33 54.215 94.59 54.475 ;
        RECT 94.33 53.455 94.59 53.715 ;
        RECT 94.33 52.695 94.59 52.955 ;
        RECT 94.33 51.935 94.59 52.195 ;
        RECT 94.33 51.175 94.59 51.435 ;
        RECT 94.33 50.415 94.59 50.675 ;
        RECT 94.33 49.655 94.59 49.915 ;
        RECT 94.33 48.895 94.59 49.155 ;
        RECT 94.33 48.135 94.59 48.395 ;
        RECT 94.33 47.375 94.59 47.635 ;
        RECT 94.33 46.615 94.59 46.875 ;
        RECT 94.33 45.855 94.59 46.115 ;
        RECT 94.33 45.095 94.59 45.355 ;
        RECT 94.33 44.335 94.59 44.595 ;
        RECT 94.33 43.575 94.59 43.835 ;
        RECT 94.33 42.815 94.59 43.075 ;
        RECT 94.33 42.055 94.59 42.315 ;
        RECT 94.33 41.295 94.59 41.555 ;
        RECT 94.33 40.535 94.59 40.795 ;
        RECT 94.33 39.775 94.59 40.035 ;
        RECT 94.33 39.015 94.59 39.275 ;
        RECT 94.33 38.255 94.59 38.515 ;
        RECT 94.33 37.495 94.59 37.755 ;
        RECT 94.33 36.735 94.59 36.995 ;
        RECT 95.09 58.775 95.35 59.035 ;
        RECT 95.09 58.015 95.35 58.275 ;
        RECT 95.09 57.255 95.35 57.515 ;
        RECT 95.09 56.495 95.35 56.755 ;
        RECT 95.09 55.735 95.35 55.995 ;
        RECT 95.09 54.975 95.35 55.235 ;
        RECT 95.09 54.215 95.35 54.475 ;
        RECT 95.09 53.455 95.35 53.715 ;
        RECT 95.09 52.695 95.35 52.955 ;
        RECT 95.09 51.935 95.35 52.195 ;
        RECT 95.09 51.175 95.35 51.435 ;
        RECT 95.09 50.415 95.35 50.675 ;
        RECT 95.09 49.655 95.35 49.915 ;
        RECT 95.09 48.895 95.35 49.155 ;
        RECT 95.09 48.135 95.35 48.395 ;
        RECT 95.09 47.375 95.35 47.635 ;
        RECT 95.09 46.615 95.35 46.875 ;
        RECT 95.09 45.855 95.35 46.115 ;
        RECT 95.09 45.095 95.35 45.355 ;
        RECT 95.09 44.335 95.35 44.595 ;
        RECT 95.09 43.575 95.35 43.835 ;
        RECT 95.09 42.815 95.35 43.075 ;
        RECT 95.09 42.055 95.35 42.315 ;
        RECT 95.09 41.295 95.35 41.555 ;
        RECT 95.09 40.535 95.35 40.795 ;
        RECT 95.09 39.775 95.35 40.035 ;
        RECT 95.09 39.015 95.35 39.275 ;
        RECT 95.09 38.255 95.35 38.515 ;
        RECT 95.09 37.495 95.35 37.755 ;
        RECT 95.09 36.735 95.35 36.995 ;
        RECT 54.81 43.575 55.07 43.835 ;
        RECT 54.81 42.815 55.07 43.075 ;
        RECT 54.81 42.055 55.07 42.315 ;
        RECT 54.81 41.295 55.07 41.555 ;
        RECT 54.81 40.535 55.07 40.795 ;
        RECT 54.81 39.775 55.07 40.035 ;
        RECT 54.81 39.015 55.07 39.275 ;
        RECT 54.81 38.255 55.07 38.515 ;
        RECT 54.81 37.495 55.07 37.755 ;
        RECT 54.81 36.735 55.07 36.995 ;
        RECT 55.57 58.775 55.83 59.035 ;
        RECT 55.57 58.015 55.83 58.275 ;
        RECT 55.57 57.255 55.83 57.515 ;
        RECT 55.57 56.495 55.83 56.755 ;
        RECT 55.57 55.735 55.83 55.995 ;
        RECT 55.57 54.975 55.83 55.235 ;
        RECT 55.57 54.215 55.83 54.475 ;
        RECT 55.57 53.455 55.83 53.715 ;
        RECT 55.57 52.695 55.83 52.955 ;
        RECT 55.57 51.935 55.83 52.195 ;
        RECT 55.57 51.175 55.83 51.435 ;
        RECT 55.57 50.415 55.83 50.675 ;
        RECT 55.57 49.655 55.83 49.915 ;
        RECT 55.57 48.895 55.83 49.155 ;
        RECT 55.57 48.135 55.83 48.395 ;
        RECT 55.57 47.375 55.83 47.635 ;
        RECT 55.57 46.615 55.83 46.875 ;
        RECT 55.57 45.855 55.83 46.115 ;
        RECT 55.57 45.095 55.83 45.355 ;
        RECT 55.57 44.335 55.83 44.595 ;
        RECT 55.57 43.575 55.83 43.835 ;
        RECT 55.57 42.815 55.83 43.075 ;
        RECT 55.57 42.055 55.83 42.315 ;
        RECT 55.57 41.295 55.83 41.555 ;
        RECT 55.57 40.535 55.83 40.795 ;
        RECT 55.57 39.775 55.83 40.035 ;
        RECT 55.57 39.015 55.83 39.275 ;
        RECT 55.57 38.255 55.83 38.515 ;
        RECT 55.57 37.495 55.83 37.755 ;
        RECT 55.57 36.735 55.83 36.995 ;
        RECT 56.33 58.775 56.59 59.035 ;
        RECT 56.33 58.015 56.59 58.275 ;
        RECT 56.33 57.255 56.59 57.515 ;
        RECT 56.33 56.495 56.59 56.755 ;
        RECT 56.33 55.735 56.59 55.995 ;
        RECT 56.33 54.975 56.59 55.235 ;
        RECT 56.33 54.215 56.59 54.475 ;
        RECT 56.33 53.455 56.59 53.715 ;
        RECT 56.33 52.695 56.59 52.955 ;
        RECT 56.33 51.935 56.59 52.195 ;
        RECT 56.33 51.175 56.59 51.435 ;
        RECT 56.33 50.415 56.59 50.675 ;
        RECT 56.33 49.655 56.59 49.915 ;
        RECT 56.33 48.895 56.59 49.155 ;
        RECT 56.33 48.135 56.59 48.395 ;
        RECT 56.33 47.375 56.59 47.635 ;
        RECT 56.33 46.615 56.59 46.875 ;
        RECT 56.33 45.855 56.59 46.115 ;
        RECT 56.33 45.095 56.59 45.355 ;
        RECT 56.33 44.335 56.59 44.595 ;
        RECT 56.33 43.575 56.59 43.835 ;
        RECT 56.33 42.815 56.59 43.075 ;
        RECT 56.33 42.055 56.59 42.315 ;
        RECT 56.33 41.295 56.59 41.555 ;
        RECT 56.33 40.535 56.59 40.795 ;
        RECT 56.33 39.775 56.59 40.035 ;
        RECT 56.33 39.015 56.59 39.275 ;
        RECT 56.33 38.255 56.59 38.515 ;
        RECT 56.33 37.495 56.59 37.755 ;
        RECT 56.33 36.735 56.59 36.995 ;
        RECT 57.09 58.775 57.35 59.035 ;
        RECT 57.09 58.015 57.35 58.275 ;
        RECT 57.09 57.255 57.35 57.515 ;
        RECT 57.09 56.495 57.35 56.755 ;
        RECT 57.09 55.735 57.35 55.995 ;
        RECT 57.09 54.975 57.35 55.235 ;
        RECT 57.09 54.215 57.35 54.475 ;
        RECT 57.09 53.455 57.35 53.715 ;
        RECT 57.09 52.695 57.35 52.955 ;
        RECT 57.09 51.935 57.35 52.195 ;
        RECT 57.09 51.175 57.35 51.435 ;
        RECT 57.09 50.415 57.35 50.675 ;
        RECT 57.09 49.655 57.35 49.915 ;
        RECT 57.09 48.895 57.35 49.155 ;
        RECT 57.09 48.135 57.35 48.395 ;
        RECT 57.09 47.375 57.35 47.635 ;
        RECT 57.09 46.615 57.35 46.875 ;
        RECT 57.09 45.855 57.35 46.115 ;
        RECT 57.09 45.095 57.35 45.355 ;
        RECT 57.09 44.335 57.35 44.595 ;
        RECT 57.09 43.575 57.35 43.835 ;
        RECT 57.09 42.815 57.35 43.075 ;
        RECT 57.09 42.055 57.35 42.315 ;
        RECT 57.09 41.295 57.35 41.555 ;
        RECT 57.09 40.535 57.35 40.795 ;
        RECT 57.09 39.775 57.35 40.035 ;
        RECT 57.09 39.015 57.35 39.275 ;
        RECT 57.09 38.255 57.35 38.515 ;
        RECT 57.09 37.495 57.35 37.755 ;
        RECT 57.09 36.735 57.35 36.995 ;
        RECT 57.85 58.775 58.11 59.035 ;
        RECT 57.85 58.015 58.11 58.275 ;
        RECT 57.85 57.255 58.11 57.515 ;
        RECT 57.85 56.495 58.11 56.755 ;
        RECT 57.85 55.735 58.11 55.995 ;
        RECT 57.85 54.975 58.11 55.235 ;
        RECT 57.85 54.215 58.11 54.475 ;
        RECT 57.85 53.455 58.11 53.715 ;
        RECT 57.85 52.695 58.11 52.955 ;
        RECT 57.85 51.935 58.11 52.195 ;
        RECT 57.85 51.175 58.11 51.435 ;
        RECT 57.85 50.415 58.11 50.675 ;
        RECT 57.85 49.655 58.11 49.915 ;
        RECT 57.85 48.895 58.11 49.155 ;
        RECT 57.85 48.135 58.11 48.395 ;
        RECT 57.85 47.375 58.11 47.635 ;
        RECT 57.85 46.615 58.11 46.875 ;
        RECT 57.85 45.855 58.11 46.115 ;
        RECT 57.85 45.095 58.11 45.355 ;
        RECT 57.85 44.335 58.11 44.595 ;
        RECT 57.85 43.575 58.11 43.835 ;
        RECT 57.85 42.815 58.11 43.075 ;
        RECT 57.85 42.055 58.11 42.315 ;
        RECT 57.85 41.295 58.11 41.555 ;
        RECT 57.85 40.535 58.11 40.795 ;
        RECT 57.85 39.775 58.11 40.035 ;
        RECT 57.85 39.015 58.11 39.275 ;
        RECT 57.85 38.255 58.11 38.515 ;
        RECT 57.85 37.495 58.11 37.755 ;
        RECT 57.85 36.735 58.11 36.995 ;
        RECT 58.61 58.775 58.87 59.035 ;
        RECT 58.61 58.015 58.87 58.275 ;
        RECT 58.61 57.255 58.87 57.515 ;
        RECT 58.61 56.495 58.87 56.755 ;
        RECT 58.61 55.735 58.87 55.995 ;
        RECT 58.61 54.975 58.87 55.235 ;
        RECT 58.61 54.215 58.87 54.475 ;
        RECT 58.61 53.455 58.87 53.715 ;
        RECT 58.61 52.695 58.87 52.955 ;
        RECT 58.61 51.935 58.87 52.195 ;
        RECT 58.61 51.175 58.87 51.435 ;
        RECT 58.61 50.415 58.87 50.675 ;
        RECT 58.61 49.655 58.87 49.915 ;
        RECT 58.61 48.895 58.87 49.155 ;
        RECT 58.61 48.135 58.87 48.395 ;
        RECT 58.61 47.375 58.87 47.635 ;
        RECT 58.61 46.615 58.87 46.875 ;
        RECT 58.61 45.855 58.87 46.115 ;
        RECT 58.61 45.095 58.87 45.355 ;
        RECT 58.61 44.335 58.87 44.595 ;
        RECT 58.61 43.575 58.87 43.835 ;
        RECT 58.61 42.815 58.87 43.075 ;
        RECT 58.61 42.055 58.87 42.315 ;
        RECT 58.61 41.295 58.87 41.555 ;
        RECT 58.61 40.535 58.87 40.795 ;
        RECT 58.61 39.775 58.87 40.035 ;
        RECT 58.61 39.015 58.87 39.275 ;
        RECT 58.61 38.255 58.87 38.515 ;
        RECT 58.61 37.495 58.87 37.755 ;
        RECT 58.61 36.735 58.87 36.995 ;
        RECT 59.37 58.775 59.63 59.035 ;
        RECT 59.37 58.015 59.63 58.275 ;
        RECT 59.37 57.255 59.63 57.515 ;
        RECT 59.37 56.495 59.63 56.755 ;
        RECT 59.37 55.735 59.63 55.995 ;
        RECT 59.37 54.975 59.63 55.235 ;
        RECT 59.37 54.215 59.63 54.475 ;
        RECT 59.37 53.455 59.63 53.715 ;
        RECT 59.37 52.695 59.63 52.955 ;
        RECT 59.37 51.935 59.63 52.195 ;
        RECT 59.37 51.175 59.63 51.435 ;
        RECT 59.37 50.415 59.63 50.675 ;
        RECT 59.37 49.655 59.63 49.915 ;
        RECT 59.37 48.895 59.63 49.155 ;
        RECT 59.37 48.135 59.63 48.395 ;
        RECT 59.37 47.375 59.63 47.635 ;
        RECT 59.37 46.615 59.63 46.875 ;
        RECT 59.37 45.855 59.63 46.115 ;
        RECT 59.37 45.095 59.63 45.355 ;
        RECT 59.37 44.335 59.63 44.595 ;
        RECT 59.37 43.575 59.63 43.835 ;
        RECT 59.37 42.815 59.63 43.075 ;
        RECT 59.37 42.055 59.63 42.315 ;
        RECT 59.37 41.295 59.63 41.555 ;
        RECT 59.37 40.535 59.63 40.795 ;
        RECT 59.37 39.775 59.63 40.035 ;
        RECT 59.37 39.015 59.63 39.275 ;
        RECT 59.37 38.255 59.63 38.515 ;
        RECT 59.37 37.495 59.63 37.755 ;
        RECT 59.37 36.735 59.63 36.995 ;
        RECT 60.13 58.775 60.39 59.035 ;
        RECT 60.13 58.015 60.39 58.275 ;
        RECT 60.13 57.255 60.39 57.515 ;
        RECT 60.13 56.495 60.39 56.755 ;
        RECT 60.13 55.735 60.39 55.995 ;
        RECT 60.13 54.975 60.39 55.235 ;
        RECT 60.13 54.215 60.39 54.475 ;
        RECT 60.13 53.455 60.39 53.715 ;
        RECT 60.13 52.695 60.39 52.955 ;
        RECT 60.13 51.935 60.39 52.195 ;
        RECT 60.13 51.175 60.39 51.435 ;
        RECT 60.13 50.415 60.39 50.675 ;
        RECT 60.13 49.655 60.39 49.915 ;
        RECT 60.13 48.895 60.39 49.155 ;
        RECT 60.13 48.135 60.39 48.395 ;
        RECT 60.13 47.375 60.39 47.635 ;
        RECT 60.13 46.615 60.39 46.875 ;
        RECT 60.13 45.855 60.39 46.115 ;
        RECT 60.13 45.095 60.39 45.355 ;
        RECT 60.13 44.335 60.39 44.595 ;
        RECT 60.13 43.575 60.39 43.835 ;
        RECT 60.13 42.815 60.39 43.075 ;
        RECT 60.13 42.055 60.39 42.315 ;
        RECT 60.13 41.295 60.39 41.555 ;
        RECT 60.13 40.535 60.39 40.795 ;
        RECT 60.13 39.775 60.39 40.035 ;
        RECT 60.13 39.015 60.39 39.275 ;
        RECT 60.13 38.255 60.39 38.515 ;
        RECT 60.13 37.495 60.39 37.755 ;
        RECT 60.13 36.735 60.39 36.995 ;
        RECT 60.89 58.775 61.15 59.035 ;
        RECT 60.89 58.015 61.15 58.275 ;
        RECT 60.89 57.255 61.15 57.515 ;
        RECT 60.89 56.495 61.15 56.755 ;
        RECT 60.89 55.735 61.15 55.995 ;
        RECT 60.89 54.975 61.15 55.235 ;
        RECT 60.89 54.215 61.15 54.475 ;
        RECT 60.89 53.455 61.15 53.715 ;
        RECT 60.89 52.695 61.15 52.955 ;
        RECT 60.89 51.935 61.15 52.195 ;
        RECT 60.89 51.175 61.15 51.435 ;
        RECT 60.89 50.415 61.15 50.675 ;
        RECT 60.89 49.655 61.15 49.915 ;
        RECT 60.89 48.895 61.15 49.155 ;
        RECT 60.89 48.135 61.15 48.395 ;
        RECT 60.89 47.375 61.15 47.635 ;
        RECT 60.89 46.615 61.15 46.875 ;
        RECT 60.89 45.855 61.15 46.115 ;
        RECT 60.89 45.095 61.15 45.355 ;
        RECT 60.89 44.335 61.15 44.595 ;
        RECT 60.89 43.575 61.15 43.835 ;
        RECT 60.89 42.815 61.15 43.075 ;
        RECT 60.89 42.055 61.15 42.315 ;
        RECT 60.89 41.295 61.15 41.555 ;
        RECT 60.89 40.535 61.15 40.795 ;
        RECT 60.89 39.775 61.15 40.035 ;
        RECT 60.89 39.015 61.15 39.275 ;
        RECT 60.89 38.255 61.15 38.515 ;
        RECT 60.89 37.495 61.15 37.755 ;
        RECT 60.89 36.735 61.15 36.995 ;
        RECT 61.65 58.775 61.91 59.035 ;
        RECT 61.65 58.015 61.91 58.275 ;
        RECT 61.65 57.255 61.91 57.515 ;
        RECT 61.65 56.495 61.91 56.755 ;
        RECT 61.65 55.735 61.91 55.995 ;
        RECT 61.65 54.975 61.91 55.235 ;
        RECT 61.65 54.215 61.91 54.475 ;
        RECT 61.65 53.455 61.91 53.715 ;
        RECT 61.65 52.695 61.91 52.955 ;
        RECT 61.65 51.935 61.91 52.195 ;
        RECT 61.65 51.175 61.91 51.435 ;
        RECT 61.65 50.415 61.91 50.675 ;
        RECT 61.65 49.655 61.91 49.915 ;
        RECT 61.65 48.895 61.91 49.155 ;
        RECT 61.65 48.135 61.91 48.395 ;
        RECT 61.65 47.375 61.91 47.635 ;
        RECT 61.65 46.615 61.91 46.875 ;
        RECT 61.65 45.855 61.91 46.115 ;
        RECT 61.65 45.095 61.91 45.355 ;
        RECT 61.65 44.335 61.91 44.595 ;
        RECT 61.65 43.575 61.91 43.835 ;
        RECT 61.65 42.815 61.91 43.075 ;
        RECT 61.65 42.055 61.91 42.315 ;
        RECT 61.65 41.295 61.91 41.555 ;
        RECT 61.65 40.535 61.91 40.795 ;
        RECT 61.65 39.775 61.91 40.035 ;
        RECT 61.65 39.015 61.91 39.275 ;
        RECT 61.65 38.255 61.91 38.515 ;
        RECT 61.65 37.495 61.91 37.755 ;
        RECT 61.65 36.735 61.91 36.995 ;
        RECT 62.41 58.775 62.67 59.035 ;
        RECT 62.41 58.015 62.67 58.275 ;
        RECT 62.41 57.255 62.67 57.515 ;
        RECT 62.41 56.495 62.67 56.755 ;
        RECT 62.41 55.735 62.67 55.995 ;
        RECT 62.41 54.975 62.67 55.235 ;
        RECT 62.41 54.215 62.67 54.475 ;
        RECT 62.41 53.455 62.67 53.715 ;
        RECT 62.41 52.695 62.67 52.955 ;
        RECT 62.41 51.935 62.67 52.195 ;
        RECT 62.41 51.175 62.67 51.435 ;
        RECT 62.41 50.415 62.67 50.675 ;
        RECT 62.41 49.655 62.67 49.915 ;
        RECT 62.41 48.895 62.67 49.155 ;
        RECT 62.41 48.135 62.67 48.395 ;
        RECT 62.41 47.375 62.67 47.635 ;
        RECT 62.41 46.615 62.67 46.875 ;
        RECT 62.41 45.855 62.67 46.115 ;
        RECT 62.41 45.095 62.67 45.355 ;
        RECT 62.41 44.335 62.67 44.595 ;
        RECT 62.41 43.575 62.67 43.835 ;
        RECT 62.41 42.815 62.67 43.075 ;
        RECT 62.41 42.055 62.67 42.315 ;
        RECT 62.41 41.295 62.67 41.555 ;
        RECT 62.41 40.535 62.67 40.795 ;
        RECT 62.41 39.775 62.67 40.035 ;
        RECT 62.41 39.015 62.67 39.275 ;
        RECT 62.41 38.255 62.67 38.515 ;
        RECT 62.41 37.495 62.67 37.755 ;
        RECT 62.41 36.735 62.67 36.995 ;
        RECT 63.17 58.775 63.43 59.035 ;
        RECT 63.17 58.015 63.43 58.275 ;
        RECT 63.17 57.255 63.43 57.515 ;
        RECT 63.17 56.495 63.43 56.755 ;
        RECT 63.17 55.735 63.43 55.995 ;
        RECT 63.17 54.975 63.43 55.235 ;
        RECT 63.17 54.215 63.43 54.475 ;
        RECT 63.17 53.455 63.43 53.715 ;
        RECT 63.17 52.695 63.43 52.955 ;
        RECT 63.17 51.935 63.43 52.195 ;
        RECT 63.17 51.175 63.43 51.435 ;
        RECT 63.17 50.415 63.43 50.675 ;
        RECT 63.17 49.655 63.43 49.915 ;
        RECT 63.17 48.895 63.43 49.155 ;
        RECT 63.17 48.135 63.43 48.395 ;
        RECT 63.17 47.375 63.43 47.635 ;
        RECT 63.17 46.615 63.43 46.875 ;
        RECT 63.17 45.855 63.43 46.115 ;
        RECT 63.17 45.095 63.43 45.355 ;
        RECT 63.17 44.335 63.43 44.595 ;
        RECT 63.17 43.575 63.43 43.835 ;
        RECT 63.17 42.815 63.43 43.075 ;
        RECT 63.17 42.055 63.43 42.315 ;
        RECT 63.17 41.295 63.43 41.555 ;
        RECT 63.17 40.535 63.43 40.795 ;
        RECT 63.17 39.775 63.43 40.035 ;
        RECT 63.17 39.015 63.43 39.275 ;
        RECT 63.17 38.255 63.43 38.515 ;
        RECT 63.17 37.495 63.43 37.755 ;
        RECT 63.17 36.735 63.43 36.995 ;
        RECT 63.93 58.775 64.19 59.035 ;
        RECT 63.93 58.015 64.19 58.275 ;
        RECT 63.93 57.255 64.19 57.515 ;
        RECT 63.93 56.495 64.19 56.755 ;
        RECT 63.93 55.735 64.19 55.995 ;
        RECT 63.93 54.975 64.19 55.235 ;
        RECT 63.93 54.215 64.19 54.475 ;
        RECT 63.93 53.455 64.19 53.715 ;
        RECT 63.93 52.695 64.19 52.955 ;
        RECT 63.93 51.935 64.19 52.195 ;
        RECT 63.93 51.175 64.19 51.435 ;
        RECT 63.93 50.415 64.19 50.675 ;
        RECT 63.93 49.655 64.19 49.915 ;
        RECT 63.93 48.895 64.19 49.155 ;
        RECT 63.93 48.135 64.19 48.395 ;
        RECT 63.93 47.375 64.19 47.635 ;
        RECT 63.93 46.615 64.19 46.875 ;
        RECT 63.93 45.855 64.19 46.115 ;
        RECT 63.93 45.095 64.19 45.355 ;
        RECT 63.93 44.335 64.19 44.595 ;
        RECT 63.93 43.575 64.19 43.835 ;
        RECT 63.93 42.815 64.19 43.075 ;
        RECT 63.93 42.055 64.19 42.315 ;
        RECT 63.93 41.295 64.19 41.555 ;
        RECT 63.93 40.535 64.19 40.795 ;
        RECT 63.93 39.775 64.19 40.035 ;
        RECT 63.93 39.015 64.19 39.275 ;
        RECT 63.93 38.255 64.19 38.515 ;
        RECT 63.93 37.495 64.19 37.755 ;
        RECT 63.93 36.735 64.19 36.995 ;
        RECT 64.69 58.775 64.95 59.035 ;
        RECT 64.69 58.015 64.95 58.275 ;
        RECT 64.69 57.255 64.95 57.515 ;
        RECT 64.69 56.495 64.95 56.755 ;
        RECT 64.69 55.735 64.95 55.995 ;
        RECT 64.69 54.975 64.95 55.235 ;
        RECT 64.69 54.215 64.95 54.475 ;
        RECT 64.69 53.455 64.95 53.715 ;
        RECT 64.69 52.695 64.95 52.955 ;
        RECT 64.69 51.935 64.95 52.195 ;
        RECT 64.69 51.175 64.95 51.435 ;
        RECT 64.69 50.415 64.95 50.675 ;
        RECT 64.69 49.655 64.95 49.915 ;
        RECT 64.69 48.895 64.95 49.155 ;
        RECT 64.69 48.135 64.95 48.395 ;
        RECT 64.69 47.375 64.95 47.635 ;
        RECT 64.69 46.615 64.95 46.875 ;
        RECT 64.69 45.855 64.95 46.115 ;
        RECT 64.69 45.095 64.95 45.355 ;
        RECT 64.69 44.335 64.95 44.595 ;
        RECT 64.69 43.575 64.95 43.835 ;
        RECT 64.69 42.815 64.95 43.075 ;
        RECT 64.69 42.055 64.95 42.315 ;
        RECT 64.69 41.295 64.95 41.555 ;
        RECT 64.69 40.535 64.95 40.795 ;
        RECT 64.69 39.775 64.95 40.035 ;
        RECT 64.69 39.015 64.95 39.275 ;
        RECT 64.69 38.255 64.95 38.515 ;
        RECT 64.69 37.495 64.95 37.755 ;
        RECT 64.69 36.735 64.95 36.995 ;
        RECT 65.45 58.775 65.71 59.035 ;
        RECT 65.45 58.015 65.71 58.275 ;
        RECT 65.45 57.255 65.71 57.515 ;
        RECT 65.45 56.495 65.71 56.755 ;
        RECT 65.45 55.735 65.71 55.995 ;
        RECT 65.45 54.975 65.71 55.235 ;
        RECT 65.45 54.215 65.71 54.475 ;
        RECT 65.45 53.455 65.71 53.715 ;
        RECT 65.45 52.695 65.71 52.955 ;
        RECT 65.45 51.935 65.71 52.195 ;
        RECT 65.45 51.175 65.71 51.435 ;
        RECT 65.45 50.415 65.71 50.675 ;
        RECT 65.45 49.655 65.71 49.915 ;
        RECT 65.45 48.895 65.71 49.155 ;
        RECT 65.45 48.135 65.71 48.395 ;
        RECT 65.45 47.375 65.71 47.635 ;
        RECT 65.45 46.615 65.71 46.875 ;
        RECT 65.45 45.855 65.71 46.115 ;
        RECT 65.45 45.095 65.71 45.355 ;
        RECT 65.45 44.335 65.71 44.595 ;
        RECT 65.45 43.575 65.71 43.835 ;
        RECT 65.45 42.815 65.71 43.075 ;
        RECT 65.45 42.055 65.71 42.315 ;
        RECT 65.45 41.295 65.71 41.555 ;
        RECT 65.45 40.535 65.71 40.795 ;
        RECT 65.45 39.775 65.71 40.035 ;
        RECT 65.45 39.015 65.71 39.275 ;
        RECT 65.45 38.255 65.71 38.515 ;
        RECT 65.45 37.495 65.71 37.755 ;
        RECT 65.45 36.735 65.71 36.995 ;
        RECT 66.21 58.775 66.47 59.035 ;
        RECT 66.21 58.015 66.47 58.275 ;
        RECT 66.21 57.255 66.47 57.515 ;
        RECT 66.21 56.495 66.47 56.755 ;
        RECT 66.21 55.735 66.47 55.995 ;
        RECT 66.21 54.975 66.47 55.235 ;
        RECT 66.21 54.215 66.47 54.475 ;
        RECT 66.21 53.455 66.47 53.715 ;
        RECT 66.21 52.695 66.47 52.955 ;
        RECT 66.21 51.935 66.47 52.195 ;
        RECT 66.21 51.175 66.47 51.435 ;
        RECT 66.21 50.415 66.47 50.675 ;
        RECT 66.21 49.655 66.47 49.915 ;
        RECT 66.21 48.895 66.47 49.155 ;
        RECT 66.21 48.135 66.47 48.395 ;
        RECT 66.21 47.375 66.47 47.635 ;
        RECT 66.21 46.615 66.47 46.875 ;
        RECT 66.21 45.855 66.47 46.115 ;
        RECT 66.21 45.095 66.47 45.355 ;
        RECT 66.21 44.335 66.47 44.595 ;
        RECT 66.21 43.575 66.47 43.835 ;
        RECT 66.21 42.815 66.47 43.075 ;
        RECT 66.21 42.055 66.47 42.315 ;
        RECT 66.21 41.295 66.47 41.555 ;
        RECT 66.21 40.535 66.47 40.795 ;
        RECT 66.21 39.775 66.47 40.035 ;
        RECT 66.21 39.015 66.47 39.275 ;
        RECT 66.21 38.255 66.47 38.515 ;
        RECT 66.21 37.495 66.47 37.755 ;
        RECT 66.21 36.735 66.47 36.995 ;
        RECT 66.97 58.775 67.23 59.035 ;
        RECT 66.97 58.015 67.23 58.275 ;
        RECT 66.97 57.255 67.23 57.515 ;
        RECT 66.97 56.495 67.23 56.755 ;
        RECT 66.97 55.735 67.23 55.995 ;
        RECT 66.97 54.975 67.23 55.235 ;
        RECT 66.97 54.215 67.23 54.475 ;
        RECT 66.97 53.455 67.23 53.715 ;
        RECT 66.97 52.695 67.23 52.955 ;
        RECT 66.97 51.935 67.23 52.195 ;
        RECT 66.97 51.175 67.23 51.435 ;
        RECT 66.97 50.415 67.23 50.675 ;
        RECT 66.97 49.655 67.23 49.915 ;
        RECT 66.97 48.895 67.23 49.155 ;
        RECT 66.97 48.135 67.23 48.395 ;
        RECT 66.97 47.375 67.23 47.635 ;
        RECT 66.97 46.615 67.23 46.875 ;
        RECT 66.97 45.855 67.23 46.115 ;
        RECT 66.97 45.095 67.23 45.355 ;
        RECT 66.97 44.335 67.23 44.595 ;
        RECT 66.97 43.575 67.23 43.835 ;
        RECT 66.97 42.815 67.23 43.075 ;
        RECT 66.97 42.055 67.23 42.315 ;
        RECT 66.97 41.295 67.23 41.555 ;
        RECT 66.97 40.535 67.23 40.795 ;
        RECT 66.97 39.775 67.23 40.035 ;
        RECT 66.97 39.015 67.23 39.275 ;
        RECT 66.97 38.255 67.23 38.515 ;
        RECT 66.97 37.495 67.23 37.755 ;
        RECT 66.97 36.735 67.23 36.995 ;
        RECT 67.73 58.775 67.99 59.035 ;
        RECT 67.73 58.015 67.99 58.275 ;
        RECT 67.73 57.255 67.99 57.515 ;
        RECT 67.73 56.495 67.99 56.755 ;
        RECT 67.73 55.735 67.99 55.995 ;
        RECT 67.73 54.975 67.99 55.235 ;
        RECT 67.73 54.215 67.99 54.475 ;
        RECT 67.73 53.455 67.99 53.715 ;
        RECT 67.73 52.695 67.99 52.955 ;
        RECT 67.73 51.935 67.99 52.195 ;
        RECT 67.73 51.175 67.99 51.435 ;
        RECT 67.73 50.415 67.99 50.675 ;
        RECT 67.73 49.655 67.99 49.915 ;
        RECT 67.73 48.895 67.99 49.155 ;
        RECT 67.73 48.135 67.99 48.395 ;
        RECT 67.73 47.375 67.99 47.635 ;
        RECT 67.73 46.615 67.99 46.875 ;
        RECT 67.73 45.855 67.99 46.115 ;
        RECT 67.73 45.095 67.99 45.355 ;
        RECT 67.73 44.335 67.99 44.595 ;
        RECT 67.73 43.575 67.99 43.835 ;
        RECT 67.73 42.815 67.99 43.075 ;
        RECT 67.73 42.055 67.99 42.315 ;
        RECT 67.73 41.295 67.99 41.555 ;
        RECT 67.73 40.535 67.99 40.795 ;
        RECT 67.73 39.775 67.99 40.035 ;
        RECT 67.73 39.015 67.99 39.275 ;
        RECT 67.73 38.255 67.99 38.515 ;
        RECT 67.73 37.495 67.99 37.755 ;
        RECT 67.73 36.735 67.99 36.995 ;
        RECT 68.49 58.775 68.75 59.035 ;
        RECT 68.49 58.015 68.75 58.275 ;
        RECT 68.49 57.255 68.75 57.515 ;
        RECT 68.49 56.495 68.75 56.755 ;
        RECT 68.49 55.735 68.75 55.995 ;
        RECT 68.49 54.975 68.75 55.235 ;
        RECT 68.49 54.215 68.75 54.475 ;
        RECT 68.49 53.455 68.75 53.715 ;
        RECT 68.49 52.695 68.75 52.955 ;
        RECT 68.49 51.935 68.75 52.195 ;
        RECT 68.49 51.175 68.75 51.435 ;
        RECT 68.49 50.415 68.75 50.675 ;
        RECT 68.49 49.655 68.75 49.915 ;
        RECT 68.49 48.895 68.75 49.155 ;
        RECT 68.49 48.135 68.75 48.395 ;
        RECT 68.49 47.375 68.75 47.635 ;
        RECT 68.49 46.615 68.75 46.875 ;
        RECT 68.49 45.855 68.75 46.115 ;
        RECT 68.49 45.095 68.75 45.355 ;
        RECT 68.49 44.335 68.75 44.595 ;
        RECT 68.49 43.575 68.75 43.835 ;
        RECT 68.49 42.815 68.75 43.075 ;
        RECT 68.49 42.055 68.75 42.315 ;
        RECT 68.49 41.295 68.75 41.555 ;
        RECT 68.49 40.535 68.75 40.795 ;
        RECT 68.49 39.775 68.75 40.035 ;
        RECT 68.49 39.015 68.75 39.275 ;
        RECT 68.49 38.255 68.75 38.515 ;
        RECT 68.49 37.495 68.75 37.755 ;
        RECT 68.49 36.735 68.75 36.995 ;
        RECT 69.25 58.775 69.51 59.035 ;
        RECT 69.25 58.015 69.51 58.275 ;
        RECT 69.25 57.255 69.51 57.515 ;
        RECT 69.25 56.495 69.51 56.755 ;
        RECT 69.25 55.735 69.51 55.995 ;
        RECT 69.25 54.975 69.51 55.235 ;
        RECT 69.25 54.215 69.51 54.475 ;
        RECT 69.25 53.455 69.51 53.715 ;
        RECT 69.25 52.695 69.51 52.955 ;
        RECT 69.25 51.935 69.51 52.195 ;
        RECT 69.25 51.175 69.51 51.435 ;
        RECT 69.25 50.415 69.51 50.675 ;
        RECT 69.25 49.655 69.51 49.915 ;
        RECT 69.25 48.895 69.51 49.155 ;
        RECT 69.25 48.135 69.51 48.395 ;
        RECT 69.25 47.375 69.51 47.635 ;
        RECT 69.25 46.615 69.51 46.875 ;
        RECT 69.25 45.855 69.51 46.115 ;
        RECT 69.25 45.095 69.51 45.355 ;
        RECT 69.25 44.335 69.51 44.595 ;
        RECT 69.25 43.575 69.51 43.835 ;
        RECT 69.25 42.815 69.51 43.075 ;
        RECT 69.25 42.055 69.51 42.315 ;
        RECT 69.25 41.295 69.51 41.555 ;
        RECT 69.25 40.535 69.51 40.795 ;
        RECT 69.25 39.775 69.51 40.035 ;
        RECT 69.25 39.015 69.51 39.275 ;
        RECT 69.25 38.255 69.51 38.515 ;
        RECT 69.25 37.495 69.51 37.755 ;
        RECT 69.25 36.735 69.51 36.995 ;
        RECT 70.01 58.775 70.27 59.035 ;
        RECT 70.01 58.015 70.27 58.275 ;
        RECT 70.01 57.255 70.27 57.515 ;
        RECT 70.01 56.495 70.27 56.755 ;
        RECT 70.01 55.735 70.27 55.995 ;
        RECT 70.01 54.975 70.27 55.235 ;
        RECT 70.01 54.215 70.27 54.475 ;
        RECT 70.01 53.455 70.27 53.715 ;
        RECT 70.01 52.695 70.27 52.955 ;
        RECT 70.01 51.935 70.27 52.195 ;
        RECT 70.01 51.175 70.27 51.435 ;
        RECT 70.01 50.415 70.27 50.675 ;
        RECT 70.01 49.655 70.27 49.915 ;
        RECT 70.01 48.895 70.27 49.155 ;
        RECT 70.01 48.135 70.27 48.395 ;
        RECT 70.01 47.375 70.27 47.635 ;
        RECT 70.01 46.615 70.27 46.875 ;
        RECT 70.01 45.855 70.27 46.115 ;
        RECT 70.01 45.095 70.27 45.355 ;
        RECT 70.01 44.335 70.27 44.595 ;
        RECT 70.01 43.575 70.27 43.835 ;
        RECT 70.01 42.815 70.27 43.075 ;
        RECT 70.01 42.055 70.27 42.315 ;
        RECT 70.01 41.295 70.27 41.555 ;
        RECT 70.01 40.535 70.27 40.795 ;
        RECT 70.01 39.775 70.27 40.035 ;
        RECT 70.01 39.015 70.27 39.275 ;
        RECT 70.01 38.255 70.27 38.515 ;
        RECT 70.01 37.495 70.27 37.755 ;
        RECT 70.01 36.735 70.27 36.995 ;
        RECT 70.77 58.775 71.03 59.035 ;
        RECT 70.77 58.015 71.03 58.275 ;
        RECT 70.77 57.255 71.03 57.515 ;
        RECT 70.77 56.495 71.03 56.755 ;
        RECT 70.77 55.735 71.03 55.995 ;
        RECT 70.77 54.975 71.03 55.235 ;
        RECT 70.77 54.215 71.03 54.475 ;
        RECT 70.77 53.455 71.03 53.715 ;
        RECT 70.77 52.695 71.03 52.955 ;
        RECT 70.77 51.935 71.03 52.195 ;
        RECT 70.77 51.175 71.03 51.435 ;
        RECT 70.77 50.415 71.03 50.675 ;
        RECT 70.77 49.655 71.03 49.915 ;
        RECT 70.77 48.895 71.03 49.155 ;
        RECT 70.77 48.135 71.03 48.395 ;
        RECT 70.77 47.375 71.03 47.635 ;
        RECT 70.77 46.615 71.03 46.875 ;
        RECT 70.77 45.855 71.03 46.115 ;
        RECT 70.77 45.095 71.03 45.355 ;
        RECT 70.77 44.335 71.03 44.595 ;
        RECT 70.77 43.575 71.03 43.835 ;
        RECT 70.77 42.815 71.03 43.075 ;
        RECT 70.77 42.055 71.03 42.315 ;
        RECT 70.77 41.295 71.03 41.555 ;
        RECT 70.77 40.535 71.03 40.795 ;
        RECT 70.77 39.775 71.03 40.035 ;
        RECT 70.77 39.015 71.03 39.275 ;
        RECT 70.77 38.255 71.03 38.515 ;
        RECT 70.77 37.495 71.03 37.755 ;
        RECT 70.77 36.735 71.03 36.995 ;
        RECT 71.53 58.775 71.79 59.035 ;
        RECT 71.53 58.015 71.79 58.275 ;
        RECT 71.53 57.255 71.79 57.515 ;
        RECT 71.53 56.495 71.79 56.755 ;
        RECT 71.53 55.735 71.79 55.995 ;
        RECT 71.53 54.975 71.79 55.235 ;
        RECT 71.53 54.215 71.79 54.475 ;
        RECT 71.53 53.455 71.79 53.715 ;
        RECT 71.53 52.695 71.79 52.955 ;
        RECT 71.53 51.935 71.79 52.195 ;
        RECT 71.53 51.175 71.79 51.435 ;
        RECT 71.53 50.415 71.79 50.675 ;
        RECT 71.53 49.655 71.79 49.915 ;
        RECT 71.53 48.895 71.79 49.155 ;
        RECT 71.53 48.135 71.79 48.395 ;
        RECT 71.53 47.375 71.79 47.635 ;
        RECT 71.53 46.615 71.79 46.875 ;
        RECT 71.53 45.855 71.79 46.115 ;
        RECT 71.53 45.095 71.79 45.355 ;
        RECT 71.53 44.335 71.79 44.595 ;
        RECT 71.53 43.575 71.79 43.835 ;
        RECT 71.53 42.815 71.79 43.075 ;
        RECT 71.53 42.055 71.79 42.315 ;
        RECT 71.53 41.295 71.79 41.555 ;
        RECT 71.53 40.535 71.79 40.795 ;
        RECT 71.53 39.775 71.79 40.035 ;
        RECT 71.53 39.015 71.79 39.275 ;
        RECT 71.53 38.255 71.79 38.515 ;
        RECT 71.53 37.495 71.79 37.755 ;
        RECT 71.53 36.735 71.79 36.995 ;
        RECT 72.29 58.775 72.55 59.035 ;
        RECT 72.29 58.015 72.55 58.275 ;
        RECT 72.29 57.255 72.55 57.515 ;
        RECT 72.29 56.495 72.55 56.755 ;
        RECT 72.29 55.735 72.55 55.995 ;
        RECT 72.29 54.975 72.55 55.235 ;
        RECT 72.29 54.215 72.55 54.475 ;
        RECT 72.29 53.455 72.55 53.715 ;
        RECT 72.29 52.695 72.55 52.955 ;
        RECT 72.29 51.935 72.55 52.195 ;
        RECT 72.29 51.175 72.55 51.435 ;
        RECT 72.29 50.415 72.55 50.675 ;
        RECT 72.29 49.655 72.55 49.915 ;
        RECT 72.29 48.895 72.55 49.155 ;
        RECT 72.29 48.135 72.55 48.395 ;
        RECT 72.29 47.375 72.55 47.635 ;
        RECT 72.29 46.615 72.55 46.875 ;
        RECT 72.29 45.855 72.55 46.115 ;
        RECT 72.29 45.095 72.55 45.355 ;
        RECT 72.29 44.335 72.55 44.595 ;
        RECT 72.29 43.575 72.55 43.835 ;
        RECT 72.29 42.815 72.55 43.075 ;
        RECT 72.29 42.055 72.55 42.315 ;
        RECT 72.29 41.295 72.55 41.555 ;
        RECT 72.29 40.535 72.55 40.795 ;
        RECT 72.29 39.775 72.55 40.035 ;
        RECT 72.29 39.015 72.55 39.275 ;
        RECT 72.29 38.255 72.55 38.515 ;
        RECT 72.29 37.495 72.55 37.755 ;
        RECT 72.29 36.735 72.55 36.995 ;
        RECT 73.05 58.775 73.31 59.035 ;
        RECT 73.05 58.015 73.31 58.275 ;
        RECT 73.05 57.255 73.31 57.515 ;
        RECT 73.05 56.495 73.31 56.755 ;
        RECT 73.05 55.735 73.31 55.995 ;
        RECT 73.05 54.975 73.31 55.235 ;
        RECT 73.05 54.215 73.31 54.475 ;
        RECT 73.05 53.455 73.31 53.715 ;
        RECT 73.05 52.695 73.31 52.955 ;
        RECT 73.05 51.935 73.31 52.195 ;
        RECT 73.05 51.175 73.31 51.435 ;
        RECT 73.05 50.415 73.31 50.675 ;
        RECT 73.05 49.655 73.31 49.915 ;
        RECT 73.05 48.895 73.31 49.155 ;
        RECT 73.05 48.135 73.31 48.395 ;
        RECT 73.05 47.375 73.31 47.635 ;
        RECT 73.05 46.615 73.31 46.875 ;
        RECT 73.05 45.855 73.31 46.115 ;
        RECT 73.05 45.095 73.31 45.355 ;
        RECT 73.05 44.335 73.31 44.595 ;
        RECT 73.05 43.575 73.31 43.835 ;
        RECT 73.05 42.815 73.31 43.075 ;
        RECT 73.05 42.055 73.31 42.315 ;
        RECT 73.05 41.295 73.31 41.555 ;
        RECT 73.05 40.535 73.31 40.795 ;
        RECT 73.05 39.775 73.31 40.035 ;
        RECT 73.05 39.015 73.31 39.275 ;
        RECT 73.05 38.255 73.31 38.515 ;
        RECT 73.05 37.495 73.31 37.755 ;
        RECT 73.05 36.735 73.31 36.995 ;
        RECT 73.81 58.775 74.07 59.035 ;
        RECT 73.81 58.015 74.07 58.275 ;
        RECT 73.81 57.255 74.07 57.515 ;
        RECT 73.81 56.495 74.07 56.755 ;
        RECT 73.81 55.735 74.07 55.995 ;
        RECT 73.81 54.975 74.07 55.235 ;
        RECT 73.81 54.215 74.07 54.475 ;
        RECT 73.81 53.455 74.07 53.715 ;
        RECT 73.81 52.695 74.07 52.955 ;
        RECT 73.81 51.935 74.07 52.195 ;
        RECT 73.81 51.175 74.07 51.435 ;
        RECT 73.81 50.415 74.07 50.675 ;
        RECT 73.81 49.655 74.07 49.915 ;
        RECT 73.81 48.895 74.07 49.155 ;
        RECT 73.81 48.135 74.07 48.395 ;
        RECT 73.81 47.375 74.07 47.635 ;
        RECT 73.81 46.615 74.07 46.875 ;
        RECT 73.81 45.855 74.07 46.115 ;
        RECT 73.81 45.095 74.07 45.355 ;
        RECT 73.81 44.335 74.07 44.595 ;
        RECT 73.81 43.575 74.07 43.835 ;
        RECT 73.81 42.815 74.07 43.075 ;
        RECT 73.81 42.055 74.07 42.315 ;
        RECT 73.81 41.295 74.07 41.555 ;
        RECT 73.81 40.535 74.07 40.795 ;
        RECT 73.81 39.775 74.07 40.035 ;
        RECT 73.81 39.015 74.07 39.275 ;
        RECT 73.81 38.255 74.07 38.515 ;
        RECT 73.81 37.495 74.07 37.755 ;
        RECT 73.81 36.735 74.07 36.995 ;
        RECT 74.57 58.775 74.83 59.035 ;
        RECT 74.57 58.015 74.83 58.275 ;
        RECT 74.57 57.255 74.83 57.515 ;
        RECT 74.57 56.495 74.83 56.755 ;
        RECT 74.57 55.735 74.83 55.995 ;
        RECT 74.57 54.975 74.83 55.235 ;
        RECT 74.57 54.215 74.83 54.475 ;
        RECT 74.57 53.455 74.83 53.715 ;
        RECT 74.57 52.695 74.83 52.955 ;
        RECT 74.57 51.935 74.83 52.195 ;
        RECT 74.57 51.175 74.83 51.435 ;
        RECT 74.57 50.415 74.83 50.675 ;
        RECT 74.57 49.655 74.83 49.915 ;
        RECT 74.57 48.895 74.83 49.155 ;
        RECT 74.57 48.135 74.83 48.395 ;
        RECT 74.57 47.375 74.83 47.635 ;
        RECT 74.57 46.615 74.83 46.875 ;
        RECT 74.57 45.855 74.83 46.115 ;
        RECT 74.57 45.095 74.83 45.355 ;
        RECT 74.57 44.335 74.83 44.595 ;
        RECT 74.57 43.575 74.83 43.835 ;
        RECT 74.57 42.815 74.83 43.075 ;
        RECT 74.57 42.055 74.83 42.315 ;
        RECT 74.57 41.295 74.83 41.555 ;
        RECT 74.57 40.535 74.83 40.795 ;
        RECT 74.57 39.775 74.83 40.035 ;
        RECT 74.57 39.015 74.83 39.275 ;
        RECT 74.57 38.255 74.83 38.515 ;
        RECT 74.57 37.495 74.83 37.755 ;
        RECT 74.57 36.735 74.83 36.995 ;
        RECT 75.33 58.775 75.59 59.035 ;
        RECT 75.33 58.015 75.59 58.275 ;
        RECT 75.33 57.255 75.59 57.515 ;
        RECT 75.33 56.495 75.59 56.755 ;
        RECT 75.33 55.735 75.59 55.995 ;
        RECT 75.33 54.975 75.59 55.235 ;
        RECT 75.33 54.215 75.59 54.475 ;
        RECT 75.33 53.455 75.59 53.715 ;
        RECT 75.33 52.695 75.59 52.955 ;
        RECT 75.33 51.935 75.59 52.195 ;
        RECT 75.33 51.175 75.59 51.435 ;
        RECT 75.33 50.415 75.59 50.675 ;
        RECT 75.33 49.655 75.59 49.915 ;
        RECT 75.33 48.895 75.59 49.155 ;
        RECT 75.33 48.135 75.59 48.395 ;
        RECT 75.33 47.375 75.59 47.635 ;
        RECT 75.33 46.615 75.59 46.875 ;
        RECT 75.33 45.855 75.59 46.115 ;
        RECT 75.33 45.095 75.59 45.355 ;
        RECT 75.33 44.335 75.59 44.595 ;
        RECT 75.33 43.575 75.59 43.835 ;
        RECT 75.33 42.815 75.59 43.075 ;
        RECT 75.33 42.055 75.59 42.315 ;
        RECT 75.33 41.295 75.59 41.555 ;
        RECT 75.33 40.535 75.59 40.795 ;
        RECT 75.33 39.775 75.59 40.035 ;
        RECT 75.33 39.015 75.59 39.275 ;
        RECT 75.33 38.255 75.59 38.515 ;
        RECT 75.33 37.495 75.59 37.755 ;
        RECT 75.33 36.735 75.59 36.995 ;
        RECT 76.09 58.775 76.35 59.035 ;
        RECT 76.09 58.015 76.35 58.275 ;
        RECT 76.09 57.255 76.35 57.515 ;
        RECT 76.09 56.495 76.35 56.755 ;
        RECT 76.09 55.735 76.35 55.995 ;
        RECT 76.09 54.975 76.35 55.235 ;
        RECT 76.09 54.215 76.35 54.475 ;
        RECT 76.09 53.455 76.35 53.715 ;
        RECT 76.09 52.695 76.35 52.955 ;
        RECT 76.09 51.935 76.35 52.195 ;
        RECT 76.09 51.175 76.35 51.435 ;
        RECT 76.09 50.415 76.35 50.675 ;
        RECT 76.09 49.655 76.35 49.915 ;
        RECT 76.09 48.895 76.35 49.155 ;
        RECT 76.09 48.135 76.35 48.395 ;
        RECT 76.09 47.375 76.35 47.635 ;
        RECT 76.09 46.615 76.35 46.875 ;
        RECT 76.09 45.855 76.35 46.115 ;
        RECT 76.09 45.095 76.35 45.355 ;
        RECT 76.09 44.335 76.35 44.595 ;
        RECT 76.09 43.575 76.35 43.835 ;
        RECT 76.09 42.815 76.35 43.075 ;
        RECT 76.09 42.055 76.35 42.315 ;
        RECT 76.09 41.295 76.35 41.555 ;
        RECT 76.09 40.535 76.35 40.795 ;
        RECT 76.09 39.775 76.35 40.035 ;
        RECT 76.09 39.015 76.35 39.275 ;
        RECT 76.09 38.255 76.35 38.515 ;
        RECT 76.09 37.495 76.35 37.755 ;
        RECT 76.09 36.735 76.35 36.995 ;
        RECT 76.85 58.775 77.11 59.035 ;
        RECT 76.85 58.015 77.11 58.275 ;
        RECT 76.85 57.255 77.11 57.515 ;
        RECT 76.85 56.495 77.11 56.755 ;
        RECT 76.85 55.735 77.11 55.995 ;
        RECT 76.85 54.975 77.11 55.235 ;
        RECT 76.85 54.215 77.11 54.475 ;
        RECT 76.85 53.455 77.11 53.715 ;
        RECT 76.85 52.695 77.11 52.955 ;
        RECT 76.85 51.935 77.11 52.195 ;
        RECT 76.85 51.175 77.11 51.435 ;
        RECT 76.85 50.415 77.11 50.675 ;
        RECT 76.85 49.655 77.11 49.915 ;
        RECT 76.85 48.895 77.11 49.155 ;
        RECT 76.85 48.135 77.11 48.395 ;
        RECT 76.85 47.375 77.11 47.635 ;
        RECT 76.85 46.615 77.11 46.875 ;
        RECT 76.85 45.855 77.11 46.115 ;
        RECT 76.85 45.095 77.11 45.355 ;
        RECT 76.85 44.335 77.11 44.595 ;
        RECT 76.85 43.575 77.11 43.835 ;
        RECT 76.85 42.815 77.11 43.075 ;
        RECT 76.85 42.055 77.11 42.315 ;
        RECT 76.85 41.295 77.11 41.555 ;
        RECT 76.85 40.535 77.11 40.795 ;
        RECT 76.85 39.775 77.11 40.035 ;
        RECT 76.85 39.015 77.11 39.275 ;
        RECT 76.85 38.255 77.11 38.515 ;
        RECT 76.85 37.495 77.11 37.755 ;
        RECT 76.85 36.735 77.11 36.995 ;
        RECT 77.61 58.775 77.87 59.035 ;
        RECT 77.61 58.015 77.87 58.275 ;
        RECT 77.61 57.255 77.87 57.515 ;
        RECT 77.61 56.495 77.87 56.755 ;
        RECT 77.61 55.735 77.87 55.995 ;
        RECT 77.61 54.975 77.87 55.235 ;
        RECT 77.61 54.215 77.87 54.475 ;
        RECT 77.61 53.455 77.87 53.715 ;
        RECT 77.61 52.695 77.87 52.955 ;
        RECT 77.61 51.935 77.87 52.195 ;
        RECT 77.61 51.175 77.87 51.435 ;
        RECT 77.61 50.415 77.87 50.675 ;
        RECT 77.61 49.655 77.87 49.915 ;
        RECT 77.61 48.895 77.87 49.155 ;
        RECT 77.61 48.135 77.87 48.395 ;
        RECT 77.61 47.375 77.87 47.635 ;
        RECT 77.61 46.615 77.87 46.875 ;
        RECT 77.61 45.855 77.87 46.115 ;
        RECT 77.61 45.095 77.87 45.355 ;
        RECT 77.61 44.335 77.87 44.595 ;
        RECT 77.61 43.575 77.87 43.835 ;
        RECT 77.61 42.815 77.87 43.075 ;
        RECT 77.61 42.055 77.87 42.315 ;
        RECT 77.61 41.295 77.87 41.555 ;
        RECT 77.61 40.535 77.87 40.795 ;
        RECT 77.61 39.775 77.87 40.035 ;
        RECT 77.61 39.015 77.87 39.275 ;
        RECT 77.61 38.255 77.87 38.515 ;
        RECT 77.61 37.495 77.87 37.755 ;
        RECT 77.61 36.735 77.87 36.995 ;
        RECT 78.37 58.775 78.63 59.035 ;
        RECT 78.37 58.015 78.63 58.275 ;
        RECT 78.37 57.255 78.63 57.515 ;
        RECT 78.37 56.495 78.63 56.755 ;
        RECT 78.37 55.735 78.63 55.995 ;
        RECT 78.37 54.975 78.63 55.235 ;
        RECT 78.37 54.215 78.63 54.475 ;
        RECT 78.37 53.455 78.63 53.715 ;
        RECT 78.37 52.695 78.63 52.955 ;
        RECT 78.37 51.935 78.63 52.195 ;
        RECT 78.37 51.175 78.63 51.435 ;
        RECT 78.37 50.415 78.63 50.675 ;
        RECT 78.37 49.655 78.63 49.915 ;
        RECT 78.37 48.895 78.63 49.155 ;
        RECT 78.37 48.135 78.63 48.395 ;
        RECT 78.37 47.375 78.63 47.635 ;
        RECT 78.37 46.615 78.63 46.875 ;
        RECT 78.37 45.855 78.63 46.115 ;
        RECT 78.37 45.095 78.63 45.355 ;
        RECT 78.37 44.335 78.63 44.595 ;
        RECT 78.37 43.575 78.63 43.835 ;
        RECT 78.37 42.815 78.63 43.075 ;
        RECT 78.37 42.055 78.63 42.315 ;
        RECT 78.37 41.295 78.63 41.555 ;
        RECT 78.37 40.535 78.63 40.795 ;
        RECT 78.37 39.775 78.63 40.035 ;
        RECT 78.37 39.015 78.63 39.275 ;
        RECT 78.37 38.255 78.63 38.515 ;
        RECT 78.37 37.495 78.63 37.755 ;
        RECT 78.37 36.735 78.63 36.995 ;
        RECT 79.13 58.775 79.39 59.035 ;
        RECT 79.13 58.015 79.39 58.275 ;
        RECT 79.13 57.255 79.39 57.515 ;
        RECT 79.13 56.495 79.39 56.755 ;
        RECT 79.13 55.735 79.39 55.995 ;
        RECT 79.13 54.975 79.39 55.235 ;
        RECT 79.13 54.215 79.39 54.475 ;
        RECT 79.13 53.455 79.39 53.715 ;
        RECT 79.13 52.695 79.39 52.955 ;
        RECT 79.13 51.935 79.39 52.195 ;
        RECT 79.13 51.175 79.39 51.435 ;
        RECT 79.13 50.415 79.39 50.675 ;
        RECT 79.13 49.655 79.39 49.915 ;
        RECT 79.13 48.895 79.39 49.155 ;
        RECT 79.13 48.135 79.39 48.395 ;
        RECT 79.13 47.375 79.39 47.635 ;
        RECT 79.13 46.615 79.39 46.875 ;
        RECT 79.13 45.855 79.39 46.115 ;
        RECT 79.13 45.095 79.39 45.355 ;
        RECT 79.13 44.335 79.39 44.595 ;
        RECT 79.13 43.575 79.39 43.835 ;
        RECT 79.13 42.815 79.39 43.075 ;
        RECT 79.13 42.055 79.39 42.315 ;
        RECT 79.13 41.295 79.39 41.555 ;
        RECT 79.13 40.535 79.39 40.795 ;
        RECT 79.13 39.775 79.39 40.035 ;
        RECT 79.13 39.015 79.39 39.275 ;
        RECT 79.13 38.255 79.39 38.515 ;
        RECT 79.13 37.495 79.39 37.755 ;
        RECT 79.13 36.735 79.39 36.995 ;
        RECT 79.89 58.775 80.15 59.035 ;
        RECT 79.89 58.015 80.15 58.275 ;
        RECT 79.89 57.255 80.15 57.515 ;
        RECT 79.89 56.495 80.15 56.755 ;
        RECT 79.89 55.735 80.15 55.995 ;
        RECT 79.89 54.975 80.15 55.235 ;
        RECT 79.89 54.215 80.15 54.475 ;
        RECT 79.89 53.455 80.15 53.715 ;
        RECT 79.89 52.695 80.15 52.955 ;
        RECT 79.89 51.935 80.15 52.195 ;
        RECT 79.89 51.175 80.15 51.435 ;
        RECT 79.89 50.415 80.15 50.675 ;
        RECT 79.89 49.655 80.15 49.915 ;
        RECT 79.89 48.895 80.15 49.155 ;
        RECT 79.89 48.135 80.15 48.395 ;
        RECT 79.89 47.375 80.15 47.635 ;
        RECT 79.89 46.615 80.15 46.875 ;
        RECT 79.89 45.855 80.15 46.115 ;
        RECT 79.89 45.095 80.15 45.355 ;
        RECT 79.89 44.335 80.15 44.595 ;
        RECT 79.89 43.575 80.15 43.835 ;
        RECT 79.89 42.815 80.15 43.075 ;
        RECT 79.89 42.055 80.15 42.315 ;
        RECT 79.89 41.295 80.15 41.555 ;
        RECT 79.89 40.535 80.15 40.795 ;
        RECT 79.89 39.775 80.15 40.035 ;
        RECT 79.89 39.015 80.15 39.275 ;
        RECT 79.89 38.255 80.15 38.515 ;
        RECT 79.89 37.495 80.15 37.755 ;
        RECT 79.89 36.735 80.15 36.995 ;
        RECT 29.73 51.175 29.99 51.435 ;
        RECT 29.73 50.415 29.99 50.675 ;
        RECT 29.73 49.655 29.99 49.915 ;
        RECT 29.73 48.895 29.99 49.155 ;
        RECT 29.73 48.135 29.99 48.395 ;
        RECT 29.73 47.375 29.99 47.635 ;
        RECT 29.73 46.615 29.99 46.875 ;
        RECT 29.73 45.855 29.99 46.115 ;
        RECT 29.73 45.095 29.99 45.355 ;
        RECT 29.73 44.335 29.99 44.595 ;
        RECT 29.73 43.575 29.99 43.835 ;
        RECT 29.73 42.815 29.99 43.075 ;
        RECT 29.73 42.055 29.99 42.315 ;
        RECT 29.73 41.295 29.99 41.555 ;
        RECT 29.73 40.535 29.99 40.795 ;
        RECT 29.73 39.775 29.99 40.035 ;
        RECT 29.73 39.015 29.99 39.275 ;
        RECT 29.73 38.255 29.99 38.515 ;
        RECT 29.73 37.495 29.99 37.755 ;
        RECT 29.73 36.735 29.99 36.995 ;
        RECT 30.49 58.775 30.75 59.035 ;
        RECT 30.49 58.015 30.75 58.275 ;
        RECT 30.49 57.255 30.75 57.515 ;
        RECT 30.49 56.495 30.75 56.755 ;
        RECT 30.49 55.735 30.75 55.995 ;
        RECT 30.49 54.975 30.75 55.235 ;
        RECT 30.49 54.215 30.75 54.475 ;
        RECT 30.49 53.455 30.75 53.715 ;
        RECT 30.49 52.695 30.75 52.955 ;
        RECT 30.49 51.935 30.75 52.195 ;
        RECT 30.49 51.175 30.75 51.435 ;
        RECT 30.49 50.415 30.75 50.675 ;
        RECT 30.49 49.655 30.75 49.915 ;
        RECT 30.49 48.895 30.75 49.155 ;
        RECT 30.49 48.135 30.75 48.395 ;
        RECT 30.49 47.375 30.75 47.635 ;
        RECT 30.49 46.615 30.75 46.875 ;
        RECT 30.49 45.855 30.75 46.115 ;
        RECT 30.49 45.095 30.75 45.355 ;
        RECT 30.49 44.335 30.75 44.595 ;
        RECT 30.49 43.575 30.75 43.835 ;
        RECT 30.49 42.815 30.75 43.075 ;
        RECT 30.49 42.055 30.75 42.315 ;
        RECT 30.49 41.295 30.75 41.555 ;
        RECT 30.49 40.535 30.75 40.795 ;
        RECT 30.49 39.775 30.75 40.035 ;
        RECT 30.49 39.015 30.75 39.275 ;
        RECT 30.49 38.255 30.75 38.515 ;
        RECT 30.49 37.495 30.75 37.755 ;
        RECT 30.49 36.735 30.75 36.995 ;
        RECT 31.25 58.775 31.51 59.035 ;
        RECT 31.25 58.015 31.51 58.275 ;
        RECT 31.25 57.255 31.51 57.515 ;
        RECT 31.25 56.495 31.51 56.755 ;
        RECT 31.25 55.735 31.51 55.995 ;
        RECT 31.25 54.975 31.51 55.235 ;
        RECT 31.25 54.215 31.51 54.475 ;
        RECT 31.25 53.455 31.51 53.715 ;
        RECT 31.25 52.695 31.51 52.955 ;
        RECT 31.25 51.935 31.51 52.195 ;
        RECT 31.25 51.175 31.51 51.435 ;
        RECT 31.25 50.415 31.51 50.675 ;
        RECT 31.25 49.655 31.51 49.915 ;
        RECT 31.25 48.895 31.51 49.155 ;
        RECT 31.25 48.135 31.51 48.395 ;
        RECT 31.25 47.375 31.51 47.635 ;
        RECT 31.25 46.615 31.51 46.875 ;
        RECT 31.25 45.855 31.51 46.115 ;
        RECT 31.25 45.095 31.51 45.355 ;
        RECT 31.25 44.335 31.51 44.595 ;
        RECT 31.25 43.575 31.51 43.835 ;
        RECT 31.25 42.815 31.51 43.075 ;
        RECT 31.25 42.055 31.51 42.315 ;
        RECT 31.25 41.295 31.51 41.555 ;
        RECT 31.25 40.535 31.51 40.795 ;
        RECT 31.25 39.775 31.51 40.035 ;
        RECT 31.25 39.015 31.51 39.275 ;
        RECT 31.25 38.255 31.51 38.515 ;
        RECT 31.25 37.495 31.51 37.755 ;
        RECT 31.25 36.735 31.51 36.995 ;
        RECT 32.01 58.775 32.27 59.035 ;
        RECT 32.01 58.015 32.27 58.275 ;
        RECT 32.01 57.255 32.27 57.515 ;
        RECT 32.01 56.495 32.27 56.755 ;
        RECT 32.01 55.735 32.27 55.995 ;
        RECT 32.01 54.975 32.27 55.235 ;
        RECT 32.01 54.215 32.27 54.475 ;
        RECT 32.01 53.455 32.27 53.715 ;
        RECT 32.01 52.695 32.27 52.955 ;
        RECT 32.01 51.935 32.27 52.195 ;
        RECT 32.01 51.175 32.27 51.435 ;
        RECT 32.01 50.415 32.27 50.675 ;
        RECT 32.01 49.655 32.27 49.915 ;
        RECT 32.01 48.895 32.27 49.155 ;
        RECT 32.01 48.135 32.27 48.395 ;
        RECT 32.01 47.375 32.27 47.635 ;
        RECT 32.01 46.615 32.27 46.875 ;
        RECT 32.01 45.855 32.27 46.115 ;
        RECT 32.01 45.095 32.27 45.355 ;
        RECT 32.01 44.335 32.27 44.595 ;
        RECT 32.01 43.575 32.27 43.835 ;
        RECT 32.01 42.815 32.27 43.075 ;
        RECT 32.01 42.055 32.27 42.315 ;
        RECT 32.01 41.295 32.27 41.555 ;
        RECT 32.01 40.535 32.27 40.795 ;
        RECT 32.01 39.775 32.27 40.035 ;
        RECT 32.01 39.015 32.27 39.275 ;
        RECT 32.01 38.255 32.27 38.515 ;
        RECT 32.01 37.495 32.27 37.755 ;
        RECT 32.01 36.735 32.27 36.995 ;
        RECT 32.77 58.775 33.03 59.035 ;
        RECT 32.77 58.015 33.03 58.275 ;
        RECT 32.77 57.255 33.03 57.515 ;
        RECT 32.77 56.495 33.03 56.755 ;
        RECT 32.77 55.735 33.03 55.995 ;
        RECT 32.77 54.975 33.03 55.235 ;
        RECT 32.77 54.215 33.03 54.475 ;
        RECT 32.77 53.455 33.03 53.715 ;
        RECT 32.77 52.695 33.03 52.955 ;
        RECT 32.77 51.935 33.03 52.195 ;
        RECT 32.77 51.175 33.03 51.435 ;
        RECT 32.77 50.415 33.03 50.675 ;
        RECT 32.77 49.655 33.03 49.915 ;
        RECT 32.77 48.895 33.03 49.155 ;
        RECT 32.77 48.135 33.03 48.395 ;
        RECT 32.77 47.375 33.03 47.635 ;
        RECT 32.77 46.615 33.03 46.875 ;
        RECT 32.77 45.855 33.03 46.115 ;
        RECT 32.77 45.095 33.03 45.355 ;
        RECT 32.77 44.335 33.03 44.595 ;
        RECT 32.77 43.575 33.03 43.835 ;
        RECT 32.77 42.815 33.03 43.075 ;
        RECT 32.77 42.055 33.03 42.315 ;
        RECT 32.77 41.295 33.03 41.555 ;
        RECT 32.77 40.535 33.03 40.795 ;
        RECT 32.77 39.775 33.03 40.035 ;
        RECT 32.77 39.015 33.03 39.275 ;
        RECT 32.77 38.255 33.03 38.515 ;
        RECT 32.77 37.495 33.03 37.755 ;
        RECT 32.77 36.735 33.03 36.995 ;
        RECT 33.53 58.775 33.79 59.035 ;
        RECT 33.53 58.015 33.79 58.275 ;
        RECT 33.53 57.255 33.79 57.515 ;
        RECT 33.53 56.495 33.79 56.755 ;
        RECT 33.53 55.735 33.79 55.995 ;
        RECT 33.53 54.975 33.79 55.235 ;
        RECT 33.53 54.215 33.79 54.475 ;
        RECT 33.53 53.455 33.79 53.715 ;
        RECT 33.53 52.695 33.79 52.955 ;
        RECT 33.53 51.935 33.79 52.195 ;
        RECT 33.53 51.175 33.79 51.435 ;
        RECT 33.53 50.415 33.79 50.675 ;
        RECT 33.53 49.655 33.79 49.915 ;
        RECT 33.53 48.895 33.79 49.155 ;
        RECT 33.53 48.135 33.79 48.395 ;
        RECT 33.53 47.375 33.79 47.635 ;
        RECT 33.53 46.615 33.79 46.875 ;
        RECT 33.53 45.855 33.79 46.115 ;
        RECT 33.53 45.095 33.79 45.355 ;
        RECT 33.53 44.335 33.79 44.595 ;
        RECT 33.53 43.575 33.79 43.835 ;
        RECT 33.53 42.815 33.79 43.075 ;
        RECT 33.53 42.055 33.79 42.315 ;
        RECT 33.53 41.295 33.79 41.555 ;
        RECT 33.53 40.535 33.79 40.795 ;
        RECT 33.53 39.775 33.79 40.035 ;
        RECT 33.53 39.015 33.79 39.275 ;
        RECT 33.53 38.255 33.79 38.515 ;
        RECT 33.53 37.495 33.79 37.755 ;
        RECT 33.53 36.735 33.79 36.995 ;
        RECT 34.29 58.775 34.55 59.035 ;
        RECT 34.29 58.015 34.55 58.275 ;
        RECT 34.29 57.255 34.55 57.515 ;
        RECT 34.29 56.495 34.55 56.755 ;
        RECT 34.29 55.735 34.55 55.995 ;
        RECT 34.29 54.975 34.55 55.235 ;
        RECT 34.29 54.215 34.55 54.475 ;
        RECT 34.29 53.455 34.55 53.715 ;
        RECT 34.29 52.695 34.55 52.955 ;
        RECT 34.29 51.935 34.55 52.195 ;
        RECT 34.29 51.175 34.55 51.435 ;
        RECT 34.29 50.415 34.55 50.675 ;
        RECT 34.29 49.655 34.55 49.915 ;
        RECT 34.29 48.895 34.55 49.155 ;
        RECT 34.29 48.135 34.55 48.395 ;
        RECT 34.29 47.375 34.55 47.635 ;
        RECT 34.29 46.615 34.55 46.875 ;
        RECT 34.29 45.855 34.55 46.115 ;
        RECT 34.29 45.095 34.55 45.355 ;
        RECT 34.29 44.335 34.55 44.595 ;
        RECT 34.29 43.575 34.55 43.835 ;
        RECT 34.29 42.815 34.55 43.075 ;
        RECT 34.29 42.055 34.55 42.315 ;
        RECT 34.29 41.295 34.55 41.555 ;
        RECT 34.29 40.535 34.55 40.795 ;
        RECT 34.29 39.775 34.55 40.035 ;
        RECT 34.29 39.015 34.55 39.275 ;
        RECT 34.29 38.255 34.55 38.515 ;
        RECT 34.29 37.495 34.55 37.755 ;
        RECT 34.29 36.735 34.55 36.995 ;
        RECT 35.05 58.775 35.31 59.035 ;
        RECT 35.05 58.015 35.31 58.275 ;
        RECT 35.05 57.255 35.31 57.515 ;
        RECT 35.05 56.495 35.31 56.755 ;
        RECT 35.05 55.735 35.31 55.995 ;
        RECT 35.05 54.975 35.31 55.235 ;
        RECT 35.05 54.215 35.31 54.475 ;
        RECT 35.05 53.455 35.31 53.715 ;
        RECT 35.05 52.695 35.31 52.955 ;
        RECT 35.05 51.935 35.31 52.195 ;
        RECT 35.05 51.175 35.31 51.435 ;
        RECT 35.05 50.415 35.31 50.675 ;
        RECT 35.05 49.655 35.31 49.915 ;
        RECT 35.05 48.895 35.31 49.155 ;
        RECT 35.05 48.135 35.31 48.395 ;
        RECT 35.05 47.375 35.31 47.635 ;
        RECT 35.05 46.615 35.31 46.875 ;
        RECT 35.05 45.855 35.31 46.115 ;
        RECT 35.05 45.095 35.31 45.355 ;
        RECT 35.05 44.335 35.31 44.595 ;
        RECT 35.05 43.575 35.31 43.835 ;
        RECT 35.05 42.815 35.31 43.075 ;
        RECT 35.05 42.055 35.31 42.315 ;
        RECT 35.05 41.295 35.31 41.555 ;
        RECT 35.05 40.535 35.31 40.795 ;
        RECT 35.05 39.775 35.31 40.035 ;
        RECT 35.05 39.015 35.31 39.275 ;
        RECT 35.05 38.255 35.31 38.515 ;
        RECT 35.05 37.495 35.31 37.755 ;
        RECT 35.05 36.735 35.31 36.995 ;
        RECT 35.81 58.775 36.07 59.035 ;
        RECT 35.81 58.015 36.07 58.275 ;
        RECT 35.81 57.255 36.07 57.515 ;
        RECT 35.81 56.495 36.07 56.755 ;
        RECT 35.81 55.735 36.07 55.995 ;
        RECT 35.81 54.975 36.07 55.235 ;
        RECT 35.81 54.215 36.07 54.475 ;
        RECT 35.81 53.455 36.07 53.715 ;
        RECT 35.81 52.695 36.07 52.955 ;
        RECT 35.81 51.935 36.07 52.195 ;
        RECT 35.81 51.175 36.07 51.435 ;
        RECT 35.81 50.415 36.07 50.675 ;
        RECT 35.81 49.655 36.07 49.915 ;
        RECT 35.81 48.895 36.07 49.155 ;
        RECT 35.81 48.135 36.07 48.395 ;
        RECT 35.81 47.375 36.07 47.635 ;
        RECT 35.81 46.615 36.07 46.875 ;
        RECT 35.81 45.855 36.07 46.115 ;
        RECT 35.81 45.095 36.07 45.355 ;
        RECT 35.81 44.335 36.07 44.595 ;
        RECT 35.81 43.575 36.07 43.835 ;
        RECT 35.81 42.815 36.07 43.075 ;
        RECT 35.81 42.055 36.07 42.315 ;
        RECT 35.81 41.295 36.07 41.555 ;
        RECT 35.81 40.535 36.07 40.795 ;
        RECT 35.81 39.775 36.07 40.035 ;
        RECT 35.81 39.015 36.07 39.275 ;
        RECT 35.81 38.255 36.07 38.515 ;
        RECT 35.81 37.495 36.07 37.755 ;
        RECT 35.81 36.735 36.07 36.995 ;
        RECT 36.57 58.775 36.83 59.035 ;
        RECT 36.57 58.015 36.83 58.275 ;
        RECT 36.57 57.255 36.83 57.515 ;
        RECT 36.57 56.495 36.83 56.755 ;
        RECT 36.57 55.735 36.83 55.995 ;
        RECT 36.57 54.975 36.83 55.235 ;
        RECT 36.57 54.215 36.83 54.475 ;
        RECT 36.57 53.455 36.83 53.715 ;
        RECT 36.57 52.695 36.83 52.955 ;
        RECT 36.57 51.935 36.83 52.195 ;
        RECT 36.57 51.175 36.83 51.435 ;
        RECT 36.57 50.415 36.83 50.675 ;
        RECT 36.57 49.655 36.83 49.915 ;
        RECT 36.57 48.895 36.83 49.155 ;
        RECT 36.57 48.135 36.83 48.395 ;
        RECT 36.57 47.375 36.83 47.635 ;
        RECT 36.57 46.615 36.83 46.875 ;
        RECT 36.57 45.855 36.83 46.115 ;
        RECT 36.57 45.095 36.83 45.355 ;
        RECT 36.57 44.335 36.83 44.595 ;
        RECT 36.57 43.575 36.83 43.835 ;
        RECT 36.57 42.815 36.83 43.075 ;
        RECT 36.57 42.055 36.83 42.315 ;
        RECT 36.57 41.295 36.83 41.555 ;
        RECT 36.57 40.535 36.83 40.795 ;
        RECT 36.57 39.775 36.83 40.035 ;
        RECT 36.57 39.015 36.83 39.275 ;
        RECT 36.57 38.255 36.83 38.515 ;
        RECT 36.57 37.495 36.83 37.755 ;
        RECT 36.57 36.735 36.83 36.995 ;
        RECT 37.33 58.775 37.59 59.035 ;
        RECT 37.33 58.015 37.59 58.275 ;
        RECT 37.33 57.255 37.59 57.515 ;
        RECT 37.33 56.495 37.59 56.755 ;
        RECT 37.33 55.735 37.59 55.995 ;
        RECT 37.33 54.975 37.59 55.235 ;
        RECT 37.33 54.215 37.59 54.475 ;
        RECT 37.33 53.455 37.59 53.715 ;
        RECT 37.33 52.695 37.59 52.955 ;
        RECT 37.33 51.935 37.59 52.195 ;
        RECT 37.33 51.175 37.59 51.435 ;
        RECT 37.33 50.415 37.59 50.675 ;
        RECT 37.33 49.655 37.59 49.915 ;
        RECT 37.33 48.895 37.59 49.155 ;
        RECT 37.33 48.135 37.59 48.395 ;
        RECT 37.33 47.375 37.59 47.635 ;
        RECT 37.33 46.615 37.59 46.875 ;
        RECT 37.33 45.855 37.59 46.115 ;
        RECT 37.33 45.095 37.59 45.355 ;
        RECT 37.33 44.335 37.59 44.595 ;
        RECT 37.33 43.575 37.59 43.835 ;
        RECT 37.33 42.815 37.59 43.075 ;
        RECT 37.33 42.055 37.59 42.315 ;
        RECT 37.33 41.295 37.59 41.555 ;
        RECT 37.33 40.535 37.59 40.795 ;
        RECT 37.33 39.775 37.59 40.035 ;
        RECT 37.33 39.015 37.59 39.275 ;
        RECT 37.33 38.255 37.59 38.515 ;
        RECT 37.33 37.495 37.59 37.755 ;
        RECT 37.33 36.735 37.59 36.995 ;
        RECT 38.09 58.775 38.35 59.035 ;
        RECT 38.09 58.015 38.35 58.275 ;
        RECT 38.09 57.255 38.35 57.515 ;
        RECT 38.09 56.495 38.35 56.755 ;
        RECT 38.09 55.735 38.35 55.995 ;
        RECT 38.09 54.975 38.35 55.235 ;
        RECT 38.09 54.215 38.35 54.475 ;
        RECT 38.09 53.455 38.35 53.715 ;
        RECT 38.09 52.695 38.35 52.955 ;
        RECT 38.09 51.935 38.35 52.195 ;
        RECT 38.09 51.175 38.35 51.435 ;
        RECT 38.09 50.415 38.35 50.675 ;
        RECT 38.09 49.655 38.35 49.915 ;
        RECT 38.09 48.895 38.35 49.155 ;
        RECT 38.09 48.135 38.35 48.395 ;
        RECT 38.09 47.375 38.35 47.635 ;
        RECT 38.09 46.615 38.35 46.875 ;
        RECT 38.09 45.855 38.35 46.115 ;
        RECT 38.09 45.095 38.35 45.355 ;
        RECT 38.09 44.335 38.35 44.595 ;
        RECT 38.09 43.575 38.35 43.835 ;
        RECT 38.09 42.815 38.35 43.075 ;
        RECT 38.09 42.055 38.35 42.315 ;
        RECT 38.09 41.295 38.35 41.555 ;
        RECT 38.09 40.535 38.35 40.795 ;
        RECT 38.09 39.775 38.35 40.035 ;
        RECT 38.09 39.015 38.35 39.275 ;
        RECT 38.09 38.255 38.35 38.515 ;
        RECT 38.09 37.495 38.35 37.755 ;
        RECT 38.09 36.735 38.35 36.995 ;
        RECT 38.85 58.775 39.11 59.035 ;
        RECT 38.85 58.015 39.11 58.275 ;
        RECT 38.85 57.255 39.11 57.515 ;
        RECT 38.85 56.495 39.11 56.755 ;
        RECT 38.85 55.735 39.11 55.995 ;
        RECT 38.85 54.975 39.11 55.235 ;
        RECT 38.85 54.215 39.11 54.475 ;
        RECT 38.85 53.455 39.11 53.715 ;
        RECT 38.85 52.695 39.11 52.955 ;
        RECT 38.85 51.935 39.11 52.195 ;
        RECT 38.85 51.175 39.11 51.435 ;
        RECT 38.85 50.415 39.11 50.675 ;
        RECT 38.85 49.655 39.11 49.915 ;
        RECT 38.85 48.895 39.11 49.155 ;
        RECT 38.85 48.135 39.11 48.395 ;
        RECT 38.85 47.375 39.11 47.635 ;
        RECT 38.85 46.615 39.11 46.875 ;
        RECT 38.85 45.855 39.11 46.115 ;
        RECT 38.85 45.095 39.11 45.355 ;
        RECT 38.85 44.335 39.11 44.595 ;
        RECT 38.85 43.575 39.11 43.835 ;
        RECT 38.85 42.815 39.11 43.075 ;
        RECT 38.85 42.055 39.11 42.315 ;
        RECT 38.85 41.295 39.11 41.555 ;
        RECT 38.85 40.535 39.11 40.795 ;
        RECT 38.85 39.775 39.11 40.035 ;
        RECT 38.85 39.015 39.11 39.275 ;
        RECT 38.85 38.255 39.11 38.515 ;
        RECT 38.85 37.495 39.11 37.755 ;
        RECT 38.85 36.735 39.11 36.995 ;
        RECT 39.61 58.775 39.87 59.035 ;
        RECT 39.61 58.015 39.87 58.275 ;
        RECT 39.61 57.255 39.87 57.515 ;
        RECT 39.61 56.495 39.87 56.755 ;
        RECT 39.61 55.735 39.87 55.995 ;
        RECT 39.61 54.975 39.87 55.235 ;
        RECT 39.61 54.215 39.87 54.475 ;
        RECT 39.61 53.455 39.87 53.715 ;
        RECT 39.61 52.695 39.87 52.955 ;
        RECT 39.61 51.935 39.87 52.195 ;
        RECT 39.61 51.175 39.87 51.435 ;
        RECT 39.61 50.415 39.87 50.675 ;
        RECT 39.61 49.655 39.87 49.915 ;
        RECT 39.61 48.895 39.87 49.155 ;
        RECT 39.61 48.135 39.87 48.395 ;
        RECT 39.61 47.375 39.87 47.635 ;
        RECT 39.61 46.615 39.87 46.875 ;
        RECT 39.61 45.855 39.87 46.115 ;
        RECT 39.61 45.095 39.87 45.355 ;
        RECT 39.61 44.335 39.87 44.595 ;
        RECT 39.61 43.575 39.87 43.835 ;
        RECT 39.61 42.815 39.87 43.075 ;
        RECT 39.61 42.055 39.87 42.315 ;
        RECT 39.61 41.295 39.87 41.555 ;
        RECT 39.61 40.535 39.87 40.795 ;
        RECT 39.61 39.775 39.87 40.035 ;
        RECT 39.61 39.015 39.87 39.275 ;
        RECT 39.61 38.255 39.87 38.515 ;
        RECT 39.61 37.495 39.87 37.755 ;
        RECT 39.61 36.735 39.87 36.995 ;
        RECT 40.37 58.775 40.63 59.035 ;
        RECT 40.37 58.015 40.63 58.275 ;
        RECT 40.37 57.255 40.63 57.515 ;
        RECT 40.37 56.495 40.63 56.755 ;
        RECT 40.37 55.735 40.63 55.995 ;
        RECT 40.37 54.975 40.63 55.235 ;
        RECT 40.37 54.215 40.63 54.475 ;
        RECT 40.37 53.455 40.63 53.715 ;
        RECT 40.37 52.695 40.63 52.955 ;
        RECT 40.37 51.935 40.63 52.195 ;
        RECT 40.37 51.175 40.63 51.435 ;
        RECT 40.37 50.415 40.63 50.675 ;
        RECT 40.37 49.655 40.63 49.915 ;
        RECT 40.37 48.895 40.63 49.155 ;
        RECT 40.37 48.135 40.63 48.395 ;
        RECT 40.37 47.375 40.63 47.635 ;
        RECT 40.37 46.615 40.63 46.875 ;
        RECT 40.37 45.855 40.63 46.115 ;
        RECT 40.37 45.095 40.63 45.355 ;
        RECT 40.37 44.335 40.63 44.595 ;
        RECT 40.37 43.575 40.63 43.835 ;
        RECT 40.37 42.815 40.63 43.075 ;
        RECT 40.37 42.055 40.63 42.315 ;
        RECT 40.37 41.295 40.63 41.555 ;
        RECT 40.37 40.535 40.63 40.795 ;
        RECT 40.37 39.775 40.63 40.035 ;
        RECT 40.37 39.015 40.63 39.275 ;
        RECT 40.37 38.255 40.63 38.515 ;
        RECT 40.37 37.495 40.63 37.755 ;
        RECT 40.37 36.735 40.63 36.995 ;
        RECT 41.13 58.775 41.39 59.035 ;
        RECT 41.13 58.015 41.39 58.275 ;
        RECT 41.13 57.255 41.39 57.515 ;
        RECT 41.13 56.495 41.39 56.755 ;
        RECT 41.13 55.735 41.39 55.995 ;
        RECT 41.13 54.975 41.39 55.235 ;
        RECT 41.13 54.215 41.39 54.475 ;
        RECT 41.13 53.455 41.39 53.715 ;
        RECT 41.13 52.695 41.39 52.955 ;
        RECT 41.13 51.935 41.39 52.195 ;
        RECT 41.13 51.175 41.39 51.435 ;
        RECT 41.13 50.415 41.39 50.675 ;
        RECT 41.13 49.655 41.39 49.915 ;
        RECT 41.13 48.895 41.39 49.155 ;
        RECT 41.13 48.135 41.39 48.395 ;
        RECT 41.13 47.375 41.39 47.635 ;
        RECT 41.13 46.615 41.39 46.875 ;
        RECT 41.13 45.855 41.39 46.115 ;
        RECT 41.13 45.095 41.39 45.355 ;
        RECT 41.13 44.335 41.39 44.595 ;
        RECT 41.13 43.575 41.39 43.835 ;
        RECT 41.13 42.815 41.39 43.075 ;
        RECT 41.13 42.055 41.39 42.315 ;
        RECT 41.13 41.295 41.39 41.555 ;
        RECT 41.13 40.535 41.39 40.795 ;
        RECT 41.13 39.775 41.39 40.035 ;
        RECT 41.13 39.015 41.39 39.275 ;
        RECT 41.13 38.255 41.39 38.515 ;
        RECT 41.13 37.495 41.39 37.755 ;
        RECT 41.13 36.735 41.39 36.995 ;
        RECT 41.89 58.775 42.15 59.035 ;
        RECT 41.89 58.015 42.15 58.275 ;
        RECT 41.89 57.255 42.15 57.515 ;
        RECT 41.89 56.495 42.15 56.755 ;
        RECT 41.89 55.735 42.15 55.995 ;
        RECT 41.89 54.975 42.15 55.235 ;
        RECT 41.89 54.215 42.15 54.475 ;
        RECT 41.89 53.455 42.15 53.715 ;
        RECT 41.89 52.695 42.15 52.955 ;
        RECT 41.89 51.935 42.15 52.195 ;
        RECT 41.89 51.175 42.15 51.435 ;
        RECT 41.89 50.415 42.15 50.675 ;
        RECT 41.89 49.655 42.15 49.915 ;
        RECT 41.89 48.895 42.15 49.155 ;
        RECT 41.89 48.135 42.15 48.395 ;
        RECT 41.89 47.375 42.15 47.635 ;
        RECT 41.89 46.615 42.15 46.875 ;
        RECT 41.89 45.855 42.15 46.115 ;
        RECT 41.89 45.095 42.15 45.355 ;
        RECT 41.89 44.335 42.15 44.595 ;
        RECT 41.89 43.575 42.15 43.835 ;
        RECT 41.89 42.815 42.15 43.075 ;
        RECT 41.89 42.055 42.15 42.315 ;
        RECT 41.89 41.295 42.15 41.555 ;
        RECT 41.89 40.535 42.15 40.795 ;
        RECT 41.89 39.775 42.15 40.035 ;
        RECT 41.89 39.015 42.15 39.275 ;
        RECT 41.89 38.255 42.15 38.515 ;
        RECT 41.89 37.495 42.15 37.755 ;
        RECT 41.89 36.735 42.15 36.995 ;
        RECT 42.65 58.775 42.91 59.035 ;
        RECT 42.65 58.015 42.91 58.275 ;
        RECT 42.65 57.255 42.91 57.515 ;
        RECT 42.65 56.495 42.91 56.755 ;
        RECT 42.65 55.735 42.91 55.995 ;
        RECT 42.65 54.975 42.91 55.235 ;
        RECT 42.65 54.215 42.91 54.475 ;
        RECT 42.65 53.455 42.91 53.715 ;
        RECT 42.65 52.695 42.91 52.955 ;
        RECT 42.65 51.935 42.91 52.195 ;
        RECT 42.65 51.175 42.91 51.435 ;
        RECT 42.65 50.415 42.91 50.675 ;
        RECT 42.65 49.655 42.91 49.915 ;
        RECT 42.65 48.895 42.91 49.155 ;
        RECT 42.65 48.135 42.91 48.395 ;
        RECT 42.65 47.375 42.91 47.635 ;
        RECT 42.65 46.615 42.91 46.875 ;
        RECT 42.65 45.855 42.91 46.115 ;
        RECT 42.65 45.095 42.91 45.355 ;
        RECT 42.65 44.335 42.91 44.595 ;
        RECT 42.65 43.575 42.91 43.835 ;
        RECT 42.65 42.815 42.91 43.075 ;
        RECT 42.65 42.055 42.91 42.315 ;
        RECT 42.65 41.295 42.91 41.555 ;
        RECT 42.65 40.535 42.91 40.795 ;
        RECT 42.65 39.775 42.91 40.035 ;
        RECT 42.65 39.015 42.91 39.275 ;
        RECT 42.65 38.255 42.91 38.515 ;
        RECT 42.65 37.495 42.91 37.755 ;
        RECT 42.65 36.735 42.91 36.995 ;
        RECT 43.41 58.775 43.67 59.035 ;
        RECT 43.41 58.015 43.67 58.275 ;
        RECT 43.41 57.255 43.67 57.515 ;
        RECT 43.41 56.495 43.67 56.755 ;
        RECT 43.41 55.735 43.67 55.995 ;
        RECT 43.41 54.975 43.67 55.235 ;
        RECT 43.41 54.215 43.67 54.475 ;
        RECT 43.41 53.455 43.67 53.715 ;
        RECT 43.41 52.695 43.67 52.955 ;
        RECT 43.41 51.935 43.67 52.195 ;
        RECT 43.41 51.175 43.67 51.435 ;
        RECT 43.41 50.415 43.67 50.675 ;
        RECT 43.41 49.655 43.67 49.915 ;
        RECT 43.41 48.895 43.67 49.155 ;
        RECT 43.41 48.135 43.67 48.395 ;
        RECT 43.41 47.375 43.67 47.635 ;
        RECT 43.41 46.615 43.67 46.875 ;
        RECT 43.41 45.855 43.67 46.115 ;
        RECT 43.41 45.095 43.67 45.355 ;
        RECT 43.41 44.335 43.67 44.595 ;
        RECT 43.41 43.575 43.67 43.835 ;
        RECT 43.41 42.815 43.67 43.075 ;
        RECT 43.41 42.055 43.67 42.315 ;
        RECT 43.41 41.295 43.67 41.555 ;
        RECT 43.41 40.535 43.67 40.795 ;
        RECT 43.41 39.775 43.67 40.035 ;
        RECT 43.41 39.015 43.67 39.275 ;
        RECT 43.41 38.255 43.67 38.515 ;
        RECT 43.41 37.495 43.67 37.755 ;
        RECT 43.41 36.735 43.67 36.995 ;
        RECT 44.17 58.775 44.43 59.035 ;
        RECT 44.17 58.015 44.43 58.275 ;
        RECT 44.17 57.255 44.43 57.515 ;
        RECT 44.17 56.495 44.43 56.755 ;
        RECT 44.17 55.735 44.43 55.995 ;
        RECT 44.17 54.975 44.43 55.235 ;
        RECT 44.17 54.215 44.43 54.475 ;
        RECT 44.17 53.455 44.43 53.715 ;
        RECT 44.17 52.695 44.43 52.955 ;
        RECT 44.17 51.935 44.43 52.195 ;
        RECT 44.17 51.175 44.43 51.435 ;
        RECT 44.17 50.415 44.43 50.675 ;
        RECT 44.17 49.655 44.43 49.915 ;
        RECT 44.17 48.895 44.43 49.155 ;
        RECT 44.17 48.135 44.43 48.395 ;
        RECT 44.17 47.375 44.43 47.635 ;
        RECT 44.17 46.615 44.43 46.875 ;
        RECT 44.17 45.855 44.43 46.115 ;
        RECT 44.17 45.095 44.43 45.355 ;
        RECT 44.17 44.335 44.43 44.595 ;
        RECT 44.17 43.575 44.43 43.835 ;
        RECT 44.17 42.815 44.43 43.075 ;
        RECT 44.17 42.055 44.43 42.315 ;
        RECT 44.17 41.295 44.43 41.555 ;
        RECT 44.17 40.535 44.43 40.795 ;
        RECT 44.17 39.775 44.43 40.035 ;
        RECT 44.17 39.015 44.43 39.275 ;
        RECT 44.17 38.255 44.43 38.515 ;
        RECT 44.17 37.495 44.43 37.755 ;
        RECT 44.17 36.735 44.43 36.995 ;
        RECT 44.93 58.775 45.19 59.035 ;
        RECT 44.93 58.015 45.19 58.275 ;
        RECT 44.93 57.255 45.19 57.515 ;
        RECT 44.93 56.495 45.19 56.755 ;
        RECT 44.93 55.735 45.19 55.995 ;
        RECT 44.93 54.975 45.19 55.235 ;
        RECT 44.93 54.215 45.19 54.475 ;
        RECT 44.93 53.455 45.19 53.715 ;
        RECT 44.93 52.695 45.19 52.955 ;
        RECT 44.93 51.935 45.19 52.195 ;
        RECT 44.93 51.175 45.19 51.435 ;
        RECT 44.93 50.415 45.19 50.675 ;
        RECT 44.93 49.655 45.19 49.915 ;
        RECT 44.93 48.895 45.19 49.155 ;
        RECT 44.93 48.135 45.19 48.395 ;
        RECT 44.93 47.375 45.19 47.635 ;
        RECT 44.93 46.615 45.19 46.875 ;
        RECT 44.93 45.855 45.19 46.115 ;
        RECT 44.93 45.095 45.19 45.355 ;
        RECT 44.93 44.335 45.19 44.595 ;
        RECT 44.93 43.575 45.19 43.835 ;
        RECT 44.93 42.815 45.19 43.075 ;
        RECT 44.93 42.055 45.19 42.315 ;
        RECT 44.93 41.295 45.19 41.555 ;
        RECT 44.93 40.535 45.19 40.795 ;
        RECT 44.93 39.775 45.19 40.035 ;
        RECT 44.93 39.015 45.19 39.275 ;
        RECT 44.93 38.255 45.19 38.515 ;
        RECT 44.93 37.495 45.19 37.755 ;
        RECT 44.93 36.735 45.19 36.995 ;
        RECT 45.69 58.775 45.95 59.035 ;
        RECT 45.69 58.015 45.95 58.275 ;
        RECT 45.69 57.255 45.95 57.515 ;
        RECT 45.69 56.495 45.95 56.755 ;
        RECT 45.69 55.735 45.95 55.995 ;
        RECT 45.69 54.975 45.95 55.235 ;
        RECT 45.69 54.215 45.95 54.475 ;
        RECT 45.69 53.455 45.95 53.715 ;
        RECT 45.69 52.695 45.95 52.955 ;
        RECT 45.69 51.935 45.95 52.195 ;
        RECT 45.69 51.175 45.95 51.435 ;
        RECT 45.69 50.415 45.95 50.675 ;
        RECT 45.69 49.655 45.95 49.915 ;
        RECT 45.69 48.895 45.95 49.155 ;
        RECT 45.69 48.135 45.95 48.395 ;
        RECT 45.69 47.375 45.95 47.635 ;
        RECT 45.69 46.615 45.95 46.875 ;
        RECT 45.69 45.855 45.95 46.115 ;
        RECT 45.69 45.095 45.95 45.355 ;
        RECT 45.69 44.335 45.95 44.595 ;
        RECT 45.69 43.575 45.95 43.835 ;
        RECT 45.69 42.815 45.95 43.075 ;
        RECT 45.69 42.055 45.95 42.315 ;
        RECT 45.69 41.295 45.95 41.555 ;
        RECT 45.69 40.535 45.95 40.795 ;
        RECT 45.69 39.775 45.95 40.035 ;
        RECT 45.69 39.015 45.95 39.275 ;
        RECT 45.69 38.255 45.95 38.515 ;
        RECT 45.69 37.495 45.95 37.755 ;
        RECT 45.69 36.735 45.95 36.995 ;
        RECT 46.45 58.775 46.71 59.035 ;
        RECT 46.45 58.015 46.71 58.275 ;
        RECT 46.45 57.255 46.71 57.515 ;
        RECT 46.45 56.495 46.71 56.755 ;
        RECT 46.45 55.735 46.71 55.995 ;
        RECT 46.45 54.975 46.71 55.235 ;
        RECT 46.45 54.215 46.71 54.475 ;
        RECT 46.45 53.455 46.71 53.715 ;
        RECT 46.45 52.695 46.71 52.955 ;
        RECT 46.45 51.935 46.71 52.195 ;
        RECT 46.45 51.175 46.71 51.435 ;
        RECT 46.45 50.415 46.71 50.675 ;
        RECT 46.45 49.655 46.71 49.915 ;
        RECT 46.45 48.895 46.71 49.155 ;
        RECT 46.45 48.135 46.71 48.395 ;
        RECT 46.45 47.375 46.71 47.635 ;
        RECT 46.45 46.615 46.71 46.875 ;
        RECT 46.45 45.855 46.71 46.115 ;
        RECT 46.45 45.095 46.71 45.355 ;
        RECT 46.45 44.335 46.71 44.595 ;
        RECT 46.45 43.575 46.71 43.835 ;
        RECT 46.45 42.815 46.71 43.075 ;
        RECT 46.45 42.055 46.71 42.315 ;
        RECT 46.45 41.295 46.71 41.555 ;
        RECT 46.45 40.535 46.71 40.795 ;
        RECT 46.45 39.775 46.71 40.035 ;
        RECT 46.45 39.015 46.71 39.275 ;
        RECT 46.45 38.255 46.71 38.515 ;
        RECT 46.45 37.495 46.71 37.755 ;
        RECT 46.45 36.735 46.71 36.995 ;
        RECT 47.21 58.775 47.47 59.035 ;
        RECT 47.21 58.015 47.47 58.275 ;
        RECT 47.21 57.255 47.47 57.515 ;
        RECT 47.21 56.495 47.47 56.755 ;
        RECT 47.21 55.735 47.47 55.995 ;
        RECT 47.21 54.975 47.47 55.235 ;
        RECT 47.21 54.215 47.47 54.475 ;
        RECT 47.21 53.455 47.47 53.715 ;
        RECT 47.21 52.695 47.47 52.955 ;
        RECT 47.21 51.935 47.47 52.195 ;
        RECT 47.21 51.175 47.47 51.435 ;
        RECT 47.21 50.415 47.47 50.675 ;
        RECT 47.21 49.655 47.47 49.915 ;
        RECT 47.21 48.895 47.47 49.155 ;
        RECT 47.21 48.135 47.47 48.395 ;
        RECT 47.21 47.375 47.47 47.635 ;
        RECT 47.21 46.615 47.47 46.875 ;
        RECT 47.21 45.855 47.47 46.115 ;
        RECT 47.21 45.095 47.47 45.355 ;
        RECT 47.21 44.335 47.47 44.595 ;
        RECT 47.21 43.575 47.47 43.835 ;
        RECT 47.21 42.815 47.47 43.075 ;
        RECT 47.21 42.055 47.47 42.315 ;
        RECT 47.21 41.295 47.47 41.555 ;
        RECT 47.21 40.535 47.47 40.795 ;
        RECT 47.21 39.775 47.47 40.035 ;
        RECT 47.21 39.015 47.47 39.275 ;
        RECT 47.21 38.255 47.47 38.515 ;
        RECT 47.21 37.495 47.47 37.755 ;
        RECT 47.21 36.735 47.47 36.995 ;
        RECT 47.97 58.775 48.23 59.035 ;
        RECT 47.97 58.015 48.23 58.275 ;
        RECT 47.97 57.255 48.23 57.515 ;
        RECT 47.97 56.495 48.23 56.755 ;
        RECT 47.97 55.735 48.23 55.995 ;
        RECT 47.97 54.975 48.23 55.235 ;
        RECT 47.97 54.215 48.23 54.475 ;
        RECT 47.97 53.455 48.23 53.715 ;
        RECT 47.97 52.695 48.23 52.955 ;
        RECT 47.97 51.935 48.23 52.195 ;
        RECT 47.97 51.175 48.23 51.435 ;
        RECT 47.97 50.415 48.23 50.675 ;
        RECT 47.97 49.655 48.23 49.915 ;
        RECT 47.97 48.895 48.23 49.155 ;
        RECT 47.97 48.135 48.23 48.395 ;
        RECT 47.97 47.375 48.23 47.635 ;
        RECT 47.97 46.615 48.23 46.875 ;
        RECT 47.97 45.855 48.23 46.115 ;
        RECT 47.97 45.095 48.23 45.355 ;
        RECT 47.97 44.335 48.23 44.595 ;
        RECT 47.97 43.575 48.23 43.835 ;
        RECT 47.97 42.815 48.23 43.075 ;
        RECT 47.97 42.055 48.23 42.315 ;
        RECT 47.97 41.295 48.23 41.555 ;
        RECT 47.97 40.535 48.23 40.795 ;
        RECT 47.97 39.775 48.23 40.035 ;
        RECT 47.97 39.015 48.23 39.275 ;
        RECT 47.97 38.255 48.23 38.515 ;
        RECT 47.97 37.495 48.23 37.755 ;
        RECT 47.97 36.735 48.23 36.995 ;
        RECT 48.73 58.775 48.99 59.035 ;
        RECT 48.73 58.015 48.99 58.275 ;
        RECT 48.73 57.255 48.99 57.515 ;
        RECT 48.73 56.495 48.99 56.755 ;
        RECT 48.73 55.735 48.99 55.995 ;
        RECT 48.73 54.975 48.99 55.235 ;
        RECT 48.73 54.215 48.99 54.475 ;
        RECT 48.73 53.455 48.99 53.715 ;
        RECT 48.73 52.695 48.99 52.955 ;
        RECT 48.73 51.935 48.99 52.195 ;
        RECT 48.73 51.175 48.99 51.435 ;
        RECT 48.73 50.415 48.99 50.675 ;
        RECT 48.73 49.655 48.99 49.915 ;
        RECT 48.73 48.895 48.99 49.155 ;
        RECT 48.73 48.135 48.99 48.395 ;
        RECT 48.73 47.375 48.99 47.635 ;
        RECT 48.73 46.615 48.99 46.875 ;
        RECT 48.73 45.855 48.99 46.115 ;
        RECT 48.73 45.095 48.99 45.355 ;
        RECT 48.73 44.335 48.99 44.595 ;
        RECT 48.73 43.575 48.99 43.835 ;
        RECT 48.73 42.815 48.99 43.075 ;
        RECT 48.73 42.055 48.99 42.315 ;
        RECT 48.73 41.295 48.99 41.555 ;
        RECT 48.73 40.535 48.99 40.795 ;
        RECT 48.73 39.775 48.99 40.035 ;
        RECT 48.73 39.015 48.99 39.275 ;
        RECT 48.73 38.255 48.99 38.515 ;
        RECT 48.73 37.495 48.99 37.755 ;
        RECT 48.73 36.735 48.99 36.995 ;
        RECT 49.49 58.775 49.75 59.035 ;
        RECT 49.49 58.015 49.75 58.275 ;
        RECT 49.49 57.255 49.75 57.515 ;
        RECT 49.49 56.495 49.75 56.755 ;
        RECT 49.49 55.735 49.75 55.995 ;
        RECT 49.49 54.975 49.75 55.235 ;
        RECT 49.49 54.215 49.75 54.475 ;
        RECT 49.49 53.455 49.75 53.715 ;
        RECT 49.49 52.695 49.75 52.955 ;
        RECT 49.49 51.935 49.75 52.195 ;
        RECT 49.49 51.175 49.75 51.435 ;
        RECT 49.49 50.415 49.75 50.675 ;
        RECT 49.49 49.655 49.75 49.915 ;
        RECT 49.49 48.895 49.75 49.155 ;
        RECT 49.49 48.135 49.75 48.395 ;
        RECT 49.49 47.375 49.75 47.635 ;
        RECT 49.49 46.615 49.75 46.875 ;
        RECT 49.49 45.855 49.75 46.115 ;
        RECT 49.49 45.095 49.75 45.355 ;
        RECT 49.49 44.335 49.75 44.595 ;
        RECT 49.49 43.575 49.75 43.835 ;
        RECT 49.49 42.815 49.75 43.075 ;
        RECT 49.49 42.055 49.75 42.315 ;
        RECT 49.49 41.295 49.75 41.555 ;
        RECT 49.49 40.535 49.75 40.795 ;
        RECT 49.49 39.775 49.75 40.035 ;
        RECT 49.49 39.015 49.75 39.275 ;
        RECT 49.49 38.255 49.75 38.515 ;
        RECT 49.49 37.495 49.75 37.755 ;
        RECT 49.49 36.735 49.75 36.995 ;
        RECT 50.25 58.775 50.51 59.035 ;
        RECT 50.25 58.015 50.51 58.275 ;
        RECT 50.25 57.255 50.51 57.515 ;
        RECT 50.25 56.495 50.51 56.755 ;
        RECT 50.25 55.735 50.51 55.995 ;
        RECT 50.25 54.975 50.51 55.235 ;
        RECT 50.25 54.215 50.51 54.475 ;
        RECT 50.25 53.455 50.51 53.715 ;
        RECT 50.25 52.695 50.51 52.955 ;
        RECT 50.25 51.935 50.51 52.195 ;
        RECT 50.25 51.175 50.51 51.435 ;
        RECT 50.25 50.415 50.51 50.675 ;
        RECT 50.25 49.655 50.51 49.915 ;
        RECT 50.25 48.895 50.51 49.155 ;
        RECT 50.25 48.135 50.51 48.395 ;
        RECT 50.25 47.375 50.51 47.635 ;
        RECT 50.25 46.615 50.51 46.875 ;
        RECT 50.25 45.855 50.51 46.115 ;
        RECT 50.25 45.095 50.51 45.355 ;
        RECT 50.25 44.335 50.51 44.595 ;
        RECT 50.25 43.575 50.51 43.835 ;
        RECT 50.25 42.815 50.51 43.075 ;
        RECT 50.25 42.055 50.51 42.315 ;
        RECT 50.25 41.295 50.51 41.555 ;
        RECT 50.25 40.535 50.51 40.795 ;
        RECT 50.25 39.775 50.51 40.035 ;
        RECT 50.25 39.015 50.51 39.275 ;
        RECT 50.25 38.255 50.51 38.515 ;
        RECT 50.25 37.495 50.51 37.755 ;
        RECT 50.25 36.735 50.51 36.995 ;
        RECT 51.01 58.775 51.27 59.035 ;
        RECT 51.01 58.015 51.27 58.275 ;
        RECT 51.01 57.255 51.27 57.515 ;
        RECT 51.01 56.495 51.27 56.755 ;
        RECT 51.01 55.735 51.27 55.995 ;
        RECT 51.01 54.975 51.27 55.235 ;
        RECT 51.01 54.215 51.27 54.475 ;
        RECT 51.01 53.455 51.27 53.715 ;
        RECT 51.01 52.695 51.27 52.955 ;
        RECT 51.01 51.935 51.27 52.195 ;
        RECT 51.01 51.175 51.27 51.435 ;
        RECT 51.01 50.415 51.27 50.675 ;
        RECT 51.01 49.655 51.27 49.915 ;
        RECT 51.01 48.895 51.27 49.155 ;
        RECT 51.01 48.135 51.27 48.395 ;
        RECT 51.01 47.375 51.27 47.635 ;
        RECT 51.01 46.615 51.27 46.875 ;
        RECT 51.01 45.855 51.27 46.115 ;
        RECT 51.01 45.095 51.27 45.355 ;
        RECT 51.01 44.335 51.27 44.595 ;
        RECT 51.01 43.575 51.27 43.835 ;
        RECT 51.01 42.815 51.27 43.075 ;
        RECT 51.01 42.055 51.27 42.315 ;
        RECT 51.01 41.295 51.27 41.555 ;
        RECT 51.01 40.535 51.27 40.795 ;
        RECT 51.01 39.775 51.27 40.035 ;
        RECT 51.01 39.015 51.27 39.275 ;
        RECT 51.01 38.255 51.27 38.515 ;
        RECT 51.01 37.495 51.27 37.755 ;
        RECT 51.01 36.735 51.27 36.995 ;
        RECT 51.77 58.775 52.03 59.035 ;
        RECT 51.77 58.015 52.03 58.275 ;
        RECT 51.77 57.255 52.03 57.515 ;
        RECT 51.77 56.495 52.03 56.755 ;
        RECT 51.77 55.735 52.03 55.995 ;
        RECT 51.77 54.975 52.03 55.235 ;
        RECT 51.77 54.215 52.03 54.475 ;
        RECT 51.77 53.455 52.03 53.715 ;
        RECT 51.77 52.695 52.03 52.955 ;
        RECT 51.77 51.935 52.03 52.195 ;
        RECT 51.77 51.175 52.03 51.435 ;
        RECT 51.77 50.415 52.03 50.675 ;
        RECT 51.77 49.655 52.03 49.915 ;
        RECT 51.77 48.895 52.03 49.155 ;
        RECT 51.77 48.135 52.03 48.395 ;
        RECT 51.77 47.375 52.03 47.635 ;
        RECT 51.77 46.615 52.03 46.875 ;
        RECT 51.77 45.855 52.03 46.115 ;
        RECT 51.77 45.095 52.03 45.355 ;
        RECT 51.77 44.335 52.03 44.595 ;
        RECT 51.77 43.575 52.03 43.835 ;
        RECT 51.77 42.815 52.03 43.075 ;
        RECT 51.77 42.055 52.03 42.315 ;
        RECT 51.77 41.295 52.03 41.555 ;
        RECT 51.77 40.535 52.03 40.795 ;
        RECT 51.77 39.775 52.03 40.035 ;
        RECT 51.77 39.015 52.03 39.275 ;
        RECT 51.77 38.255 52.03 38.515 ;
        RECT 51.77 37.495 52.03 37.755 ;
        RECT 51.77 36.735 52.03 36.995 ;
        RECT 52.53 58.775 52.79 59.035 ;
        RECT 52.53 58.015 52.79 58.275 ;
        RECT 52.53 57.255 52.79 57.515 ;
        RECT 52.53 56.495 52.79 56.755 ;
        RECT 52.53 55.735 52.79 55.995 ;
        RECT 52.53 54.975 52.79 55.235 ;
        RECT 52.53 54.215 52.79 54.475 ;
        RECT 52.53 53.455 52.79 53.715 ;
        RECT 52.53 52.695 52.79 52.955 ;
        RECT 52.53 51.935 52.79 52.195 ;
        RECT 52.53 51.175 52.79 51.435 ;
        RECT 52.53 50.415 52.79 50.675 ;
        RECT 52.53 49.655 52.79 49.915 ;
        RECT 52.53 48.895 52.79 49.155 ;
        RECT 52.53 48.135 52.79 48.395 ;
        RECT 52.53 47.375 52.79 47.635 ;
        RECT 52.53 46.615 52.79 46.875 ;
        RECT 52.53 45.855 52.79 46.115 ;
        RECT 52.53 45.095 52.79 45.355 ;
        RECT 52.53 44.335 52.79 44.595 ;
        RECT 52.53 43.575 52.79 43.835 ;
        RECT 52.53 42.815 52.79 43.075 ;
        RECT 52.53 42.055 52.79 42.315 ;
        RECT 52.53 41.295 52.79 41.555 ;
        RECT 52.53 40.535 52.79 40.795 ;
        RECT 52.53 39.775 52.79 40.035 ;
        RECT 52.53 39.015 52.79 39.275 ;
        RECT 52.53 38.255 52.79 38.515 ;
        RECT 52.53 37.495 52.79 37.755 ;
        RECT 52.53 36.735 52.79 36.995 ;
        RECT 53.29 58.775 53.55 59.035 ;
        RECT 53.29 58.015 53.55 58.275 ;
        RECT 53.29 57.255 53.55 57.515 ;
        RECT 53.29 56.495 53.55 56.755 ;
        RECT 53.29 55.735 53.55 55.995 ;
        RECT 53.29 54.975 53.55 55.235 ;
        RECT 53.29 54.215 53.55 54.475 ;
        RECT 53.29 53.455 53.55 53.715 ;
        RECT 53.29 52.695 53.55 52.955 ;
        RECT 53.29 51.935 53.55 52.195 ;
        RECT 53.29 51.175 53.55 51.435 ;
        RECT 53.29 50.415 53.55 50.675 ;
        RECT 53.29 49.655 53.55 49.915 ;
        RECT 53.29 48.895 53.55 49.155 ;
        RECT 53.29 48.135 53.55 48.395 ;
        RECT 53.29 47.375 53.55 47.635 ;
        RECT 53.29 46.615 53.55 46.875 ;
        RECT 53.29 45.855 53.55 46.115 ;
        RECT 53.29 45.095 53.55 45.355 ;
        RECT 53.29 44.335 53.55 44.595 ;
        RECT 53.29 43.575 53.55 43.835 ;
        RECT 53.29 42.815 53.55 43.075 ;
        RECT 53.29 42.055 53.55 42.315 ;
        RECT 53.29 41.295 53.55 41.555 ;
        RECT 53.29 40.535 53.55 40.795 ;
        RECT 53.29 39.775 53.55 40.035 ;
        RECT 53.29 39.015 53.55 39.275 ;
        RECT 53.29 38.255 53.55 38.515 ;
        RECT 53.29 37.495 53.55 37.755 ;
        RECT 53.29 36.735 53.55 36.995 ;
        RECT 54.05 58.775 54.31 59.035 ;
        RECT 54.05 58.015 54.31 58.275 ;
        RECT 54.05 57.255 54.31 57.515 ;
        RECT 54.05 56.495 54.31 56.755 ;
        RECT 54.05 55.735 54.31 55.995 ;
        RECT 54.05 54.975 54.31 55.235 ;
        RECT 54.05 54.215 54.31 54.475 ;
        RECT 54.05 53.455 54.31 53.715 ;
        RECT 54.05 52.695 54.31 52.955 ;
        RECT 54.05 51.935 54.31 52.195 ;
        RECT 54.05 51.175 54.31 51.435 ;
        RECT 54.05 50.415 54.31 50.675 ;
        RECT 54.05 49.655 54.31 49.915 ;
        RECT 54.05 48.895 54.31 49.155 ;
        RECT 54.05 48.135 54.31 48.395 ;
        RECT 54.05 47.375 54.31 47.635 ;
        RECT 54.05 46.615 54.31 46.875 ;
        RECT 54.05 45.855 54.31 46.115 ;
        RECT 54.05 45.095 54.31 45.355 ;
        RECT 54.05 44.335 54.31 44.595 ;
        RECT 54.05 43.575 54.31 43.835 ;
        RECT 54.05 42.815 54.31 43.075 ;
        RECT 54.05 42.055 54.31 42.315 ;
        RECT 54.05 41.295 54.31 41.555 ;
        RECT 54.05 40.535 54.31 40.795 ;
        RECT 54.05 39.775 54.31 40.035 ;
        RECT 54.05 39.015 54.31 39.275 ;
        RECT 54.05 38.255 54.31 38.515 ;
        RECT 54.05 37.495 54.31 37.755 ;
        RECT 54.05 36.735 54.31 36.995 ;
        RECT 54.81 58.775 55.07 59.035 ;
        RECT 54.81 58.015 55.07 58.275 ;
        RECT 54.81 57.255 55.07 57.515 ;
        RECT 54.81 56.495 55.07 56.755 ;
        RECT 54.81 55.735 55.07 55.995 ;
        RECT 54.81 54.975 55.07 55.235 ;
        RECT 54.81 54.215 55.07 54.475 ;
        RECT 54.81 53.455 55.07 53.715 ;
        RECT 54.81 52.695 55.07 52.955 ;
        RECT 54.81 51.935 55.07 52.195 ;
        RECT 54.81 51.175 55.07 51.435 ;
        RECT 54.81 50.415 55.07 50.675 ;
        RECT 54.81 49.655 55.07 49.915 ;
        RECT 54.81 48.895 55.07 49.155 ;
        RECT 54.81 48.135 55.07 48.395 ;
        RECT 54.81 47.375 55.07 47.635 ;
        RECT 54.81 46.615 55.07 46.875 ;
        RECT 54.81 45.855 55.07 46.115 ;
        RECT 54.81 45.095 55.07 45.355 ;
        RECT 54.81 44.335 55.07 44.595 ;
        RECT 4.65 58.775 4.91 59.035 ;
        RECT 4.65 58.015 4.91 58.275 ;
        RECT 4.65 57.255 4.91 57.515 ;
        RECT 4.65 56.495 4.91 56.755 ;
        RECT 4.65 55.735 4.91 55.995 ;
        RECT 4.65 54.975 4.91 55.235 ;
        RECT 4.65 54.215 4.91 54.475 ;
        RECT 4.65 53.455 4.91 53.715 ;
        RECT 4.65 52.695 4.91 52.955 ;
        RECT 4.65 51.935 4.91 52.195 ;
        RECT 4.65 51.175 4.91 51.435 ;
        RECT 4.65 50.415 4.91 50.675 ;
        RECT 4.65 49.655 4.91 49.915 ;
        RECT 4.65 48.895 4.91 49.155 ;
        RECT 4.65 48.135 4.91 48.395 ;
        RECT 4.65 47.375 4.91 47.635 ;
        RECT 4.65 46.615 4.91 46.875 ;
        RECT 4.65 45.855 4.91 46.115 ;
        RECT 4.65 45.095 4.91 45.355 ;
        RECT 4.65 44.335 4.91 44.595 ;
        RECT 4.65 43.575 4.91 43.835 ;
        RECT 4.65 42.815 4.91 43.075 ;
        RECT 4.65 42.055 4.91 42.315 ;
        RECT 4.65 41.295 4.91 41.555 ;
        RECT 4.65 40.535 4.91 40.795 ;
        RECT 4.65 39.775 4.91 40.035 ;
        RECT 4.65 39.015 4.91 39.275 ;
        RECT 4.65 38.255 4.91 38.515 ;
        RECT 4.65 37.495 4.91 37.755 ;
        RECT 4.65 36.735 4.91 36.995 ;
        RECT 5.41 58.775 5.67 59.035 ;
        RECT 5.41 58.015 5.67 58.275 ;
        RECT 5.41 57.255 5.67 57.515 ;
        RECT 5.41 56.495 5.67 56.755 ;
        RECT 5.41 55.735 5.67 55.995 ;
        RECT 5.41 54.975 5.67 55.235 ;
        RECT 5.41 54.215 5.67 54.475 ;
        RECT 5.41 53.455 5.67 53.715 ;
        RECT 5.41 52.695 5.67 52.955 ;
        RECT 5.41 51.935 5.67 52.195 ;
        RECT 5.41 51.175 5.67 51.435 ;
        RECT 5.41 50.415 5.67 50.675 ;
        RECT 5.41 49.655 5.67 49.915 ;
        RECT 5.41 48.895 5.67 49.155 ;
        RECT 5.41 48.135 5.67 48.395 ;
        RECT 5.41 47.375 5.67 47.635 ;
        RECT 5.41 46.615 5.67 46.875 ;
        RECT 5.41 45.855 5.67 46.115 ;
        RECT 5.41 45.095 5.67 45.355 ;
        RECT 5.41 44.335 5.67 44.595 ;
        RECT 5.41 43.575 5.67 43.835 ;
        RECT 5.41 42.815 5.67 43.075 ;
        RECT 5.41 42.055 5.67 42.315 ;
        RECT 5.41 41.295 5.67 41.555 ;
        RECT 5.41 40.535 5.67 40.795 ;
        RECT 5.41 39.775 5.67 40.035 ;
        RECT 5.41 39.015 5.67 39.275 ;
        RECT 5.41 38.255 5.67 38.515 ;
        RECT 5.41 37.495 5.67 37.755 ;
        RECT 5.41 36.735 5.67 36.995 ;
        RECT 6.17 58.775 6.43 59.035 ;
        RECT 6.17 58.015 6.43 58.275 ;
        RECT 6.17 57.255 6.43 57.515 ;
        RECT 6.17 56.495 6.43 56.755 ;
        RECT 6.17 55.735 6.43 55.995 ;
        RECT 6.17 54.975 6.43 55.235 ;
        RECT 6.17 54.215 6.43 54.475 ;
        RECT 6.17 53.455 6.43 53.715 ;
        RECT 6.17 52.695 6.43 52.955 ;
        RECT 6.17 51.935 6.43 52.195 ;
        RECT 6.17 51.175 6.43 51.435 ;
        RECT 6.17 50.415 6.43 50.675 ;
        RECT 6.17 49.655 6.43 49.915 ;
        RECT 6.17 48.895 6.43 49.155 ;
        RECT 6.17 48.135 6.43 48.395 ;
        RECT 6.17 47.375 6.43 47.635 ;
        RECT 6.17 46.615 6.43 46.875 ;
        RECT 6.17 45.855 6.43 46.115 ;
        RECT 6.17 45.095 6.43 45.355 ;
        RECT 6.17 44.335 6.43 44.595 ;
        RECT 6.17 43.575 6.43 43.835 ;
        RECT 6.17 42.815 6.43 43.075 ;
        RECT 6.17 42.055 6.43 42.315 ;
        RECT 6.17 41.295 6.43 41.555 ;
        RECT 6.17 40.535 6.43 40.795 ;
        RECT 6.17 39.775 6.43 40.035 ;
        RECT 6.17 39.015 6.43 39.275 ;
        RECT 6.17 38.255 6.43 38.515 ;
        RECT 6.17 37.495 6.43 37.755 ;
        RECT 6.17 36.735 6.43 36.995 ;
        RECT 6.93 58.775 7.19 59.035 ;
        RECT 6.93 58.015 7.19 58.275 ;
        RECT 6.93 57.255 7.19 57.515 ;
        RECT 6.93 56.495 7.19 56.755 ;
        RECT 6.93 55.735 7.19 55.995 ;
        RECT 6.93 54.975 7.19 55.235 ;
        RECT 6.93 54.215 7.19 54.475 ;
        RECT 6.93 53.455 7.19 53.715 ;
        RECT 6.93 52.695 7.19 52.955 ;
        RECT 6.93 51.935 7.19 52.195 ;
        RECT 6.93 51.175 7.19 51.435 ;
        RECT 6.93 50.415 7.19 50.675 ;
        RECT 6.93 49.655 7.19 49.915 ;
        RECT 6.93 48.895 7.19 49.155 ;
        RECT 6.93 48.135 7.19 48.395 ;
        RECT 6.93 47.375 7.19 47.635 ;
        RECT 6.93 46.615 7.19 46.875 ;
        RECT 6.93 45.855 7.19 46.115 ;
        RECT 6.93 45.095 7.19 45.355 ;
        RECT 6.93 44.335 7.19 44.595 ;
        RECT 6.93 43.575 7.19 43.835 ;
        RECT 6.93 42.815 7.19 43.075 ;
        RECT 6.93 42.055 7.19 42.315 ;
        RECT 6.93 41.295 7.19 41.555 ;
        RECT 6.93 40.535 7.19 40.795 ;
        RECT 6.93 39.775 7.19 40.035 ;
        RECT 6.93 39.015 7.19 39.275 ;
        RECT 6.93 38.255 7.19 38.515 ;
        RECT 6.93 37.495 7.19 37.755 ;
        RECT 6.93 36.735 7.19 36.995 ;
        RECT 7.69 58.775 7.95 59.035 ;
        RECT 7.69 58.015 7.95 58.275 ;
        RECT 7.69 57.255 7.95 57.515 ;
        RECT 7.69 56.495 7.95 56.755 ;
        RECT 7.69 55.735 7.95 55.995 ;
        RECT 7.69 54.975 7.95 55.235 ;
        RECT 7.69 54.215 7.95 54.475 ;
        RECT 7.69 53.455 7.95 53.715 ;
        RECT 7.69 52.695 7.95 52.955 ;
        RECT 7.69 51.935 7.95 52.195 ;
        RECT 7.69 51.175 7.95 51.435 ;
        RECT 7.69 50.415 7.95 50.675 ;
        RECT 7.69 49.655 7.95 49.915 ;
        RECT 7.69 48.895 7.95 49.155 ;
        RECT 7.69 48.135 7.95 48.395 ;
        RECT 7.69 47.375 7.95 47.635 ;
        RECT 7.69 46.615 7.95 46.875 ;
        RECT 7.69 45.855 7.95 46.115 ;
        RECT 7.69 45.095 7.95 45.355 ;
        RECT 7.69 44.335 7.95 44.595 ;
        RECT 7.69 43.575 7.95 43.835 ;
        RECT 7.69 42.815 7.95 43.075 ;
        RECT 7.69 42.055 7.95 42.315 ;
        RECT 7.69 41.295 7.95 41.555 ;
        RECT 7.69 40.535 7.95 40.795 ;
        RECT 7.69 39.775 7.95 40.035 ;
        RECT 7.69 39.015 7.95 39.275 ;
        RECT 7.69 38.255 7.95 38.515 ;
        RECT 7.69 37.495 7.95 37.755 ;
        RECT 7.69 36.735 7.95 36.995 ;
        RECT 8.45 58.775 8.71 59.035 ;
        RECT 8.45 58.015 8.71 58.275 ;
        RECT 8.45 57.255 8.71 57.515 ;
        RECT 8.45 56.495 8.71 56.755 ;
        RECT 8.45 55.735 8.71 55.995 ;
        RECT 8.45 54.975 8.71 55.235 ;
        RECT 8.45 54.215 8.71 54.475 ;
        RECT 8.45 53.455 8.71 53.715 ;
        RECT 8.45 52.695 8.71 52.955 ;
        RECT 8.45 51.935 8.71 52.195 ;
        RECT 8.45 51.175 8.71 51.435 ;
        RECT 8.45 50.415 8.71 50.675 ;
        RECT 8.45 49.655 8.71 49.915 ;
        RECT 8.45 48.895 8.71 49.155 ;
        RECT 8.45 48.135 8.71 48.395 ;
        RECT 8.45 47.375 8.71 47.635 ;
        RECT 8.45 46.615 8.71 46.875 ;
        RECT 8.45 45.855 8.71 46.115 ;
        RECT 8.45 45.095 8.71 45.355 ;
        RECT 8.45 44.335 8.71 44.595 ;
        RECT 8.45 43.575 8.71 43.835 ;
        RECT 8.45 42.815 8.71 43.075 ;
        RECT 8.45 42.055 8.71 42.315 ;
        RECT 8.45 41.295 8.71 41.555 ;
        RECT 8.45 40.535 8.71 40.795 ;
        RECT 8.45 39.775 8.71 40.035 ;
        RECT 8.45 39.015 8.71 39.275 ;
        RECT 8.45 38.255 8.71 38.515 ;
        RECT 8.45 37.495 8.71 37.755 ;
        RECT 8.45 36.735 8.71 36.995 ;
        RECT 9.21 58.775 9.47 59.035 ;
        RECT 9.21 58.015 9.47 58.275 ;
        RECT 9.21 57.255 9.47 57.515 ;
        RECT 9.21 56.495 9.47 56.755 ;
        RECT 9.21 55.735 9.47 55.995 ;
        RECT 9.21 54.975 9.47 55.235 ;
        RECT 9.21 54.215 9.47 54.475 ;
        RECT 9.21 53.455 9.47 53.715 ;
        RECT 9.21 52.695 9.47 52.955 ;
        RECT 9.21 51.935 9.47 52.195 ;
        RECT 9.21 51.175 9.47 51.435 ;
        RECT 9.21 50.415 9.47 50.675 ;
        RECT 9.21 49.655 9.47 49.915 ;
        RECT 9.21 48.895 9.47 49.155 ;
        RECT 9.21 48.135 9.47 48.395 ;
        RECT 9.21 47.375 9.47 47.635 ;
        RECT 9.21 46.615 9.47 46.875 ;
        RECT 9.21 45.855 9.47 46.115 ;
        RECT 9.21 45.095 9.47 45.355 ;
        RECT 9.21 44.335 9.47 44.595 ;
        RECT 9.21 43.575 9.47 43.835 ;
        RECT 9.21 42.815 9.47 43.075 ;
        RECT 9.21 42.055 9.47 42.315 ;
        RECT 9.21 41.295 9.47 41.555 ;
        RECT 9.21 40.535 9.47 40.795 ;
        RECT 9.21 39.775 9.47 40.035 ;
        RECT 9.21 39.015 9.47 39.275 ;
        RECT 9.21 38.255 9.47 38.515 ;
        RECT 9.21 37.495 9.47 37.755 ;
        RECT 9.21 36.735 9.47 36.995 ;
        RECT 9.97 58.775 10.23 59.035 ;
        RECT 9.97 58.015 10.23 58.275 ;
        RECT 9.97 57.255 10.23 57.515 ;
        RECT 9.97 56.495 10.23 56.755 ;
        RECT 9.97 55.735 10.23 55.995 ;
        RECT 9.97 54.975 10.23 55.235 ;
        RECT 9.97 54.215 10.23 54.475 ;
        RECT 9.97 53.455 10.23 53.715 ;
        RECT 9.97 52.695 10.23 52.955 ;
        RECT 9.97 51.935 10.23 52.195 ;
        RECT 9.97 51.175 10.23 51.435 ;
        RECT 9.97 50.415 10.23 50.675 ;
        RECT 9.97 49.655 10.23 49.915 ;
        RECT 9.97 48.895 10.23 49.155 ;
        RECT 9.97 48.135 10.23 48.395 ;
        RECT 9.97 47.375 10.23 47.635 ;
        RECT 9.97 46.615 10.23 46.875 ;
        RECT 9.97 45.855 10.23 46.115 ;
        RECT 9.97 45.095 10.23 45.355 ;
        RECT 9.97 44.335 10.23 44.595 ;
        RECT 9.97 43.575 10.23 43.835 ;
        RECT 9.97 42.815 10.23 43.075 ;
        RECT 9.97 42.055 10.23 42.315 ;
        RECT 9.97 41.295 10.23 41.555 ;
        RECT 9.97 40.535 10.23 40.795 ;
        RECT 9.97 39.775 10.23 40.035 ;
        RECT 9.97 39.015 10.23 39.275 ;
        RECT 9.97 38.255 10.23 38.515 ;
        RECT 9.97 37.495 10.23 37.755 ;
        RECT 9.97 36.735 10.23 36.995 ;
        RECT 10.73 58.775 10.99 59.035 ;
        RECT 10.73 58.015 10.99 58.275 ;
        RECT 10.73 57.255 10.99 57.515 ;
        RECT 10.73 56.495 10.99 56.755 ;
        RECT 10.73 55.735 10.99 55.995 ;
        RECT 10.73 54.975 10.99 55.235 ;
        RECT 10.73 54.215 10.99 54.475 ;
        RECT 10.73 53.455 10.99 53.715 ;
        RECT 10.73 52.695 10.99 52.955 ;
        RECT 10.73 51.935 10.99 52.195 ;
        RECT 10.73 51.175 10.99 51.435 ;
        RECT 10.73 50.415 10.99 50.675 ;
        RECT 10.73 49.655 10.99 49.915 ;
        RECT 10.73 48.895 10.99 49.155 ;
        RECT 10.73 48.135 10.99 48.395 ;
        RECT 10.73 47.375 10.99 47.635 ;
        RECT 10.73 46.615 10.99 46.875 ;
        RECT 10.73 45.855 10.99 46.115 ;
        RECT 10.73 45.095 10.99 45.355 ;
        RECT 10.73 44.335 10.99 44.595 ;
        RECT 10.73 43.575 10.99 43.835 ;
        RECT 10.73 42.815 10.99 43.075 ;
        RECT 10.73 42.055 10.99 42.315 ;
        RECT 10.73 41.295 10.99 41.555 ;
        RECT 10.73 40.535 10.99 40.795 ;
        RECT 10.73 39.775 10.99 40.035 ;
        RECT 10.73 39.015 10.99 39.275 ;
        RECT 10.73 38.255 10.99 38.515 ;
        RECT 10.73 37.495 10.99 37.755 ;
        RECT 10.73 36.735 10.99 36.995 ;
        RECT 11.49 58.775 11.75 59.035 ;
        RECT 11.49 58.015 11.75 58.275 ;
        RECT 11.49 57.255 11.75 57.515 ;
        RECT 11.49 56.495 11.75 56.755 ;
        RECT 11.49 55.735 11.75 55.995 ;
        RECT 11.49 54.975 11.75 55.235 ;
        RECT 11.49 54.215 11.75 54.475 ;
        RECT 11.49 53.455 11.75 53.715 ;
        RECT 11.49 52.695 11.75 52.955 ;
        RECT 11.49 51.935 11.75 52.195 ;
        RECT 11.49 51.175 11.75 51.435 ;
        RECT 11.49 50.415 11.75 50.675 ;
        RECT 11.49 49.655 11.75 49.915 ;
        RECT 11.49 48.895 11.75 49.155 ;
        RECT 11.49 48.135 11.75 48.395 ;
        RECT 11.49 47.375 11.75 47.635 ;
        RECT 11.49 46.615 11.75 46.875 ;
        RECT 11.49 45.855 11.75 46.115 ;
        RECT 11.49 45.095 11.75 45.355 ;
        RECT 11.49 44.335 11.75 44.595 ;
        RECT 11.49 43.575 11.75 43.835 ;
        RECT 11.49 42.815 11.75 43.075 ;
        RECT 11.49 42.055 11.75 42.315 ;
        RECT 11.49 41.295 11.75 41.555 ;
        RECT 11.49 40.535 11.75 40.795 ;
        RECT 11.49 39.775 11.75 40.035 ;
        RECT 11.49 39.015 11.75 39.275 ;
        RECT 11.49 38.255 11.75 38.515 ;
        RECT 11.49 37.495 11.75 37.755 ;
        RECT 11.49 36.735 11.75 36.995 ;
        RECT 12.25 58.775 12.51 59.035 ;
        RECT 12.25 58.015 12.51 58.275 ;
        RECT 12.25 57.255 12.51 57.515 ;
        RECT 12.25 56.495 12.51 56.755 ;
        RECT 12.25 55.735 12.51 55.995 ;
        RECT 12.25 54.975 12.51 55.235 ;
        RECT 12.25 54.215 12.51 54.475 ;
        RECT 12.25 53.455 12.51 53.715 ;
        RECT 12.25 52.695 12.51 52.955 ;
        RECT 12.25 51.935 12.51 52.195 ;
        RECT 12.25 51.175 12.51 51.435 ;
        RECT 12.25 50.415 12.51 50.675 ;
        RECT 12.25 49.655 12.51 49.915 ;
        RECT 12.25 48.895 12.51 49.155 ;
        RECT 12.25 48.135 12.51 48.395 ;
        RECT 12.25 47.375 12.51 47.635 ;
        RECT 12.25 46.615 12.51 46.875 ;
        RECT 12.25 45.855 12.51 46.115 ;
        RECT 12.25 45.095 12.51 45.355 ;
        RECT 12.25 44.335 12.51 44.595 ;
        RECT 12.25 43.575 12.51 43.835 ;
        RECT 12.25 42.815 12.51 43.075 ;
        RECT 12.25 42.055 12.51 42.315 ;
        RECT 12.25 41.295 12.51 41.555 ;
        RECT 12.25 40.535 12.51 40.795 ;
        RECT 12.25 39.775 12.51 40.035 ;
        RECT 12.25 39.015 12.51 39.275 ;
        RECT 12.25 38.255 12.51 38.515 ;
        RECT 12.25 37.495 12.51 37.755 ;
        RECT 12.25 36.735 12.51 36.995 ;
        RECT 13.01 58.775 13.27 59.035 ;
        RECT 13.01 58.015 13.27 58.275 ;
        RECT 13.01 57.255 13.27 57.515 ;
        RECT 13.01 56.495 13.27 56.755 ;
        RECT 13.01 55.735 13.27 55.995 ;
        RECT 13.01 54.975 13.27 55.235 ;
        RECT 13.01 54.215 13.27 54.475 ;
        RECT 13.01 53.455 13.27 53.715 ;
        RECT 13.01 52.695 13.27 52.955 ;
        RECT 13.01 51.935 13.27 52.195 ;
        RECT 13.01 51.175 13.27 51.435 ;
        RECT 13.01 50.415 13.27 50.675 ;
        RECT 13.01 49.655 13.27 49.915 ;
        RECT 13.01 48.895 13.27 49.155 ;
        RECT 13.01 48.135 13.27 48.395 ;
        RECT 13.01 47.375 13.27 47.635 ;
        RECT 13.01 46.615 13.27 46.875 ;
        RECT 13.01 45.855 13.27 46.115 ;
        RECT 13.01 45.095 13.27 45.355 ;
        RECT 13.01 44.335 13.27 44.595 ;
        RECT 13.01 43.575 13.27 43.835 ;
        RECT 13.01 42.815 13.27 43.075 ;
        RECT 13.01 42.055 13.27 42.315 ;
        RECT 13.01 41.295 13.27 41.555 ;
        RECT 13.01 40.535 13.27 40.795 ;
        RECT 13.01 39.775 13.27 40.035 ;
        RECT 13.01 39.015 13.27 39.275 ;
        RECT 13.01 38.255 13.27 38.515 ;
        RECT 13.01 37.495 13.27 37.755 ;
        RECT 13.01 36.735 13.27 36.995 ;
        RECT 13.77 58.775 14.03 59.035 ;
        RECT 13.77 58.015 14.03 58.275 ;
        RECT 13.77 57.255 14.03 57.515 ;
        RECT 13.77 56.495 14.03 56.755 ;
        RECT 13.77 55.735 14.03 55.995 ;
        RECT 13.77 54.975 14.03 55.235 ;
        RECT 13.77 54.215 14.03 54.475 ;
        RECT 13.77 53.455 14.03 53.715 ;
        RECT 13.77 52.695 14.03 52.955 ;
        RECT 13.77 51.935 14.03 52.195 ;
        RECT 13.77 51.175 14.03 51.435 ;
        RECT 13.77 50.415 14.03 50.675 ;
        RECT 13.77 49.655 14.03 49.915 ;
        RECT 13.77 48.895 14.03 49.155 ;
        RECT 13.77 48.135 14.03 48.395 ;
        RECT 13.77 47.375 14.03 47.635 ;
        RECT 13.77 46.615 14.03 46.875 ;
        RECT 13.77 45.855 14.03 46.115 ;
        RECT 13.77 45.095 14.03 45.355 ;
        RECT 13.77 44.335 14.03 44.595 ;
        RECT 13.77 43.575 14.03 43.835 ;
        RECT 13.77 42.815 14.03 43.075 ;
        RECT 13.77 42.055 14.03 42.315 ;
        RECT 13.77 41.295 14.03 41.555 ;
        RECT 13.77 40.535 14.03 40.795 ;
        RECT 13.77 39.775 14.03 40.035 ;
        RECT 13.77 39.015 14.03 39.275 ;
        RECT 13.77 38.255 14.03 38.515 ;
        RECT 13.77 37.495 14.03 37.755 ;
        RECT 13.77 36.735 14.03 36.995 ;
        RECT 14.53 58.775 14.79 59.035 ;
        RECT 14.53 58.015 14.79 58.275 ;
        RECT 14.53 57.255 14.79 57.515 ;
        RECT 14.53 56.495 14.79 56.755 ;
        RECT 14.53 55.735 14.79 55.995 ;
        RECT 14.53 54.975 14.79 55.235 ;
        RECT 14.53 54.215 14.79 54.475 ;
        RECT 14.53 53.455 14.79 53.715 ;
        RECT 14.53 52.695 14.79 52.955 ;
        RECT 14.53 51.935 14.79 52.195 ;
        RECT 14.53 51.175 14.79 51.435 ;
        RECT 14.53 50.415 14.79 50.675 ;
        RECT 14.53 49.655 14.79 49.915 ;
        RECT 14.53 48.895 14.79 49.155 ;
        RECT 14.53 48.135 14.79 48.395 ;
        RECT 14.53 47.375 14.79 47.635 ;
        RECT 14.53 46.615 14.79 46.875 ;
        RECT 14.53 45.855 14.79 46.115 ;
        RECT 14.53 45.095 14.79 45.355 ;
        RECT 14.53 44.335 14.79 44.595 ;
        RECT 14.53 43.575 14.79 43.835 ;
        RECT 14.53 42.815 14.79 43.075 ;
        RECT 14.53 42.055 14.79 42.315 ;
        RECT 14.53 41.295 14.79 41.555 ;
        RECT 14.53 40.535 14.79 40.795 ;
        RECT 14.53 39.775 14.79 40.035 ;
        RECT 14.53 39.015 14.79 39.275 ;
        RECT 14.53 38.255 14.79 38.515 ;
        RECT 14.53 37.495 14.79 37.755 ;
        RECT 14.53 36.735 14.79 36.995 ;
        RECT 15.29 58.775 15.55 59.035 ;
        RECT 15.29 58.015 15.55 58.275 ;
        RECT 15.29 57.255 15.55 57.515 ;
        RECT 15.29 56.495 15.55 56.755 ;
        RECT 15.29 55.735 15.55 55.995 ;
        RECT 15.29 54.975 15.55 55.235 ;
        RECT 15.29 54.215 15.55 54.475 ;
        RECT 15.29 53.455 15.55 53.715 ;
        RECT 15.29 52.695 15.55 52.955 ;
        RECT 15.29 51.935 15.55 52.195 ;
        RECT 15.29 51.175 15.55 51.435 ;
        RECT 15.29 50.415 15.55 50.675 ;
        RECT 15.29 49.655 15.55 49.915 ;
        RECT 15.29 48.895 15.55 49.155 ;
        RECT 15.29 48.135 15.55 48.395 ;
        RECT 15.29 47.375 15.55 47.635 ;
        RECT 15.29 46.615 15.55 46.875 ;
        RECT 15.29 45.855 15.55 46.115 ;
        RECT 15.29 45.095 15.55 45.355 ;
        RECT 15.29 44.335 15.55 44.595 ;
        RECT 15.29 43.575 15.55 43.835 ;
        RECT 15.29 42.815 15.55 43.075 ;
        RECT 15.29 42.055 15.55 42.315 ;
        RECT 15.29 41.295 15.55 41.555 ;
        RECT 15.29 40.535 15.55 40.795 ;
        RECT 15.29 39.775 15.55 40.035 ;
        RECT 15.29 39.015 15.55 39.275 ;
        RECT 15.29 38.255 15.55 38.515 ;
        RECT 15.29 37.495 15.55 37.755 ;
        RECT 15.29 36.735 15.55 36.995 ;
        RECT 16.05 58.775 16.31 59.035 ;
        RECT 16.05 58.015 16.31 58.275 ;
        RECT 16.05 57.255 16.31 57.515 ;
        RECT 16.05 56.495 16.31 56.755 ;
        RECT 16.05 55.735 16.31 55.995 ;
        RECT 16.05 54.975 16.31 55.235 ;
        RECT 16.05 54.215 16.31 54.475 ;
        RECT 16.05 53.455 16.31 53.715 ;
        RECT 16.05 52.695 16.31 52.955 ;
        RECT 16.05 51.935 16.31 52.195 ;
        RECT 16.05 51.175 16.31 51.435 ;
        RECT 16.05 50.415 16.31 50.675 ;
        RECT 16.05 49.655 16.31 49.915 ;
        RECT 16.05 48.895 16.31 49.155 ;
        RECT 16.05 48.135 16.31 48.395 ;
        RECT 16.05 47.375 16.31 47.635 ;
        RECT 16.05 46.615 16.31 46.875 ;
        RECT 16.05 45.855 16.31 46.115 ;
        RECT 16.05 45.095 16.31 45.355 ;
        RECT 16.05 44.335 16.31 44.595 ;
        RECT 16.05 43.575 16.31 43.835 ;
        RECT 16.05 42.815 16.31 43.075 ;
        RECT 16.05 42.055 16.31 42.315 ;
        RECT 16.05 41.295 16.31 41.555 ;
        RECT 16.05 40.535 16.31 40.795 ;
        RECT 16.05 39.775 16.31 40.035 ;
        RECT 16.05 39.015 16.31 39.275 ;
        RECT 16.05 38.255 16.31 38.515 ;
        RECT 16.05 37.495 16.31 37.755 ;
        RECT 16.05 36.735 16.31 36.995 ;
        RECT 16.81 58.775 17.07 59.035 ;
        RECT 16.81 58.015 17.07 58.275 ;
        RECT 16.81 57.255 17.07 57.515 ;
        RECT 16.81 56.495 17.07 56.755 ;
        RECT 16.81 55.735 17.07 55.995 ;
        RECT 16.81 54.975 17.07 55.235 ;
        RECT 16.81 54.215 17.07 54.475 ;
        RECT 16.81 53.455 17.07 53.715 ;
        RECT 16.81 52.695 17.07 52.955 ;
        RECT 16.81 51.935 17.07 52.195 ;
        RECT 16.81 51.175 17.07 51.435 ;
        RECT 16.81 50.415 17.07 50.675 ;
        RECT 16.81 49.655 17.07 49.915 ;
        RECT 16.81 48.895 17.07 49.155 ;
        RECT 16.81 48.135 17.07 48.395 ;
        RECT 16.81 47.375 17.07 47.635 ;
        RECT 16.81 46.615 17.07 46.875 ;
        RECT 16.81 45.855 17.07 46.115 ;
        RECT 16.81 45.095 17.07 45.355 ;
        RECT 16.81 44.335 17.07 44.595 ;
        RECT 16.81 43.575 17.07 43.835 ;
        RECT 16.81 42.815 17.07 43.075 ;
        RECT 16.81 42.055 17.07 42.315 ;
        RECT 16.81 41.295 17.07 41.555 ;
        RECT 16.81 40.535 17.07 40.795 ;
        RECT 16.81 39.775 17.07 40.035 ;
        RECT 16.81 39.015 17.07 39.275 ;
        RECT 16.81 38.255 17.07 38.515 ;
        RECT 16.81 37.495 17.07 37.755 ;
        RECT 16.81 36.735 17.07 36.995 ;
        RECT 17.57 58.775 17.83 59.035 ;
        RECT 17.57 58.015 17.83 58.275 ;
        RECT 17.57 57.255 17.83 57.515 ;
        RECT 17.57 56.495 17.83 56.755 ;
        RECT 17.57 55.735 17.83 55.995 ;
        RECT 17.57 54.975 17.83 55.235 ;
        RECT 17.57 54.215 17.83 54.475 ;
        RECT 17.57 53.455 17.83 53.715 ;
        RECT 17.57 52.695 17.83 52.955 ;
        RECT 17.57 51.935 17.83 52.195 ;
        RECT 17.57 51.175 17.83 51.435 ;
        RECT 17.57 50.415 17.83 50.675 ;
        RECT 17.57 49.655 17.83 49.915 ;
        RECT 17.57 48.895 17.83 49.155 ;
        RECT 17.57 48.135 17.83 48.395 ;
        RECT 17.57 47.375 17.83 47.635 ;
        RECT 17.57 46.615 17.83 46.875 ;
        RECT 17.57 45.855 17.83 46.115 ;
        RECT 17.57 45.095 17.83 45.355 ;
        RECT 17.57 44.335 17.83 44.595 ;
        RECT 17.57 43.575 17.83 43.835 ;
        RECT 17.57 42.815 17.83 43.075 ;
        RECT 17.57 42.055 17.83 42.315 ;
        RECT 17.57 41.295 17.83 41.555 ;
        RECT 17.57 40.535 17.83 40.795 ;
        RECT 17.57 39.775 17.83 40.035 ;
        RECT 17.57 39.015 17.83 39.275 ;
        RECT 17.57 38.255 17.83 38.515 ;
        RECT 17.57 37.495 17.83 37.755 ;
        RECT 17.57 36.735 17.83 36.995 ;
        RECT 18.33 58.775 18.59 59.035 ;
        RECT 18.33 58.015 18.59 58.275 ;
        RECT 18.33 57.255 18.59 57.515 ;
        RECT 18.33 56.495 18.59 56.755 ;
        RECT 18.33 55.735 18.59 55.995 ;
        RECT 18.33 54.975 18.59 55.235 ;
        RECT 18.33 54.215 18.59 54.475 ;
        RECT 18.33 53.455 18.59 53.715 ;
        RECT 18.33 52.695 18.59 52.955 ;
        RECT 18.33 51.935 18.59 52.195 ;
        RECT 18.33 51.175 18.59 51.435 ;
        RECT 18.33 50.415 18.59 50.675 ;
        RECT 18.33 49.655 18.59 49.915 ;
        RECT 18.33 48.895 18.59 49.155 ;
        RECT 18.33 48.135 18.59 48.395 ;
        RECT 18.33 47.375 18.59 47.635 ;
        RECT 18.33 46.615 18.59 46.875 ;
        RECT 18.33 45.855 18.59 46.115 ;
        RECT 18.33 45.095 18.59 45.355 ;
        RECT 18.33 44.335 18.59 44.595 ;
        RECT 18.33 43.575 18.59 43.835 ;
        RECT 18.33 42.815 18.59 43.075 ;
        RECT 18.33 42.055 18.59 42.315 ;
        RECT 18.33 41.295 18.59 41.555 ;
        RECT 18.33 40.535 18.59 40.795 ;
        RECT 18.33 39.775 18.59 40.035 ;
        RECT 18.33 39.015 18.59 39.275 ;
        RECT 18.33 38.255 18.59 38.515 ;
        RECT 18.33 37.495 18.59 37.755 ;
        RECT 18.33 36.735 18.59 36.995 ;
        RECT 19.09 58.775 19.35 59.035 ;
        RECT 19.09 58.015 19.35 58.275 ;
        RECT 19.09 57.255 19.35 57.515 ;
        RECT 19.09 56.495 19.35 56.755 ;
        RECT 19.09 55.735 19.35 55.995 ;
        RECT 19.09 54.975 19.35 55.235 ;
        RECT 19.09 54.215 19.35 54.475 ;
        RECT 19.09 53.455 19.35 53.715 ;
        RECT 19.09 52.695 19.35 52.955 ;
        RECT 19.09 51.935 19.35 52.195 ;
        RECT 19.09 51.175 19.35 51.435 ;
        RECT 19.09 50.415 19.35 50.675 ;
        RECT 19.09 49.655 19.35 49.915 ;
        RECT 19.09 48.895 19.35 49.155 ;
        RECT 19.09 48.135 19.35 48.395 ;
        RECT 19.09 47.375 19.35 47.635 ;
        RECT 19.09 46.615 19.35 46.875 ;
        RECT 19.09 45.855 19.35 46.115 ;
        RECT 19.09 45.095 19.35 45.355 ;
        RECT 19.09 44.335 19.35 44.595 ;
        RECT 19.09 43.575 19.35 43.835 ;
        RECT 19.09 42.815 19.35 43.075 ;
        RECT 19.09 42.055 19.35 42.315 ;
        RECT 19.09 41.295 19.35 41.555 ;
        RECT 19.09 40.535 19.35 40.795 ;
        RECT 19.09 39.775 19.35 40.035 ;
        RECT 19.09 39.015 19.35 39.275 ;
        RECT 19.09 38.255 19.35 38.515 ;
        RECT 19.09 37.495 19.35 37.755 ;
        RECT 19.09 36.735 19.35 36.995 ;
        RECT 19.85 58.775 20.11 59.035 ;
        RECT 19.85 58.015 20.11 58.275 ;
        RECT 19.85 57.255 20.11 57.515 ;
        RECT 19.85 56.495 20.11 56.755 ;
        RECT 19.85 55.735 20.11 55.995 ;
        RECT 19.85 54.975 20.11 55.235 ;
        RECT 19.85 54.215 20.11 54.475 ;
        RECT 19.85 53.455 20.11 53.715 ;
        RECT 19.85 52.695 20.11 52.955 ;
        RECT 19.85 51.935 20.11 52.195 ;
        RECT 19.85 51.175 20.11 51.435 ;
        RECT 19.85 50.415 20.11 50.675 ;
        RECT 19.85 49.655 20.11 49.915 ;
        RECT 19.85 48.895 20.11 49.155 ;
        RECT 19.85 48.135 20.11 48.395 ;
        RECT 19.85 47.375 20.11 47.635 ;
        RECT 19.85 46.615 20.11 46.875 ;
        RECT 19.85 45.855 20.11 46.115 ;
        RECT 19.85 45.095 20.11 45.355 ;
        RECT 19.85 44.335 20.11 44.595 ;
        RECT 19.85 43.575 20.11 43.835 ;
        RECT 19.85 42.815 20.11 43.075 ;
        RECT 19.85 42.055 20.11 42.315 ;
        RECT 19.85 41.295 20.11 41.555 ;
        RECT 19.85 40.535 20.11 40.795 ;
        RECT 19.85 39.775 20.11 40.035 ;
        RECT 19.85 39.015 20.11 39.275 ;
        RECT 19.85 38.255 20.11 38.515 ;
        RECT 19.85 37.495 20.11 37.755 ;
        RECT 19.85 36.735 20.11 36.995 ;
        RECT 20.61 58.775 20.87 59.035 ;
        RECT 20.61 58.015 20.87 58.275 ;
        RECT 20.61 57.255 20.87 57.515 ;
        RECT 20.61 56.495 20.87 56.755 ;
        RECT 20.61 55.735 20.87 55.995 ;
        RECT 20.61 54.975 20.87 55.235 ;
        RECT 20.61 54.215 20.87 54.475 ;
        RECT 20.61 53.455 20.87 53.715 ;
        RECT 20.61 52.695 20.87 52.955 ;
        RECT 20.61 51.935 20.87 52.195 ;
        RECT 20.61 51.175 20.87 51.435 ;
        RECT 20.61 50.415 20.87 50.675 ;
        RECT 20.61 49.655 20.87 49.915 ;
        RECT 20.61 48.895 20.87 49.155 ;
        RECT 20.61 48.135 20.87 48.395 ;
        RECT 20.61 47.375 20.87 47.635 ;
        RECT 20.61 46.615 20.87 46.875 ;
        RECT 20.61 45.855 20.87 46.115 ;
        RECT 20.61 45.095 20.87 45.355 ;
        RECT 20.61 44.335 20.87 44.595 ;
        RECT 20.61 43.575 20.87 43.835 ;
        RECT 20.61 42.815 20.87 43.075 ;
        RECT 20.61 42.055 20.87 42.315 ;
        RECT 20.61 41.295 20.87 41.555 ;
        RECT 20.61 40.535 20.87 40.795 ;
        RECT 20.61 39.775 20.87 40.035 ;
        RECT 20.61 39.015 20.87 39.275 ;
        RECT 20.61 38.255 20.87 38.515 ;
        RECT 20.61 37.495 20.87 37.755 ;
        RECT 20.61 36.735 20.87 36.995 ;
        RECT 21.37 58.775 21.63 59.035 ;
        RECT 21.37 58.015 21.63 58.275 ;
        RECT 21.37 57.255 21.63 57.515 ;
        RECT 21.37 56.495 21.63 56.755 ;
        RECT 21.37 55.735 21.63 55.995 ;
        RECT 21.37 54.975 21.63 55.235 ;
        RECT 21.37 54.215 21.63 54.475 ;
        RECT 21.37 53.455 21.63 53.715 ;
        RECT 21.37 52.695 21.63 52.955 ;
        RECT 21.37 51.935 21.63 52.195 ;
        RECT 21.37 51.175 21.63 51.435 ;
        RECT 21.37 50.415 21.63 50.675 ;
        RECT 21.37 49.655 21.63 49.915 ;
        RECT 21.37 48.895 21.63 49.155 ;
        RECT 21.37 48.135 21.63 48.395 ;
        RECT 21.37 47.375 21.63 47.635 ;
        RECT 21.37 46.615 21.63 46.875 ;
        RECT 21.37 45.855 21.63 46.115 ;
        RECT 21.37 45.095 21.63 45.355 ;
        RECT 21.37 44.335 21.63 44.595 ;
        RECT 21.37 43.575 21.63 43.835 ;
        RECT 21.37 42.815 21.63 43.075 ;
        RECT 21.37 42.055 21.63 42.315 ;
        RECT 21.37 41.295 21.63 41.555 ;
        RECT 21.37 40.535 21.63 40.795 ;
        RECT 21.37 39.775 21.63 40.035 ;
        RECT 21.37 39.015 21.63 39.275 ;
        RECT 21.37 38.255 21.63 38.515 ;
        RECT 21.37 37.495 21.63 37.755 ;
        RECT 21.37 36.735 21.63 36.995 ;
        RECT 22.13 58.775 22.39 59.035 ;
        RECT 22.13 58.015 22.39 58.275 ;
        RECT 22.13 57.255 22.39 57.515 ;
        RECT 22.13 56.495 22.39 56.755 ;
        RECT 22.13 55.735 22.39 55.995 ;
        RECT 22.13 54.975 22.39 55.235 ;
        RECT 22.13 54.215 22.39 54.475 ;
        RECT 22.13 53.455 22.39 53.715 ;
        RECT 22.13 52.695 22.39 52.955 ;
        RECT 22.13 51.935 22.39 52.195 ;
        RECT 22.13 51.175 22.39 51.435 ;
        RECT 22.13 50.415 22.39 50.675 ;
        RECT 22.13 49.655 22.39 49.915 ;
        RECT 22.13 48.895 22.39 49.155 ;
        RECT 22.13 48.135 22.39 48.395 ;
        RECT 22.13 47.375 22.39 47.635 ;
        RECT 22.13 46.615 22.39 46.875 ;
        RECT 22.13 45.855 22.39 46.115 ;
        RECT 22.13 45.095 22.39 45.355 ;
        RECT 22.13 44.335 22.39 44.595 ;
        RECT 22.13 43.575 22.39 43.835 ;
        RECT 22.13 42.815 22.39 43.075 ;
        RECT 22.13 42.055 22.39 42.315 ;
        RECT 22.13 41.295 22.39 41.555 ;
        RECT 22.13 40.535 22.39 40.795 ;
        RECT 22.13 39.775 22.39 40.035 ;
        RECT 22.13 39.015 22.39 39.275 ;
        RECT 22.13 38.255 22.39 38.515 ;
        RECT 22.13 37.495 22.39 37.755 ;
        RECT 22.13 36.735 22.39 36.995 ;
        RECT 22.89 58.775 23.15 59.035 ;
        RECT 22.89 58.015 23.15 58.275 ;
        RECT 22.89 57.255 23.15 57.515 ;
        RECT 22.89 56.495 23.15 56.755 ;
        RECT 22.89 55.735 23.15 55.995 ;
        RECT 22.89 54.975 23.15 55.235 ;
        RECT 22.89 54.215 23.15 54.475 ;
        RECT 22.89 53.455 23.15 53.715 ;
        RECT 22.89 52.695 23.15 52.955 ;
        RECT 22.89 51.935 23.15 52.195 ;
        RECT 22.89 51.175 23.15 51.435 ;
        RECT 22.89 50.415 23.15 50.675 ;
        RECT 22.89 49.655 23.15 49.915 ;
        RECT 22.89 48.895 23.15 49.155 ;
        RECT 22.89 48.135 23.15 48.395 ;
        RECT 22.89 47.375 23.15 47.635 ;
        RECT 22.89 46.615 23.15 46.875 ;
        RECT 22.89 45.855 23.15 46.115 ;
        RECT 22.89 45.095 23.15 45.355 ;
        RECT 22.89 44.335 23.15 44.595 ;
        RECT 22.89 43.575 23.15 43.835 ;
        RECT 22.89 42.815 23.15 43.075 ;
        RECT 22.89 42.055 23.15 42.315 ;
        RECT 22.89 41.295 23.15 41.555 ;
        RECT 22.89 40.535 23.15 40.795 ;
        RECT 22.89 39.775 23.15 40.035 ;
        RECT 22.89 39.015 23.15 39.275 ;
        RECT 22.89 38.255 23.15 38.515 ;
        RECT 22.89 37.495 23.15 37.755 ;
        RECT 22.89 36.735 23.15 36.995 ;
        RECT 23.65 58.775 23.91 59.035 ;
        RECT 23.65 58.015 23.91 58.275 ;
        RECT 23.65 57.255 23.91 57.515 ;
        RECT 23.65 56.495 23.91 56.755 ;
        RECT 23.65 55.735 23.91 55.995 ;
        RECT 23.65 54.975 23.91 55.235 ;
        RECT 23.65 54.215 23.91 54.475 ;
        RECT 23.65 53.455 23.91 53.715 ;
        RECT 23.65 52.695 23.91 52.955 ;
        RECT 23.65 51.935 23.91 52.195 ;
        RECT 23.65 51.175 23.91 51.435 ;
        RECT 23.65 50.415 23.91 50.675 ;
        RECT 23.65 49.655 23.91 49.915 ;
        RECT 23.65 48.895 23.91 49.155 ;
        RECT 23.65 48.135 23.91 48.395 ;
        RECT 23.65 47.375 23.91 47.635 ;
        RECT 23.65 46.615 23.91 46.875 ;
        RECT 23.65 45.855 23.91 46.115 ;
        RECT 23.65 45.095 23.91 45.355 ;
        RECT 23.65 44.335 23.91 44.595 ;
        RECT 23.65 43.575 23.91 43.835 ;
        RECT 23.65 42.815 23.91 43.075 ;
        RECT 23.65 42.055 23.91 42.315 ;
        RECT 23.65 41.295 23.91 41.555 ;
        RECT 23.65 40.535 23.91 40.795 ;
        RECT 23.65 39.775 23.91 40.035 ;
        RECT 23.65 39.015 23.91 39.275 ;
        RECT 23.65 38.255 23.91 38.515 ;
        RECT 23.65 37.495 23.91 37.755 ;
        RECT 23.65 36.735 23.91 36.995 ;
        RECT 24.41 58.775 24.67 59.035 ;
        RECT 24.41 58.015 24.67 58.275 ;
        RECT 24.41 57.255 24.67 57.515 ;
        RECT 24.41 56.495 24.67 56.755 ;
        RECT 24.41 55.735 24.67 55.995 ;
        RECT 24.41 54.975 24.67 55.235 ;
        RECT 24.41 54.215 24.67 54.475 ;
        RECT 24.41 53.455 24.67 53.715 ;
        RECT 24.41 52.695 24.67 52.955 ;
        RECT 24.41 51.935 24.67 52.195 ;
        RECT 24.41 51.175 24.67 51.435 ;
        RECT 24.41 50.415 24.67 50.675 ;
        RECT 24.41 49.655 24.67 49.915 ;
        RECT 24.41 48.895 24.67 49.155 ;
        RECT 24.41 48.135 24.67 48.395 ;
        RECT 24.41 47.375 24.67 47.635 ;
        RECT 24.41 46.615 24.67 46.875 ;
        RECT 24.41 45.855 24.67 46.115 ;
        RECT 24.41 45.095 24.67 45.355 ;
        RECT 24.41 44.335 24.67 44.595 ;
        RECT 24.41 43.575 24.67 43.835 ;
        RECT 24.41 42.815 24.67 43.075 ;
        RECT 24.41 42.055 24.67 42.315 ;
        RECT 24.41 41.295 24.67 41.555 ;
        RECT 24.41 40.535 24.67 40.795 ;
        RECT 24.41 39.775 24.67 40.035 ;
        RECT 24.41 39.015 24.67 39.275 ;
        RECT 24.41 38.255 24.67 38.515 ;
        RECT 24.41 37.495 24.67 37.755 ;
        RECT 24.41 36.735 24.67 36.995 ;
        RECT 25.17 58.775 25.43 59.035 ;
        RECT 25.17 58.015 25.43 58.275 ;
        RECT 25.17 57.255 25.43 57.515 ;
        RECT 25.17 56.495 25.43 56.755 ;
        RECT 25.17 55.735 25.43 55.995 ;
        RECT 25.17 54.975 25.43 55.235 ;
        RECT 25.17 54.215 25.43 54.475 ;
        RECT 25.17 53.455 25.43 53.715 ;
        RECT 25.17 52.695 25.43 52.955 ;
        RECT 25.17 51.935 25.43 52.195 ;
        RECT 25.17 51.175 25.43 51.435 ;
        RECT 25.17 50.415 25.43 50.675 ;
        RECT 25.17 49.655 25.43 49.915 ;
        RECT 25.17 48.895 25.43 49.155 ;
        RECT 25.17 48.135 25.43 48.395 ;
        RECT 25.17 47.375 25.43 47.635 ;
        RECT 25.17 46.615 25.43 46.875 ;
        RECT 25.17 45.855 25.43 46.115 ;
        RECT 25.17 45.095 25.43 45.355 ;
        RECT 25.17 44.335 25.43 44.595 ;
        RECT 25.17 43.575 25.43 43.835 ;
        RECT 25.17 42.815 25.43 43.075 ;
        RECT 25.17 42.055 25.43 42.315 ;
        RECT 25.17 41.295 25.43 41.555 ;
        RECT 25.17 40.535 25.43 40.795 ;
        RECT 25.17 39.775 25.43 40.035 ;
        RECT 25.17 39.015 25.43 39.275 ;
        RECT 25.17 38.255 25.43 38.515 ;
        RECT 25.17 37.495 25.43 37.755 ;
        RECT 25.17 36.735 25.43 36.995 ;
        RECT 25.93 58.775 26.19 59.035 ;
        RECT 25.93 58.015 26.19 58.275 ;
        RECT 25.93 57.255 26.19 57.515 ;
        RECT 25.93 56.495 26.19 56.755 ;
        RECT 25.93 55.735 26.19 55.995 ;
        RECT 25.93 54.975 26.19 55.235 ;
        RECT 25.93 54.215 26.19 54.475 ;
        RECT 25.93 53.455 26.19 53.715 ;
        RECT 25.93 52.695 26.19 52.955 ;
        RECT 25.93 51.935 26.19 52.195 ;
        RECT 25.93 51.175 26.19 51.435 ;
        RECT 25.93 50.415 26.19 50.675 ;
        RECT 25.93 49.655 26.19 49.915 ;
        RECT 25.93 48.895 26.19 49.155 ;
        RECT 25.93 48.135 26.19 48.395 ;
        RECT 25.93 47.375 26.19 47.635 ;
        RECT 25.93 46.615 26.19 46.875 ;
        RECT 25.93 45.855 26.19 46.115 ;
        RECT 25.93 45.095 26.19 45.355 ;
        RECT 25.93 44.335 26.19 44.595 ;
        RECT 25.93 43.575 26.19 43.835 ;
        RECT 25.93 42.815 26.19 43.075 ;
        RECT 25.93 42.055 26.19 42.315 ;
        RECT 25.93 41.295 26.19 41.555 ;
        RECT 25.93 40.535 26.19 40.795 ;
        RECT 25.93 39.775 26.19 40.035 ;
        RECT 25.93 39.015 26.19 39.275 ;
        RECT 25.93 38.255 26.19 38.515 ;
        RECT 25.93 37.495 26.19 37.755 ;
        RECT 25.93 36.735 26.19 36.995 ;
        RECT 26.69 58.775 26.95 59.035 ;
        RECT 26.69 58.015 26.95 58.275 ;
        RECT 26.69 57.255 26.95 57.515 ;
        RECT 26.69 56.495 26.95 56.755 ;
        RECT 26.69 55.735 26.95 55.995 ;
        RECT 26.69 54.975 26.95 55.235 ;
        RECT 26.69 54.215 26.95 54.475 ;
        RECT 26.69 53.455 26.95 53.715 ;
        RECT 26.69 52.695 26.95 52.955 ;
        RECT 26.69 51.935 26.95 52.195 ;
        RECT 26.69 51.175 26.95 51.435 ;
        RECT 26.69 50.415 26.95 50.675 ;
        RECT 26.69 49.655 26.95 49.915 ;
        RECT 26.69 48.895 26.95 49.155 ;
        RECT 26.69 48.135 26.95 48.395 ;
        RECT 26.69 47.375 26.95 47.635 ;
        RECT 26.69 46.615 26.95 46.875 ;
        RECT 26.69 45.855 26.95 46.115 ;
        RECT 26.69 45.095 26.95 45.355 ;
        RECT 26.69 44.335 26.95 44.595 ;
        RECT 26.69 43.575 26.95 43.835 ;
        RECT 26.69 42.815 26.95 43.075 ;
        RECT 26.69 42.055 26.95 42.315 ;
        RECT 26.69 41.295 26.95 41.555 ;
        RECT 26.69 40.535 26.95 40.795 ;
        RECT 26.69 39.775 26.95 40.035 ;
        RECT 26.69 39.015 26.95 39.275 ;
        RECT 26.69 38.255 26.95 38.515 ;
        RECT 26.69 37.495 26.95 37.755 ;
        RECT 26.69 36.735 26.95 36.995 ;
        RECT 27.45 58.775 27.71 59.035 ;
        RECT 27.45 58.015 27.71 58.275 ;
        RECT 27.45 57.255 27.71 57.515 ;
        RECT 27.45 56.495 27.71 56.755 ;
        RECT 27.45 55.735 27.71 55.995 ;
        RECT 27.45 54.975 27.71 55.235 ;
        RECT 27.45 54.215 27.71 54.475 ;
        RECT 27.45 53.455 27.71 53.715 ;
        RECT 27.45 52.695 27.71 52.955 ;
        RECT 27.45 51.935 27.71 52.195 ;
        RECT 27.45 51.175 27.71 51.435 ;
        RECT 27.45 50.415 27.71 50.675 ;
        RECT 27.45 49.655 27.71 49.915 ;
        RECT 27.45 48.895 27.71 49.155 ;
        RECT 27.45 48.135 27.71 48.395 ;
        RECT 27.45 47.375 27.71 47.635 ;
        RECT 27.45 46.615 27.71 46.875 ;
        RECT 27.45 45.855 27.71 46.115 ;
        RECT 27.45 45.095 27.71 45.355 ;
        RECT 27.45 44.335 27.71 44.595 ;
        RECT 27.45 43.575 27.71 43.835 ;
        RECT 27.45 42.815 27.71 43.075 ;
        RECT 27.45 42.055 27.71 42.315 ;
        RECT 27.45 41.295 27.71 41.555 ;
        RECT 27.45 40.535 27.71 40.795 ;
        RECT 27.45 39.775 27.71 40.035 ;
        RECT 27.45 39.015 27.71 39.275 ;
        RECT 27.45 38.255 27.71 38.515 ;
        RECT 27.45 37.495 27.71 37.755 ;
        RECT 27.45 36.735 27.71 36.995 ;
        RECT 28.21 58.775 28.47 59.035 ;
        RECT 28.21 58.015 28.47 58.275 ;
        RECT 28.21 57.255 28.47 57.515 ;
        RECT 28.21 56.495 28.47 56.755 ;
        RECT 28.21 55.735 28.47 55.995 ;
        RECT 28.21 54.975 28.47 55.235 ;
        RECT 28.21 54.215 28.47 54.475 ;
        RECT 28.21 53.455 28.47 53.715 ;
        RECT 28.21 52.695 28.47 52.955 ;
        RECT 28.21 51.935 28.47 52.195 ;
        RECT 28.21 51.175 28.47 51.435 ;
        RECT 28.21 50.415 28.47 50.675 ;
        RECT 28.21 49.655 28.47 49.915 ;
        RECT 28.21 48.895 28.47 49.155 ;
        RECT 28.21 48.135 28.47 48.395 ;
        RECT 28.21 47.375 28.47 47.635 ;
        RECT 28.21 46.615 28.47 46.875 ;
        RECT 28.21 45.855 28.47 46.115 ;
        RECT 28.21 45.095 28.47 45.355 ;
        RECT 28.21 44.335 28.47 44.595 ;
        RECT 28.21 43.575 28.47 43.835 ;
        RECT 28.21 42.815 28.47 43.075 ;
        RECT 28.21 42.055 28.47 42.315 ;
        RECT 28.21 41.295 28.47 41.555 ;
        RECT 28.21 40.535 28.47 40.795 ;
        RECT 28.21 39.775 28.47 40.035 ;
        RECT 28.21 39.015 28.47 39.275 ;
        RECT 28.21 38.255 28.47 38.515 ;
        RECT 28.21 37.495 28.47 37.755 ;
        RECT 28.21 36.735 28.47 36.995 ;
        RECT 28.97 58.775 29.23 59.035 ;
        RECT 28.97 58.015 29.23 58.275 ;
        RECT 28.97 57.255 29.23 57.515 ;
        RECT 28.97 56.495 29.23 56.755 ;
        RECT 28.97 55.735 29.23 55.995 ;
        RECT 28.97 54.975 29.23 55.235 ;
        RECT 28.97 54.215 29.23 54.475 ;
        RECT 28.97 53.455 29.23 53.715 ;
        RECT 28.97 52.695 29.23 52.955 ;
        RECT 28.97 51.935 29.23 52.195 ;
        RECT 28.97 51.175 29.23 51.435 ;
        RECT 28.97 50.415 29.23 50.675 ;
        RECT 28.97 49.655 29.23 49.915 ;
        RECT 28.97 48.895 29.23 49.155 ;
        RECT 28.97 48.135 29.23 48.395 ;
        RECT 28.97 47.375 29.23 47.635 ;
        RECT 28.97 46.615 29.23 46.875 ;
        RECT 28.97 45.855 29.23 46.115 ;
        RECT 28.97 45.095 29.23 45.355 ;
        RECT 28.97 44.335 29.23 44.595 ;
        RECT 28.97 43.575 29.23 43.835 ;
        RECT 28.97 42.815 29.23 43.075 ;
        RECT 28.97 42.055 29.23 42.315 ;
        RECT 28.97 41.295 29.23 41.555 ;
        RECT 28.97 40.535 29.23 40.795 ;
        RECT 28.97 39.775 29.23 40.035 ;
        RECT 28.97 39.015 29.23 39.275 ;
        RECT 28.97 38.255 29.23 38.515 ;
        RECT 28.97 37.495 29.23 37.755 ;
        RECT 28.97 36.735 29.23 36.995 ;
        RECT 29.73 58.775 29.99 59.035 ;
        RECT 29.73 58.015 29.99 58.275 ;
        RECT 29.73 57.255 29.99 57.515 ;
        RECT 29.73 56.495 29.99 56.755 ;
        RECT 29.73 55.735 29.99 55.995 ;
        RECT 29.73 54.975 29.99 55.235 ;
        RECT 29.73 54.215 29.99 54.475 ;
        RECT 29.73 53.455 29.99 53.715 ;
        RECT 29.73 52.695 29.99 52.955 ;
        RECT 29.73 51.935 29.99 52.195 ;
      LAYER M5 ;
        RECT 4 4 96 96 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M3 ;
        RECT 0 66 100 96 ;
      LAYER M4 ;
        RECT 0 66 100 96 ;
      LAYER V4 ;
        RECT 80.65 91.2 80.91 91.46 ;
        RECT 80.65 90.44 80.91 90.7 ;
        RECT 80.65 89.68 80.91 89.94 ;
        RECT 80.65 88.92 80.91 89.18 ;
        RECT 80.65 88.16 80.91 88.42 ;
        RECT 80.65 87.4 80.91 87.66 ;
        RECT 80.65 86.64 80.91 86.9 ;
        RECT 80.65 85.88 80.91 86.14 ;
        RECT 80.65 85.12 80.91 85.38 ;
        RECT 80.65 84.36 80.91 84.62 ;
        RECT 80.65 83.6 80.91 83.86 ;
        RECT 80.65 82.84 80.91 83.1 ;
        RECT 80.65 82.08 80.91 82.34 ;
        RECT 80.65 81.32 80.91 81.58 ;
        RECT 80.65 80.56 80.91 80.82 ;
        RECT 80.65 79.8 80.91 80.06 ;
        RECT 80.65 79.04 80.91 79.3 ;
        RECT 80.65 78.28 80.91 78.54 ;
        RECT 80.65 77.52 80.91 77.78 ;
        RECT 80.65 76.76 80.91 77.02 ;
        RECT 80.65 76 80.91 76.26 ;
        RECT 80.65 75.24 80.91 75.5 ;
        RECT 80.65 74.48 80.91 74.74 ;
        RECT 80.65 73.72 80.91 73.98 ;
        RECT 80.65 72.96 80.91 73.22 ;
        RECT 80.65 72.2 80.91 72.46 ;
        RECT 80.65 71.44 80.91 71.7 ;
        RECT 80.65 70.68 80.91 70.94 ;
        RECT 80.65 69.92 80.91 70.18 ;
        RECT 80.65 69.16 80.91 69.42 ;
        RECT 81.41 91.2 81.67 91.46 ;
        RECT 81.41 90.44 81.67 90.7 ;
        RECT 81.41 89.68 81.67 89.94 ;
        RECT 81.41 88.92 81.67 89.18 ;
        RECT 81.41 88.16 81.67 88.42 ;
        RECT 81.41 87.4 81.67 87.66 ;
        RECT 81.41 86.64 81.67 86.9 ;
        RECT 81.41 85.88 81.67 86.14 ;
        RECT 81.41 85.12 81.67 85.38 ;
        RECT 81.41 84.36 81.67 84.62 ;
        RECT 81.41 83.6 81.67 83.86 ;
        RECT 81.41 82.84 81.67 83.1 ;
        RECT 81.41 82.08 81.67 82.34 ;
        RECT 81.41 81.32 81.67 81.58 ;
        RECT 81.41 80.56 81.67 80.82 ;
        RECT 81.41 79.8 81.67 80.06 ;
        RECT 81.41 79.04 81.67 79.3 ;
        RECT 81.41 78.28 81.67 78.54 ;
        RECT 81.41 77.52 81.67 77.78 ;
        RECT 81.41 76.76 81.67 77.02 ;
        RECT 81.41 76 81.67 76.26 ;
        RECT 81.41 75.24 81.67 75.5 ;
        RECT 81.41 74.48 81.67 74.74 ;
        RECT 81.41 73.72 81.67 73.98 ;
        RECT 81.41 72.96 81.67 73.22 ;
        RECT 81.41 72.2 81.67 72.46 ;
        RECT 81.41 71.44 81.67 71.7 ;
        RECT 81.41 70.68 81.67 70.94 ;
        RECT 81.41 69.92 81.67 70.18 ;
        RECT 81.41 69.16 81.67 69.42 ;
        RECT 82.17 91.2 82.43 91.46 ;
        RECT 82.17 90.44 82.43 90.7 ;
        RECT 82.17 89.68 82.43 89.94 ;
        RECT 82.17 88.92 82.43 89.18 ;
        RECT 82.17 88.16 82.43 88.42 ;
        RECT 82.17 87.4 82.43 87.66 ;
        RECT 82.17 86.64 82.43 86.9 ;
        RECT 82.17 85.88 82.43 86.14 ;
        RECT 82.17 85.12 82.43 85.38 ;
        RECT 82.17 84.36 82.43 84.62 ;
        RECT 82.17 83.6 82.43 83.86 ;
        RECT 82.17 82.84 82.43 83.1 ;
        RECT 82.17 82.08 82.43 82.34 ;
        RECT 82.17 81.32 82.43 81.58 ;
        RECT 82.17 80.56 82.43 80.82 ;
        RECT 82.17 79.8 82.43 80.06 ;
        RECT 82.17 79.04 82.43 79.3 ;
        RECT 82.17 78.28 82.43 78.54 ;
        RECT 82.17 77.52 82.43 77.78 ;
        RECT 82.17 76.76 82.43 77.02 ;
        RECT 82.17 76 82.43 76.26 ;
        RECT 82.17 75.24 82.43 75.5 ;
        RECT 82.17 74.48 82.43 74.74 ;
        RECT 82.17 73.72 82.43 73.98 ;
        RECT 82.17 72.96 82.43 73.22 ;
        RECT 82.17 72.2 82.43 72.46 ;
        RECT 82.17 71.44 82.43 71.7 ;
        RECT 82.17 70.68 82.43 70.94 ;
        RECT 82.17 69.92 82.43 70.18 ;
        RECT 82.17 69.16 82.43 69.42 ;
        RECT 82.93 91.2 83.19 91.46 ;
        RECT 82.93 90.44 83.19 90.7 ;
        RECT 82.93 89.68 83.19 89.94 ;
        RECT 82.93 88.92 83.19 89.18 ;
        RECT 82.93 88.16 83.19 88.42 ;
        RECT 82.93 87.4 83.19 87.66 ;
        RECT 82.93 86.64 83.19 86.9 ;
        RECT 82.93 85.88 83.19 86.14 ;
        RECT 82.93 85.12 83.19 85.38 ;
        RECT 82.93 84.36 83.19 84.62 ;
        RECT 82.93 83.6 83.19 83.86 ;
        RECT 82.93 82.84 83.19 83.1 ;
        RECT 82.93 82.08 83.19 82.34 ;
        RECT 82.93 81.32 83.19 81.58 ;
        RECT 82.93 80.56 83.19 80.82 ;
        RECT 82.93 79.8 83.19 80.06 ;
        RECT 82.93 79.04 83.19 79.3 ;
        RECT 82.93 78.28 83.19 78.54 ;
        RECT 82.93 77.52 83.19 77.78 ;
        RECT 82.93 76.76 83.19 77.02 ;
        RECT 82.93 76 83.19 76.26 ;
        RECT 82.93 75.24 83.19 75.5 ;
        RECT 82.93 74.48 83.19 74.74 ;
        RECT 82.93 73.72 83.19 73.98 ;
        RECT 82.93 72.96 83.19 73.22 ;
        RECT 82.93 72.2 83.19 72.46 ;
        RECT 82.93 71.44 83.19 71.7 ;
        RECT 82.93 70.68 83.19 70.94 ;
        RECT 82.93 69.92 83.19 70.18 ;
        RECT 82.93 69.16 83.19 69.42 ;
        RECT 83.69 91.2 83.95 91.46 ;
        RECT 83.69 90.44 83.95 90.7 ;
        RECT 83.69 89.68 83.95 89.94 ;
        RECT 83.69 88.92 83.95 89.18 ;
        RECT 83.69 88.16 83.95 88.42 ;
        RECT 83.69 87.4 83.95 87.66 ;
        RECT 83.69 86.64 83.95 86.9 ;
        RECT 83.69 85.88 83.95 86.14 ;
        RECT 83.69 85.12 83.95 85.38 ;
        RECT 83.69 84.36 83.95 84.62 ;
        RECT 83.69 83.6 83.95 83.86 ;
        RECT 83.69 82.84 83.95 83.1 ;
        RECT 83.69 82.08 83.95 82.34 ;
        RECT 83.69 81.32 83.95 81.58 ;
        RECT 83.69 80.56 83.95 80.82 ;
        RECT 83.69 79.8 83.95 80.06 ;
        RECT 83.69 79.04 83.95 79.3 ;
        RECT 83.69 78.28 83.95 78.54 ;
        RECT 83.69 77.52 83.95 77.78 ;
        RECT 83.69 76.76 83.95 77.02 ;
        RECT 83.69 76 83.95 76.26 ;
        RECT 83.69 75.24 83.95 75.5 ;
        RECT 83.69 74.48 83.95 74.74 ;
        RECT 83.69 73.72 83.95 73.98 ;
        RECT 83.69 72.96 83.95 73.22 ;
        RECT 83.69 72.2 83.95 72.46 ;
        RECT 83.69 71.44 83.95 71.7 ;
        RECT 83.69 70.68 83.95 70.94 ;
        RECT 83.69 69.92 83.95 70.18 ;
        RECT 83.69 69.16 83.95 69.42 ;
        RECT 84.45 91.2 84.71 91.46 ;
        RECT 84.45 90.44 84.71 90.7 ;
        RECT 84.45 89.68 84.71 89.94 ;
        RECT 84.45 88.92 84.71 89.18 ;
        RECT 84.45 88.16 84.71 88.42 ;
        RECT 84.45 87.4 84.71 87.66 ;
        RECT 84.45 86.64 84.71 86.9 ;
        RECT 84.45 85.88 84.71 86.14 ;
        RECT 84.45 85.12 84.71 85.38 ;
        RECT 84.45 84.36 84.71 84.62 ;
        RECT 84.45 83.6 84.71 83.86 ;
        RECT 84.45 82.84 84.71 83.1 ;
        RECT 84.45 82.08 84.71 82.34 ;
        RECT 84.45 81.32 84.71 81.58 ;
        RECT 84.45 80.56 84.71 80.82 ;
        RECT 84.45 79.8 84.71 80.06 ;
        RECT 84.45 79.04 84.71 79.3 ;
        RECT 84.45 78.28 84.71 78.54 ;
        RECT 84.45 77.52 84.71 77.78 ;
        RECT 84.45 76.76 84.71 77.02 ;
        RECT 84.45 76 84.71 76.26 ;
        RECT 84.45 75.24 84.71 75.5 ;
        RECT 84.45 74.48 84.71 74.74 ;
        RECT 84.45 73.72 84.71 73.98 ;
        RECT 84.45 72.96 84.71 73.22 ;
        RECT 84.45 72.2 84.71 72.46 ;
        RECT 84.45 71.44 84.71 71.7 ;
        RECT 84.45 70.68 84.71 70.94 ;
        RECT 84.45 69.92 84.71 70.18 ;
        RECT 84.45 69.16 84.71 69.42 ;
        RECT 85.21 91.2 85.47 91.46 ;
        RECT 85.21 90.44 85.47 90.7 ;
        RECT 85.21 89.68 85.47 89.94 ;
        RECT 85.21 88.92 85.47 89.18 ;
        RECT 85.21 88.16 85.47 88.42 ;
        RECT 85.21 87.4 85.47 87.66 ;
        RECT 85.21 86.64 85.47 86.9 ;
        RECT 85.21 85.88 85.47 86.14 ;
        RECT 85.21 85.12 85.47 85.38 ;
        RECT 85.21 84.36 85.47 84.62 ;
        RECT 85.21 83.6 85.47 83.86 ;
        RECT 85.21 82.84 85.47 83.1 ;
        RECT 85.21 82.08 85.47 82.34 ;
        RECT 85.21 81.32 85.47 81.58 ;
        RECT 85.21 80.56 85.47 80.82 ;
        RECT 85.21 79.8 85.47 80.06 ;
        RECT 85.21 79.04 85.47 79.3 ;
        RECT 85.21 78.28 85.47 78.54 ;
        RECT 85.21 77.52 85.47 77.78 ;
        RECT 85.21 76.76 85.47 77.02 ;
        RECT 85.21 76 85.47 76.26 ;
        RECT 85.21 75.24 85.47 75.5 ;
        RECT 85.21 74.48 85.47 74.74 ;
        RECT 85.21 73.72 85.47 73.98 ;
        RECT 85.21 72.96 85.47 73.22 ;
        RECT 85.21 72.2 85.47 72.46 ;
        RECT 85.21 71.44 85.47 71.7 ;
        RECT 85.21 70.68 85.47 70.94 ;
        RECT 85.21 69.92 85.47 70.18 ;
        RECT 85.21 69.16 85.47 69.42 ;
        RECT 85.97 91.2 86.23 91.46 ;
        RECT 85.97 90.44 86.23 90.7 ;
        RECT 85.97 89.68 86.23 89.94 ;
        RECT 85.97 88.92 86.23 89.18 ;
        RECT 85.97 88.16 86.23 88.42 ;
        RECT 85.97 87.4 86.23 87.66 ;
        RECT 85.97 86.64 86.23 86.9 ;
        RECT 85.97 85.88 86.23 86.14 ;
        RECT 85.97 85.12 86.23 85.38 ;
        RECT 85.97 84.36 86.23 84.62 ;
        RECT 85.97 83.6 86.23 83.86 ;
        RECT 85.97 82.84 86.23 83.1 ;
        RECT 85.97 82.08 86.23 82.34 ;
        RECT 85.97 81.32 86.23 81.58 ;
        RECT 85.97 80.56 86.23 80.82 ;
        RECT 85.97 79.8 86.23 80.06 ;
        RECT 85.97 79.04 86.23 79.3 ;
        RECT 85.97 78.28 86.23 78.54 ;
        RECT 85.97 77.52 86.23 77.78 ;
        RECT 85.97 76.76 86.23 77.02 ;
        RECT 85.97 76 86.23 76.26 ;
        RECT 85.97 75.24 86.23 75.5 ;
        RECT 85.97 74.48 86.23 74.74 ;
        RECT 85.97 73.72 86.23 73.98 ;
        RECT 85.97 72.96 86.23 73.22 ;
        RECT 85.97 72.2 86.23 72.46 ;
        RECT 85.97 71.44 86.23 71.7 ;
        RECT 85.97 70.68 86.23 70.94 ;
        RECT 85.97 69.92 86.23 70.18 ;
        RECT 85.97 69.16 86.23 69.42 ;
        RECT 86.73 91.2 86.99 91.46 ;
        RECT 86.73 90.44 86.99 90.7 ;
        RECT 86.73 89.68 86.99 89.94 ;
        RECT 86.73 88.92 86.99 89.18 ;
        RECT 86.73 88.16 86.99 88.42 ;
        RECT 86.73 87.4 86.99 87.66 ;
        RECT 86.73 86.64 86.99 86.9 ;
        RECT 86.73 85.88 86.99 86.14 ;
        RECT 86.73 85.12 86.99 85.38 ;
        RECT 86.73 84.36 86.99 84.62 ;
        RECT 86.73 83.6 86.99 83.86 ;
        RECT 86.73 82.84 86.99 83.1 ;
        RECT 86.73 82.08 86.99 82.34 ;
        RECT 86.73 81.32 86.99 81.58 ;
        RECT 86.73 80.56 86.99 80.82 ;
        RECT 86.73 79.8 86.99 80.06 ;
        RECT 86.73 79.04 86.99 79.3 ;
        RECT 86.73 78.28 86.99 78.54 ;
        RECT 86.73 77.52 86.99 77.78 ;
        RECT 86.73 76.76 86.99 77.02 ;
        RECT 86.73 76 86.99 76.26 ;
        RECT 86.73 75.24 86.99 75.5 ;
        RECT 86.73 74.48 86.99 74.74 ;
        RECT 86.73 73.72 86.99 73.98 ;
        RECT 86.73 72.96 86.99 73.22 ;
        RECT 86.73 72.2 86.99 72.46 ;
        RECT 86.73 71.44 86.99 71.7 ;
        RECT 86.73 70.68 86.99 70.94 ;
        RECT 86.73 69.92 86.99 70.18 ;
        RECT 86.73 69.16 86.99 69.42 ;
        RECT 87.49 91.2 87.75 91.46 ;
        RECT 87.49 90.44 87.75 90.7 ;
        RECT 87.49 89.68 87.75 89.94 ;
        RECT 87.49 88.92 87.75 89.18 ;
        RECT 87.49 88.16 87.75 88.42 ;
        RECT 87.49 87.4 87.75 87.66 ;
        RECT 87.49 86.64 87.75 86.9 ;
        RECT 87.49 85.88 87.75 86.14 ;
        RECT 87.49 85.12 87.75 85.38 ;
        RECT 87.49 84.36 87.75 84.62 ;
        RECT 87.49 83.6 87.75 83.86 ;
        RECT 87.49 82.84 87.75 83.1 ;
        RECT 87.49 82.08 87.75 82.34 ;
        RECT 87.49 81.32 87.75 81.58 ;
        RECT 87.49 80.56 87.75 80.82 ;
        RECT 87.49 79.8 87.75 80.06 ;
        RECT 87.49 79.04 87.75 79.3 ;
        RECT 87.49 78.28 87.75 78.54 ;
        RECT 87.49 77.52 87.75 77.78 ;
        RECT 87.49 76.76 87.75 77.02 ;
        RECT 87.49 76 87.75 76.26 ;
        RECT 87.49 75.24 87.75 75.5 ;
        RECT 87.49 74.48 87.75 74.74 ;
        RECT 87.49 73.72 87.75 73.98 ;
        RECT 87.49 72.96 87.75 73.22 ;
        RECT 87.49 72.2 87.75 72.46 ;
        RECT 87.49 71.44 87.75 71.7 ;
        RECT 87.49 70.68 87.75 70.94 ;
        RECT 87.49 69.92 87.75 70.18 ;
        RECT 87.49 69.16 87.75 69.42 ;
        RECT 88.25 91.2 88.51 91.46 ;
        RECT 88.25 90.44 88.51 90.7 ;
        RECT 88.25 89.68 88.51 89.94 ;
        RECT 88.25 88.92 88.51 89.18 ;
        RECT 88.25 88.16 88.51 88.42 ;
        RECT 88.25 87.4 88.51 87.66 ;
        RECT 88.25 86.64 88.51 86.9 ;
        RECT 88.25 85.88 88.51 86.14 ;
        RECT 88.25 85.12 88.51 85.38 ;
        RECT 88.25 84.36 88.51 84.62 ;
        RECT 88.25 83.6 88.51 83.86 ;
        RECT 88.25 82.84 88.51 83.1 ;
        RECT 88.25 82.08 88.51 82.34 ;
        RECT 88.25 81.32 88.51 81.58 ;
        RECT 88.25 80.56 88.51 80.82 ;
        RECT 88.25 79.8 88.51 80.06 ;
        RECT 88.25 79.04 88.51 79.3 ;
        RECT 88.25 78.28 88.51 78.54 ;
        RECT 88.25 77.52 88.51 77.78 ;
        RECT 88.25 76.76 88.51 77.02 ;
        RECT 88.25 76 88.51 76.26 ;
        RECT 88.25 75.24 88.51 75.5 ;
        RECT 88.25 74.48 88.51 74.74 ;
        RECT 88.25 73.72 88.51 73.98 ;
        RECT 88.25 72.96 88.51 73.22 ;
        RECT 88.25 72.2 88.51 72.46 ;
        RECT 88.25 71.44 88.51 71.7 ;
        RECT 88.25 70.68 88.51 70.94 ;
        RECT 88.25 69.92 88.51 70.18 ;
        RECT 88.25 69.16 88.51 69.42 ;
        RECT 89.01 91.2 89.27 91.46 ;
        RECT 89.01 90.44 89.27 90.7 ;
        RECT 89.01 89.68 89.27 89.94 ;
        RECT 89.01 88.92 89.27 89.18 ;
        RECT 89.01 88.16 89.27 88.42 ;
        RECT 89.01 87.4 89.27 87.66 ;
        RECT 89.01 86.64 89.27 86.9 ;
        RECT 89.01 85.88 89.27 86.14 ;
        RECT 89.01 85.12 89.27 85.38 ;
        RECT 89.01 84.36 89.27 84.62 ;
        RECT 89.01 83.6 89.27 83.86 ;
        RECT 89.01 82.84 89.27 83.1 ;
        RECT 89.01 82.08 89.27 82.34 ;
        RECT 89.01 81.32 89.27 81.58 ;
        RECT 89.01 80.56 89.27 80.82 ;
        RECT 89.01 79.8 89.27 80.06 ;
        RECT 89.01 79.04 89.27 79.3 ;
        RECT 89.01 78.28 89.27 78.54 ;
        RECT 89.01 77.52 89.27 77.78 ;
        RECT 89.01 76.76 89.27 77.02 ;
        RECT 89.01 76 89.27 76.26 ;
        RECT 89.01 75.24 89.27 75.5 ;
        RECT 89.01 74.48 89.27 74.74 ;
        RECT 89.01 73.72 89.27 73.98 ;
        RECT 89.01 72.96 89.27 73.22 ;
        RECT 89.01 72.2 89.27 72.46 ;
        RECT 89.01 71.44 89.27 71.7 ;
        RECT 89.01 70.68 89.27 70.94 ;
        RECT 89.01 69.92 89.27 70.18 ;
        RECT 89.01 69.16 89.27 69.42 ;
        RECT 89.77 91.2 90.03 91.46 ;
        RECT 89.77 90.44 90.03 90.7 ;
        RECT 89.77 89.68 90.03 89.94 ;
        RECT 89.77 88.92 90.03 89.18 ;
        RECT 89.77 88.16 90.03 88.42 ;
        RECT 89.77 87.4 90.03 87.66 ;
        RECT 89.77 86.64 90.03 86.9 ;
        RECT 89.77 85.88 90.03 86.14 ;
        RECT 89.77 85.12 90.03 85.38 ;
        RECT 89.77 84.36 90.03 84.62 ;
        RECT 89.77 83.6 90.03 83.86 ;
        RECT 89.77 82.84 90.03 83.1 ;
        RECT 89.77 82.08 90.03 82.34 ;
        RECT 89.77 81.32 90.03 81.58 ;
        RECT 89.77 80.56 90.03 80.82 ;
        RECT 89.77 79.8 90.03 80.06 ;
        RECT 89.77 79.04 90.03 79.3 ;
        RECT 89.77 78.28 90.03 78.54 ;
        RECT 89.77 77.52 90.03 77.78 ;
        RECT 89.77 76.76 90.03 77.02 ;
        RECT 89.77 76 90.03 76.26 ;
        RECT 89.77 75.24 90.03 75.5 ;
        RECT 89.77 74.48 90.03 74.74 ;
        RECT 89.77 73.72 90.03 73.98 ;
        RECT 89.77 72.96 90.03 73.22 ;
        RECT 89.77 72.2 90.03 72.46 ;
        RECT 89.77 71.44 90.03 71.7 ;
        RECT 89.77 70.68 90.03 70.94 ;
        RECT 89.77 69.92 90.03 70.18 ;
        RECT 89.77 69.16 90.03 69.42 ;
        RECT 90.53 91.2 90.79 91.46 ;
        RECT 90.53 90.44 90.79 90.7 ;
        RECT 90.53 89.68 90.79 89.94 ;
        RECT 90.53 88.92 90.79 89.18 ;
        RECT 90.53 88.16 90.79 88.42 ;
        RECT 90.53 87.4 90.79 87.66 ;
        RECT 90.53 86.64 90.79 86.9 ;
        RECT 90.53 85.88 90.79 86.14 ;
        RECT 90.53 85.12 90.79 85.38 ;
        RECT 90.53 84.36 90.79 84.62 ;
        RECT 90.53 83.6 90.79 83.86 ;
        RECT 90.53 82.84 90.79 83.1 ;
        RECT 90.53 82.08 90.79 82.34 ;
        RECT 90.53 81.32 90.79 81.58 ;
        RECT 90.53 80.56 90.79 80.82 ;
        RECT 90.53 79.8 90.79 80.06 ;
        RECT 90.53 79.04 90.79 79.3 ;
        RECT 90.53 78.28 90.79 78.54 ;
        RECT 90.53 77.52 90.79 77.78 ;
        RECT 90.53 76.76 90.79 77.02 ;
        RECT 90.53 76 90.79 76.26 ;
        RECT 90.53 75.24 90.79 75.5 ;
        RECT 90.53 74.48 90.79 74.74 ;
        RECT 90.53 73.72 90.79 73.98 ;
        RECT 90.53 72.96 90.79 73.22 ;
        RECT 90.53 72.2 90.79 72.46 ;
        RECT 90.53 71.44 90.79 71.7 ;
        RECT 90.53 70.68 90.79 70.94 ;
        RECT 90.53 69.92 90.79 70.18 ;
        RECT 90.53 69.16 90.79 69.42 ;
        RECT 91.29 91.2 91.55 91.46 ;
        RECT 91.29 90.44 91.55 90.7 ;
        RECT 91.29 89.68 91.55 89.94 ;
        RECT 91.29 88.92 91.55 89.18 ;
        RECT 91.29 88.16 91.55 88.42 ;
        RECT 91.29 87.4 91.55 87.66 ;
        RECT 91.29 86.64 91.55 86.9 ;
        RECT 91.29 85.88 91.55 86.14 ;
        RECT 91.29 85.12 91.55 85.38 ;
        RECT 91.29 84.36 91.55 84.62 ;
        RECT 91.29 83.6 91.55 83.86 ;
        RECT 91.29 82.84 91.55 83.1 ;
        RECT 91.29 82.08 91.55 82.34 ;
        RECT 91.29 81.32 91.55 81.58 ;
        RECT 91.29 80.56 91.55 80.82 ;
        RECT 91.29 79.8 91.55 80.06 ;
        RECT 91.29 79.04 91.55 79.3 ;
        RECT 91.29 78.28 91.55 78.54 ;
        RECT 91.29 77.52 91.55 77.78 ;
        RECT 91.29 76.76 91.55 77.02 ;
        RECT 91.29 76 91.55 76.26 ;
        RECT 91.29 75.24 91.55 75.5 ;
        RECT 91.29 74.48 91.55 74.74 ;
        RECT 91.29 73.72 91.55 73.98 ;
        RECT 91.29 72.96 91.55 73.22 ;
        RECT 91.29 72.2 91.55 72.46 ;
        RECT 91.29 71.44 91.55 71.7 ;
        RECT 91.29 70.68 91.55 70.94 ;
        RECT 91.29 69.92 91.55 70.18 ;
        RECT 91.29 69.16 91.55 69.42 ;
        RECT 92.05 91.2 92.31 91.46 ;
        RECT 92.05 90.44 92.31 90.7 ;
        RECT 92.05 89.68 92.31 89.94 ;
        RECT 92.05 88.92 92.31 89.18 ;
        RECT 92.05 88.16 92.31 88.42 ;
        RECT 92.05 87.4 92.31 87.66 ;
        RECT 92.05 86.64 92.31 86.9 ;
        RECT 92.05 85.88 92.31 86.14 ;
        RECT 92.05 85.12 92.31 85.38 ;
        RECT 92.05 84.36 92.31 84.62 ;
        RECT 92.05 83.6 92.31 83.86 ;
        RECT 92.05 82.84 92.31 83.1 ;
        RECT 92.05 82.08 92.31 82.34 ;
        RECT 92.05 81.32 92.31 81.58 ;
        RECT 92.05 80.56 92.31 80.82 ;
        RECT 92.05 79.8 92.31 80.06 ;
        RECT 92.05 79.04 92.31 79.3 ;
        RECT 92.05 78.28 92.31 78.54 ;
        RECT 92.05 77.52 92.31 77.78 ;
        RECT 92.05 76.76 92.31 77.02 ;
        RECT 92.05 76 92.31 76.26 ;
        RECT 92.05 75.24 92.31 75.5 ;
        RECT 92.05 74.48 92.31 74.74 ;
        RECT 92.05 73.72 92.31 73.98 ;
        RECT 92.05 72.96 92.31 73.22 ;
        RECT 92.05 72.2 92.31 72.46 ;
        RECT 92.05 71.44 92.31 71.7 ;
        RECT 92.05 70.68 92.31 70.94 ;
        RECT 92.05 69.92 92.31 70.18 ;
        RECT 92.05 69.16 92.31 69.42 ;
        RECT 92.81 91.2 93.07 91.46 ;
        RECT 92.81 90.44 93.07 90.7 ;
        RECT 92.81 89.68 93.07 89.94 ;
        RECT 92.81 88.92 93.07 89.18 ;
        RECT 92.81 88.16 93.07 88.42 ;
        RECT 92.81 87.4 93.07 87.66 ;
        RECT 92.81 86.64 93.07 86.9 ;
        RECT 92.81 85.88 93.07 86.14 ;
        RECT 92.81 85.12 93.07 85.38 ;
        RECT 92.81 84.36 93.07 84.62 ;
        RECT 92.81 83.6 93.07 83.86 ;
        RECT 92.81 82.84 93.07 83.1 ;
        RECT 92.81 82.08 93.07 82.34 ;
        RECT 92.81 81.32 93.07 81.58 ;
        RECT 92.81 80.56 93.07 80.82 ;
        RECT 92.81 79.8 93.07 80.06 ;
        RECT 92.81 79.04 93.07 79.3 ;
        RECT 92.81 78.28 93.07 78.54 ;
        RECT 92.81 77.52 93.07 77.78 ;
        RECT 92.81 76.76 93.07 77.02 ;
        RECT 92.81 76 93.07 76.26 ;
        RECT 92.81 75.24 93.07 75.5 ;
        RECT 92.81 74.48 93.07 74.74 ;
        RECT 92.81 73.72 93.07 73.98 ;
        RECT 92.81 72.96 93.07 73.22 ;
        RECT 92.81 72.2 93.07 72.46 ;
        RECT 92.81 71.44 93.07 71.7 ;
        RECT 92.81 70.68 93.07 70.94 ;
        RECT 92.81 69.92 93.07 70.18 ;
        RECT 92.81 69.16 93.07 69.42 ;
        RECT 93.57 91.2 93.83 91.46 ;
        RECT 93.57 90.44 93.83 90.7 ;
        RECT 93.57 89.68 93.83 89.94 ;
        RECT 93.57 88.92 93.83 89.18 ;
        RECT 93.57 88.16 93.83 88.42 ;
        RECT 93.57 87.4 93.83 87.66 ;
        RECT 93.57 86.64 93.83 86.9 ;
        RECT 93.57 85.88 93.83 86.14 ;
        RECT 93.57 85.12 93.83 85.38 ;
        RECT 93.57 84.36 93.83 84.62 ;
        RECT 93.57 83.6 93.83 83.86 ;
        RECT 93.57 82.84 93.83 83.1 ;
        RECT 93.57 82.08 93.83 82.34 ;
        RECT 93.57 81.32 93.83 81.58 ;
        RECT 93.57 80.56 93.83 80.82 ;
        RECT 93.57 79.8 93.83 80.06 ;
        RECT 93.57 79.04 93.83 79.3 ;
        RECT 93.57 78.28 93.83 78.54 ;
        RECT 93.57 77.52 93.83 77.78 ;
        RECT 93.57 76.76 93.83 77.02 ;
        RECT 93.57 76 93.83 76.26 ;
        RECT 93.57 75.24 93.83 75.5 ;
        RECT 93.57 74.48 93.83 74.74 ;
        RECT 93.57 73.72 93.83 73.98 ;
        RECT 93.57 72.96 93.83 73.22 ;
        RECT 93.57 72.2 93.83 72.46 ;
        RECT 93.57 71.44 93.83 71.7 ;
        RECT 93.57 70.68 93.83 70.94 ;
        RECT 93.57 69.92 93.83 70.18 ;
        RECT 93.57 69.16 93.83 69.42 ;
        RECT 94.33 91.2 94.59 91.46 ;
        RECT 94.33 90.44 94.59 90.7 ;
        RECT 94.33 89.68 94.59 89.94 ;
        RECT 94.33 88.92 94.59 89.18 ;
        RECT 94.33 88.16 94.59 88.42 ;
        RECT 94.33 87.4 94.59 87.66 ;
        RECT 94.33 86.64 94.59 86.9 ;
        RECT 94.33 85.88 94.59 86.14 ;
        RECT 94.33 85.12 94.59 85.38 ;
        RECT 94.33 84.36 94.59 84.62 ;
        RECT 94.33 83.6 94.59 83.86 ;
        RECT 94.33 82.84 94.59 83.1 ;
        RECT 94.33 82.08 94.59 82.34 ;
        RECT 94.33 81.32 94.59 81.58 ;
        RECT 94.33 80.56 94.59 80.82 ;
        RECT 94.33 79.8 94.59 80.06 ;
        RECT 94.33 79.04 94.59 79.3 ;
        RECT 94.33 78.28 94.59 78.54 ;
        RECT 94.33 77.52 94.59 77.78 ;
        RECT 94.33 76.76 94.59 77.02 ;
        RECT 94.33 76 94.59 76.26 ;
        RECT 94.33 75.24 94.59 75.5 ;
        RECT 94.33 74.48 94.59 74.74 ;
        RECT 94.33 73.72 94.59 73.98 ;
        RECT 94.33 72.96 94.59 73.22 ;
        RECT 94.33 72.2 94.59 72.46 ;
        RECT 94.33 71.44 94.59 71.7 ;
        RECT 94.33 70.68 94.59 70.94 ;
        RECT 94.33 69.92 94.59 70.18 ;
        RECT 94.33 69.16 94.59 69.42 ;
        RECT 95.09 91.2 95.35 91.46 ;
        RECT 95.09 90.44 95.35 90.7 ;
        RECT 95.09 89.68 95.35 89.94 ;
        RECT 95.09 88.92 95.35 89.18 ;
        RECT 95.09 88.16 95.35 88.42 ;
        RECT 95.09 87.4 95.35 87.66 ;
        RECT 95.09 86.64 95.35 86.9 ;
        RECT 95.09 85.88 95.35 86.14 ;
        RECT 95.09 85.12 95.35 85.38 ;
        RECT 95.09 84.36 95.35 84.62 ;
        RECT 95.09 83.6 95.35 83.86 ;
        RECT 95.09 82.84 95.35 83.1 ;
        RECT 95.09 82.08 95.35 82.34 ;
        RECT 95.09 81.32 95.35 81.58 ;
        RECT 95.09 80.56 95.35 80.82 ;
        RECT 95.09 79.8 95.35 80.06 ;
        RECT 95.09 79.04 95.35 79.3 ;
        RECT 95.09 78.28 95.35 78.54 ;
        RECT 95.09 77.52 95.35 77.78 ;
        RECT 95.09 76.76 95.35 77.02 ;
        RECT 95.09 76 95.35 76.26 ;
        RECT 95.09 75.24 95.35 75.5 ;
        RECT 95.09 74.48 95.35 74.74 ;
        RECT 95.09 73.72 95.35 73.98 ;
        RECT 95.09 72.96 95.35 73.22 ;
        RECT 95.09 72.2 95.35 72.46 ;
        RECT 95.09 71.44 95.35 71.7 ;
        RECT 95.09 70.68 95.35 70.94 ;
        RECT 95.09 69.92 95.35 70.18 ;
        RECT 95.09 69.16 95.35 69.42 ;
        RECT 54.81 76 55.07 76.26 ;
        RECT 54.81 75.24 55.07 75.5 ;
        RECT 54.81 74.48 55.07 74.74 ;
        RECT 54.81 73.72 55.07 73.98 ;
        RECT 54.81 72.96 55.07 73.22 ;
        RECT 54.81 72.2 55.07 72.46 ;
        RECT 54.81 71.44 55.07 71.7 ;
        RECT 54.81 70.68 55.07 70.94 ;
        RECT 54.81 69.92 55.07 70.18 ;
        RECT 54.81 69.16 55.07 69.42 ;
        RECT 55.57 91.2 55.83 91.46 ;
        RECT 55.57 90.44 55.83 90.7 ;
        RECT 55.57 89.68 55.83 89.94 ;
        RECT 55.57 88.92 55.83 89.18 ;
        RECT 55.57 88.16 55.83 88.42 ;
        RECT 55.57 87.4 55.83 87.66 ;
        RECT 55.57 86.64 55.83 86.9 ;
        RECT 55.57 85.88 55.83 86.14 ;
        RECT 55.57 85.12 55.83 85.38 ;
        RECT 55.57 84.36 55.83 84.62 ;
        RECT 55.57 83.6 55.83 83.86 ;
        RECT 55.57 82.84 55.83 83.1 ;
        RECT 55.57 82.08 55.83 82.34 ;
        RECT 55.57 81.32 55.83 81.58 ;
        RECT 55.57 80.56 55.83 80.82 ;
        RECT 55.57 79.8 55.83 80.06 ;
        RECT 55.57 79.04 55.83 79.3 ;
        RECT 55.57 78.28 55.83 78.54 ;
        RECT 55.57 77.52 55.83 77.78 ;
        RECT 55.57 76.76 55.83 77.02 ;
        RECT 55.57 76 55.83 76.26 ;
        RECT 55.57 75.24 55.83 75.5 ;
        RECT 55.57 74.48 55.83 74.74 ;
        RECT 55.57 73.72 55.83 73.98 ;
        RECT 55.57 72.96 55.83 73.22 ;
        RECT 55.57 72.2 55.83 72.46 ;
        RECT 55.57 71.44 55.83 71.7 ;
        RECT 55.57 70.68 55.83 70.94 ;
        RECT 55.57 69.92 55.83 70.18 ;
        RECT 55.57 69.16 55.83 69.42 ;
        RECT 56.33 91.2 56.59 91.46 ;
        RECT 56.33 90.44 56.59 90.7 ;
        RECT 56.33 89.68 56.59 89.94 ;
        RECT 56.33 88.92 56.59 89.18 ;
        RECT 56.33 88.16 56.59 88.42 ;
        RECT 56.33 87.4 56.59 87.66 ;
        RECT 56.33 86.64 56.59 86.9 ;
        RECT 56.33 85.88 56.59 86.14 ;
        RECT 56.33 85.12 56.59 85.38 ;
        RECT 56.33 84.36 56.59 84.62 ;
        RECT 56.33 83.6 56.59 83.86 ;
        RECT 56.33 82.84 56.59 83.1 ;
        RECT 56.33 82.08 56.59 82.34 ;
        RECT 56.33 81.32 56.59 81.58 ;
        RECT 56.33 80.56 56.59 80.82 ;
        RECT 56.33 79.8 56.59 80.06 ;
        RECT 56.33 79.04 56.59 79.3 ;
        RECT 56.33 78.28 56.59 78.54 ;
        RECT 56.33 77.52 56.59 77.78 ;
        RECT 56.33 76.76 56.59 77.02 ;
        RECT 56.33 76 56.59 76.26 ;
        RECT 56.33 75.24 56.59 75.5 ;
        RECT 56.33 74.48 56.59 74.74 ;
        RECT 56.33 73.72 56.59 73.98 ;
        RECT 56.33 72.96 56.59 73.22 ;
        RECT 56.33 72.2 56.59 72.46 ;
        RECT 56.33 71.44 56.59 71.7 ;
        RECT 56.33 70.68 56.59 70.94 ;
        RECT 56.33 69.92 56.59 70.18 ;
        RECT 56.33 69.16 56.59 69.42 ;
        RECT 57.09 91.2 57.35 91.46 ;
        RECT 57.09 90.44 57.35 90.7 ;
        RECT 57.09 89.68 57.35 89.94 ;
        RECT 57.09 88.92 57.35 89.18 ;
        RECT 57.09 88.16 57.35 88.42 ;
        RECT 57.09 87.4 57.35 87.66 ;
        RECT 57.09 86.64 57.35 86.9 ;
        RECT 57.09 85.88 57.35 86.14 ;
        RECT 57.09 85.12 57.35 85.38 ;
        RECT 57.09 84.36 57.35 84.62 ;
        RECT 57.09 83.6 57.35 83.86 ;
        RECT 57.09 82.84 57.35 83.1 ;
        RECT 57.09 82.08 57.35 82.34 ;
        RECT 57.09 81.32 57.35 81.58 ;
        RECT 57.09 80.56 57.35 80.82 ;
        RECT 57.09 79.8 57.35 80.06 ;
        RECT 57.09 79.04 57.35 79.3 ;
        RECT 57.09 78.28 57.35 78.54 ;
        RECT 57.09 77.52 57.35 77.78 ;
        RECT 57.09 76.76 57.35 77.02 ;
        RECT 57.09 76 57.35 76.26 ;
        RECT 57.09 75.24 57.35 75.5 ;
        RECT 57.09 74.48 57.35 74.74 ;
        RECT 57.09 73.72 57.35 73.98 ;
        RECT 57.09 72.96 57.35 73.22 ;
        RECT 57.09 72.2 57.35 72.46 ;
        RECT 57.09 71.44 57.35 71.7 ;
        RECT 57.09 70.68 57.35 70.94 ;
        RECT 57.09 69.92 57.35 70.18 ;
        RECT 57.09 69.16 57.35 69.42 ;
        RECT 57.85 91.2 58.11 91.46 ;
        RECT 57.85 90.44 58.11 90.7 ;
        RECT 57.85 89.68 58.11 89.94 ;
        RECT 57.85 88.92 58.11 89.18 ;
        RECT 57.85 88.16 58.11 88.42 ;
        RECT 57.85 87.4 58.11 87.66 ;
        RECT 57.85 86.64 58.11 86.9 ;
        RECT 57.85 85.88 58.11 86.14 ;
        RECT 57.85 85.12 58.11 85.38 ;
        RECT 57.85 84.36 58.11 84.62 ;
        RECT 57.85 83.6 58.11 83.86 ;
        RECT 57.85 82.84 58.11 83.1 ;
        RECT 57.85 82.08 58.11 82.34 ;
        RECT 57.85 81.32 58.11 81.58 ;
        RECT 57.85 80.56 58.11 80.82 ;
        RECT 57.85 79.8 58.11 80.06 ;
        RECT 57.85 79.04 58.11 79.3 ;
        RECT 57.85 78.28 58.11 78.54 ;
        RECT 57.85 77.52 58.11 77.78 ;
        RECT 57.85 76.76 58.11 77.02 ;
        RECT 57.85 76 58.11 76.26 ;
        RECT 57.85 75.24 58.11 75.5 ;
        RECT 57.85 74.48 58.11 74.74 ;
        RECT 57.85 73.72 58.11 73.98 ;
        RECT 57.85 72.96 58.11 73.22 ;
        RECT 57.85 72.2 58.11 72.46 ;
        RECT 57.85 71.44 58.11 71.7 ;
        RECT 57.85 70.68 58.11 70.94 ;
        RECT 57.85 69.92 58.11 70.18 ;
        RECT 57.85 69.16 58.11 69.42 ;
        RECT 58.61 91.2 58.87 91.46 ;
        RECT 58.61 90.44 58.87 90.7 ;
        RECT 58.61 89.68 58.87 89.94 ;
        RECT 58.61 88.92 58.87 89.18 ;
        RECT 58.61 88.16 58.87 88.42 ;
        RECT 58.61 87.4 58.87 87.66 ;
        RECT 58.61 86.64 58.87 86.9 ;
        RECT 58.61 85.88 58.87 86.14 ;
        RECT 58.61 85.12 58.87 85.38 ;
        RECT 58.61 84.36 58.87 84.62 ;
        RECT 58.61 83.6 58.87 83.86 ;
        RECT 58.61 82.84 58.87 83.1 ;
        RECT 58.61 82.08 58.87 82.34 ;
        RECT 58.61 81.32 58.87 81.58 ;
        RECT 58.61 80.56 58.87 80.82 ;
        RECT 58.61 79.8 58.87 80.06 ;
        RECT 58.61 79.04 58.87 79.3 ;
        RECT 58.61 78.28 58.87 78.54 ;
        RECT 58.61 77.52 58.87 77.78 ;
        RECT 58.61 76.76 58.87 77.02 ;
        RECT 58.61 76 58.87 76.26 ;
        RECT 58.61 75.24 58.87 75.5 ;
        RECT 58.61 74.48 58.87 74.74 ;
        RECT 58.61 73.72 58.87 73.98 ;
        RECT 58.61 72.96 58.87 73.22 ;
        RECT 58.61 72.2 58.87 72.46 ;
        RECT 58.61 71.44 58.87 71.7 ;
        RECT 58.61 70.68 58.87 70.94 ;
        RECT 58.61 69.92 58.87 70.18 ;
        RECT 58.61 69.16 58.87 69.42 ;
        RECT 59.37 91.2 59.63 91.46 ;
        RECT 59.37 90.44 59.63 90.7 ;
        RECT 59.37 89.68 59.63 89.94 ;
        RECT 59.37 88.92 59.63 89.18 ;
        RECT 59.37 88.16 59.63 88.42 ;
        RECT 59.37 87.4 59.63 87.66 ;
        RECT 59.37 86.64 59.63 86.9 ;
        RECT 59.37 85.88 59.63 86.14 ;
        RECT 59.37 85.12 59.63 85.38 ;
        RECT 59.37 84.36 59.63 84.62 ;
        RECT 59.37 83.6 59.63 83.86 ;
        RECT 59.37 82.84 59.63 83.1 ;
        RECT 59.37 82.08 59.63 82.34 ;
        RECT 59.37 81.32 59.63 81.58 ;
        RECT 59.37 80.56 59.63 80.82 ;
        RECT 59.37 79.8 59.63 80.06 ;
        RECT 59.37 79.04 59.63 79.3 ;
        RECT 59.37 78.28 59.63 78.54 ;
        RECT 59.37 77.52 59.63 77.78 ;
        RECT 59.37 76.76 59.63 77.02 ;
        RECT 59.37 76 59.63 76.26 ;
        RECT 59.37 75.24 59.63 75.5 ;
        RECT 59.37 74.48 59.63 74.74 ;
        RECT 59.37 73.72 59.63 73.98 ;
        RECT 59.37 72.96 59.63 73.22 ;
        RECT 59.37 72.2 59.63 72.46 ;
        RECT 59.37 71.44 59.63 71.7 ;
        RECT 59.37 70.68 59.63 70.94 ;
        RECT 59.37 69.92 59.63 70.18 ;
        RECT 59.37 69.16 59.63 69.42 ;
        RECT 60.13 91.2 60.39 91.46 ;
        RECT 60.13 90.44 60.39 90.7 ;
        RECT 60.13 89.68 60.39 89.94 ;
        RECT 60.13 88.92 60.39 89.18 ;
        RECT 60.13 88.16 60.39 88.42 ;
        RECT 60.13 87.4 60.39 87.66 ;
        RECT 60.13 86.64 60.39 86.9 ;
        RECT 60.13 85.88 60.39 86.14 ;
        RECT 60.13 85.12 60.39 85.38 ;
        RECT 60.13 84.36 60.39 84.62 ;
        RECT 60.13 83.6 60.39 83.86 ;
        RECT 60.13 82.84 60.39 83.1 ;
        RECT 60.13 82.08 60.39 82.34 ;
        RECT 60.13 81.32 60.39 81.58 ;
        RECT 60.13 80.56 60.39 80.82 ;
        RECT 60.13 79.8 60.39 80.06 ;
        RECT 60.13 79.04 60.39 79.3 ;
        RECT 60.13 78.28 60.39 78.54 ;
        RECT 60.13 77.52 60.39 77.78 ;
        RECT 60.13 76.76 60.39 77.02 ;
        RECT 60.13 76 60.39 76.26 ;
        RECT 60.13 75.24 60.39 75.5 ;
        RECT 60.13 74.48 60.39 74.74 ;
        RECT 60.13 73.72 60.39 73.98 ;
        RECT 60.13 72.96 60.39 73.22 ;
        RECT 60.13 72.2 60.39 72.46 ;
        RECT 60.13 71.44 60.39 71.7 ;
        RECT 60.13 70.68 60.39 70.94 ;
        RECT 60.13 69.92 60.39 70.18 ;
        RECT 60.13 69.16 60.39 69.42 ;
        RECT 60.89 91.2 61.15 91.46 ;
        RECT 60.89 90.44 61.15 90.7 ;
        RECT 60.89 89.68 61.15 89.94 ;
        RECT 60.89 88.92 61.15 89.18 ;
        RECT 60.89 88.16 61.15 88.42 ;
        RECT 60.89 87.4 61.15 87.66 ;
        RECT 60.89 86.64 61.15 86.9 ;
        RECT 60.89 85.88 61.15 86.14 ;
        RECT 60.89 85.12 61.15 85.38 ;
        RECT 60.89 84.36 61.15 84.62 ;
        RECT 60.89 83.6 61.15 83.86 ;
        RECT 60.89 82.84 61.15 83.1 ;
        RECT 60.89 82.08 61.15 82.34 ;
        RECT 60.89 81.32 61.15 81.58 ;
        RECT 60.89 80.56 61.15 80.82 ;
        RECT 60.89 79.8 61.15 80.06 ;
        RECT 60.89 79.04 61.15 79.3 ;
        RECT 60.89 78.28 61.15 78.54 ;
        RECT 60.89 77.52 61.15 77.78 ;
        RECT 60.89 76.76 61.15 77.02 ;
        RECT 60.89 76 61.15 76.26 ;
        RECT 60.89 75.24 61.15 75.5 ;
        RECT 60.89 74.48 61.15 74.74 ;
        RECT 60.89 73.72 61.15 73.98 ;
        RECT 60.89 72.96 61.15 73.22 ;
        RECT 60.89 72.2 61.15 72.46 ;
        RECT 60.89 71.44 61.15 71.7 ;
        RECT 60.89 70.68 61.15 70.94 ;
        RECT 60.89 69.92 61.15 70.18 ;
        RECT 60.89 69.16 61.15 69.42 ;
        RECT 61.65 91.2 61.91 91.46 ;
        RECT 61.65 90.44 61.91 90.7 ;
        RECT 61.65 89.68 61.91 89.94 ;
        RECT 61.65 88.92 61.91 89.18 ;
        RECT 61.65 88.16 61.91 88.42 ;
        RECT 61.65 87.4 61.91 87.66 ;
        RECT 61.65 86.64 61.91 86.9 ;
        RECT 61.65 85.88 61.91 86.14 ;
        RECT 61.65 85.12 61.91 85.38 ;
        RECT 61.65 84.36 61.91 84.62 ;
        RECT 61.65 83.6 61.91 83.86 ;
        RECT 61.65 82.84 61.91 83.1 ;
        RECT 61.65 82.08 61.91 82.34 ;
        RECT 61.65 81.32 61.91 81.58 ;
        RECT 61.65 80.56 61.91 80.82 ;
        RECT 61.65 79.8 61.91 80.06 ;
        RECT 61.65 79.04 61.91 79.3 ;
        RECT 61.65 78.28 61.91 78.54 ;
        RECT 61.65 77.52 61.91 77.78 ;
        RECT 61.65 76.76 61.91 77.02 ;
        RECT 61.65 76 61.91 76.26 ;
        RECT 61.65 75.24 61.91 75.5 ;
        RECT 61.65 74.48 61.91 74.74 ;
        RECT 61.65 73.72 61.91 73.98 ;
        RECT 61.65 72.96 61.91 73.22 ;
        RECT 61.65 72.2 61.91 72.46 ;
        RECT 61.65 71.44 61.91 71.7 ;
        RECT 61.65 70.68 61.91 70.94 ;
        RECT 61.65 69.92 61.91 70.18 ;
        RECT 61.65 69.16 61.91 69.42 ;
        RECT 62.41 91.2 62.67 91.46 ;
        RECT 62.41 90.44 62.67 90.7 ;
        RECT 62.41 89.68 62.67 89.94 ;
        RECT 62.41 88.92 62.67 89.18 ;
        RECT 62.41 88.16 62.67 88.42 ;
        RECT 62.41 87.4 62.67 87.66 ;
        RECT 62.41 86.64 62.67 86.9 ;
        RECT 62.41 85.88 62.67 86.14 ;
        RECT 62.41 85.12 62.67 85.38 ;
        RECT 62.41 84.36 62.67 84.62 ;
        RECT 62.41 83.6 62.67 83.86 ;
        RECT 62.41 82.84 62.67 83.1 ;
        RECT 62.41 82.08 62.67 82.34 ;
        RECT 62.41 81.32 62.67 81.58 ;
        RECT 62.41 80.56 62.67 80.82 ;
        RECT 62.41 79.8 62.67 80.06 ;
        RECT 62.41 79.04 62.67 79.3 ;
        RECT 62.41 78.28 62.67 78.54 ;
        RECT 62.41 77.52 62.67 77.78 ;
        RECT 62.41 76.76 62.67 77.02 ;
        RECT 62.41 76 62.67 76.26 ;
        RECT 62.41 75.24 62.67 75.5 ;
        RECT 62.41 74.48 62.67 74.74 ;
        RECT 62.41 73.72 62.67 73.98 ;
        RECT 62.41 72.96 62.67 73.22 ;
        RECT 62.41 72.2 62.67 72.46 ;
        RECT 62.41 71.44 62.67 71.7 ;
        RECT 62.41 70.68 62.67 70.94 ;
        RECT 62.41 69.92 62.67 70.18 ;
        RECT 62.41 69.16 62.67 69.42 ;
        RECT 63.17 91.2 63.43 91.46 ;
        RECT 63.17 90.44 63.43 90.7 ;
        RECT 63.17 89.68 63.43 89.94 ;
        RECT 63.17 88.92 63.43 89.18 ;
        RECT 63.17 88.16 63.43 88.42 ;
        RECT 63.17 87.4 63.43 87.66 ;
        RECT 63.17 86.64 63.43 86.9 ;
        RECT 63.17 85.88 63.43 86.14 ;
        RECT 63.17 85.12 63.43 85.38 ;
        RECT 63.17 84.36 63.43 84.62 ;
        RECT 63.17 83.6 63.43 83.86 ;
        RECT 63.17 82.84 63.43 83.1 ;
        RECT 63.17 82.08 63.43 82.34 ;
        RECT 63.17 81.32 63.43 81.58 ;
        RECT 63.17 80.56 63.43 80.82 ;
        RECT 63.17 79.8 63.43 80.06 ;
        RECT 63.17 79.04 63.43 79.3 ;
        RECT 63.17 78.28 63.43 78.54 ;
        RECT 63.17 77.52 63.43 77.78 ;
        RECT 63.17 76.76 63.43 77.02 ;
        RECT 63.17 76 63.43 76.26 ;
        RECT 63.17 75.24 63.43 75.5 ;
        RECT 63.17 74.48 63.43 74.74 ;
        RECT 63.17 73.72 63.43 73.98 ;
        RECT 63.17 72.96 63.43 73.22 ;
        RECT 63.17 72.2 63.43 72.46 ;
        RECT 63.17 71.44 63.43 71.7 ;
        RECT 63.17 70.68 63.43 70.94 ;
        RECT 63.17 69.92 63.43 70.18 ;
        RECT 63.17 69.16 63.43 69.42 ;
        RECT 63.93 91.2 64.19 91.46 ;
        RECT 63.93 90.44 64.19 90.7 ;
        RECT 63.93 89.68 64.19 89.94 ;
        RECT 63.93 88.92 64.19 89.18 ;
        RECT 63.93 88.16 64.19 88.42 ;
        RECT 63.93 87.4 64.19 87.66 ;
        RECT 63.93 86.64 64.19 86.9 ;
        RECT 63.93 85.88 64.19 86.14 ;
        RECT 63.93 85.12 64.19 85.38 ;
        RECT 63.93 84.36 64.19 84.62 ;
        RECT 63.93 83.6 64.19 83.86 ;
        RECT 63.93 82.84 64.19 83.1 ;
        RECT 63.93 82.08 64.19 82.34 ;
        RECT 63.93 81.32 64.19 81.58 ;
        RECT 63.93 80.56 64.19 80.82 ;
        RECT 63.93 79.8 64.19 80.06 ;
        RECT 63.93 79.04 64.19 79.3 ;
        RECT 63.93 78.28 64.19 78.54 ;
        RECT 63.93 77.52 64.19 77.78 ;
        RECT 63.93 76.76 64.19 77.02 ;
        RECT 63.93 76 64.19 76.26 ;
        RECT 63.93 75.24 64.19 75.5 ;
        RECT 63.93 74.48 64.19 74.74 ;
        RECT 63.93 73.72 64.19 73.98 ;
        RECT 63.93 72.96 64.19 73.22 ;
        RECT 63.93 72.2 64.19 72.46 ;
        RECT 63.93 71.44 64.19 71.7 ;
        RECT 63.93 70.68 64.19 70.94 ;
        RECT 63.93 69.92 64.19 70.18 ;
        RECT 63.93 69.16 64.19 69.42 ;
        RECT 64.69 91.2 64.95 91.46 ;
        RECT 64.69 90.44 64.95 90.7 ;
        RECT 64.69 89.68 64.95 89.94 ;
        RECT 64.69 88.92 64.95 89.18 ;
        RECT 64.69 88.16 64.95 88.42 ;
        RECT 64.69 87.4 64.95 87.66 ;
        RECT 64.69 86.64 64.95 86.9 ;
        RECT 64.69 85.88 64.95 86.14 ;
        RECT 64.69 85.12 64.95 85.38 ;
        RECT 64.69 84.36 64.95 84.62 ;
        RECT 64.69 83.6 64.95 83.86 ;
        RECT 64.69 82.84 64.95 83.1 ;
        RECT 64.69 82.08 64.95 82.34 ;
        RECT 64.69 81.32 64.95 81.58 ;
        RECT 64.69 80.56 64.95 80.82 ;
        RECT 64.69 79.8 64.95 80.06 ;
        RECT 64.69 79.04 64.95 79.3 ;
        RECT 64.69 78.28 64.95 78.54 ;
        RECT 64.69 77.52 64.95 77.78 ;
        RECT 64.69 76.76 64.95 77.02 ;
        RECT 64.69 76 64.95 76.26 ;
        RECT 64.69 75.24 64.95 75.5 ;
        RECT 64.69 74.48 64.95 74.74 ;
        RECT 64.69 73.72 64.95 73.98 ;
        RECT 64.69 72.96 64.95 73.22 ;
        RECT 64.69 72.2 64.95 72.46 ;
        RECT 64.69 71.44 64.95 71.7 ;
        RECT 64.69 70.68 64.95 70.94 ;
        RECT 64.69 69.92 64.95 70.18 ;
        RECT 64.69 69.16 64.95 69.42 ;
        RECT 65.45 91.2 65.71 91.46 ;
        RECT 65.45 90.44 65.71 90.7 ;
        RECT 65.45 89.68 65.71 89.94 ;
        RECT 65.45 88.92 65.71 89.18 ;
        RECT 65.45 88.16 65.71 88.42 ;
        RECT 65.45 87.4 65.71 87.66 ;
        RECT 65.45 86.64 65.71 86.9 ;
        RECT 65.45 85.88 65.71 86.14 ;
        RECT 65.45 85.12 65.71 85.38 ;
        RECT 65.45 84.36 65.71 84.62 ;
        RECT 65.45 83.6 65.71 83.86 ;
        RECT 65.45 82.84 65.71 83.1 ;
        RECT 65.45 82.08 65.71 82.34 ;
        RECT 65.45 81.32 65.71 81.58 ;
        RECT 65.45 80.56 65.71 80.82 ;
        RECT 65.45 79.8 65.71 80.06 ;
        RECT 65.45 79.04 65.71 79.3 ;
        RECT 65.45 78.28 65.71 78.54 ;
        RECT 65.45 77.52 65.71 77.78 ;
        RECT 65.45 76.76 65.71 77.02 ;
        RECT 65.45 76 65.71 76.26 ;
        RECT 65.45 75.24 65.71 75.5 ;
        RECT 65.45 74.48 65.71 74.74 ;
        RECT 65.45 73.72 65.71 73.98 ;
        RECT 65.45 72.96 65.71 73.22 ;
        RECT 65.45 72.2 65.71 72.46 ;
        RECT 65.45 71.44 65.71 71.7 ;
        RECT 65.45 70.68 65.71 70.94 ;
        RECT 65.45 69.92 65.71 70.18 ;
        RECT 65.45 69.16 65.71 69.42 ;
        RECT 66.21 91.2 66.47 91.46 ;
        RECT 66.21 90.44 66.47 90.7 ;
        RECT 66.21 89.68 66.47 89.94 ;
        RECT 66.21 88.92 66.47 89.18 ;
        RECT 66.21 88.16 66.47 88.42 ;
        RECT 66.21 87.4 66.47 87.66 ;
        RECT 66.21 86.64 66.47 86.9 ;
        RECT 66.21 85.88 66.47 86.14 ;
        RECT 66.21 85.12 66.47 85.38 ;
        RECT 66.21 84.36 66.47 84.62 ;
        RECT 66.21 83.6 66.47 83.86 ;
        RECT 66.21 82.84 66.47 83.1 ;
        RECT 66.21 82.08 66.47 82.34 ;
        RECT 66.21 81.32 66.47 81.58 ;
        RECT 66.21 80.56 66.47 80.82 ;
        RECT 66.21 79.8 66.47 80.06 ;
        RECT 66.21 79.04 66.47 79.3 ;
        RECT 66.21 78.28 66.47 78.54 ;
        RECT 66.21 77.52 66.47 77.78 ;
        RECT 66.21 76.76 66.47 77.02 ;
        RECT 66.21 76 66.47 76.26 ;
        RECT 66.21 75.24 66.47 75.5 ;
        RECT 66.21 74.48 66.47 74.74 ;
        RECT 66.21 73.72 66.47 73.98 ;
        RECT 66.21 72.96 66.47 73.22 ;
        RECT 66.21 72.2 66.47 72.46 ;
        RECT 66.21 71.44 66.47 71.7 ;
        RECT 66.21 70.68 66.47 70.94 ;
        RECT 66.21 69.92 66.47 70.18 ;
        RECT 66.21 69.16 66.47 69.42 ;
        RECT 66.97 91.2 67.23 91.46 ;
        RECT 66.97 90.44 67.23 90.7 ;
        RECT 66.97 89.68 67.23 89.94 ;
        RECT 66.97 88.92 67.23 89.18 ;
        RECT 66.97 88.16 67.23 88.42 ;
        RECT 66.97 87.4 67.23 87.66 ;
        RECT 66.97 86.64 67.23 86.9 ;
        RECT 66.97 85.88 67.23 86.14 ;
        RECT 66.97 85.12 67.23 85.38 ;
        RECT 66.97 84.36 67.23 84.62 ;
        RECT 66.97 83.6 67.23 83.86 ;
        RECT 66.97 82.84 67.23 83.1 ;
        RECT 66.97 82.08 67.23 82.34 ;
        RECT 66.97 81.32 67.23 81.58 ;
        RECT 66.97 80.56 67.23 80.82 ;
        RECT 66.97 79.8 67.23 80.06 ;
        RECT 66.97 79.04 67.23 79.3 ;
        RECT 66.97 78.28 67.23 78.54 ;
        RECT 66.97 77.52 67.23 77.78 ;
        RECT 66.97 76.76 67.23 77.02 ;
        RECT 66.97 76 67.23 76.26 ;
        RECT 66.97 75.24 67.23 75.5 ;
        RECT 66.97 74.48 67.23 74.74 ;
        RECT 66.97 73.72 67.23 73.98 ;
        RECT 66.97 72.96 67.23 73.22 ;
        RECT 66.97 72.2 67.23 72.46 ;
        RECT 66.97 71.44 67.23 71.7 ;
        RECT 66.97 70.68 67.23 70.94 ;
        RECT 66.97 69.92 67.23 70.18 ;
        RECT 66.97 69.16 67.23 69.42 ;
        RECT 67.73 91.2 67.99 91.46 ;
        RECT 67.73 90.44 67.99 90.7 ;
        RECT 67.73 89.68 67.99 89.94 ;
        RECT 67.73 88.92 67.99 89.18 ;
        RECT 67.73 88.16 67.99 88.42 ;
        RECT 67.73 87.4 67.99 87.66 ;
        RECT 67.73 86.64 67.99 86.9 ;
        RECT 67.73 85.88 67.99 86.14 ;
        RECT 67.73 85.12 67.99 85.38 ;
        RECT 67.73 84.36 67.99 84.62 ;
        RECT 67.73 83.6 67.99 83.86 ;
        RECT 67.73 82.84 67.99 83.1 ;
        RECT 67.73 82.08 67.99 82.34 ;
        RECT 67.73 81.32 67.99 81.58 ;
        RECT 67.73 80.56 67.99 80.82 ;
        RECT 67.73 79.8 67.99 80.06 ;
        RECT 67.73 79.04 67.99 79.3 ;
        RECT 67.73 78.28 67.99 78.54 ;
        RECT 67.73 77.52 67.99 77.78 ;
        RECT 67.73 76.76 67.99 77.02 ;
        RECT 67.73 76 67.99 76.26 ;
        RECT 67.73 75.24 67.99 75.5 ;
        RECT 67.73 74.48 67.99 74.74 ;
        RECT 67.73 73.72 67.99 73.98 ;
        RECT 67.73 72.96 67.99 73.22 ;
        RECT 67.73 72.2 67.99 72.46 ;
        RECT 67.73 71.44 67.99 71.7 ;
        RECT 67.73 70.68 67.99 70.94 ;
        RECT 67.73 69.92 67.99 70.18 ;
        RECT 67.73 69.16 67.99 69.42 ;
        RECT 68.49 91.2 68.75 91.46 ;
        RECT 68.49 90.44 68.75 90.7 ;
        RECT 68.49 89.68 68.75 89.94 ;
        RECT 68.49 88.92 68.75 89.18 ;
        RECT 68.49 88.16 68.75 88.42 ;
        RECT 68.49 87.4 68.75 87.66 ;
        RECT 68.49 86.64 68.75 86.9 ;
        RECT 68.49 85.88 68.75 86.14 ;
        RECT 68.49 85.12 68.75 85.38 ;
        RECT 68.49 84.36 68.75 84.62 ;
        RECT 68.49 83.6 68.75 83.86 ;
        RECT 68.49 82.84 68.75 83.1 ;
        RECT 68.49 82.08 68.75 82.34 ;
        RECT 68.49 81.32 68.75 81.58 ;
        RECT 68.49 80.56 68.75 80.82 ;
        RECT 68.49 79.8 68.75 80.06 ;
        RECT 68.49 79.04 68.75 79.3 ;
        RECT 68.49 78.28 68.75 78.54 ;
        RECT 68.49 77.52 68.75 77.78 ;
        RECT 68.49 76.76 68.75 77.02 ;
        RECT 68.49 76 68.75 76.26 ;
        RECT 68.49 75.24 68.75 75.5 ;
        RECT 68.49 74.48 68.75 74.74 ;
        RECT 68.49 73.72 68.75 73.98 ;
        RECT 68.49 72.96 68.75 73.22 ;
        RECT 68.49 72.2 68.75 72.46 ;
        RECT 68.49 71.44 68.75 71.7 ;
        RECT 68.49 70.68 68.75 70.94 ;
        RECT 68.49 69.92 68.75 70.18 ;
        RECT 68.49 69.16 68.75 69.42 ;
        RECT 69.25 91.2 69.51 91.46 ;
        RECT 69.25 90.44 69.51 90.7 ;
        RECT 69.25 89.68 69.51 89.94 ;
        RECT 69.25 88.92 69.51 89.18 ;
        RECT 69.25 88.16 69.51 88.42 ;
        RECT 69.25 87.4 69.51 87.66 ;
        RECT 69.25 86.64 69.51 86.9 ;
        RECT 69.25 85.88 69.51 86.14 ;
        RECT 69.25 85.12 69.51 85.38 ;
        RECT 69.25 84.36 69.51 84.62 ;
        RECT 69.25 83.6 69.51 83.86 ;
        RECT 69.25 82.84 69.51 83.1 ;
        RECT 69.25 82.08 69.51 82.34 ;
        RECT 69.25 81.32 69.51 81.58 ;
        RECT 69.25 80.56 69.51 80.82 ;
        RECT 69.25 79.8 69.51 80.06 ;
        RECT 69.25 79.04 69.51 79.3 ;
        RECT 69.25 78.28 69.51 78.54 ;
        RECT 69.25 77.52 69.51 77.78 ;
        RECT 69.25 76.76 69.51 77.02 ;
        RECT 69.25 76 69.51 76.26 ;
        RECT 69.25 75.24 69.51 75.5 ;
        RECT 69.25 74.48 69.51 74.74 ;
        RECT 69.25 73.72 69.51 73.98 ;
        RECT 69.25 72.96 69.51 73.22 ;
        RECT 69.25 72.2 69.51 72.46 ;
        RECT 69.25 71.44 69.51 71.7 ;
        RECT 69.25 70.68 69.51 70.94 ;
        RECT 69.25 69.92 69.51 70.18 ;
        RECT 69.25 69.16 69.51 69.42 ;
        RECT 70.01 91.2 70.27 91.46 ;
        RECT 70.01 90.44 70.27 90.7 ;
        RECT 70.01 89.68 70.27 89.94 ;
        RECT 70.01 88.92 70.27 89.18 ;
        RECT 70.01 88.16 70.27 88.42 ;
        RECT 70.01 87.4 70.27 87.66 ;
        RECT 70.01 86.64 70.27 86.9 ;
        RECT 70.01 85.88 70.27 86.14 ;
        RECT 70.01 85.12 70.27 85.38 ;
        RECT 70.01 84.36 70.27 84.62 ;
        RECT 70.01 83.6 70.27 83.86 ;
        RECT 70.01 82.84 70.27 83.1 ;
        RECT 70.01 82.08 70.27 82.34 ;
        RECT 70.01 81.32 70.27 81.58 ;
        RECT 70.01 80.56 70.27 80.82 ;
        RECT 70.01 79.8 70.27 80.06 ;
        RECT 70.01 79.04 70.27 79.3 ;
        RECT 70.01 78.28 70.27 78.54 ;
        RECT 70.01 77.52 70.27 77.78 ;
        RECT 70.01 76.76 70.27 77.02 ;
        RECT 70.01 76 70.27 76.26 ;
        RECT 70.01 75.24 70.27 75.5 ;
        RECT 70.01 74.48 70.27 74.74 ;
        RECT 70.01 73.72 70.27 73.98 ;
        RECT 70.01 72.96 70.27 73.22 ;
        RECT 70.01 72.2 70.27 72.46 ;
        RECT 70.01 71.44 70.27 71.7 ;
        RECT 70.01 70.68 70.27 70.94 ;
        RECT 70.01 69.92 70.27 70.18 ;
        RECT 70.01 69.16 70.27 69.42 ;
        RECT 70.77 91.2 71.03 91.46 ;
        RECT 70.77 90.44 71.03 90.7 ;
        RECT 70.77 89.68 71.03 89.94 ;
        RECT 70.77 88.92 71.03 89.18 ;
        RECT 70.77 88.16 71.03 88.42 ;
        RECT 70.77 87.4 71.03 87.66 ;
        RECT 70.77 86.64 71.03 86.9 ;
        RECT 70.77 85.88 71.03 86.14 ;
        RECT 70.77 85.12 71.03 85.38 ;
        RECT 70.77 84.36 71.03 84.62 ;
        RECT 70.77 83.6 71.03 83.86 ;
        RECT 70.77 82.84 71.03 83.1 ;
        RECT 70.77 82.08 71.03 82.34 ;
        RECT 70.77 81.32 71.03 81.58 ;
        RECT 70.77 80.56 71.03 80.82 ;
        RECT 70.77 79.8 71.03 80.06 ;
        RECT 70.77 79.04 71.03 79.3 ;
        RECT 70.77 78.28 71.03 78.54 ;
        RECT 70.77 77.52 71.03 77.78 ;
        RECT 70.77 76.76 71.03 77.02 ;
        RECT 70.77 76 71.03 76.26 ;
        RECT 70.77 75.24 71.03 75.5 ;
        RECT 70.77 74.48 71.03 74.74 ;
        RECT 70.77 73.72 71.03 73.98 ;
        RECT 70.77 72.96 71.03 73.22 ;
        RECT 70.77 72.2 71.03 72.46 ;
        RECT 70.77 71.44 71.03 71.7 ;
        RECT 70.77 70.68 71.03 70.94 ;
        RECT 70.77 69.92 71.03 70.18 ;
        RECT 70.77 69.16 71.03 69.42 ;
        RECT 71.53 91.2 71.79 91.46 ;
        RECT 71.53 90.44 71.79 90.7 ;
        RECT 71.53 89.68 71.79 89.94 ;
        RECT 71.53 88.92 71.79 89.18 ;
        RECT 71.53 88.16 71.79 88.42 ;
        RECT 71.53 87.4 71.79 87.66 ;
        RECT 71.53 86.64 71.79 86.9 ;
        RECT 71.53 85.88 71.79 86.14 ;
        RECT 71.53 85.12 71.79 85.38 ;
        RECT 71.53 84.36 71.79 84.62 ;
        RECT 71.53 83.6 71.79 83.86 ;
        RECT 71.53 82.84 71.79 83.1 ;
        RECT 71.53 82.08 71.79 82.34 ;
        RECT 71.53 81.32 71.79 81.58 ;
        RECT 71.53 80.56 71.79 80.82 ;
        RECT 71.53 79.8 71.79 80.06 ;
        RECT 71.53 79.04 71.79 79.3 ;
        RECT 71.53 78.28 71.79 78.54 ;
        RECT 71.53 77.52 71.79 77.78 ;
        RECT 71.53 76.76 71.79 77.02 ;
        RECT 71.53 76 71.79 76.26 ;
        RECT 71.53 75.24 71.79 75.5 ;
        RECT 71.53 74.48 71.79 74.74 ;
        RECT 71.53 73.72 71.79 73.98 ;
        RECT 71.53 72.96 71.79 73.22 ;
        RECT 71.53 72.2 71.79 72.46 ;
        RECT 71.53 71.44 71.79 71.7 ;
        RECT 71.53 70.68 71.79 70.94 ;
        RECT 71.53 69.92 71.79 70.18 ;
        RECT 71.53 69.16 71.79 69.42 ;
        RECT 72.29 91.2 72.55 91.46 ;
        RECT 72.29 90.44 72.55 90.7 ;
        RECT 72.29 89.68 72.55 89.94 ;
        RECT 72.29 88.92 72.55 89.18 ;
        RECT 72.29 88.16 72.55 88.42 ;
        RECT 72.29 87.4 72.55 87.66 ;
        RECT 72.29 86.64 72.55 86.9 ;
        RECT 72.29 85.88 72.55 86.14 ;
        RECT 72.29 85.12 72.55 85.38 ;
        RECT 72.29 84.36 72.55 84.62 ;
        RECT 72.29 83.6 72.55 83.86 ;
        RECT 72.29 82.84 72.55 83.1 ;
        RECT 72.29 82.08 72.55 82.34 ;
        RECT 72.29 81.32 72.55 81.58 ;
        RECT 72.29 80.56 72.55 80.82 ;
        RECT 72.29 79.8 72.55 80.06 ;
        RECT 72.29 79.04 72.55 79.3 ;
        RECT 72.29 78.28 72.55 78.54 ;
        RECT 72.29 77.52 72.55 77.78 ;
        RECT 72.29 76.76 72.55 77.02 ;
        RECT 72.29 76 72.55 76.26 ;
        RECT 72.29 75.24 72.55 75.5 ;
        RECT 72.29 74.48 72.55 74.74 ;
        RECT 72.29 73.72 72.55 73.98 ;
        RECT 72.29 72.96 72.55 73.22 ;
        RECT 72.29 72.2 72.55 72.46 ;
        RECT 72.29 71.44 72.55 71.7 ;
        RECT 72.29 70.68 72.55 70.94 ;
        RECT 72.29 69.92 72.55 70.18 ;
        RECT 72.29 69.16 72.55 69.42 ;
        RECT 73.05 91.2 73.31 91.46 ;
        RECT 73.05 90.44 73.31 90.7 ;
        RECT 73.05 89.68 73.31 89.94 ;
        RECT 73.05 88.92 73.31 89.18 ;
        RECT 73.05 88.16 73.31 88.42 ;
        RECT 73.05 87.4 73.31 87.66 ;
        RECT 73.05 86.64 73.31 86.9 ;
        RECT 73.05 85.88 73.31 86.14 ;
        RECT 73.05 85.12 73.31 85.38 ;
        RECT 73.05 84.36 73.31 84.62 ;
        RECT 73.05 83.6 73.31 83.86 ;
        RECT 73.05 82.84 73.31 83.1 ;
        RECT 73.05 82.08 73.31 82.34 ;
        RECT 73.05 81.32 73.31 81.58 ;
        RECT 73.05 80.56 73.31 80.82 ;
        RECT 73.05 79.8 73.31 80.06 ;
        RECT 73.05 79.04 73.31 79.3 ;
        RECT 73.05 78.28 73.31 78.54 ;
        RECT 73.05 77.52 73.31 77.78 ;
        RECT 73.05 76.76 73.31 77.02 ;
        RECT 73.05 76 73.31 76.26 ;
        RECT 73.05 75.24 73.31 75.5 ;
        RECT 73.05 74.48 73.31 74.74 ;
        RECT 73.05 73.72 73.31 73.98 ;
        RECT 73.05 72.96 73.31 73.22 ;
        RECT 73.05 72.2 73.31 72.46 ;
        RECT 73.05 71.44 73.31 71.7 ;
        RECT 73.05 70.68 73.31 70.94 ;
        RECT 73.05 69.92 73.31 70.18 ;
        RECT 73.05 69.16 73.31 69.42 ;
        RECT 73.81 91.2 74.07 91.46 ;
        RECT 73.81 90.44 74.07 90.7 ;
        RECT 73.81 89.68 74.07 89.94 ;
        RECT 73.81 88.92 74.07 89.18 ;
        RECT 73.81 88.16 74.07 88.42 ;
        RECT 73.81 87.4 74.07 87.66 ;
        RECT 73.81 86.64 74.07 86.9 ;
        RECT 73.81 85.88 74.07 86.14 ;
        RECT 73.81 85.12 74.07 85.38 ;
        RECT 73.81 84.36 74.07 84.62 ;
        RECT 73.81 83.6 74.07 83.86 ;
        RECT 73.81 82.84 74.07 83.1 ;
        RECT 73.81 82.08 74.07 82.34 ;
        RECT 73.81 81.32 74.07 81.58 ;
        RECT 73.81 80.56 74.07 80.82 ;
        RECT 73.81 79.8 74.07 80.06 ;
        RECT 73.81 79.04 74.07 79.3 ;
        RECT 73.81 78.28 74.07 78.54 ;
        RECT 73.81 77.52 74.07 77.78 ;
        RECT 73.81 76.76 74.07 77.02 ;
        RECT 73.81 76 74.07 76.26 ;
        RECT 73.81 75.24 74.07 75.5 ;
        RECT 73.81 74.48 74.07 74.74 ;
        RECT 73.81 73.72 74.07 73.98 ;
        RECT 73.81 72.96 74.07 73.22 ;
        RECT 73.81 72.2 74.07 72.46 ;
        RECT 73.81 71.44 74.07 71.7 ;
        RECT 73.81 70.68 74.07 70.94 ;
        RECT 73.81 69.92 74.07 70.18 ;
        RECT 73.81 69.16 74.07 69.42 ;
        RECT 74.57 91.2 74.83 91.46 ;
        RECT 74.57 90.44 74.83 90.7 ;
        RECT 74.57 89.68 74.83 89.94 ;
        RECT 74.57 88.92 74.83 89.18 ;
        RECT 74.57 88.16 74.83 88.42 ;
        RECT 74.57 87.4 74.83 87.66 ;
        RECT 74.57 86.64 74.83 86.9 ;
        RECT 74.57 85.88 74.83 86.14 ;
        RECT 74.57 85.12 74.83 85.38 ;
        RECT 74.57 84.36 74.83 84.62 ;
        RECT 74.57 83.6 74.83 83.86 ;
        RECT 74.57 82.84 74.83 83.1 ;
        RECT 74.57 82.08 74.83 82.34 ;
        RECT 74.57 81.32 74.83 81.58 ;
        RECT 74.57 80.56 74.83 80.82 ;
        RECT 74.57 79.8 74.83 80.06 ;
        RECT 74.57 79.04 74.83 79.3 ;
        RECT 74.57 78.28 74.83 78.54 ;
        RECT 74.57 77.52 74.83 77.78 ;
        RECT 74.57 76.76 74.83 77.02 ;
        RECT 74.57 76 74.83 76.26 ;
        RECT 74.57 75.24 74.83 75.5 ;
        RECT 74.57 74.48 74.83 74.74 ;
        RECT 74.57 73.72 74.83 73.98 ;
        RECT 74.57 72.96 74.83 73.22 ;
        RECT 74.57 72.2 74.83 72.46 ;
        RECT 74.57 71.44 74.83 71.7 ;
        RECT 74.57 70.68 74.83 70.94 ;
        RECT 74.57 69.92 74.83 70.18 ;
        RECT 74.57 69.16 74.83 69.42 ;
        RECT 75.33 91.2 75.59 91.46 ;
        RECT 75.33 90.44 75.59 90.7 ;
        RECT 75.33 89.68 75.59 89.94 ;
        RECT 75.33 88.92 75.59 89.18 ;
        RECT 75.33 88.16 75.59 88.42 ;
        RECT 75.33 87.4 75.59 87.66 ;
        RECT 75.33 86.64 75.59 86.9 ;
        RECT 75.33 85.88 75.59 86.14 ;
        RECT 75.33 85.12 75.59 85.38 ;
        RECT 75.33 84.36 75.59 84.62 ;
        RECT 75.33 83.6 75.59 83.86 ;
        RECT 75.33 82.84 75.59 83.1 ;
        RECT 75.33 82.08 75.59 82.34 ;
        RECT 75.33 81.32 75.59 81.58 ;
        RECT 75.33 80.56 75.59 80.82 ;
        RECT 75.33 79.8 75.59 80.06 ;
        RECT 75.33 79.04 75.59 79.3 ;
        RECT 75.33 78.28 75.59 78.54 ;
        RECT 75.33 77.52 75.59 77.78 ;
        RECT 75.33 76.76 75.59 77.02 ;
        RECT 75.33 76 75.59 76.26 ;
        RECT 75.33 75.24 75.59 75.5 ;
        RECT 75.33 74.48 75.59 74.74 ;
        RECT 75.33 73.72 75.59 73.98 ;
        RECT 75.33 72.96 75.59 73.22 ;
        RECT 75.33 72.2 75.59 72.46 ;
        RECT 75.33 71.44 75.59 71.7 ;
        RECT 75.33 70.68 75.59 70.94 ;
        RECT 75.33 69.92 75.59 70.18 ;
        RECT 75.33 69.16 75.59 69.42 ;
        RECT 76.09 91.2 76.35 91.46 ;
        RECT 76.09 90.44 76.35 90.7 ;
        RECT 76.09 89.68 76.35 89.94 ;
        RECT 76.09 88.92 76.35 89.18 ;
        RECT 76.09 88.16 76.35 88.42 ;
        RECT 76.09 87.4 76.35 87.66 ;
        RECT 76.09 86.64 76.35 86.9 ;
        RECT 76.09 85.88 76.35 86.14 ;
        RECT 76.09 85.12 76.35 85.38 ;
        RECT 76.09 84.36 76.35 84.62 ;
        RECT 76.09 83.6 76.35 83.86 ;
        RECT 76.09 82.84 76.35 83.1 ;
        RECT 76.09 82.08 76.35 82.34 ;
        RECT 76.09 81.32 76.35 81.58 ;
        RECT 76.09 80.56 76.35 80.82 ;
        RECT 76.09 79.8 76.35 80.06 ;
        RECT 76.09 79.04 76.35 79.3 ;
        RECT 76.09 78.28 76.35 78.54 ;
        RECT 76.09 77.52 76.35 77.78 ;
        RECT 76.09 76.76 76.35 77.02 ;
        RECT 76.09 76 76.35 76.26 ;
        RECT 76.09 75.24 76.35 75.5 ;
        RECT 76.09 74.48 76.35 74.74 ;
        RECT 76.09 73.72 76.35 73.98 ;
        RECT 76.09 72.96 76.35 73.22 ;
        RECT 76.09 72.2 76.35 72.46 ;
        RECT 76.09 71.44 76.35 71.7 ;
        RECT 76.09 70.68 76.35 70.94 ;
        RECT 76.09 69.92 76.35 70.18 ;
        RECT 76.09 69.16 76.35 69.42 ;
        RECT 76.85 91.2 77.11 91.46 ;
        RECT 76.85 90.44 77.11 90.7 ;
        RECT 76.85 89.68 77.11 89.94 ;
        RECT 76.85 88.92 77.11 89.18 ;
        RECT 76.85 88.16 77.11 88.42 ;
        RECT 76.85 87.4 77.11 87.66 ;
        RECT 76.85 86.64 77.11 86.9 ;
        RECT 76.85 85.88 77.11 86.14 ;
        RECT 76.85 85.12 77.11 85.38 ;
        RECT 76.85 84.36 77.11 84.62 ;
        RECT 76.85 83.6 77.11 83.86 ;
        RECT 76.85 82.84 77.11 83.1 ;
        RECT 76.85 82.08 77.11 82.34 ;
        RECT 76.85 81.32 77.11 81.58 ;
        RECT 76.85 80.56 77.11 80.82 ;
        RECT 76.85 79.8 77.11 80.06 ;
        RECT 76.85 79.04 77.11 79.3 ;
        RECT 76.85 78.28 77.11 78.54 ;
        RECT 76.85 77.52 77.11 77.78 ;
        RECT 76.85 76.76 77.11 77.02 ;
        RECT 76.85 76 77.11 76.26 ;
        RECT 76.85 75.24 77.11 75.5 ;
        RECT 76.85 74.48 77.11 74.74 ;
        RECT 76.85 73.72 77.11 73.98 ;
        RECT 76.85 72.96 77.11 73.22 ;
        RECT 76.85 72.2 77.11 72.46 ;
        RECT 76.85 71.44 77.11 71.7 ;
        RECT 76.85 70.68 77.11 70.94 ;
        RECT 76.85 69.92 77.11 70.18 ;
        RECT 76.85 69.16 77.11 69.42 ;
        RECT 77.61 91.2 77.87 91.46 ;
        RECT 77.61 90.44 77.87 90.7 ;
        RECT 77.61 89.68 77.87 89.94 ;
        RECT 77.61 88.92 77.87 89.18 ;
        RECT 77.61 88.16 77.87 88.42 ;
        RECT 77.61 87.4 77.87 87.66 ;
        RECT 77.61 86.64 77.87 86.9 ;
        RECT 77.61 85.88 77.87 86.14 ;
        RECT 77.61 85.12 77.87 85.38 ;
        RECT 77.61 84.36 77.87 84.62 ;
        RECT 77.61 83.6 77.87 83.86 ;
        RECT 77.61 82.84 77.87 83.1 ;
        RECT 77.61 82.08 77.87 82.34 ;
        RECT 77.61 81.32 77.87 81.58 ;
        RECT 77.61 80.56 77.87 80.82 ;
        RECT 77.61 79.8 77.87 80.06 ;
        RECT 77.61 79.04 77.87 79.3 ;
        RECT 77.61 78.28 77.87 78.54 ;
        RECT 77.61 77.52 77.87 77.78 ;
        RECT 77.61 76.76 77.87 77.02 ;
        RECT 77.61 76 77.87 76.26 ;
        RECT 77.61 75.24 77.87 75.5 ;
        RECT 77.61 74.48 77.87 74.74 ;
        RECT 77.61 73.72 77.87 73.98 ;
        RECT 77.61 72.96 77.87 73.22 ;
        RECT 77.61 72.2 77.87 72.46 ;
        RECT 77.61 71.44 77.87 71.7 ;
        RECT 77.61 70.68 77.87 70.94 ;
        RECT 77.61 69.92 77.87 70.18 ;
        RECT 77.61 69.16 77.87 69.42 ;
        RECT 78.37 91.2 78.63 91.46 ;
        RECT 78.37 90.44 78.63 90.7 ;
        RECT 78.37 89.68 78.63 89.94 ;
        RECT 78.37 88.92 78.63 89.18 ;
        RECT 78.37 88.16 78.63 88.42 ;
        RECT 78.37 87.4 78.63 87.66 ;
        RECT 78.37 86.64 78.63 86.9 ;
        RECT 78.37 85.88 78.63 86.14 ;
        RECT 78.37 85.12 78.63 85.38 ;
        RECT 78.37 84.36 78.63 84.62 ;
        RECT 78.37 83.6 78.63 83.86 ;
        RECT 78.37 82.84 78.63 83.1 ;
        RECT 78.37 82.08 78.63 82.34 ;
        RECT 78.37 81.32 78.63 81.58 ;
        RECT 78.37 80.56 78.63 80.82 ;
        RECT 78.37 79.8 78.63 80.06 ;
        RECT 78.37 79.04 78.63 79.3 ;
        RECT 78.37 78.28 78.63 78.54 ;
        RECT 78.37 77.52 78.63 77.78 ;
        RECT 78.37 76.76 78.63 77.02 ;
        RECT 78.37 76 78.63 76.26 ;
        RECT 78.37 75.24 78.63 75.5 ;
        RECT 78.37 74.48 78.63 74.74 ;
        RECT 78.37 73.72 78.63 73.98 ;
        RECT 78.37 72.96 78.63 73.22 ;
        RECT 78.37 72.2 78.63 72.46 ;
        RECT 78.37 71.44 78.63 71.7 ;
        RECT 78.37 70.68 78.63 70.94 ;
        RECT 78.37 69.92 78.63 70.18 ;
        RECT 78.37 69.16 78.63 69.42 ;
        RECT 79.13 91.2 79.39 91.46 ;
        RECT 79.13 90.44 79.39 90.7 ;
        RECT 79.13 89.68 79.39 89.94 ;
        RECT 79.13 88.92 79.39 89.18 ;
        RECT 79.13 88.16 79.39 88.42 ;
        RECT 79.13 87.4 79.39 87.66 ;
        RECT 79.13 86.64 79.39 86.9 ;
        RECT 79.13 85.88 79.39 86.14 ;
        RECT 79.13 85.12 79.39 85.38 ;
        RECT 79.13 84.36 79.39 84.62 ;
        RECT 79.13 83.6 79.39 83.86 ;
        RECT 79.13 82.84 79.39 83.1 ;
        RECT 79.13 82.08 79.39 82.34 ;
        RECT 79.13 81.32 79.39 81.58 ;
        RECT 79.13 80.56 79.39 80.82 ;
        RECT 79.13 79.8 79.39 80.06 ;
        RECT 79.13 79.04 79.39 79.3 ;
        RECT 79.13 78.28 79.39 78.54 ;
        RECT 79.13 77.52 79.39 77.78 ;
        RECT 79.13 76.76 79.39 77.02 ;
        RECT 79.13 76 79.39 76.26 ;
        RECT 79.13 75.24 79.39 75.5 ;
        RECT 79.13 74.48 79.39 74.74 ;
        RECT 79.13 73.72 79.39 73.98 ;
        RECT 79.13 72.96 79.39 73.22 ;
        RECT 79.13 72.2 79.39 72.46 ;
        RECT 79.13 71.44 79.39 71.7 ;
        RECT 79.13 70.68 79.39 70.94 ;
        RECT 79.13 69.92 79.39 70.18 ;
        RECT 79.13 69.16 79.39 69.42 ;
        RECT 79.89 91.2 80.15 91.46 ;
        RECT 79.89 90.44 80.15 90.7 ;
        RECT 79.89 89.68 80.15 89.94 ;
        RECT 79.89 88.92 80.15 89.18 ;
        RECT 79.89 88.16 80.15 88.42 ;
        RECT 79.89 87.4 80.15 87.66 ;
        RECT 79.89 86.64 80.15 86.9 ;
        RECT 79.89 85.88 80.15 86.14 ;
        RECT 79.89 85.12 80.15 85.38 ;
        RECT 79.89 84.36 80.15 84.62 ;
        RECT 79.89 83.6 80.15 83.86 ;
        RECT 79.89 82.84 80.15 83.1 ;
        RECT 79.89 82.08 80.15 82.34 ;
        RECT 79.89 81.32 80.15 81.58 ;
        RECT 79.89 80.56 80.15 80.82 ;
        RECT 79.89 79.8 80.15 80.06 ;
        RECT 79.89 79.04 80.15 79.3 ;
        RECT 79.89 78.28 80.15 78.54 ;
        RECT 79.89 77.52 80.15 77.78 ;
        RECT 79.89 76.76 80.15 77.02 ;
        RECT 79.89 76 80.15 76.26 ;
        RECT 79.89 75.24 80.15 75.5 ;
        RECT 79.89 74.48 80.15 74.74 ;
        RECT 79.89 73.72 80.15 73.98 ;
        RECT 79.89 72.96 80.15 73.22 ;
        RECT 79.89 72.2 80.15 72.46 ;
        RECT 79.89 71.44 80.15 71.7 ;
        RECT 79.89 70.68 80.15 70.94 ;
        RECT 79.89 69.92 80.15 70.18 ;
        RECT 79.89 69.16 80.15 69.42 ;
        RECT 29.73 83.6 29.99 83.86 ;
        RECT 29.73 82.84 29.99 83.1 ;
        RECT 29.73 82.08 29.99 82.34 ;
        RECT 29.73 81.32 29.99 81.58 ;
        RECT 29.73 80.56 29.99 80.82 ;
        RECT 29.73 79.8 29.99 80.06 ;
        RECT 29.73 79.04 29.99 79.3 ;
        RECT 29.73 78.28 29.99 78.54 ;
        RECT 29.73 77.52 29.99 77.78 ;
        RECT 29.73 76.76 29.99 77.02 ;
        RECT 29.73 76 29.99 76.26 ;
        RECT 29.73 75.24 29.99 75.5 ;
        RECT 29.73 74.48 29.99 74.74 ;
        RECT 29.73 73.72 29.99 73.98 ;
        RECT 29.73 72.96 29.99 73.22 ;
        RECT 29.73 72.2 29.99 72.46 ;
        RECT 29.73 71.44 29.99 71.7 ;
        RECT 29.73 70.68 29.99 70.94 ;
        RECT 29.73 69.92 29.99 70.18 ;
        RECT 29.73 69.16 29.99 69.42 ;
        RECT 30.49 91.2 30.75 91.46 ;
        RECT 30.49 90.44 30.75 90.7 ;
        RECT 30.49 89.68 30.75 89.94 ;
        RECT 30.49 88.92 30.75 89.18 ;
        RECT 30.49 88.16 30.75 88.42 ;
        RECT 30.49 87.4 30.75 87.66 ;
        RECT 30.49 86.64 30.75 86.9 ;
        RECT 30.49 85.88 30.75 86.14 ;
        RECT 30.49 85.12 30.75 85.38 ;
        RECT 30.49 84.36 30.75 84.62 ;
        RECT 30.49 83.6 30.75 83.86 ;
        RECT 30.49 82.84 30.75 83.1 ;
        RECT 30.49 82.08 30.75 82.34 ;
        RECT 30.49 81.32 30.75 81.58 ;
        RECT 30.49 80.56 30.75 80.82 ;
        RECT 30.49 79.8 30.75 80.06 ;
        RECT 30.49 79.04 30.75 79.3 ;
        RECT 30.49 78.28 30.75 78.54 ;
        RECT 30.49 77.52 30.75 77.78 ;
        RECT 30.49 76.76 30.75 77.02 ;
        RECT 30.49 76 30.75 76.26 ;
        RECT 30.49 75.24 30.75 75.5 ;
        RECT 30.49 74.48 30.75 74.74 ;
        RECT 30.49 73.72 30.75 73.98 ;
        RECT 30.49 72.96 30.75 73.22 ;
        RECT 30.49 72.2 30.75 72.46 ;
        RECT 30.49 71.44 30.75 71.7 ;
        RECT 30.49 70.68 30.75 70.94 ;
        RECT 30.49 69.92 30.75 70.18 ;
        RECT 30.49 69.16 30.75 69.42 ;
        RECT 31.25 91.2 31.51 91.46 ;
        RECT 31.25 90.44 31.51 90.7 ;
        RECT 31.25 89.68 31.51 89.94 ;
        RECT 31.25 88.92 31.51 89.18 ;
        RECT 31.25 88.16 31.51 88.42 ;
        RECT 31.25 87.4 31.51 87.66 ;
        RECT 31.25 86.64 31.51 86.9 ;
        RECT 31.25 85.88 31.51 86.14 ;
        RECT 31.25 85.12 31.51 85.38 ;
        RECT 31.25 84.36 31.51 84.62 ;
        RECT 31.25 83.6 31.51 83.86 ;
        RECT 31.25 82.84 31.51 83.1 ;
        RECT 31.25 82.08 31.51 82.34 ;
        RECT 31.25 81.32 31.51 81.58 ;
        RECT 31.25 80.56 31.51 80.82 ;
        RECT 31.25 79.8 31.51 80.06 ;
        RECT 31.25 79.04 31.51 79.3 ;
        RECT 31.25 78.28 31.51 78.54 ;
        RECT 31.25 77.52 31.51 77.78 ;
        RECT 31.25 76.76 31.51 77.02 ;
        RECT 31.25 76 31.51 76.26 ;
        RECT 31.25 75.24 31.51 75.5 ;
        RECT 31.25 74.48 31.51 74.74 ;
        RECT 31.25 73.72 31.51 73.98 ;
        RECT 31.25 72.96 31.51 73.22 ;
        RECT 31.25 72.2 31.51 72.46 ;
        RECT 31.25 71.44 31.51 71.7 ;
        RECT 31.25 70.68 31.51 70.94 ;
        RECT 31.25 69.92 31.51 70.18 ;
        RECT 31.25 69.16 31.51 69.42 ;
        RECT 32.01 91.2 32.27 91.46 ;
        RECT 32.01 90.44 32.27 90.7 ;
        RECT 32.01 89.68 32.27 89.94 ;
        RECT 32.01 88.92 32.27 89.18 ;
        RECT 32.01 88.16 32.27 88.42 ;
        RECT 32.01 87.4 32.27 87.66 ;
        RECT 32.01 86.64 32.27 86.9 ;
        RECT 32.01 85.88 32.27 86.14 ;
        RECT 32.01 85.12 32.27 85.38 ;
        RECT 32.01 84.36 32.27 84.62 ;
        RECT 32.01 83.6 32.27 83.86 ;
        RECT 32.01 82.84 32.27 83.1 ;
        RECT 32.01 82.08 32.27 82.34 ;
        RECT 32.01 81.32 32.27 81.58 ;
        RECT 32.01 80.56 32.27 80.82 ;
        RECT 32.01 79.8 32.27 80.06 ;
        RECT 32.01 79.04 32.27 79.3 ;
        RECT 32.01 78.28 32.27 78.54 ;
        RECT 32.01 77.52 32.27 77.78 ;
        RECT 32.01 76.76 32.27 77.02 ;
        RECT 32.01 76 32.27 76.26 ;
        RECT 32.01 75.24 32.27 75.5 ;
        RECT 32.01 74.48 32.27 74.74 ;
        RECT 32.01 73.72 32.27 73.98 ;
        RECT 32.01 72.96 32.27 73.22 ;
        RECT 32.01 72.2 32.27 72.46 ;
        RECT 32.01 71.44 32.27 71.7 ;
        RECT 32.01 70.68 32.27 70.94 ;
        RECT 32.01 69.92 32.27 70.18 ;
        RECT 32.01 69.16 32.27 69.42 ;
        RECT 32.77 91.2 33.03 91.46 ;
        RECT 32.77 90.44 33.03 90.7 ;
        RECT 32.77 89.68 33.03 89.94 ;
        RECT 32.77 88.92 33.03 89.18 ;
        RECT 32.77 88.16 33.03 88.42 ;
        RECT 32.77 87.4 33.03 87.66 ;
        RECT 32.77 86.64 33.03 86.9 ;
        RECT 32.77 85.88 33.03 86.14 ;
        RECT 32.77 85.12 33.03 85.38 ;
        RECT 32.77 84.36 33.03 84.62 ;
        RECT 32.77 83.6 33.03 83.86 ;
        RECT 32.77 82.84 33.03 83.1 ;
        RECT 32.77 82.08 33.03 82.34 ;
        RECT 32.77 81.32 33.03 81.58 ;
        RECT 32.77 80.56 33.03 80.82 ;
        RECT 32.77 79.8 33.03 80.06 ;
        RECT 32.77 79.04 33.03 79.3 ;
        RECT 32.77 78.28 33.03 78.54 ;
        RECT 32.77 77.52 33.03 77.78 ;
        RECT 32.77 76.76 33.03 77.02 ;
        RECT 32.77 76 33.03 76.26 ;
        RECT 32.77 75.24 33.03 75.5 ;
        RECT 32.77 74.48 33.03 74.74 ;
        RECT 32.77 73.72 33.03 73.98 ;
        RECT 32.77 72.96 33.03 73.22 ;
        RECT 32.77 72.2 33.03 72.46 ;
        RECT 32.77 71.44 33.03 71.7 ;
        RECT 32.77 70.68 33.03 70.94 ;
        RECT 32.77 69.92 33.03 70.18 ;
        RECT 32.77 69.16 33.03 69.42 ;
        RECT 33.53 91.2 33.79 91.46 ;
        RECT 33.53 90.44 33.79 90.7 ;
        RECT 33.53 89.68 33.79 89.94 ;
        RECT 33.53 88.92 33.79 89.18 ;
        RECT 33.53 88.16 33.79 88.42 ;
        RECT 33.53 87.4 33.79 87.66 ;
        RECT 33.53 86.64 33.79 86.9 ;
        RECT 33.53 85.88 33.79 86.14 ;
        RECT 33.53 85.12 33.79 85.38 ;
        RECT 33.53 84.36 33.79 84.62 ;
        RECT 33.53 83.6 33.79 83.86 ;
        RECT 33.53 82.84 33.79 83.1 ;
        RECT 33.53 82.08 33.79 82.34 ;
        RECT 33.53 81.32 33.79 81.58 ;
        RECT 33.53 80.56 33.79 80.82 ;
        RECT 33.53 79.8 33.79 80.06 ;
        RECT 33.53 79.04 33.79 79.3 ;
        RECT 33.53 78.28 33.79 78.54 ;
        RECT 33.53 77.52 33.79 77.78 ;
        RECT 33.53 76.76 33.79 77.02 ;
        RECT 33.53 76 33.79 76.26 ;
        RECT 33.53 75.24 33.79 75.5 ;
        RECT 33.53 74.48 33.79 74.74 ;
        RECT 33.53 73.72 33.79 73.98 ;
        RECT 33.53 72.96 33.79 73.22 ;
        RECT 33.53 72.2 33.79 72.46 ;
        RECT 33.53 71.44 33.79 71.7 ;
        RECT 33.53 70.68 33.79 70.94 ;
        RECT 33.53 69.92 33.79 70.18 ;
        RECT 33.53 69.16 33.79 69.42 ;
        RECT 34.29 91.2 34.55 91.46 ;
        RECT 34.29 90.44 34.55 90.7 ;
        RECT 34.29 89.68 34.55 89.94 ;
        RECT 34.29 88.92 34.55 89.18 ;
        RECT 34.29 88.16 34.55 88.42 ;
        RECT 34.29 87.4 34.55 87.66 ;
        RECT 34.29 86.64 34.55 86.9 ;
        RECT 34.29 85.88 34.55 86.14 ;
        RECT 34.29 85.12 34.55 85.38 ;
        RECT 34.29 84.36 34.55 84.62 ;
        RECT 34.29 83.6 34.55 83.86 ;
        RECT 34.29 82.84 34.55 83.1 ;
        RECT 34.29 82.08 34.55 82.34 ;
        RECT 34.29 81.32 34.55 81.58 ;
        RECT 34.29 80.56 34.55 80.82 ;
        RECT 34.29 79.8 34.55 80.06 ;
        RECT 34.29 79.04 34.55 79.3 ;
        RECT 34.29 78.28 34.55 78.54 ;
        RECT 34.29 77.52 34.55 77.78 ;
        RECT 34.29 76.76 34.55 77.02 ;
        RECT 34.29 76 34.55 76.26 ;
        RECT 34.29 75.24 34.55 75.5 ;
        RECT 34.29 74.48 34.55 74.74 ;
        RECT 34.29 73.72 34.55 73.98 ;
        RECT 34.29 72.96 34.55 73.22 ;
        RECT 34.29 72.2 34.55 72.46 ;
        RECT 34.29 71.44 34.55 71.7 ;
        RECT 34.29 70.68 34.55 70.94 ;
        RECT 34.29 69.92 34.55 70.18 ;
        RECT 34.29 69.16 34.55 69.42 ;
        RECT 35.05 91.2 35.31 91.46 ;
        RECT 35.05 90.44 35.31 90.7 ;
        RECT 35.05 89.68 35.31 89.94 ;
        RECT 35.05 88.92 35.31 89.18 ;
        RECT 35.05 88.16 35.31 88.42 ;
        RECT 35.05 87.4 35.31 87.66 ;
        RECT 35.05 86.64 35.31 86.9 ;
        RECT 35.05 85.88 35.31 86.14 ;
        RECT 35.05 85.12 35.31 85.38 ;
        RECT 35.05 84.36 35.31 84.62 ;
        RECT 35.05 83.6 35.31 83.86 ;
        RECT 35.05 82.84 35.31 83.1 ;
        RECT 35.05 82.08 35.31 82.34 ;
        RECT 35.05 81.32 35.31 81.58 ;
        RECT 35.05 80.56 35.31 80.82 ;
        RECT 35.05 79.8 35.31 80.06 ;
        RECT 35.05 79.04 35.31 79.3 ;
        RECT 35.05 78.28 35.31 78.54 ;
        RECT 35.05 77.52 35.31 77.78 ;
        RECT 35.05 76.76 35.31 77.02 ;
        RECT 35.05 76 35.31 76.26 ;
        RECT 35.05 75.24 35.31 75.5 ;
        RECT 35.05 74.48 35.31 74.74 ;
        RECT 35.05 73.72 35.31 73.98 ;
        RECT 35.05 72.96 35.31 73.22 ;
        RECT 35.05 72.2 35.31 72.46 ;
        RECT 35.05 71.44 35.31 71.7 ;
        RECT 35.05 70.68 35.31 70.94 ;
        RECT 35.05 69.92 35.31 70.18 ;
        RECT 35.05 69.16 35.31 69.42 ;
        RECT 35.81 91.2 36.07 91.46 ;
        RECT 35.81 90.44 36.07 90.7 ;
        RECT 35.81 89.68 36.07 89.94 ;
        RECT 35.81 88.92 36.07 89.18 ;
        RECT 35.81 88.16 36.07 88.42 ;
        RECT 35.81 87.4 36.07 87.66 ;
        RECT 35.81 86.64 36.07 86.9 ;
        RECT 35.81 85.88 36.07 86.14 ;
        RECT 35.81 85.12 36.07 85.38 ;
        RECT 35.81 84.36 36.07 84.62 ;
        RECT 35.81 83.6 36.07 83.86 ;
        RECT 35.81 82.84 36.07 83.1 ;
        RECT 35.81 82.08 36.07 82.34 ;
        RECT 35.81 81.32 36.07 81.58 ;
        RECT 35.81 80.56 36.07 80.82 ;
        RECT 35.81 79.8 36.07 80.06 ;
        RECT 35.81 79.04 36.07 79.3 ;
        RECT 35.81 78.28 36.07 78.54 ;
        RECT 35.81 77.52 36.07 77.78 ;
        RECT 35.81 76.76 36.07 77.02 ;
        RECT 35.81 76 36.07 76.26 ;
        RECT 35.81 75.24 36.07 75.5 ;
        RECT 35.81 74.48 36.07 74.74 ;
        RECT 35.81 73.72 36.07 73.98 ;
        RECT 35.81 72.96 36.07 73.22 ;
        RECT 35.81 72.2 36.07 72.46 ;
        RECT 35.81 71.44 36.07 71.7 ;
        RECT 35.81 70.68 36.07 70.94 ;
        RECT 35.81 69.92 36.07 70.18 ;
        RECT 35.81 69.16 36.07 69.42 ;
        RECT 36.57 91.2 36.83 91.46 ;
        RECT 36.57 90.44 36.83 90.7 ;
        RECT 36.57 89.68 36.83 89.94 ;
        RECT 36.57 88.92 36.83 89.18 ;
        RECT 36.57 88.16 36.83 88.42 ;
        RECT 36.57 87.4 36.83 87.66 ;
        RECT 36.57 86.64 36.83 86.9 ;
        RECT 36.57 85.88 36.83 86.14 ;
        RECT 36.57 85.12 36.83 85.38 ;
        RECT 36.57 84.36 36.83 84.62 ;
        RECT 36.57 83.6 36.83 83.86 ;
        RECT 36.57 82.84 36.83 83.1 ;
        RECT 36.57 82.08 36.83 82.34 ;
        RECT 36.57 81.32 36.83 81.58 ;
        RECT 36.57 80.56 36.83 80.82 ;
        RECT 36.57 79.8 36.83 80.06 ;
        RECT 36.57 79.04 36.83 79.3 ;
        RECT 36.57 78.28 36.83 78.54 ;
        RECT 36.57 77.52 36.83 77.78 ;
        RECT 36.57 76.76 36.83 77.02 ;
        RECT 36.57 76 36.83 76.26 ;
        RECT 36.57 75.24 36.83 75.5 ;
        RECT 36.57 74.48 36.83 74.74 ;
        RECT 36.57 73.72 36.83 73.98 ;
        RECT 36.57 72.96 36.83 73.22 ;
        RECT 36.57 72.2 36.83 72.46 ;
        RECT 36.57 71.44 36.83 71.7 ;
        RECT 36.57 70.68 36.83 70.94 ;
        RECT 36.57 69.92 36.83 70.18 ;
        RECT 36.57 69.16 36.83 69.42 ;
        RECT 37.33 91.2 37.59 91.46 ;
        RECT 37.33 90.44 37.59 90.7 ;
        RECT 37.33 89.68 37.59 89.94 ;
        RECT 37.33 88.92 37.59 89.18 ;
        RECT 37.33 88.16 37.59 88.42 ;
        RECT 37.33 87.4 37.59 87.66 ;
        RECT 37.33 86.64 37.59 86.9 ;
        RECT 37.33 85.88 37.59 86.14 ;
        RECT 37.33 85.12 37.59 85.38 ;
        RECT 37.33 84.36 37.59 84.62 ;
        RECT 37.33 83.6 37.59 83.86 ;
        RECT 37.33 82.84 37.59 83.1 ;
        RECT 37.33 82.08 37.59 82.34 ;
        RECT 37.33 81.32 37.59 81.58 ;
        RECT 37.33 80.56 37.59 80.82 ;
        RECT 37.33 79.8 37.59 80.06 ;
        RECT 37.33 79.04 37.59 79.3 ;
        RECT 37.33 78.28 37.59 78.54 ;
        RECT 37.33 77.52 37.59 77.78 ;
        RECT 37.33 76.76 37.59 77.02 ;
        RECT 37.33 76 37.59 76.26 ;
        RECT 37.33 75.24 37.59 75.5 ;
        RECT 37.33 74.48 37.59 74.74 ;
        RECT 37.33 73.72 37.59 73.98 ;
        RECT 37.33 72.96 37.59 73.22 ;
        RECT 37.33 72.2 37.59 72.46 ;
        RECT 37.33 71.44 37.59 71.7 ;
        RECT 37.33 70.68 37.59 70.94 ;
        RECT 37.33 69.92 37.59 70.18 ;
        RECT 37.33 69.16 37.59 69.42 ;
        RECT 38.09 91.2 38.35 91.46 ;
        RECT 38.09 90.44 38.35 90.7 ;
        RECT 38.09 89.68 38.35 89.94 ;
        RECT 38.09 88.92 38.35 89.18 ;
        RECT 38.09 88.16 38.35 88.42 ;
        RECT 38.09 87.4 38.35 87.66 ;
        RECT 38.09 86.64 38.35 86.9 ;
        RECT 38.09 85.88 38.35 86.14 ;
        RECT 38.09 85.12 38.35 85.38 ;
        RECT 38.09 84.36 38.35 84.62 ;
        RECT 38.09 83.6 38.35 83.86 ;
        RECT 38.09 82.84 38.35 83.1 ;
        RECT 38.09 82.08 38.35 82.34 ;
        RECT 38.09 81.32 38.35 81.58 ;
        RECT 38.09 80.56 38.35 80.82 ;
        RECT 38.09 79.8 38.35 80.06 ;
        RECT 38.09 79.04 38.35 79.3 ;
        RECT 38.09 78.28 38.35 78.54 ;
        RECT 38.09 77.52 38.35 77.78 ;
        RECT 38.09 76.76 38.35 77.02 ;
        RECT 38.09 76 38.35 76.26 ;
        RECT 38.09 75.24 38.35 75.5 ;
        RECT 38.09 74.48 38.35 74.74 ;
        RECT 38.09 73.72 38.35 73.98 ;
        RECT 38.09 72.96 38.35 73.22 ;
        RECT 38.09 72.2 38.35 72.46 ;
        RECT 38.09 71.44 38.35 71.7 ;
        RECT 38.09 70.68 38.35 70.94 ;
        RECT 38.09 69.92 38.35 70.18 ;
        RECT 38.09 69.16 38.35 69.42 ;
        RECT 38.85 91.2 39.11 91.46 ;
        RECT 38.85 90.44 39.11 90.7 ;
        RECT 38.85 89.68 39.11 89.94 ;
        RECT 38.85 88.92 39.11 89.18 ;
        RECT 38.85 88.16 39.11 88.42 ;
        RECT 38.85 87.4 39.11 87.66 ;
        RECT 38.85 86.64 39.11 86.9 ;
        RECT 38.85 85.88 39.11 86.14 ;
        RECT 38.85 85.12 39.11 85.38 ;
        RECT 38.85 84.36 39.11 84.62 ;
        RECT 38.85 83.6 39.11 83.86 ;
        RECT 38.85 82.84 39.11 83.1 ;
        RECT 38.85 82.08 39.11 82.34 ;
        RECT 38.85 81.32 39.11 81.58 ;
        RECT 38.85 80.56 39.11 80.82 ;
        RECT 38.85 79.8 39.11 80.06 ;
        RECT 38.85 79.04 39.11 79.3 ;
        RECT 38.85 78.28 39.11 78.54 ;
        RECT 38.85 77.52 39.11 77.78 ;
        RECT 38.85 76.76 39.11 77.02 ;
        RECT 38.85 76 39.11 76.26 ;
        RECT 38.85 75.24 39.11 75.5 ;
        RECT 38.85 74.48 39.11 74.74 ;
        RECT 38.85 73.72 39.11 73.98 ;
        RECT 38.85 72.96 39.11 73.22 ;
        RECT 38.85 72.2 39.11 72.46 ;
        RECT 38.85 71.44 39.11 71.7 ;
        RECT 38.85 70.68 39.11 70.94 ;
        RECT 38.85 69.92 39.11 70.18 ;
        RECT 38.85 69.16 39.11 69.42 ;
        RECT 39.61 91.2 39.87 91.46 ;
        RECT 39.61 90.44 39.87 90.7 ;
        RECT 39.61 89.68 39.87 89.94 ;
        RECT 39.61 88.92 39.87 89.18 ;
        RECT 39.61 88.16 39.87 88.42 ;
        RECT 39.61 87.4 39.87 87.66 ;
        RECT 39.61 86.64 39.87 86.9 ;
        RECT 39.61 85.88 39.87 86.14 ;
        RECT 39.61 85.12 39.87 85.38 ;
        RECT 39.61 84.36 39.87 84.62 ;
        RECT 39.61 83.6 39.87 83.86 ;
        RECT 39.61 82.84 39.87 83.1 ;
        RECT 39.61 82.08 39.87 82.34 ;
        RECT 39.61 81.32 39.87 81.58 ;
        RECT 39.61 80.56 39.87 80.82 ;
        RECT 39.61 79.8 39.87 80.06 ;
        RECT 39.61 79.04 39.87 79.3 ;
        RECT 39.61 78.28 39.87 78.54 ;
        RECT 39.61 77.52 39.87 77.78 ;
        RECT 39.61 76.76 39.87 77.02 ;
        RECT 39.61 76 39.87 76.26 ;
        RECT 39.61 75.24 39.87 75.5 ;
        RECT 39.61 74.48 39.87 74.74 ;
        RECT 39.61 73.72 39.87 73.98 ;
        RECT 39.61 72.96 39.87 73.22 ;
        RECT 39.61 72.2 39.87 72.46 ;
        RECT 39.61 71.44 39.87 71.7 ;
        RECT 39.61 70.68 39.87 70.94 ;
        RECT 39.61 69.92 39.87 70.18 ;
        RECT 39.61 69.16 39.87 69.42 ;
        RECT 40.37 91.2 40.63 91.46 ;
        RECT 40.37 90.44 40.63 90.7 ;
        RECT 40.37 89.68 40.63 89.94 ;
        RECT 40.37 88.92 40.63 89.18 ;
        RECT 40.37 88.16 40.63 88.42 ;
        RECT 40.37 87.4 40.63 87.66 ;
        RECT 40.37 86.64 40.63 86.9 ;
        RECT 40.37 85.88 40.63 86.14 ;
        RECT 40.37 85.12 40.63 85.38 ;
        RECT 40.37 84.36 40.63 84.62 ;
        RECT 40.37 83.6 40.63 83.86 ;
        RECT 40.37 82.84 40.63 83.1 ;
        RECT 40.37 82.08 40.63 82.34 ;
        RECT 40.37 81.32 40.63 81.58 ;
        RECT 40.37 80.56 40.63 80.82 ;
        RECT 40.37 79.8 40.63 80.06 ;
        RECT 40.37 79.04 40.63 79.3 ;
        RECT 40.37 78.28 40.63 78.54 ;
        RECT 40.37 77.52 40.63 77.78 ;
        RECT 40.37 76.76 40.63 77.02 ;
        RECT 40.37 76 40.63 76.26 ;
        RECT 40.37 75.24 40.63 75.5 ;
        RECT 40.37 74.48 40.63 74.74 ;
        RECT 40.37 73.72 40.63 73.98 ;
        RECT 40.37 72.96 40.63 73.22 ;
        RECT 40.37 72.2 40.63 72.46 ;
        RECT 40.37 71.44 40.63 71.7 ;
        RECT 40.37 70.68 40.63 70.94 ;
        RECT 40.37 69.92 40.63 70.18 ;
        RECT 40.37 69.16 40.63 69.42 ;
        RECT 41.13 91.2 41.39 91.46 ;
        RECT 41.13 90.44 41.39 90.7 ;
        RECT 41.13 89.68 41.39 89.94 ;
        RECT 41.13 88.92 41.39 89.18 ;
        RECT 41.13 88.16 41.39 88.42 ;
        RECT 41.13 87.4 41.39 87.66 ;
        RECT 41.13 86.64 41.39 86.9 ;
        RECT 41.13 85.88 41.39 86.14 ;
        RECT 41.13 85.12 41.39 85.38 ;
        RECT 41.13 84.36 41.39 84.62 ;
        RECT 41.13 83.6 41.39 83.86 ;
        RECT 41.13 82.84 41.39 83.1 ;
        RECT 41.13 82.08 41.39 82.34 ;
        RECT 41.13 81.32 41.39 81.58 ;
        RECT 41.13 80.56 41.39 80.82 ;
        RECT 41.13 79.8 41.39 80.06 ;
        RECT 41.13 79.04 41.39 79.3 ;
        RECT 41.13 78.28 41.39 78.54 ;
        RECT 41.13 77.52 41.39 77.78 ;
        RECT 41.13 76.76 41.39 77.02 ;
        RECT 41.13 76 41.39 76.26 ;
        RECT 41.13 75.24 41.39 75.5 ;
        RECT 41.13 74.48 41.39 74.74 ;
        RECT 41.13 73.72 41.39 73.98 ;
        RECT 41.13 72.96 41.39 73.22 ;
        RECT 41.13 72.2 41.39 72.46 ;
        RECT 41.13 71.44 41.39 71.7 ;
        RECT 41.13 70.68 41.39 70.94 ;
        RECT 41.13 69.92 41.39 70.18 ;
        RECT 41.13 69.16 41.39 69.42 ;
        RECT 41.89 91.2 42.15 91.46 ;
        RECT 41.89 90.44 42.15 90.7 ;
        RECT 41.89 89.68 42.15 89.94 ;
        RECT 41.89 88.92 42.15 89.18 ;
        RECT 41.89 88.16 42.15 88.42 ;
        RECT 41.89 87.4 42.15 87.66 ;
        RECT 41.89 86.64 42.15 86.9 ;
        RECT 41.89 85.88 42.15 86.14 ;
        RECT 41.89 85.12 42.15 85.38 ;
        RECT 41.89 84.36 42.15 84.62 ;
        RECT 41.89 83.6 42.15 83.86 ;
        RECT 41.89 82.84 42.15 83.1 ;
        RECT 41.89 82.08 42.15 82.34 ;
        RECT 41.89 81.32 42.15 81.58 ;
        RECT 41.89 80.56 42.15 80.82 ;
        RECT 41.89 79.8 42.15 80.06 ;
        RECT 41.89 79.04 42.15 79.3 ;
        RECT 41.89 78.28 42.15 78.54 ;
        RECT 41.89 77.52 42.15 77.78 ;
        RECT 41.89 76.76 42.15 77.02 ;
        RECT 41.89 76 42.15 76.26 ;
        RECT 41.89 75.24 42.15 75.5 ;
        RECT 41.89 74.48 42.15 74.74 ;
        RECT 41.89 73.72 42.15 73.98 ;
        RECT 41.89 72.96 42.15 73.22 ;
        RECT 41.89 72.2 42.15 72.46 ;
        RECT 41.89 71.44 42.15 71.7 ;
        RECT 41.89 70.68 42.15 70.94 ;
        RECT 41.89 69.92 42.15 70.18 ;
        RECT 41.89 69.16 42.15 69.42 ;
        RECT 42.65 91.2 42.91 91.46 ;
        RECT 42.65 90.44 42.91 90.7 ;
        RECT 42.65 89.68 42.91 89.94 ;
        RECT 42.65 88.92 42.91 89.18 ;
        RECT 42.65 88.16 42.91 88.42 ;
        RECT 42.65 87.4 42.91 87.66 ;
        RECT 42.65 86.64 42.91 86.9 ;
        RECT 42.65 85.88 42.91 86.14 ;
        RECT 42.65 85.12 42.91 85.38 ;
        RECT 42.65 84.36 42.91 84.62 ;
        RECT 42.65 83.6 42.91 83.86 ;
        RECT 42.65 82.84 42.91 83.1 ;
        RECT 42.65 82.08 42.91 82.34 ;
        RECT 42.65 81.32 42.91 81.58 ;
        RECT 42.65 80.56 42.91 80.82 ;
        RECT 42.65 79.8 42.91 80.06 ;
        RECT 42.65 79.04 42.91 79.3 ;
        RECT 42.65 78.28 42.91 78.54 ;
        RECT 42.65 77.52 42.91 77.78 ;
        RECT 42.65 76.76 42.91 77.02 ;
        RECT 42.65 76 42.91 76.26 ;
        RECT 42.65 75.24 42.91 75.5 ;
        RECT 42.65 74.48 42.91 74.74 ;
        RECT 42.65 73.72 42.91 73.98 ;
        RECT 42.65 72.96 42.91 73.22 ;
        RECT 42.65 72.2 42.91 72.46 ;
        RECT 42.65 71.44 42.91 71.7 ;
        RECT 42.65 70.68 42.91 70.94 ;
        RECT 42.65 69.92 42.91 70.18 ;
        RECT 42.65 69.16 42.91 69.42 ;
        RECT 43.41 91.2 43.67 91.46 ;
        RECT 43.41 90.44 43.67 90.7 ;
        RECT 43.41 89.68 43.67 89.94 ;
        RECT 43.41 88.92 43.67 89.18 ;
        RECT 43.41 88.16 43.67 88.42 ;
        RECT 43.41 87.4 43.67 87.66 ;
        RECT 43.41 86.64 43.67 86.9 ;
        RECT 43.41 85.88 43.67 86.14 ;
        RECT 43.41 85.12 43.67 85.38 ;
        RECT 43.41 84.36 43.67 84.62 ;
        RECT 43.41 83.6 43.67 83.86 ;
        RECT 43.41 82.84 43.67 83.1 ;
        RECT 43.41 82.08 43.67 82.34 ;
        RECT 43.41 81.32 43.67 81.58 ;
        RECT 43.41 80.56 43.67 80.82 ;
        RECT 43.41 79.8 43.67 80.06 ;
        RECT 43.41 79.04 43.67 79.3 ;
        RECT 43.41 78.28 43.67 78.54 ;
        RECT 43.41 77.52 43.67 77.78 ;
        RECT 43.41 76.76 43.67 77.02 ;
        RECT 43.41 76 43.67 76.26 ;
        RECT 43.41 75.24 43.67 75.5 ;
        RECT 43.41 74.48 43.67 74.74 ;
        RECT 43.41 73.72 43.67 73.98 ;
        RECT 43.41 72.96 43.67 73.22 ;
        RECT 43.41 72.2 43.67 72.46 ;
        RECT 43.41 71.44 43.67 71.7 ;
        RECT 43.41 70.68 43.67 70.94 ;
        RECT 43.41 69.92 43.67 70.18 ;
        RECT 43.41 69.16 43.67 69.42 ;
        RECT 44.17 91.2 44.43 91.46 ;
        RECT 44.17 90.44 44.43 90.7 ;
        RECT 44.17 89.68 44.43 89.94 ;
        RECT 44.17 88.92 44.43 89.18 ;
        RECT 44.17 88.16 44.43 88.42 ;
        RECT 44.17 87.4 44.43 87.66 ;
        RECT 44.17 86.64 44.43 86.9 ;
        RECT 44.17 85.88 44.43 86.14 ;
        RECT 44.17 85.12 44.43 85.38 ;
        RECT 44.17 84.36 44.43 84.62 ;
        RECT 44.17 83.6 44.43 83.86 ;
        RECT 44.17 82.84 44.43 83.1 ;
        RECT 44.17 82.08 44.43 82.34 ;
        RECT 44.17 81.32 44.43 81.58 ;
        RECT 44.17 80.56 44.43 80.82 ;
        RECT 44.17 79.8 44.43 80.06 ;
        RECT 44.17 79.04 44.43 79.3 ;
        RECT 44.17 78.28 44.43 78.54 ;
        RECT 44.17 77.52 44.43 77.78 ;
        RECT 44.17 76.76 44.43 77.02 ;
        RECT 44.17 76 44.43 76.26 ;
        RECT 44.17 75.24 44.43 75.5 ;
        RECT 44.17 74.48 44.43 74.74 ;
        RECT 44.17 73.72 44.43 73.98 ;
        RECT 44.17 72.96 44.43 73.22 ;
        RECT 44.17 72.2 44.43 72.46 ;
        RECT 44.17 71.44 44.43 71.7 ;
        RECT 44.17 70.68 44.43 70.94 ;
        RECT 44.17 69.92 44.43 70.18 ;
        RECT 44.17 69.16 44.43 69.42 ;
        RECT 44.93 91.2 45.19 91.46 ;
        RECT 44.93 90.44 45.19 90.7 ;
        RECT 44.93 89.68 45.19 89.94 ;
        RECT 44.93 88.92 45.19 89.18 ;
        RECT 44.93 88.16 45.19 88.42 ;
        RECT 44.93 87.4 45.19 87.66 ;
        RECT 44.93 86.64 45.19 86.9 ;
        RECT 44.93 85.88 45.19 86.14 ;
        RECT 44.93 85.12 45.19 85.38 ;
        RECT 44.93 84.36 45.19 84.62 ;
        RECT 44.93 83.6 45.19 83.86 ;
        RECT 44.93 82.84 45.19 83.1 ;
        RECT 44.93 82.08 45.19 82.34 ;
        RECT 44.93 81.32 45.19 81.58 ;
        RECT 44.93 80.56 45.19 80.82 ;
        RECT 44.93 79.8 45.19 80.06 ;
        RECT 44.93 79.04 45.19 79.3 ;
        RECT 44.93 78.28 45.19 78.54 ;
        RECT 44.93 77.52 45.19 77.78 ;
        RECT 44.93 76.76 45.19 77.02 ;
        RECT 44.93 76 45.19 76.26 ;
        RECT 44.93 75.24 45.19 75.5 ;
        RECT 44.93 74.48 45.19 74.74 ;
        RECT 44.93 73.72 45.19 73.98 ;
        RECT 44.93 72.96 45.19 73.22 ;
        RECT 44.93 72.2 45.19 72.46 ;
        RECT 44.93 71.44 45.19 71.7 ;
        RECT 44.93 70.68 45.19 70.94 ;
        RECT 44.93 69.92 45.19 70.18 ;
        RECT 44.93 69.16 45.19 69.42 ;
        RECT 45.69 91.2 45.95 91.46 ;
        RECT 45.69 90.44 45.95 90.7 ;
        RECT 45.69 89.68 45.95 89.94 ;
        RECT 45.69 88.92 45.95 89.18 ;
        RECT 45.69 88.16 45.95 88.42 ;
        RECT 45.69 87.4 45.95 87.66 ;
        RECT 45.69 86.64 45.95 86.9 ;
        RECT 45.69 85.88 45.95 86.14 ;
        RECT 45.69 85.12 45.95 85.38 ;
        RECT 45.69 84.36 45.95 84.62 ;
        RECT 45.69 83.6 45.95 83.86 ;
        RECT 45.69 82.84 45.95 83.1 ;
        RECT 45.69 82.08 45.95 82.34 ;
        RECT 45.69 81.32 45.95 81.58 ;
        RECT 45.69 80.56 45.95 80.82 ;
        RECT 45.69 79.8 45.95 80.06 ;
        RECT 45.69 79.04 45.95 79.3 ;
        RECT 45.69 78.28 45.95 78.54 ;
        RECT 45.69 77.52 45.95 77.78 ;
        RECT 45.69 76.76 45.95 77.02 ;
        RECT 45.69 76 45.95 76.26 ;
        RECT 45.69 75.24 45.95 75.5 ;
        RECT 45.69 74.48 45.95 74.74 ;
        RECT 45.69 73.72 45.95 73.98 ;
        RECT 45.69 72.96 45.95 73.22 ;
        RECT 45.69 72.2 45.95 72.46 ;
        RECT 45.69 71.44 45.95 71.7 ;
        RECT 45.69 70.68 45.95 70.94 ;
        RECT 45.69 69.92 45.95 70.18 ;
        RECT 45.69 69.16 45.95 69.42 ;
        RECT 46.45 91.2 46.71 91.46 ;
        RECT 46.45 90.44 46.71 90.7 ;
        RECT 46.45 89.68 46.71 89.94 ;
        RECT 46.45 88.92 46.71 89.18 ;
        RECT 46.45 88.16 46.71 88.42 ;
        RECT 46.45 87.4 46.71 87.66 ;
        RECT 46.45 86.64 46.71 86.9 ;
        RECT 46.45 85.88 46.71 86.14 ;
        RECT 46.45 85.12 46.71 85.38 ;
        RECT 46.45 84.36 46.71 84.62 ;
        RECT 46.45 83.6 46.71 83.86 ;
        RECT 46.45 82.84 46.71 83.1 ;
        RECT 46.45 82.08 46.71 82.34 ;
        RECT 46.45 81.32 46.71 81.58 ;
        RECT 46.45 80.56 46.71 80.82 ;
        RECT 46.45 79.8 46.71 80.06 ;
        RECT 46.45 79.04 46.71 79.3 ;
        RECT 46.45 78.28 46.71 78.54 ;
        RECT 46.45 77.52 46.71 77.78 ;
        RECT 46.45 76.76 46.71 77.02 ;
        RECT 46.45 76 46.71 76.26 ;
        RECT 46.45 75.24 46.71 75.5 ;
        RECT 46.45 74.48 46.71 74.74 ;
        RECT 46.45 73.72 46.71 73.98 ;
        RECT 46.45 72.96 46.71 73.22 ;
        RECT 46.45 72.2 46.71 72.46 ;
        RECT 46.45 71.44 46.71 71.7 ;
        RECT 46.45 70.68 46.71 70.94 ;
        RECT 46.45 69.92 46.71 70.18 ;
        RECT 46.45 69.16 46.71 69.42 ;
        RECT 47.21 91.2 47.47 91.46 ;
        RECT 47.21 90.44 47.47 90.7 ;
        RECT 47.21 89.68 47.47 89.94 ;
        RECT 47.21 88.92 47.47 89.18 ;
        RECT 47.21 88.16 47.47 88.42 ;
        RECT 47.21 87.4 47.47 87.66 ;
        RECT 47.21 86.64 47.47 86.9 ;
        RECT 47.21 85.88 47.47 86.14 ;
        RECT 47.21 85.12 47.47 85.38 ;
        RECT 47.21 84.36 47.47 84.62 ;
        RECT 47.21 83.6 47.47 83.86 ;
        RECT 47.21 82.84 47.47 83.1 ;
        RECT 47.21 82.08 47.47 82.34 ;
        RECT 47.21 81.32 47.47 81.58 ;
        RECT 47.21 80.56 47.47 80.82 ;
        RECT 47.21 79.8 47.47 80.06 ;
        RECT 47.21 79.04 47.47 79.3 ;
        RECT 47.21 78.28 47.47 78.54 ;
        RECT 47.21 77.52 47.47 77.78 ;
        RECT 47.21 76.76 47.47 77.02 ;
        RECT 47.21 76 47.47 76.26 ;
        RECT 47.21 75.24 47.47 75.5 ;
        RECT 47.21 74.48 47.47 74.74 ;
        RECT 47.21 73.72 47.47 73.98 ;
        RECT 47.21 72.96 47.47 73.22 ;
        RECT 47.21 72.2 47.47 72.46 ;
        RECT 47.21 71.44 47.47 71.7 ;
        RECT 47.21 70.68 47.47 70.94 ;
        RECT 47.21 69.92 47.47 70.18 ;
        RECT 47.21 69.16 47.47 69.42 ;
        RECT 47.97 91.2 48.23 91.46 ;
        RECT 47.97 90.44 48.23 90.7 ;
        RECT 47.97 89.68 48.23 89.94 ;
        RECT 47.97 88.92 48.23 89.18 ;
        RECT 47.97 88.16 48.23 88.42 ;
        RECT 47.97 87.4 48.23 87.66 ;
        RECT 47.97 86.64 48.23 86.9 ;
        RECT 47.97 85.88 48.23 86.14 ;
        RECT 47.97 85.12 48.23 85.38 ;
        RECT 47.97 84.36 48.23 84.62 ;
        RECT 47.97 83.6 48.23 83.86 ;
        RECT 47.97 82.84 48.23 83.1 ;
        RECT 47.97 82.08 48.23 82.34 ;
        RECT 47.97 81.32 48.23 81.58 ;
        RECT 47.97 80.56 48.23 80.82 ;
        RECT 47.97 79.8 48.23 80.06 ;
        RECT 47.97 79.04 48.23 79.3 ;
        RECT 47.97 78.28 48.23 78.54 ;
        RECT 47.97 77.52 48.23 77.78 ;
        RECT 47.97 76.76 48.23 77.02 ;
        RECT 47.97 76 48.23 76.26 ;
        RECT 47.97 75.24 48.23 75.5 ;
        RECT 47.97 74.48 48.23 74.74 ;
        RECT 47.97 73.72 48.23 73.98 ;
        RECT 47.97 72.96 48.23 73.22 ;
        RECT 47.97 72.2 48.23 72.46 ;
        RECT 47.97 71.44 48.23 71.7 ;
        RECT 47.97 70.68 48.23 70.94 ;
        RECT 47.97 69.92 48.23 70.18 ;
        RECT 47.97 69.16 48.23 69.42 ;
        RECT 48.73 91.2 48.99 91.46 ;
        RECT 48.73 90.44 48.99 90.7 ;
        RECT 48.73 89.68 48.99 89.94 ;
        RECT 48.73 88.92 48.99 89.18 ;
        RECT 48.73 88.16 48.99 88.42 ;
        RECT 48.73 87.4 48.99 87.66 ;
        RECT 48.73 86.64 48.99 86.9 ;
        RECT 48.73 85.88 48.99 86.14 ;
        RECT 48.73 85.12 48.99 85.38 ;
        RECT 48.73 84.36 48.99 84.62 ;
        RECT 48.73 83.6 48.99 83.86 ;
        RECT 48.73 82.84 48.99 83.1 ;
        RECT 48.73 82.08 48.99 82.34 ;
        RECT 48.73 81.32 48.99 81.58 ;
        RECT 48.73 80.56 48.99 80.82 ;
        RECT 48.73 79.8 48.99 80.06 ;
        RECT 48.73 79.04 48.99 79.3 ;
        RECT 48.73 78.28 48.99 78.54 ;
        RECT 48.73 77.52 48.99 77.78 ;
        RECT 48.73 76.76 48.99 77.02 ;
        RECT 48.73 76 48.99 76.26 ;
        RECT 48.73 75.24 48.99 75.5 ;
        RECT 48.73 74.48 48.99 74.74 ;
        RECT 48.73 73.72 48.99 73.98 ;
        RECT 48.73 72.96 48.99 73.22 ;
        RECT 48.73 72.2 48.99 72.46 ;
        RECT 48.73 71.44 48.99 71.7 ;
        RECT 48.73 70.68 48.99 70.94 ;
        RECT 48.73 69.92 48.99 70.18 ;
        RECT 48.73 69.16 48.99 69.42 ;
        RECT 49.49 91.2 49.75 91.46 ;
        RECT 49.49 90.44 49.75 90.7 ;
        RECT 49.49 89.68 49.75 89.94 ;
        RECT 49.49 88.92 49.75 89.18 ;
        RECT 49.49 88.16 49.75 88.42 ;
        RECT 49.49 87.4 49.75 87.66 ;
        RECT 49.49 86.64 49.75 86.9 ;
        RECT 49.49 85.88 49.75 86.14 ;
        RECT 49.49 85.12 49.75 85.38 ;
        RECT 49.49 84.36 49.75 84.62 ;
        RECT 49.49 83.6 49.75 83.86 ;
        RECT 49.49 82.84 49.75 83.1 ;
        RECT 49.49 82.08 49.75 82.34 ;
        RECT 49.49 81.32 49.75 81.58 ;
        RECT 49.49 80.56 49.75 80.82 ;
        RECT 49.49 79.8 49.75 80.06 ;
        RECT 49.49 79.04 49.75 79.3 ;
        RECT 49.49 78.28 49.75 78.54 ;
        RECT 49.49 77.52 49.75 77.78 ;
        RECT 49.49 76.76 49.75 77.02 ;
        RECT 49.49 76 49.75 76.26 ;
        RECT 49.49 75.24 49.75 75.5 ;
        RECT 49.49 74.48 49.75 74.74 ;
        RECT 49.49 73.72 49.75 73.98 ;
        RECT 49.49 72.96 49.75 73.22 ;
        RECT 49.49 72.2 49.75 72.46 ;
        RECT 49.49 71.44 49.75 71.7 ;
        RECT 49.49 70.68 49.75 70.94 ;
        RECT 49.49 69.92 49.75 70.18 ;
        RECT 49.49 69.16 49.75 69.42 ;
        RECT 50.25 91.2 50.51 91.46 ;
        RECT 50.25 90.44 50.51 90.7 ;
        RECT 50.25 89.68 50.51 89.94 ;
        RECT 50.25 88.92 50.51 89.18 ;
        RECT 50.25 88.16 50.51 88.42 ;
        RECT 50.25 87.4 50.51 87.66 ;
        RECT 50.25 86.64 50.51 86.9 ;
        RECT 50.25 85.88 50.51 86.14 ;
        RECT 50.25 85.12 50.51 85.38 ;
        RECT 50.25 84.36 50.51 84.62 ;
        RECT 50.25 83.6 50.51 83.86 ;
        RECT 50.25 82.84 50.51 83.1 ;
        RECT 50.25 82.08 50.51 82.34 ;
        RECT 50.25 81.32 50.51 81.58 ;
        RECT 50.25 80.56 50.51 80.82 ;
        RECT 50.25 79.8 50.51 80.06 ;
        RECT 50.25 79.04 50.51 79.3 ;
        RECT 50.25 78.28 50.51 78.54 ;
        RECT 50.25 77.52 50.51 77.78 ;
        RECT 50.25 76.76 50.51 77.02 ;
        RECT 50.25 76 50.51 76.26 ;
        RECT 50.25 75.24 50.51 75.5 ;
        RECT 50.25 74.48 50.51 74.74 ;
        RECT 50.25 73.72 50.51 73.98 ;
        RECT 50.25 72.96 50.51 73.22 ;
        RECT 50.25 72.2 50.51 72.46 ;
        RECT 50.25 71.44 50.51 71.7 ;
        RECT 50.25 70.68 50.51 70.94 ;
        RECT 50.25 69.92 50.51 70.18 ;
        RECT 50.25 69.16 50.51 69.42 ;
        RECT 51.01 91.2 51.27 91.46 ;
        RECT 51.01 90.44 51.27 90.7 ;
        RECT 51.01 89.68 51.27 89.94 ;
        RECT 51.01 88.92 51.27 89.18 ;
        RECT 51.01 88.16 51.27 88.42 ;
        RECT 51.01 87.4 51.27 87.66 ;
        RECT 51.01 86.64 51.27 86.9 ;
        RECT 51.01 85.88 51.27 86.14 ;
        RECT 51.01 85.12 51.27 85.38 ;
        RECT 51.01 84.36 51.27 84.62 ;
        RECT 51.01 83.6 51.27 83.86 ;
        RECT 51.01 82.84 51.27 83.1 ;
        RECT 51.01 82.08 51.27 82.34 ;
        RECT 51.01 81.32 51.27 81.58 ;
        RECT 51.01 80.56 51.27 80.82 ;
        RECT 51.01 79.8 51.27 80.06 ;
        RECT 51.01 79.04 51.27 79.3 ;
        RECT 51.01 78.28 51.27 78.54 ;
        RECT 51.01 77.52 51.27 77.78 ;
        RECT 51.01 76.76 51.27 77.02 ;
        RECT 51.01 76 51.27 76.26 ;
        RECT 51.01 75.24 51.27 75.5 ;
        RECT 51.01 74.48 51.27 74.74 ;
        RECT 51.01 73.72 51.27 73.98 ;
        RECT 51.01 72.96 51.27 73.22 ;
        RECT 51.01 72.2 51.27 72.46 ;
        RECT 51.01 71.44 51.27 71.7 ;
        RECT 51.01 70.68 51.27 70.94 ;
        RECT 51.01 69.92 51.27 70.18 ;
        RECT 51.01 69.16 51.27 69.42 ;
        RECT 51.77 91.2 52.03 91.46 ;
        RECT 51.77 90.44 52.03 90.7 ;
        RECT 51.77 89.68 52.03 89.94 ;
        RECT 51.77 88.92 52.03 89.18 ;
        RECT 51.77 88.16 52.03 88.42 ;
        RECT 51.77 87.4 52.03 87.66 ;
        RECT 51.77 86.64 52.03 86.9 ;
        RECT 51.77 85.88 52.03 86.14 ;
        RECT 51.77 85.12 52.03 85.38 ;
        RECT 51.77 84.36 52.03 84.62 ;
        RECT 51.77 83.6 52.03 83.86 ;
        RECT 51.77 82.84 52.03 83.1 ;
        RECT 51.77 82.08 52.03 82.34 ;
        RECT 51.77 81.32 52.03 81.58 ;
        RECT 51.77 80.56 52.03 80.82 ;
        RECT 51.77 79.8 52.03 80.06 ;
        RECT 51.77 79.04 52.03 79.3 ;
        RECT 51.77 78.28 52.03 78.54 ;
        RECT 51.77 77.52 52.03 77.78 ;
        RECT 51.77 76.76 52.03 77.02 ;
        RECT 51.77 76 52.03 76.26 ;
        RECT 51.77 75.24 52.03 75.5 ;
        RECT 51.77 74.48 52.03 74.74 ;
        RECT 51.77 73.72 52.03 73.98 ;
        RECT 51.77 72.96 52.03 73.22 ;
        RECT 51.77 72.2 52.03 72.46 ;
        RECT 51.77 71.44 52.03 71.7 ;
        RECT 51.77 70.68 52.03 70.94 ;
        RECT 51.77 69.92 52.03 70.18 ;
        RECT 51.77 69.16 52.03 69.42 ;
        RECT 52.53 91.2 52.79 91.46 ;
        RECT 52.53 90.44 52.79 90.7 ;
        RECT 52.53 89.68 52.79 89.94 ;
        RECT 52.53 88.92 52.79 89.18 ;
        RECT 52.53 88.16 52.79 88.42 ;
        RECT 52.53 87.4 52.79 87.66 ;
        RECT 52.53 86.64 52.79 86.9 ;
        RECT 52.53 85.88 52.79 86.14 ;
        RECT 52.53 85.12 52.79 85.38 ;
        RECT 52.53 84.36 52.79 84.62 ;
        RECT 52.53 83.6 52.79 83.86 ;
        RECT 52.53 82.84 52.79 83.1 ;
        RECT 52.53 82.08 52.79 82.34 ;
        RECT 52.53 81.32 52.79 81.58 ;
        RECT 52.53 80.56 52.79 80.82 ;
        RECT 52.53 79.8 52.79 80.06 ;
        RECT 52.53 79.04 52.79 79.3 ;
        RECT 52.53 78.28 52.79 78.54 ;
        RECT 52.53 77.52 52.79 77.78 ;
        RECT 52.53 76.76 52.79 77.02 ;
        RECT 52.53 76 52.79 76.26 ;
        RECT 52.53 75.24 52.79 75.5 ;
        RECT 52.53 74.48 52.79 74.74 ;
        RECT 52.53 73.72 52.79 73.98 ;
        RECT 52.53 72.96 52.79 73.22 ;
        RECT 52.53 72.2 52.79 72.46 ;
        RECT 52.53 71.44 52.79 71.7 ;
        RECT 52.53 70.68 52.79 70.94 ;
        RECT 52.53 69.92 52.79 70.18 ;
        RECT 52.53 69.16 52.79 69.42 ;
        RECT 53.29 91.2 53.55 91.46 ;
        RECT 53.29 90.44 53.55 90.7 ;
        RECT 53.29 89.68 53.55 89.94 ;
        RECT 53.29 88.92 53.55 89.18 ;
        RECT 53.29 88.16 53.55 88.42 ;
        RECT 53.29 87.4 53.55 87.66 ;
        RECT 53.29 86.64 53.55 86.9 ;
        RECT 53.29 85.88 53.55 86.14 ;
        RECT 53.29 85.12 53.55 85.38 ;
        RECT 53.29 84.36 53.55 84.62 ;
        RECT 53.29 83.6 53.55 83.86 ;
        RECT 53.29 82.84 53.55 83.1 ;
        RECT 53.29 82.08 53.55 82.34 ;
        RECT 53.29 81.32 53.55 81.58 ;
        RECT 53.29 80.56 53.55 80.82 ;
        RECT 53.29 79.8 53.55 80.06 ;
        RECT 53.29 79.04 53.55 79.3 ;
        RECT 53.29 78.28 53.55 78.54 ;
        RECT 53.29 77.52 53.55 77.78 ;
        RECT 53.29 76.76 53.55 77.02 ;
        RECT 53.29 76 53.55 76.26 ;
        RECT 53.29 75.24 53.55 75.5 ;
        RECT 53.29 74.48 53.55 74.74 ;
        RECT 53.29 73.72 53.55 73.98 ;
        RECT 53.29 72.96 53.55 73.22 ;
        RECT 53.29 72.2 53.55 72.46 ;
        RECT 53.29 71.44 53.55 71.7 ;
        RECT 53.29 70.68 53.55 70.94 ;
        RECT 53.29 69.92 53.55 70.18 ;
        RECT 53.29 69.16 53.55 69.42 ;
        RECT 54.05 91.2 54.31 91.46 ;
        RECT 54.05 90.44 54.31 90.7 ;
        RECT 54.05 89.68 54.31 89.94 ;
        RECT 54.05 88.92 54.31 89.18 ;
        RECT 54.05 88.16 54.31 88.42 ;
        RECT 54.05 87.4 54.31 87.66 ;
        RECT 54.05 86.64 54.31 86.9 ;
        RECT 54.05 85.88 54.31 86.14 ;
        RECT 54.05 85.12 54.31 85.38 ;
        RECT 54.05 84.36 54.31 84.62 ;
        RECT 54.05 83.6 54.31 83.86 ;
        RECT 54.05 82.84 54.31 83.1 ;
        RECT 54.05 82.08 54.31 82.34 ;
        RECT 54.05 81.32 54.31 81.58 ;
        RECT 54.05 80.56 54.31 80.82 ;
        RECT 54.05 79.8 54.31 80.06 ;
        RECT 54.05 79.04 54.31 79.3 ;
        RECT 54.05 78.28 54.31 78.54 ;
        RECT 54.05 77.52 54.31 77.78 ;
        RECT 54.05 76.76 54.31 77.02 ;
        RECT 54.05 76 54.31 76.26 ;
        RECT 54.05 75.24 54.31 75.5 ;
        RECT 54.05 74.48 54.31 74.74 ;
        RECT 54.05 73.72 54.31 73.98 ;
        RECT 54.05 72.96 54.31 73.22 ;
        RECT 54.05 72.2 54.31 72.46 ;
        RECT 54.05 71.44 54.31 71.7 ;
        RECT 54.05 70.68 54.31 70.94 ;
        RECT 54.05 69.92 54.31 70.18 ;
        RECT 54.05 69.16 54.31 69.42 ;
        RECT 54.81 91.2 55.07 91.46 ;
        RECT 54.81 90.44 55.07 90.7 ;
        RECT 54.81 89.68 55.07 89.94 ;
        RECT 54.81 88.92 55.07 89.18 ;
        RECT 54.81 88.16 55.07 88.42 ;
        RECT 54.81 87.4 55.07 87.66 ;
        RECT 54.81 86.64 55.07 86.9 ;
        RECT 54.81 85.88 55.07 86.14 ;
        RECT 54.81 85.12 55.07 85.38 ;
        RECT 54.81 84.36 55.07 84.62 ;
        RECT 54.81 83.6 55.07 83.86 ;
        RECT 54.81 82.84 55.07 83.1 ;
        RECT 54.81 82.08 55.07 82.34 ;
        RECT 54.81 81.32 55.07 81.58 ;
        RECT 54.81 80.56 55.07 80.82 ;
        RECT 54.81 79.8 55.07 80.06 ;
        RECT 54.81 79.04 55.07 79.3 ;
        RECT 54.81 78.28 55.07 78.54 ;
        RECT 54.81 77.52 55.07 77.78 ;
        RECT 54.81 76.76 55.07 77.02 ;
        RECT 4.65 91.2 4.91 91.46 ;
        RECT 4.65 90.44 4.91 90.7 ;
        RECT 4.65 89.68 4.91 89.94 ;
        RECT 4.65 88.92 4.91 89.18 ;
        RECT 4.65 88.16 4.91 88.42 ;
        RECT 4.65 87.4 4.91 87.66 ;
        RECT 4.65 86.64 4.91 86.9 ;
        RECT 4.65 85.88 4.91 86.14 ;
        RECT 4.65 85.12 4.91 85.38 ;
        RECT 4.65 84.36 4.91 84.62 ;
        RECT 4.65 83.6 4.91 83.86 ;
        RECT 4.65 82.84 4.91 83.1 ;
        RECT 4.65 82.08 4.91 82.34 ;
        RECT 4.65 81.32 4.91 81.58 ;
        RECT 4.65 80.56 4.91 80.82 ;
        RECT 4.65 79.8 4.91 80.06 ;
        RECT 4.65 79.04 4.91 79.3 ;
        RECT 4.65 78.28 4.91 78.54 ;
        RECT 4.65 77.52 4.91 77.78 ;
        RECT 4.65 76.76 4.91 77.02 ;
        RECT 4.65 76 4.91 76.26 ;
        RECT 4.65 75.24 4.91 75.5 ;
        RECT 4.65 74.48 4.91 74.74 ;
        RECT 4.65 73.72 4.91 73.98 ;
        RECT 4.65 72.96 4.91 73.22 ;
        RECT 4.65 72.2 4.91 72.46 ;
        RECT 4.65 71.44 4.91 71.7 ;
        RECT 4.65 70.68 4.91 70.94 ;
        RECT 4.65 69.92 4.91 70.18 ;
        RECT 4.65 69.16 4.91 69.42 ;
        RECT 5.41 91.2 5.67 91.46 ;
        RECT 5.41 90.44 5.67 90.7 ;
        RECT 5.41 89.68 5.67 89.94 ;
        RECT 5.41 88.92 5.67 89.18 ;
        RECT 5.41 88.16 5.67 88.42 ;
        RECT 5.41 87.4 5.67 87.66 ;
        RECT 5.41 86.64 5.67 86.9 ;
        RECT 5.41 85.88 5.67 86.14 ;
        RECT 5.41 85.12 5.67 85.38 ;
        RECT 5.41 84.36 5.67 84.62 ;
        RECT 5.41 83.6 5.67 83.86 ;
        RECT 5.41 82.84 5.67 83.1 ;
        RECT 5.41 82.08 5.67 82.34 ;
        RECT 5.41 81.32 5.67 81.58 ;
        RECT 5.41 80.56 5.67 80.82 ;
        RECT 5.41 79.8 5.67 80.06 ;
        RECT 5.41 79.04 5.67 79.3 ;
        RECT 5.41 78.28 5.67 78.54 ;
        RECT 5.41 77.52 5.67 77.78 ;
        RECT 5.41 76.76 5.67 77.02 ;
        RECT 5.41 76 5.67 76.26 ;
        RECT 5.41 75.24 5.67 75.5 ;
        RECT 5.41 74.48 5.67 74.74 ;
        RECT 5.41 73.72 5.67 73.98 ;
        RECT 5.41 72.96 5.67 73.22 ;
        RECT 5.41 72.2 5.67 72.46 ;
        RECT 5.41 71.44 5.67 71.7 ;
        RECT 5.41 70.68 5.67 70.94 ;
        RECT 5.41 69.92 5.67 70.18 ;
        RECT 5.41 69.16 5.67 69.42 ;
        RECT 6.17 91.2 6.43 91.46 ;
        RECT 6.17 90.44 6.43 90.7 ;
        RECT 6.17 89.68 6.43 89.94 ;
        RECT 6.17 88.92 6.43 89.18 ;
        RECT 6.17 88.16 6.43 88.42 ;
        RECT 6.17 87.4 6.43 87.66 ;
        RECT 6.17 86.64 6.43 86.9 ;
        RECT 6.17 85.88 6.43 86.14 ;
        RECT 6.17 85.12 6.43 85.38 ;
        RECT 6.17 84.36 6.43 84.62 ;
        RECT 6.17 83.6 6.43 83.86 ;
        RECT 6.17 82.84 6.43 83.1 ;
        RECT 6.17 82.08 6.43 82.34 ;
        RECT 6.17 81.32 6.43 81.58 ;
        RECT 6.17 80.56 6.43 80.82 ;
        RECT 6.17 79.8 6.43 80.06 ;
        RECT 6.17 79.04 6.43 79.3 ;
        RECT 6.17 78.28 6.43 78.54 ;
        RECT 6.17 77.52 6.43 77.78 ;
        RECT 6.17 76.76 6.43 77.02 ;
        RECT 6.17 76 6.43 76.26 ;
        RECT 6.17 75.24 6.43 75.5 ;
        RECT 6.17 74.48 6.43 74.74 ;
        RECT 6.17 73.72 6.43 73.98 ;
        RECT 6.17 72.96 6.43 73.22 ;
        RECT 6.17 72.2 6.43 72.46 ;
        RECT 6.17 71.44 6.43 71.7 ;
        RECT 6.17 70.68 6.43 70.94 ;
        RECT 6.17 69.92 6.43 70.18 ;
        RECT 6.17 69.16 6.43 69.42 ;
        RECT 6.93 91.2 7.19 91.46 ;
        RECT 6.93 90.44 7.19 90.7 ;
        RECT 6.93 89.68 7.19 89.94 ;
        RECT 6.93 88.92 7.19 89.18 ;
        RECT 6.93 88.16 7.19 88.42 ;
        RECT 6.93 87.4 7.19 87.66 ;
        RECT 6.93 86.64 7.19 86.9 ;
        RECT 6.93 85.88 7.19 86.14 ;
        RECT 6.93 85.12 7.19 85.38 ;
        RECT 6.93 84.36 7.19 84.62 ;
        RECT 6.93 83.6 7.19 83.86 ;
        RECT 6.93 82.84 7.19 83.1 ;
        RECT 6.93 82.08 7.19 82.34 ;
        RECT 6.93 81.32 7.19 81.58 ;
        RECT 6.93 80.56 7.19 80.82 ;
        RECT 6.93 79.8 7.19 80.06 ;
        RECT 6.93 79.04 7.19 79.3 ;
        RECT 6.93 78.28 7.19 78.54 ;
        RECT 6.93 77.52 7.19 77.78 ;
        RECT 6.93 76.76 7.19 77.02 ;
        RECT 6.93 76 7.19 76.26 ;
        RECT 6.93 75.24 7.19 75.5 ;
        RECT 6.93 74.48 7.19 74.74 ;
        RECT 6.93 73.72 7.19 73.98 ;
        RECT 6.93 72.96 7.19 73.22 ;
        RECT 6.93 72.2 7.19 72.46 ;
        RECT 6.93 71.44 7.19 71.7 ;
        RECT 6.93 70.68 7.19 70.94 ;
        RECT 6.93 69.92 7.19 70.18 ;
        RECT 6.93 69.16 7.19 69.42 ;
        RECT 7.69 91.2 7.95 91.46 ;
        RECT 7.69 90.44 7.95 90.7 ;
        RECT 7.69 89.68 7.95 89.94 ;
        RECT 7.69 88.92 7.95 89.18 ;
        RECT 7.69 88.16 7.95 88.42 ;
        RECT 7.69 87.4 7.95 87.66 ;
        RECT 7.69 86.64 7.95 86.9 ;
        RECT 7.69 85.88 7.95 86.14 ;
        RECT 7.69 85.12 7.95 85.38 ;
        RECT 7.69 84.36 7.95 84.62 ;
        RECT 7.69 83.6 7.95 83.86 ;
        RECT 7.69 82.84 7.95 83.1 ;
        RECT 7.69 82.08 7.95 82.34 ;
        RECT 7.69 81.32 7.95 81.58 ;
        RECT 7.69 80.56 7.95 80.82 ;
        RECT 7.69 79.8 7.95 80.06 ;
        RECT 7.69 79.04 7.95 79.3 ;
        RECT 7.69 78.28 7.95 78.54 ;
        RECT 7.69 77.52 7.95 77.78 ;
        RECT 7.69 76.76 7.95 77.02 ;
        RECT 7.69 76 7.95 76.26 ;
        RECT 7.69 75.24 7.95 75.5 ;
        RECT 7.69 74.48 7.95 74.74 ;
        RECT 7.69 73.72 7.95 73.98 ;
        RECT 7.69 72.96 7.95 73.22 ;
        RECT 7.69 72.2 7.95 72.46 ;
        RECT 7.69 71.44 7.95 71.7 ;
        RECT 7.69 70.68 7.95 70.94 ;
        RECT 7.69 69.92 7.95 70.18 ;
        RECT 7.69 69.16 7.95 69.42 ;
        RECT 8.45 91.2 8.71 91.46 ;
        RECT 8.45 90.44 8.71 90.7 ;
        RECT 8.45 89.68 8.71 89.94 ;
        RECT 8.45 88.92 8.71 89.18 ;
        RECT 8.45 88.16 8.71 88.42 ;
        RECT 8.45 87.4 8.71 87.66 ;
        RECT 8.45 86.64 8.71 86.9 ;
        RECT 8.45 85.88 8.71 86.14 ;
        RECT 8.45 85.12 8.71 85.38 ;
        RECT 8.45 84.36 8.71 84.62 ;
        RECT 8.45 83.6 8.71 83.86 ;
        RECT 8.45 82.84 8.71 83.1 ;
        RECT 8.45 82.08 8.71 82.34 ;
        RECT 8.45 81.32 8.71 81.58 ;
        RECT 8.45 80.56 8.71 80.82 ;
        RECT 8.45 79.8 8.71 80.06 ;
        RECT 8.45 79.04 8.71 79.3 ;
        RECT 8.45 78.28 8.71 78.54 ;
        RECT 8.45 77.52 8.71 77.78 ;
        RECT 8.45 76.76 8.71 77.02 ;
        RECT 8.45 76 8.71 76.26 ;
        RECT 8.45 75.24 8.71 75.5 ;
        RECT 8.45 74.48 8.71 74.74 ;
        RECT 8.45 73.72 8.71 73.98 ;
        RECT 8.45 72.96 8.71 73.22 ;
        RECT 8.45 72.2 8.71 72.46 ;
        RECT 8.45 71.44 8.71 71.7 ;
        RECT 8.45 70.68 8.71 70.94 ;
        RECT 8.45 69.92 8.71 70.18 ;
        RECT 8.45 69.16 8.71 69.42 ;
        RECT 9.21 91.2 9.47 91.46 ;
        RECT 9.21 90.44 9.47 90.7 ;
        RECT 9.21 89.68 9.47 89.94 ;
        RECT 9.21 88.92 9.47 89.18 ;
        RECT 9.21 88.16 9.47 88.42 ;
        RECT 9.21 87.4 9.47 87.66 ;
        RECT 9.21 86.64 9.47 86.9 ;
        RECT 9.21 85.88 9.47 86.14 ;
        RECT 9.21 85.12 9.47 85.38 ;
        RECT 9.21 84.36 9.47 84.62 ;
        RECT 9.21 83.6 9.47 83.86 ;
        RECT 9.21 82.84 9.47 83.1 ;
        RECT 9.21 82.08 9.47 82.34 ;
        RECT 9.21 81.32 9.47 81.58 ;
        RECT 9.21 80.56 9.47 80.82 ;
        RECT 9.21 79.8 9.47 80.06 ;
        RECT 9.21 79.04 9.47 79.3 ;
        RECT 9.21 78.28 9.47 78.54 ;
        RECT 9.21 77.52 9.47 77.78 ;
        RECT 9.21 76.76 9.47 77.02 ;
        RECT 9.21 76 9.47 76.26 ;
        RECT 9.21 75.24 9.47 75.5 ;
        RECT 9.21 74.48 9.47 74.74 ;
        RECT 9.21 73.72 9.47 73.98 ;
        RECT 9.21 72.96 9.47 73.22 ;
        RECT 9.21 72.2 9.47 72.46 ;
        RECT 9.21 71.44 9.47 71.7 ;
        RECT 9.21 70.68 9.47 70.94 ;
        RECT 9.21 69.92 9.47 70.18 ;
        RECT 9.21 69.16 9.47 69.42 ;
        RECT 9.97 91.2 10.23 91.46 ;
        RECT 9.97 90.44 10.23 90.7 ;
        RECT 9.97 89.68 10.23 89.94 ;
        RECT 9.97 88.92 10.23 89.18 ;
        RECT 9.97 88.16 10.23 88.42 ;
        RECT 9.97 87.4 10.23 87.66 ;
        RECT 9.97 86.64 10.23 86.9 ;
        RECT 9.97 85.88 10.23 86.14 ;
        RECT 9.97 85.12 10.23 85.38 ;
        RECT 9.97 84.36 10.23 84.62 ;
        RECT 9.97 83.6 10.23 83.86 ;
        RECT 9.97 82.84 10.23 83.1 ;
        RECT 9.97 82.08 10.23 82.34 ;
        RECT 9.97 81.32 10.23 81.58 ;
        RECT 9.97 80.56 10.23 80.82 ;
        RECT 9.97 79.8 10.23 80.06 ;
        RECT 9.97 79.04 10.23 79.3 ;
        RECT 9.97 78.28 10.23 78.54 ;
        RECT 9.97 77.52 10.23 77.78 ;
        RECT 9.97 76.76 10.23 77.02 ;
        RECT 9.97 76 10.23 76.26 ;
        RECT 9.97 75.24 10.23 75.5 ;
        RECT 9.97 74.48 10.23 74.74 ;
        RECT 9.97 73.72 10.23 73.98 ;
        RECT 9.97 72.96 10.23 73.22 ;
        RECT 9.97 72.2 10.23 72.46 ;
        RECT 9.97 71.44 10.23 71.7 ;
        RECT 9.97 70.68 10.23 70.94 ;
        RECT 9.97 69.92 10.23 70.18 ;
        RECT 9.97 69.16 10.23 69.42 ;
        RECT 10.73 91.2 10.99 91.46 ;
        RECT 10.73 90.44 10.99 90.7 ;
        RECT 10.73 89.68 10.99 89.94 ;
        RECT 10.73 88.92 10.99 89.18 ;
        RECT 10.73 88.16 10.99 88.42 ;
        RECT 10.73 87.4 10.99 87.66 ;
        RECT 10.73 86.64 10.99 86.9 ;
        RECT 10.73 85.88 10.99 86.14 ;
        RECT 10.73 85.12 10.99 85.38 ;
        RECT 10.73 84.36 10.99 84.62 ;
        RECT 10.73 83.6 10.99 83.86 ;
        RECT 10.73 82.84 10.99 83.1 ;
        RECT 10.73 82.08 10.99 82.34 ;
        RECT 10.73 81.32 10.99 81.58 ;
        RECT 10.73 80.56 10.99 80.82 ;
        RECT 10.73 79.8 10.99 80.06 ;
        RECT 10.73 79.04 10.99 79.3 ;
        RECT 10.73 78.28 10.99 78.54 ;
        RECT 10.73 77.52 10.99 77.78 ;
        RECT 10.73 76.76 10.99 77.02 ;
        RECT 10.73 76 10.99 76.26 ;
        RECT 10.73 75.24 10.99 75.5 ;
        RECT 10.73 74.48 10.99 74.74 ;
        RECT 10.73 73.72 10.99 73.98 ;
        RECT 10.73 72.96 10.99 73.22 ;
        RECT 10.73 72.2 10.99 72.46 ;
        RECT 10.73 71.44 10.99 71.7 ;
        RECT 10.73 70.68 10.99 70.94 ;
        RECT 10.73 69.92 10.99 70.18 ;
        RECT 10.73 69.16 10.99 69.42 ;
        RECT 11.49 91.2 11.75 91.46 ;
        RECT 11.49 90.44 11.75 90.7 ;
        RECT 11.49 89.68 11.75 89.94 ;
        RECT 11.49 88.92 11.75 89.18 ;
        RECT 11.49 88.16 11.75 88.42 ;
        RECT 11.49 87.4 11.75 87.66 ;
        RECT 11.49 86.64 11.75 86.9 ;
        RECT 11.49 85.88 11.75 86.14 ;
        RECT 11.49 85.12 11.75 85.38 ;
        RECT 11.49 84.36 11.75 84.62 ;
        RECT 11.49 83.6 11.75 83.86 ;
        RECT 11.49 82.84 11.75 83.1 ;
        RECT 11.49 82.08 11.75 82.34 ;
        RECT 11.49 81.32 11.75 81.58 ;
        RECT 11.49 80.56 11.75 80.82 ;
        RECT 11.49 79.8 11.75 80.06 ;
        RECT 11.49 79.04 11.75 79.3 ;
        RECT 11.49 78.28 11.75 78.54 ;
        RECT 11.49 77.52 11.75 77.78 ;
        RECT 11.49 76.76 11.75 77.02 ;
        RECT 11.49 76 11.75 76.26 ;
        RECT 11.49 75.24 11.75 75.5 ;
        RECT 11.49 74.48 11.75 74.74 ;
        RECT 11.49 73.72 11.75 73.98 ;
        RECT 11.49 72.96 11.75 73.22 ;
        RECT 11.49 72.2 11.75 72.46 ;
        RECT 11.49 71.44 11.75 71.7 ;
        RECT 11.49 70.68 11.75 70.94 ;
        RECT 11.49 69.92 11.75 70.18 ;
        RECT 11.49 69.16 11.75 69.42 ;
        RECT 12.25 91.2 12.51 91.46 ;
        RECT 12.25 90.44 12.51 90.7 ;
        RECT 12.25 89.68 12.51 89.94 ;
        RECT 12.25 88.92 12.51 89.18 ;
        RECT 12.25 88.16 12.51 88.42 ;
        RECT 12.25 87.4 12.51 87.66 ;
        RECT 12.25 86.64 12.51 86.9 ;
        RECT 12.25 85.88 12.51 86.14 ;
        RECT 12.25 85.12 12.51 85.38 ;
        RECT 12.25 84.36 12.51 84.62 ;
        RECT 12.25 83.6 12.51 83.86 ;
        RECT 12.25 82.84 12.51 83.1 ;
        RECT 12.25 82.08 12.51 82.34 ;
        RECT 12.25 81.32 12.51 81.58 ;
        RECT 12.25 80.56 12.51 80.82 ;
        RECT 12.25 79.8 12.51 80.06 ;
        RECT 12.25 79.04 12.51 79.3 ;
        RECT 12.25 78.28 12.51 78.54 ;
        RECT 12.25 77.52 12.51 77.78 ;
        RECT 12.25 76.76 12.51 77.02 ;
        RECT 12.25 76 12.51 76.26 ;
        RECT 12.25 75.24 12.51 75.5 ;
        RECT 12.25 74.48 12.51 74.74 ;
        RECT 12.25 73.72 12.51 73.98 ;
        RECT 12.25 72.96 12.51 73.22 ;
        RECT 12.25 72.2 12.51 72.46 ;
        RECT 12.25 71.44 12.51 71.7 ;
        RECT 12.25 70.68 12.51 70.94 ;
        RECT 12.25 69.92 12.51 70.18 ;
        RECT 12.25 69.16 12.51 69.42 ;
        RECT 13.01 91.2 13.27 91.46 ;
        RECT 13.01 90.44 13.27 90.7 ;
        RECT 13.01 89.68 13.27 89.94 ;
        RECT 13.01 88.92 13.27 89.18 ;
        RECT 13.01 88.16 13.27 88.42 ;
        RECT 13.01 87.4 13.27 87.66 ;
        RECT 13.01 86.64 13.27 86.9 ;
        RECT 13.01 85.88 13.27 86.14 ;
        RECT 13.01 85.12 13.27 85.38 ;
        RECT 13.01 84.36 13.27 84.62 ;
        RECT 13.01 83.6 13.27 83.86 ;
        RECT 13.01 82.84 13.27 83.1 ;
        RECT 13.01 82.08 13.27 82.34 ;
        RECT 13.01 81.32 13.27 81.58 ;
        RECT 13.01 80.56 13.27 80.82 ;
        RECT 13.01 79.8 13.27 80.06 ;
        RECT 13.01 79.04 13.27 79.3 ;
        RECT 13.01 78.28 13.27 78.54 ;
        RECT 13.01 77.52 13.27 77.78 ;
        RECT 13.01 76.76 13.27 77.02 ;
        RECT 13.01 76 13.27 76.26 ;
        RECT 13.01 75.24 13.27 75.5 ;
        RECT 13.01 74.48 13.27 74.74 ;
        RECT 13.01 73.72 13.27 73.98 ;
        RECT 13.01 72.96 13.27 73.22 ;
        RECT 13.01 72.2 13.27 72.46 ;
        RECT 13.01 71.44 13.27 71.7 ;
        RECT 13.01 70.68 13.27 70.94 ;
        RECT 13.01 69.92 13.27 70.18 ;
        RECT 13.01 69.16 13.27 69.42 ;
        RECT 13.77 91.2 14.03 91.46 ;
        RECT 13.77 90.44 14.03 90.7 ;
        RECT 13.77 89.68 14.03 89.94 ;
        RECT 13.77 88.92 14.03 89.18 ;
        RECT 13.77 88.16 14.03 88.42 ;
        RECT 13.77 87.4 14.03 87.66 ;
        RECT 13.77 86.64 14.03 86.9 ;
        RECT 13.77 85.88 14.03 86.14 ;
        RECT 13.77 85.12 14.03 85.38 ;
        RECT 13.77 84.36 14.03 84.62 ;
        RECT 13.77 83.6 14.03 83.86 ;
        RECT 13.77 82.84 14.03 83.1 ;
        RECT 13.77 82.08 14.03 82.34 ;
        RECT 13.77 81.32 14.03 81.58 ;
        RECT 13.77 80.56 14.03 80.82 ;
        RECT 13.77 79.8 14.03 80.06 ;
        RECT 13.77 79.04 14.03 79.3 ;
        RECT 13.77 78.28 14.03 78.54 ;
        RECT 13.77 77.52 14.03 77.78 ;
        RECT 13.77 76.76 14.03 77.02 ;
        RECT 13.77 76 14.03 76.26 ;
        RECT 13.77 75.24 14.03 75.5 ;
        RECT 13.77 74.48 14.03 74.74 ;
        RECT 13.77 73.72 14.03 73.98 ;
        RECT 13.77 72.96 14.03 73.22 ;
        RECT 13.77 72.2 14.03 72.46 ;
        RECT 13.77 71.44 14.03 71.7 ;
        RECT 13.77 70.68 14.03 70.94 ;
        RECT 13.77 69.92 14.03 70.18 ;
        RECT 13.77 69.16 14.03 69.42 ;
        RECT 14.53 91.2 14.79 91.46 ;
        RECT 14.53 90.44 14.79 90.7 ;
        RECT 14.53 89.68 14.79 89.94 ;
        RECT 14.53 88.92 14.79 89.18 ;
        RECT 14.53 88.16 14.79 88.42 ;
        RECT 14.53 87.4 14.79 87.66 ;
        RECT 14.53 86.64 14.79 86.9 ;
        RECT 14.53 85.88 14.79 86.14 ;
        RECT 14.53 85.12 14.79 85.38 ;
        RECT 14.53 84.36 14.79 84.62 ;
        RECT 14.53 83.6 14.79 83.86 ;
        RECT 14.53 82.84 14.79 83.1 ;
        RECT 14.53 82.08 14.79 82.34 ;
        RECT 14.53 81.32 14.79 81.58 ;
        RECT 14.53 80.56 14.79 80.82 ;
        RECT 14.53 79.8 14.79 80.06 ;
        RECT 14.53 79.04 14.79 79.3 ;
        RECT 14.53 78.28 14.79 78.54 ;
        RECT 14.53 77.52 14.79 77.78 ;
        RECT 14.53 76.76 14.79 77.02 ;
        RECT 14.53 76 14.79 76.26 ;
        RECT 14.53 75.24 14.79 75.5 ;
        RECT 14.53 74.48 14.79 74.74 ;
        RECT 14.53 73.72 14.79 73.98 ;
        RECT 14.53 72.96 14.79 73.22 ;
        RECT 14.53 72.2 14.79 72.46 ;
        RECT 14.53 71.44 14.79 71.7 ;
        RECT 14.53 70.68 14.79 70.94 ;
        RECT 14.53 69.92 14.79 70.18 ;
        RECT 14.53 69.16 14.79 69.42 ;
        RECT 15.29 91.2 15.55 91.46 ;
        RECT 15.29 90.44 15.55 90.7 ;
        RECT 15.29 89.68 15.55 89.94 ;
        RECT 15.29 88.92 15.55 89.18 ;
        RECT 15.29 88.16 15.55 88.42 ;
        RECT 15.29 87.4 15.55 87.66 ;
        RECT 15.29 86.64 15.55 86.9 ;
        RECT 15.29 85.88 15.55 86.14 ;
        RECT 15.29 85.12 15.55 85.38 ;
        RECT 15.29 84.36 15.55 84.62 ;
        RECT 15.29 83.6 15.55 83.86 ;
        RECT 15.29 82.84 15.55 83.1 ;
        RECT 15.29 82.08 15.55 82.34 ;
        RECT 15.29 81.32 15.55 81.58 ;
        RECT 15.29 80.56 15.55 80.82 ;
        RECT 15.29 79.8 15.55 80.06 ;
        RECT 15.29 79.04 15.55 79.3 ;
        RECT 15.29 78.28 15.55 78.54 ;
        RECT 15.29 77.52 15.55 77.78 ;
        RECT 15.29 76.76 15.55 77.02 ;
        RECT 15.29 76 15.55 76.26 ;
        RECT 15.29 75.24 15.55 75.5 ;
        RECT 15.29 74.48 15.55 74.74 ;
        RECT 15.29 73.72 15.55 73.98 ;
        RECT 15.29 72.96 15.55 73.22 ;
        RECT 15.29 72.2 15.55 72.46 ;
        RECT 15.29 71.44 15.55 71.7 ;
        RECT 15.29 70.68 15.55 70.94 ;
        RECT 15.29 69.92 15.55 70.18 ;
        RECT 15.29 69.16 15.55 69.42 ;
        RECT 16.05 91.2 16.31 91.46 ;
        RECT 16.05 90.44 16.31 90.7 ;
        RECT 16.05 89.68 16.31 89.94 ;
        RECT 16.05 88.92 16.31 89.18 ;
        RECT 16.05 88.16 16.31 88.42 ;
        RECT 16.05 87.4 16.31 87.66 ;
        RECT 16.05 86.64 16.31 86.9 ;
        RECT 16.05 85.88 16.31 86.14 ;
        RECT 16.05 85.12 16.31 85.38 ;
        RECT 16.05 84.36 16.31 84.62 ;
        RECT 16.05 83.6 16.31 83.86 ;
        RECT 16.05 82.84 16.31 83.1 ;
        RECT 16.05 82.08 16.31 82.34 ;
        RECT 16.05 81.32 16.31 81.58 ;
        RECT 16.05 80.56 16.31 80.82 ;
        RECT 16.05 79.8 16.31 80.06 ;
        RECT 16.05 79.04 16.31 79.3 ;
        RECT 16.05 78.28 16.31 78.54 ;
        RECT 16.05 77.52 16.31 77.78 ;
        RECT 16.05 76.76 16.31 77.02 ;
        RECT 16.05 76 16.31 76.26 ;
        RECT 16.05 75.24 16.31 75.5 ;
        RECT 16.05 74.48 16.31 74.74 ;
        RECT 16.05 73.72 16.31 73.98 ;
        RECT 16.05 72.96 16.31 73.22 ;
        RECT 16.05 72.2 16.31 72.46 ;
        RECT 16.05 71.44 16.31 71.7 ;
        RECT 16.05 70.68 16.31 70.94 ;
        RECT 16.05 69.92 16.31 70.18 ;
        RECT 16.05 69.16 16.31 69.42 ;
        RECT 16.81 91.2 17.07 91.46 ;
        RECT 16.81 90.44 17.07 90.7 ;
        RECT 16.81 89.68 17.07 89.94 ;
        RECT 16.81 88.92 17.07 89.18 ;
        RECT 16.81 88.16 17.07 88.42 ;
        RECT 16.81 87.4 17.07 87.66 ;
        RECT 16.81 86.64 17.07 86.9 ;
        RECT 16.81 85.88 17.07 86.14 ;
        RECT 16.81 85.12 17.07 85.38 ;
        RECT 16.81 84.36 17.07 84.62 ;
        RECT 16.81 83.6 17.07 83.86 ;
        RECT 16.81 82.84 17.07 83.1 ;
        RECT 16.81 82.08 17.07 82.34 ;
        RECT 16.81 81.32 17.07 81.58 ;
        RECT 16.81 80.56 17.07 80.82 ;
        RECT 16.81 79.8 17.07 80.06 ;
        RECT 16.81 79.04 17.07 79.3 ;
        RECT 16.81 78.28 17.07 78.54 ;
        RECT 16.81 77.52 17.07 77.78 ;
        RECT 16.81 76.76 17.07 77.02 ;
        RECT 16.81 76 17.07 76.26 ;
        RECT 16.81 75.24 17.07 75.5 ;
        RECT 16.81 74.48 17.07 74.74 ;
        RECT 16.81 73.72 17.07 73.98 ;
        RECT 16.81 72.96 17.07 73.22 ;
        RECT 16.81 72.2 17.07 72.46 ;
        RECT 16.81 71.44 17.07 71.7 ;
        RECT 16.81 70.68 17.07 70.94 ;
        RECT 16.81 69.92 17.07 70.18 ;
        RECT 16.81 69.16 17.07 69.42 ;
        RECT 17.57 91.2 17.83 91.46 ;
        RECT 17.57 90.44 17.83 90.7 ;
        RECT 17.57 89.68 17.83 89.94 ;
        RECT 17.57 88.92 17.83 89.18 ;
        RECT 17.57 88.16 17.83 88.42 ;
        RECT 17.57 87.4 17.83 87.66 ;
        RECT 17.57 86.64 17.83 86.9 ;
        RECT 17.57 85.88 17.83 86.14 ;
        RECT 17.57 85.12 17.83 85.38 ;
        RECT 17.57 84.36 17.83 84.62 ;
        RECT 17.57 83.6 17.83 83.86 ;
        RECT 17.57 82.84 17.83 83.1 ;
        RECT 17.57 82.08 17.83 82.34 ;
        RECT 17.57 81.32 17.83 81.58 ;
        RECT 17.57 80.56 17.83 80.82 ;
        RECT 17.57 79.8 17.83 80.06 ;
        RECT 17.57 79.04 17.83 79.3 ;
        RECT 17.57 78.28 17.83 78.54 ;
        RECT 17.57 77.52 17.83 77.78 ;
        RECT 17.57 76.76 17.83 77.02 ;
        RECT 17.57 76 17.83 76.26 ;
        RECT 17.57 75.24 17.83 75.5 ;
        RECT 17.57 74.48 17.83 74.74 ;
        RECT 17.57 73.72 17.83 73.98 ;
        RECT 17.57 72.96 17.83 73.22 ;
        RECT 17.57 72.2 17.83 72.46 ;
        RECT 17.57 71.44 17.83 71.7 ;
        RECT 17.57 70.68 17.83 70.94 ;
        RECT 17.57 69.92 17.83 70.18 ;
        RECT 17.57 69.16 17.83 69.42 ;
        RECT 18.33 91.2 18.59 91.46 ;
        RECT 18.33 90.44 18.59 90.7 ;
        RECT 18.33 89.68 18.59 89.94 ;
        RECT 18.33 88.92 18.59 89.18 ;
        RECT 18.33 88.16 18.59 88.42 ;
        RECT 18.33 87.4 18.59 87.66 ;
        RECT 18.33 86.64 18.59 86.9 ;
        RECT 18.33 85.88 18.59 86.14 ;
        RECT 18.33 85.12 18.59 85.38 ;
        RECT 18.33 84.36 18.59 84.62 ;
        RECT 18.33 83.6 18.59 83.86 ;
        RECT 18.33 82.84 18.59 83.1 ;
        RECT 18.33 82.08 18.59 82.34 ;
        RECT 18.33 81.32 18.59 81.58 ;
        RECT 18.33 80.56 18.59 80.82 ;
        RECT 18.33 79.8 18.59 80.06 ;
        RECT 18.33 79.04 18.59 79.3 ;
        RECT 18.33 78.28 18.59 78.54 ;
        RECT 18.33 77.52 18.59 77.78 ;
        RECT 18.33 76.76 18.59 77.02 ;
        RECT 18.33 76 18.59 76.26 ;
        RECT 18.33 75.24 18.59 75.5 ;
        RECT 18.33 74.48 18.59 74.74 ;
        RECT 18.33 73.72 18.59 73.98 ;
        RECT 18.33 72.96 18.59 73.22 ;
        RECT 18.33 72.2 18.59 72.46 ;
        RECT 18.33 71.44 18.59 71.7 ;
        RECT 18.33 70.68 18.59 70.94 ;
        RECT 18.33 69.92 18.59 70.18 ;
        RECT 18.33 69.16 18.59 69.42 ;
        RECT 19.09 91.2 19.35 91.46 ;
        RECT 19.09 90.44 19.35 90.7 ;
        RECT 19.09 89.68 19.35 89.94 ;
        RECT 19.09 88.92 19.35 89.18 ;
        RECT 19.09 88.16 19.35 88.42 ;
        RECT 19.09 87.4 19.35 87.66 ;
        RECT 19.09 86.64 19.35 86.9 ;
        RECT 19.09 85.88 19.35 86.14 ;
        RECT 19.09 85.12 19.35 85.38 ;
        RECT 19.09 84.36 19.35 84.62 ;
        RECT 19.09 83.6 19.35 83.86 ;
        RECT 19.09 82.84 19.35 83.1 ;
        RECT 19.09 82.08 19.35 82.34 ;
        RECT 19.09 81.32 19.35 81.58 ;
        RECT 19.09 80.56 19.35 80.82 ;
        RECT 19.09 79.8 19.35 80.06 ;
        RECT 19.09 79.04 19.35 79.3 ;
        RECT 19.09 78.28 19.35 78.54 ;
        RECT 19.09 77.52 19.35 77.78 ;
        RECT 19.09 76.76 19.35 77.02 ;
        RECT 19.09 76 19.35 76.26 ;
        RECT 19.09 75.24 19.35 75.5 ;
        RECT 19.09 74.48 19.35 74.74 ;
        RECT 19.09 73.72 19.35 73.98 ;
        RECT 19.09 72.96 19.35 73.22 ;
        RECT 19.09 72.2 19.35 72.46 ;
        RECT 19.09 71.44 19.35 71.7 ;
        RECT 19.09 70.68 19.35 70.94 ;
        RECT 19.09 69.92 19.35 70.18 ;
        RECT 19.09 69.16 19.35 69.42 ;
        RECT 19.85 91.2 20.11 91.46 ;
        RECT 19.85 90.44 20.11 90.7 ;
        RECT 19.85 89.68 20.11 89.94 ;
        RECT 19.85 88.92 20.11 89.18 ;
        RECT 19.85 88.16 20.11 88.42 ;
        RECT 19.85 87.4 20.11 87.66 ;
        RECT 19.85 86.64 20.11 86.9 ;
        RECT 19.85 85.88 20.11 86.14 ;
        RECT 19.85 85.12 20.11 85.38 ;
        RECT 19.85 84.36 20.11 84.62 ;
        RECT 19.85 83.6 20.11 83.86 ;
        RECT 19.85 82.84 20.11 83.1 ;
        RECT 19.85 82.08 20.11 82.34 ;
        RECT 19.85 81.32 20.11 81.58 ;
        RECT 19.85 80.56 20.11 80.82 ;
        RECT 19.85 79.8 20.11 80.06 ;
        RECT 19.85 79.04 20.11 79.3 ;
        RECT 19.85 78.28 20.11 78.54 ;
        RECT 19.85 77.52 20.11 77.78 ;
        RECT 19.85 76.76 20.11 77.02 ;
        RECT 19.85 76 20.11 76.26 ;
        RECT 19.85 75.24 20.11 75.5 ;
        RECT 19.85 74.48 20.11 74.74 ;
        RECT 19.85 73.72 20.11 73.98 ;
        RECT 19.85 72.96 20.11 73.22 ;
        RECT 19.85 72.2 20.11 72.46 ;
        RECT 19.85 71.44 20.11 71.7 ;
        RECT 19.85 70.68 20.11 70.94 ;
        RECT 19.85 69.92 20.11 70.18 ;
        RECT 19.85 69.16 20.11 69.42 ;
        RECT 20.61 91.2 20.87 91.46 ;
        RECT 20.61 90.44 20.87 90.7 ;
        RECT 20.61 89.68 20.87 89.94 ;
        RECT 20.61 88.92 20.87 89.18 ;
        RECT 20.61 88.16 20.87 88.42 ;
        RECT 20.61 87.4 20.87 87.66 ;
        RECT 20.61 86.64 20.87 86.9 ;
        RECT 20.61 85.88 20.87 86.14 ;
        RECT 20.61 85.12 20.87 85.38 ;
        RECT 20.61 84.36 20.87 84.62 ;
        RECT 20.61 83.6 20.87 83.86 ;
        RECT 20.61 82.84 20.87 83.1 ;
        RECT 20.61 82.08 20.87 82.34 ;
        RECT 20.61 81.32 20.87 81.58 ;
        RECT 20.61 80.56 20.87 80.82 ;
        RECT 20.61 79.8 20.87 80.06 ;
        RECT 20.61 79.04 20.87 79.3 ;
        RECT 20.61 78.28 20.87 78.54 ;
        RECT 20.61 77.52 20.87 77.78 ;
        RECT 20.61 76.76 20.87 77.02 ;
        RECT 20.61 76 20.87 76.26 ;
        RECT 20.61 75.24 20.87 75.5 ;
        RECT 20.61 74.48 20.87 74.74 ;
        RECT 20.61 73.72 20.87 73.98 ;
        RECT 20.61 72.96 20.87 73.22 ;
        RECT 20.61 72.2 20.87 72.46 ;
        RECT 20.61 71.44 20.87 71.7 ;
        RECT 20.61 70.68 20.87 70.94 ;
        RECT 20.61 69.92 20.87 70.18 ;
        RECT 20.61 69.16 20.87 69.42 ;
        RECT 21.37 91.2 21.63 91.46 ;
        RECT 21.37 90.44 21.63 90.7 ;
        RECT 21.37 89.68 21.63 89.94 ;
        RECT 21.37 88.92 21.63 89.18 ;
        RECT 21.37 88.16 21.63 88.42 ;
        RECT 21.37 87.4 21.63 87.66 ;
        RECT 21.37 86.64 21.63 86.9 ;
        RECT 21.37 85.88 21.63 86.14 ;
        RECT 21.37 85.12 21.63 85.38 ;
        RECT 21.37 84.36 21.63 84.62 ;
        RECT 21.37 83.6 21.63 83.86 ;
        RECT 21.37 82.84 21.63 83.1 ;
        RECT 21.37 82.08 21.63 82.34 ;
        RECT 21.37 81.32 21.63 81.58 ;
        RECT 21.37 80.56 21.63 80.82 ;
        RECT 21.37 79.8 21.63 80.06 ;
        RECT 21.37 79.04 21.63 79.3 ;
        RECT 21.37 78.28 21.63 78.54 ;
        RECT 21.37 77.52 21.63 77.78 ;
        RECT 21.37 76.76 21.63 77.02 ;
        RECT 21.37 76 21.63 76.26 ;
        RECT 21.37 75.24 21.63 75.5 ;
        RECT 21.37 74.48 21.63 74.74 ;
        RECT 21.37 73.72 21.63 73.98 ;
        RECT 21.37 72.96 21.63 73.22 ;
        RECT 21.37 72.2 21.63 72.46 ;
        RECT 21.37 71.44 21.63 71.7 ;
        RECT 21.37 70.68 21.63 70.94 ;
        RECT 21.37 69.92 21.63 70.18 ;
        RECT 21.37 69.16 21.63 69.42 ;
        RECT 22.13 91.2 22.39 91.46 ;
        RECT 22.13 90.44 22.39 90.7 ;
        RECT 22.13 89.68 22.39 89.94 ;
        RECT 22.13 88.92 22.39 89.18 ;
        RECT 22.13 88.16 22.39 88.42 ;
        RECT 22.13 87.4 22.39 87.66 ;
        RECT 22.13 86.64 22.39 86.9 ;
        RECT 22.13 85.88 22.39 86.14 ;
        RECT 22.13 85.12 22.39 85.38 ;
        RECT 22.13 84.36 22.39 84.62 ;
        RECT 22.13 83.6 22.39 83.86 ;
        RECT 22.13 82.84 22.39 83.1 ;
        RECT 22.13 82.08 22.39 82.34 ;
        RECT 22.13 81.32 22.39 81.58 ;
        RECT 22.13 80.56 22.39 80.82 ;
        RECT 22.13 79.8 22.39 80.06 ;
        RECT 22.13 79.04 22.39 79.3 ;
        RECT 22.13 78.28 22.39 78.54 ;
        RECT 22.13 77.52 22.39 77.78 ;
        RECT 22.13 76.76 22.39 77.02 ;
        RECT 22.13 76 22.39 76.26 ;
        RECT 22.13 75.24 22.39 75.5 ;
        RECT 22.13 74.48 22.39 74.74 ;
        RECT 22.13 73.72 22.39 73.98 ;
        RECT 22.13 72.96 22.39 73.22 ;
        RECT 22.13 72.2 22.39 72.46 ;
        RECT 22.13 71.44 22.39 71.7 ;
        RECT 22.13 70.68 22.39 70.94 ;
        RECT 22.13 69.92 22.39 70.18 ;
        RECT 22.13 69.16 22.39 69.42 ;
        RECT 22.89 91.2 23.15 91.46 ;
        RECT 22.89 90.44 23.15 90.7 ;
        RECT 22.89 89.68 23.15 89.94 ;
        RECT 22.89 88.92 23.15 89.18 ;
        RECT 22.89 88.16 23.15 88.42 ;
        RECT 22.89 87.4 23.15 87.66 ;
        RECT 22.89 86.64 23.15 86.9 ;
        RECT 22.89 85.88 23.15 86.14 ;
        RECT 22.89 85.12 23.15 85.38 ;
        RECT 22.89 84.36 23.15 84.62 ;
        RECT 22.89 83.6 23.15 83.86 ;
        RECT 22.89 82.84 23.15 83.1 ;
        RECT 22.89 82.08 23.15 82.34 ;
        RECT 22.89 81.32 23.15 81.58 ;
        RECT 22.89 80.56 23.15 80.82 ;
        RECT 22.89 79.8 23.15 80.06 ;
        RECT 22.89 79.04 23.15 79.3 ;
        RECT 22.89 78.28 23.15 78.54 ;
        RECT 22.89 77.52 23.15 77.78 ;
        RECT 22.89 76.76 23.15 77.02 ;
        RECT 22.89 76 23.15 76.26 ;
        RECT 22.89 75.24 23.15 75.5 ;
        RECT 22.89 74.48 23.15 74.74 ;
        RECT 22.89 73.72 23.15 73.98 ;
        RECT 22.89 72.96 23.15 73.22 ;
        RECT 22.89 72.2 23.15 72.46 ;
        RECT 22.89 71.44 23.15 71.7 ;
        RECT 22.89 70.68 23.15 70.94 ;
        RECT 22.89 69.92 23.15 70.18 ;
        RECT 22.89 69.16 23.15 69.42 ;
        RECT 23.65 91.2 23.91 91.46 ;
        RECT 23.65 90.44 23.91 90.7 ;
        RECT 23.65 89.68 23.91 89.94 ;
        RECT 23.65 88.92 23.91 89.18 ;
        RECT 23.65 88.16 23.91 88.42 ;
        RECT 23.65 87.4 23.91 87.66 ;
        RECT 23.65 86.64 23.91 86.9 ;
        RECT 23.65 85.88 23.91 86.14 ;
        RECT 23.65 85.12 23.91 85.38 ;
        RECT 23.65 84.36 23.91 84.62 ;
        RECT 23.65 83.6 23.91 83.86 ;
        RECT 23.65 82.84 23.91 83.1 ;
        RECT 23.65 82.08 23.91 82.34 ;
        RECT 23.65 81.32 23.91 81.58 ;
        RECT 23.65 80.56 23.91 80.82 ;
        RECT 23.65 79.8 23.91 80.06 ;
        RECT 23.65 79.04 23.91 79.3 ;
        RECT 23.65 78.28 23.91 78.54 ;
        RECT 23.65 77.52 23.91 77.78 ;
        RECT 23.65 76.76 23.91 77.02 ;
        RECT 23.65 76 23.91 76.26 ;
        RECT 23.65 75.24 23.91 75.5 ;
        RECT 23.65 74.48 23.91 74.74 ;
        RECT 23.65 73.72 23.91 73.98 ;
        RECT 23.65 72.96 23.91 73.22 ;
        RECT 23.65 72.2 23.91 72.46 ;
        RECT 23.65 71.44 23.91 71.7 ;
        RECT 23.65 70.68 23.91 70.94 ;
        RECT 23.65 69.92 23.91 70.18 ;
        RECT 23.65 69.16 23.91 69.42 ;
        RECT 24.41 91.2 24.67 91.46 ;
        RECT 24.41 90.44 24.67 90.7 ;
        RECT 24.41 89.68 24.67 89.94 ;
        RECT 24.41 88.92 24.67 89.18 ;
        RECT 24.41 88.16 24.67 88.42 ;
        RECT 24.41 87.4 24.67 87.66 ;
        RECT 24.41 86.64 24.67 86.9 ;
        RECT 24.41 85.88 24.67 86.14 ;
        RECT 24.41 85.12 24.67 85.38 ;
        RECT 24.41 84.36 24.67 84.62 ;
        RECT 24.41 83.6 24.67 83.86 ;
        RECT 24.41 82.84 24.67 83.1 ;
        RECT 24.41 82.08 24.67 82.34 ;
        RECT 24.41 81.32 24.67 81.58 ;
        RECT 24.41 80.56 24.67 80.82 ;
        RECT 24.41 79.8 24.67 80.06 ;
        RECT 24.41 79.04 24.67 79.3 ;
        RECT 24.41 78.28 24.67 78.54 ;
        RECT 24.41 77.52 24.67 77.78 ;
        RECT 24.41 76.76 24.67 77.02 ;
        RECT 24.41 76 24.67 76.26 ;
        RECT 24.41 75.24 24.67 75.5 ;
        RECT 24.41 74.48 24.67 74.74 ;
        RECT 24.41 73.72 24.67 73.98 ;
        RECT 24.41 72.96 24.67 73.22 ;
        RECT 24.41 72.2 24.67 72.46 ;
        RECT 24.41 71.44 24.67 71.7 ;
        RECT 24.41 70.68 24.67 70.94 ;
        RECT 24.41 69.92 24.67 70.18 ;
        RECT 24.41 69.16 24.67 69.42 ;
        RECT 25.17 91.2 25.43 91.46 ;
        RECT 25.17 90.44 25.43 90.7 ;
        RECT 25.17 89.68 25.43 89.94 ;
        RECT 25.17 88.92 25.43 89.18 ;
        RECT 25.17 88.16 25.43 88.42 ;
        RECT 25.17 87.4 25.43 87.66 ;
        RECT 25.17 86.64 25.43 86.9 ;
        RECT 25.17 85.88 25.43 86.14 ;
        RECT 25.17 85.12 25.43 85.38 ;
        RECT 25.17 84.36 25.43 84.62 ;
        RECT 25.17 83.6 25.43 83.86 ;
        RECT 25.17 82.84 25.43 83.1 ;
        RECT 25.17 82.08 25.43 82.34 ;
        RECT 25.17 81.32 25.43 81.58 ;
        RECT 25.17 80.56 25.43 80.82 ;
        RECT 25.17 79.8 25.43 80.06 ;
        RECT 25.17 79.04 25.43 79.3 ;
        RECT 25.17 78.28 25.43 78.54 ;
        RECT 25.17 77.52 25.43 77.78 ;
        RECT 25.17 76.76 25.43 77.02 ;
        RECT 25.17 76 25.43 76.26 ;
        RECT 25.17 75.24 25.43 75.5 ;
        RECT 25.17 74.48 25.43 74.74 ;
        RECT 25.17 73.72 25.43 73.98 ;
        RECT 25.17 72.96 25.43 73.22 ;
        RECT 25.17 72.2 25.43 72.46 ;
        RECT 25.17 71.44 25.43 71.7 ;
        RECT 25.17 70.68 25.43 70.94 ;
        RECT 25.17 69.92 25.43 70.18 ;
        RECT 25.17 69.16 25.43 69.42 ;
        RECT 25.93 91.2 26.19 91.46 ;
        RECT 25.93 90.44 26.19 90.7 ;
        RECT 25.93 89.68 26.19 89.94 ;
        RECT 25.93 88.92 26.19 89.18 ;
        RECT 25.93 88.16 26.19 88.42 ;
        RECT 25.93 87.4 26.19 87.66 ;
        RECT 25.93 86.64 26.19 86.9 ;
        RECT 25.93 85.88 26.19 86.14 ;
        RECT 25.93 85.12 26.19 85.38 ;
        RECT 25.93 84.36 26.19 84.62 ;
        RECT 25.93 83.6 26.19 83.86 ;
        RECT 25.93 82.84 26.19 83.1 ;
        RECT 25.93 82.08 26.19 82.34 ;
        RECT 25.93 81.32 26.19 81.58 ;
        RECT 25.93 80.56 26.19 80.82 ;
        RECT 25.93 79.8 26.19 80.06 ;
        RECT 25.93 79.04 26.19 79.3 ;
        RECT 25.93 78.28 26.19 78.54 ;
        RECT 25.93 77.52 26.19 77.78 ;
        RECT 25.93 76.76 26.19 77.02 ;
        RECT 25.93 76 26.19 76.26 ;
        RECT 25.93 75.24 26.19 75.5 ;
        RECT 25.93 74.48 26.19 74.74 ;
        RECT 25.93 73.72 26.19 73.98 ;
        RECT 25.93 72.96 26.19 73.22 ;
        RECT 25.93 72.2 26.19 72.46 ;
        RECT 25.93 71.44 26.19 71.7 ;
        RECT 25.93 70.68 26.19 70.94 ;
        RECT 25.93 69.92 26.19 70.18 ;
        RECT 25.93 69.16 26.19 69.42 ;
        RECT 26.69 91.2 26.95 91.46 ;
        RECT 26.69 90.44 26.95 90.7 ;
        RECT 26.69 89.68 26.95 89.94 ;
        RECT 26.69 88.92 26.95 89.18 ;
        RECT 26.69 88.16 26.95 88.42 ;
        RECT 26.69 87.4 26.95 87.66 ;
        RECT 26.69 86.64 26.95 86.9 ;
        RECT 26.69 85.88 26.95 86.14 ;
        RECT 26.69 85.12 26.95 85.38 ;
        RECT 26.69 84.36 26.95 84.62 ;
        RECT 26.69 83.6 26.95 83.86 ;
        RECT 26.69 82.84 26.95 83.1 ;
        RECT 26.69 82.08 26.95 82.34 ;
        RECT 26.69 81.32 26.95 81.58 ;
        RECT 26.69 80.56 26.95 80.82 ;
        RECT 26.69 79.8 26.95 80.06 ;
        RECT 26.69 79.04 26.95 79.3 ;
        RECT 26.69 78.28 26.95 78.54 ;
        RECT 26.69 77.52 26.95 77.78 ;
        RECT 26.69 76.76 26.95 77.02 ;
        RECT 26.69 76 26.95 76.26 ;
        RECT 26.69 75.24 26.95 75.5 ;
        RECT 26.69 74.48 26.95 74.74 ;
        RECT 26.69 73.72 26.95 73.98 ;
        RECT 26.69 72.96 26.95 73.22 ;
        RECT 26.69 72.2 26.95 72.46 ;
        RECT 26.69 71.44 26.95 71.7 ;
        RECT 26.69 70.68 26.95 70.94 ;
        RECT 26.69 69.92 26.95 70.18 ;
        RECT 26.69 69.16 26.95 69.42 ;
        RECT 27.45 91.2 27.71 91.46 ;
        RECT 27.45 90.44 27.71 90.7 ;
        RECT 27.45 89.68 27.71 89.94 ;
        RECT 27.45 88.92 27.71 89.18 ;
        RECT 27.45 88.16 27.71 88.42 ;
        RECT 27.45 87.4 27.71 87.66 ;
        RECT 27.45 86.64 27.71 86.9 ;
        RECT 27.45 85.88 27.71 86.14 ;
        RECT 27.45 85.12 27.71 85.38 ;
        RECT 27.45 84.36 27.71 84.62 ;
        RECT 27.45 83.6 27.71 83.86 ;
        RECT 27.45 82.84 27.71 83.1 ;
        RECT 27.45 82.08 27.71 82.34 ;
        RECT 27.45 81.32 27.71 81.58 ;
        RECT 27.45 80.56 27.71 80.82 ;
        RECT 27.45 79.8 27.71 80.06 ;
        RECT 27.45 79.04 27.71 79.3 ;
        RECT 27.45 78.28 27.71 78.54 ;
        RECT 27.45 77.52 27.71 77.78 ;
        RECT 27.45 76.76 27.71 77.02 ;
        RECT 27.45 76 27.71 76.26 ;
        RECT 27.45 75.24 27.71 75.5 ;
        RECT 27.45 74.48 27.71 74.74 ;
        RECT 27.45 73.72 27.71 73.98 ;
        RECT 27.45 72.96 27.71 73.22 ;
        RECT 27.45 72.2 27.71 72.46 ;
        RECT 27.45 71.44 27.71 71.7 ;
        RECT 27.45 70.68 27.71 70.94 ;
        RECT 27.45 69.92 27.71 70.18 ;
        RECT 27.45 69.16 27.71 69.42 ;
        RECT 28.21 91.2 28.47 91.46 ;
        RECT 28.21 90.44 28.47 90.7 ;
        RECT 28.21 89.68 28.47 89.94 ;
        RECT 28.21 88.92 28.47 89.18 ;
        RECT 28.21 88.16 28.47 88.42 ;
        RECT 28.21 87.4 28.47 87.66 ;
        RECT 28.21 86.64 28.47 86.9 ;
        RECT 28.21 85.88 28.47 86.14 ;
        RECT 28.21 85.12 28.47 85.38 ;
        RECT 28.21 84.36 28.47 84.62 ;
        RECT 28.21 83.6 28.47 83.86 ;
        RECT 28.21 82.84 28.47 83.1 ;
        RECT 28.21 82.08 28.47 82.34 ;
        RECT 28.21 81.32 28.47 81.58 ;
        RECT 28.21 80.56 28.47 80.82 ;
        RECT 28.21 79.8 28.47 80.06 ;
        RECT 28.21 79.04 28.47 79.3 ;
        RECT 28.21 78.28 28.47 78.54 ;
        RECT 28.21 77.52 28.47 77.78 ;
        RECT 28.21 76.76 28.47 77.02 ;
        RECT 28.21 76 28.47 76.26 ;
        RECT 28.21 75.24 28.47 75.5 ;
        RECT 28.21 74.48 28.47 74.74 ;
        RECT 28.21 73.72 28.47 73.98 ;
        RECT 28.21 72.96 28.47 73.22 ;
        RECT 28.21 72.2 28.47 72.46 ;
        RECT 28.21 71.44 28.47 71.7 ;
        RECT 28.21 70.68 28.47 70.94 ;
        RECT 28.21 69.92 28.47 70.18 ;
        RECT 28.21 69.16 28.47 69.42 ;
        RECT 28.97 91.2 29.23 91.46 ;
        RECT 28.97 90.44 29.23 90.7 ;
        RECT 28.97 89.68 29.23 89.94 ;
        RECT 28.97 88.92 29.23 89.18 ;
        RECT 28.97 88.16 29.23 88.42 ;
        RECT 28.97 87.4 29.23 87.66 ;
        RECT 28.97 86.64 29.23 86.9 ;
        RECT 28.97 85.88 29.23 86.14 ;
        RECT 28.97 85.12 29.23 85.38 ;
        RECT 28.97 84.36 29.23 84.62 ;
        RECT 28.97 83.6 29.23 83.86 ;
        RECT 28.97 82.84 29.23 83.1 ;
        RECT 28.97 82.08 29.23 82.34 ;
        RECT 28.97 81.32 29.23 81.58 ;
        RECT 28.97 80.56 29.23 80.82 ;
        RECT 28.97 79.8 29.23 80.06 ;
        RECT 28.97 79.04 29.23 79.3 ;
        RECT 28.97 78.28 29.23 78.54 ;
        RECT 28.97 77.52 29.23 77.78 ;
        RECT 28.97 76.76 29.23 77.02 ;
        RECT 28.97 76 29.23 76.26 ;
        RECT 28.97 75.24 29.23 75.5 ;
        RECT 28.97 74.48 29.23 74.74 ;
        RECT 28.97 73.72 29.23 73.98 ;
        RECT 28.97 72.96 29.23 73.22 ;
        RECT 28.97 72.2 29.23 72.46 ;
        RECT 28.97 71.44 29.23 71.7 ;
        RECT 28.97 70.68 29.23 70.94 ;
        RECT 28.97 69.92 29.23 70.18 ;
        RECT 28.97 69.16 29.23 69.42 ;
        RECT 29.73 91.2 29.99 91.46 ;
        RECT 29.73 90.44 29.99 90.7 ;
        RECT 29.73 89.68 29.99 89.94 ;
        RECT 29.73 88.92 29.99 89.18 ;
        RECT 29.73 88.16 29.99 88.42 ;
        RECT 29.73 87.4 29.99 87.66 ;
        RECT 29.73 86.64 29.99 86.9 ;
        RECT 29.73 85.88 29.99 86.14 ;
        RECT 29.73 85.12 29.99 85.38 ;
        RECT 29.73 84.36 29.99 84.62 ;
    END
  END DVSS
  PIN AVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M3 ;
        RECT 0 22 100 32 ;
      LAYER M4 ;
        RECT 0 22 100 32 ;
      LAYER V4 ;
        RECT 80.65 30.215 80.91 30.475 ;
        RECT 80.65 29.455 80.91 29.715 ;
        RECT 80.65 28.695 80.91 28.955 ;
        RECT 80.65 27.935 80.91 28.195 ;
        RECT 80.65 27.175 80.91 27.435 ;
        RECT 80.65 26.415 80.91 26.675 ;
        RECT 80.65 25.655 80.91 25.915 ;
        RECT 80.65 24.895 80.91 25.155 ;
        RECT 80.65 24.135 80.91 24.395 ;
        RECT 80.65 23.375 80.91 23.635 ;
        RECT 81.41 30.215 81.67 30.475 ;
        RECT 81.41 29.455 81.67 29.715 ;
        RECT 81.41 28.695 81.67 28.955 ;
        RECT 81.41 27.935 81.67 28.195 ;
        RECT 81.41 27.175 81.67 27.435 ;
        RECT 81.41 26.415 81.67 26.675 ;
        RECT 81.41 25.655 81.67 25.915 ;
        RECT 81.41 24.895 81.67 25.155 ;
        RECT 81.41 24.135 81.67 24.395 ;
        RECT 81.41 23.375 81.67 23.635 ;
        RECT 82.17 30.215 82.43 30.475 ;
        RECT 82.17 29.455 82.43 29.715 ;
        RECT 82.17 28.695 82.43 28.955 ;
        RECT 82.17 27.935 82.43 28.195 ;
        RECT 82.17 27.175 82.43 27.435 ;
        RECT 82.17 26.415 82.43 26.675 ;
        RECT 82.17 25.655 82.43 25.915 ;
        RECT 82.17 24.895 82.43 25.155 ;
        RECT 82.17 24.135 82.43 24.395 ;
        RECT 82.17 23.375 82.43 23.635 ;
        RECT 82.93 30.215 83.19 30.475 ;
        RECT 82.93 29.455 83.19 29.715 ;
        RECT 82.93 28.695 83.19 28.955 ;
        RECT 82.93 27.935 83.19 28.195 ;
        RECT 82.93 27.175 83.19 27.435 ;
        RECT 82.93 26.415 83.19 26.675 ;
        RECT 82.93 25.655 83.19 25.915 ;
        RECT 82.93 24.895 83.19 25.155 ;
        RECT 82.93 24.135 83.19 24.395 ;
        RECT 82.93 23.375 83.19 23.635 ;
        RECT 83.69 30.215 83.95 30.475 ;
        RECT 83.69 29.455 83.95 29.715 ;
        RECT 83.69 28.695 83.95 28.955 ;
        RECT 83.69 27.935 83.95 28.195 ;
        RECT 83.69 27.175 83.95 27.435 ;
        RECT 83.69 26.415 83.95 26.675 ;
        RECT 83.69 25.655 83.95 25.915 ;
        RECT 83.69 24.895 83.95 25.155 ;
        RECT 83.69 24.135 83.95 24.395 ;
        RECT 83.69 23.375 83.95 23.635 ;
        RECT 84.45 30.215 84.71 30.475 ;
        RECT 84.45 29.455 84.71 29.715 ;
        RECT 84.45 28.695 84.71 28.955 ;
        RECT 84.45 27.935 84.71 28.195 ;
        RECT 84.45 27.175 84.71 27.435 ;
        RECT 84.45 26.415 84.71 26.675 ;
        RECT 84.45 25.655 84.71 25.915 ;
        RECT 84.45 24.895 84.71 25.155 ;
        RECT 84.45 24.135 84.71 24.395 ;
        RECT 84.45 23.375 84.71 23.635 ;
        RECT 85.21 30.215 85.47 30.475 ;
        RECT 85.21 29.455 85.47 29.715 ;
        RECT 85.21 28.695 85.47 28.955 ;
        RECT 85.21 27.935 85.47 28.195 ;
        RECT 85.21 27.175 85.47 27.435 ;
        RECT 85.21 26.415 85.47 26.675 ;
        RECT 85.21 25.655 85.47 25.915 ;
        RECT 85.21 24.895 85.47 25.155 ;
        RECT 85.21 24.135 85.47 24.395 ;
        RECT 85.21 23.375 85.47 23.635 ;
        RECT 85.97 30.215 86.23 30.475 ;
        RECT 85.97 29.455 86.23 29.715 ;
        RECT 85.97 28.695 86.23 28.955 ;
        RECT 85.97 27.935 86.23 28.195 ;
        RECT 85.97 27.175 86.23 27.435 ;
        RECT 85.97 26.415 86.23 26.675 ;
        RECT 85.97 25.655 86.23 25.915 ;
        RECT 85.97 24.895 86.23 25.155 ;
        RECT 85.97 24.135 86.23 24.395 ;
        RECT 85.97 23.375 86.23 23.635 ;
        RECT 86.73 30.215 86.99 30.475 ;
        RECT 86.73 29.455 86.99 29.715 ;
        RECT 86.73 28.695 86.99 28.955 ;
        RECT 86.73 27.935 86.99 28.195 ;
        RECT 86.73 27.175 86.99 27.435 ;
        RECT 86.73 26.415 86.99 26.675 ;
        RECT 86.73 25.655 86.99 25.915 ;
        RECT 86.73 24.895 86.99 25.155 ;
        RECT 86.73 24.135 86.99 24.395 ;
        RECT 86.73 23.375 86.99 23.635 ;
        RECT 87.49 30.215 87.75 30.475 ;
        RECT 87.49 29.455 87.75 29.715 ;
        RECT 87.49 28.695 87.75 28.955 ;
        RECT 87.49 27.935 87.75 28.195 ;
        RECT 87.49 27.175 87.75 27.435 ;
        RECT 87.49 26.415 87.75 26.675 ;
        RECT 87.49 25.655 87.75 25.915 ;
        RECT 87.49 24.895 87.75 25.155 ;
        RECT 87.49 24.135 87.75 24.395 ;
        RECT 87.49 23.375 87.75 23.635 ;
        RECT 88.25 30.215 88.51 30.475 ;
        RECT 88.25 29.455 88.51 29.715 ;
        RECT 88.25 28.695 88.51 28.955 ;
        RECT 88.25 27.935 88.51 28.195 ;
        RECT 88.25 27.175 88.51 27.435 ;
        RECT 88.25 26.415 88.51 26.675 ;
        RECT 88.25 25.655 88.51 25.915 ;
        RECT 88.25 24.895 88.51 25.155 ;
        RECT 88.25 24.135 88.51 24.395 ;
        RECT 88.25 23.375 88.51 23.635 ;
        RECT 89.01 30.215 89.27 30.475 ;
        RECT 89.01 29.455 89.27 29.715 ;
        RECT 89.01 28.695 89.27 28.955 ;
        RECT 89.01 27.935 89.27 28.195 ;
        RECT 89.01 27.175 89.27 27.435 ;
        RECT 89.01 26.415 89.27 26.675 ;
        RECT 89.01 25.655 89.27 25.915 ;
        RECT 89.01 24.895 89.27 25.155 ;
        RECT 89.01 24.135 89.27 24.395 ;
        RECT 89.01 23.375 89.27 23.635 ;
        RECT 89.77 30.215 90.03 30.475 ;
        RECT 89.77 29.455 90.03 29.715 ;
        RECT 89.77 28.695 90.03 28.955 ;
        RECT 89.77 27.935 90.03 28.195 ;
        RECT 89.77 27.175 90.03 27.435 ;
        RECT 89.77 26.415 90.03 26.675 ;
        RECT 89.77 25.655 90.03 25.915 ;
        RECT 89.77 24.895 90.03 25.155 ;
        RECT 89.77 24.135 90.03 24.395 ;
        RECT 89.77 23.375 90.03 23.635 ;
        RECT 90.53 30.215 90.79 30.475 ;
        RECT 90.53 29.455 90.79 29.715 ;
        RECT 90.53 28.695 90.79 28.955 ;
        RECT 90.53 27.935 90.79 28.195 ;
        RECT 90.53 27.175 90.79 27.435 ;
        RECT 90.53 26.415 90.79 26.675 ;
        RECT 90.53 25.655 90.79 25.915 ;
        RECT 90.53 24.895 90.79 25.155 ;
        RECT 90.53 24.135 90.79 24.395 ;
        RECT 90.53 23.375 90.79 23.635 ;
        RECT 91.29 30.215 91.55 30.475 ;
        RECT 91.29 29.455 91.55 29.715 ;
        RECT 91.29 28.695 91.55 28.955 ;
        RECT 91.29 27.935 91.55 28.195 ;
        RECT 91.29 27.175 91.55 27.435 ;
        RECT 91.29 26.415 91.55 26.675 ;
        RECT 91.29 25.655 91.55 25.915 ;
        RECT 91.29 24.895 91.55 25.155 ;
        RECT 91.29 24.135 91.55 24.395 ;
        RECT 91.29 23.375 91.55 23.635 ;
        RECT 92.05 30.215 92.31 30.475 ;
        RECT 92.05 29.455 92.31 29.715 ;
        RECT 92.05 28.695 92.31 28.955 ;
        RECT 92.05 27.935 92.31 28.195 ;
        RECT 92.05 27.175 92.31 27.435 ;
        RECT 92.05 26.415 92.31 26.675 ;
        RECT 92.05 25.655 92.31 25.915 ;
        RECT 92.05 24.895 92.31 25.155 ;
        RECT 92.05 24.135 92.31 24.395 ;
        RECT 92.05 23.375 92.31 23.635 ;
        RECT 92.81 30.215 93.07 30.475 ;
        RECT 92.81 29.455 93.07 29.715 ;
        RECT 92.81 28.695 93.07 28.955 ;
        RECT 92.81 27.935 93.07 28.195 ;
        RECT 92.81 27.175 93.07 27.435 ;
        RECT 92.81 26.415 93.07 26.675 ;
        RECT 92.81 25.655 93.07 25.915 ;
        RECT 92.81 24.895 93.07 25.155 ;
        RECT 92.81 24.135 93.07 24.395 ;
        RECT 92.81 23.375 93.07 23.635 ;
        RECT 93.57 30.215 93.83 30.475 ;
        RECT 93.57 29.455 93.83 29.715 ;
        RECT 93.57 28.695 93.83 28.955 ;
        RECT 93.57 27.935 93.83 28.195 ;
        RECT 93.57 27.175 93.83 27.435 ;
        RECT 93.57 26.415 93.83 26.675 ;
        RECT 93.57 25.655 93.83 25.915 ;
        RECT 93.57 24.895 93.83 25.155 ;
        RECT 93.57 24.135 93.83 24.395 ;
        RECT 93.57 23.375 93.83 23.635 ;
        RECT 94.33 30.215 94.59 30.475 ;
        RECT 94.33 29.455 94.59 29.715 ;
        RECT 94.33 28.695 94.59 28.955 ;
        RECT 94.33 27.935 94.59 28.195 ;
        RECT 94.33 27.175 94.59 27.435 ;
        RECT 94.33 26.415 94.59 26.675 ;
        RECT 94.33 25.655 94.59 25.915 ;
        RECT 94.33 24.895 94.59 25.155 ;
        RECT 94.33 24.135 94.59 24.395 ;
        RECT 94.33 23.375 94.59 23.635 ;
        RECT 95.09 30.215 95.35 30.475 ;
        RECT 95.09 29.455 95.35 29.715 ;
        RECT 95.09 28.695 95.35 28.955 ;
        RECT 95.09 27.935 95.35 28.195 ;
        RECT 95.09 27.175 95.35 27.435 ;
        RECT 95.09 26.415 95.35 26.675 ;
        RECT 95.09 25.655 95.35 25.915 ;
        RECT 95.09 24.895 95.35 25.155 ;
        RECT 95.09 24.135 95.35 24.395 ;
        RECT 95.09 23.375 95.35 23.635 ;
        RECT 4.65 30.215 4.91 30.475 ;
        RECT 4.65 29.455 4.91 29.715 ;
        RECT 4.65 28.695 4.91 28.955 ;
        RECT 4.65 27.935 4.91 28.195 ;
        RECT 4.65 27.175 4.91 27.435 ;
        RECT 4.65 26.415 4.91 26.675 ;
        RECT 4.65 25.655 4.91 25.915 ;
        RECT 4.65 24.895 4.91 25.155 ;
        RECT 4.65 24.135 4.91 24.395 ;
        RECT 4.65 23.375 4.91 23.635 ;
        RECT 5.41 30.215 5.67 30.475 ;
        RECT 5.41 29.455 5.67 29.715 ;
        RECT 5.41 28.695 5.67 28.955 ;
        RECT 5.41 27.935 5.67 28.195 ;
        RECT 5.41 27.175 5.67 27.435 ;
        RECT 5.41 26.415 5.67 26.675 ;
        RECT 5.41 25.655 5.67 25.915 ;
        RECT 5.41 24.895 5.67 25.155 ;
        RECT 5.41 24.135 5.67 24.395 ;
        RECT 5.41 23.375 5.67 23.635 ;
        RECT 6.17 30.215 6.43 30.475 ;
        RECT 6.17 29.455 6.43 29.715 ;
        RECT 6.17 28.695 6.43 28.955 ;
        RECT 6.17 27.935 6.43 28.195 ;
        RECT 6.17 27.175 6.43 27.435 ;
        RECT 6.17 26.415 6.43 26.675 ;
        RECT 6.17 25.655 6.43 25.915 ;
        RECT 6.17 24.895 6.43 25.155 ;
        RECT 6.17 24.135 6.43 24.395 ;
        RECT 6.17 23.375 6.43 23.635 ;
        RECT 6.93 30.215 7.19 30.475 ;
        RECT 6.93 29.455 7.19 29.715 ;
        RECT 6.93 28.695 7.19 28.955 ;
        RECT 6.93 27.935 7.19 28.195 ;
        RECT 6.93 27.175 7.19 27.435 ;
        RECT 6.93 26.415 7.19 26.675 ;
        RECT 6.93 25.655 7.19 25.915 ;
        RECT 6.93 24.895 7.19 25.155 ;
        RECT 6.93 24.135 7.19 24.395 ;
        RECT 6.93 23.375 7.19 23.635 ;
        RECT 7.69 30.215 7.95 30.475 ;
        RECT 7.69 29.455 7.95 29.715 ;
        RECT 7.69 28.695 7.95 28.955 ;
        RECT 7.69 27.935 7.95 28.195 ;
        RECT 7.69 27.175 7.95 27.435 ;
        RECT 7.69 26.415 7.95 26.675 ;
        RECT 7.69 25.655 7.95 25.915 ;
        RECT 7.69 24.895 7.95 25.155 ;
        RECT 7.69 24.135 7.95 24.395 ;
        RECT 7.69 23.375 7.95 23.635 ;
        RECT 8.45 30.215 8.71 30.475 ;
        RECT 8.45 29.455 8.71 29.715 ;
        RECT 8.45 28.695 8.71 28.955 ;
        RECT 8.45 27.935 8.71 28.195 ;
        RECT 8.45 27.175 8.71 27.435 ;
        RECT 8.45 26.415 8.71 26.675 ;
        RECT 8.45 25.655 8.71 25.915 ;
        RECT 8.45 24.895 8.71 25.155 ;
        RECT 8.45 24.135 8.71 24.395 ;
        RECT 8.45 23.375 8.71 23.635 ;
        RECT 9.21 30.215 9.47 30.475 ;
        RECT 9.21 29.455 9.47 29.715 ;
        RECT 9.21 28.695 9.47 28.955 ;
        RECT 9.21 27.935 9.47 28.195 ;
        RECT 9.21 27.175 9.47 27.435 ;
        RECT 9.21 26.415 9.47 26.675 ;
        RECT 9.21 25.655 9.47 25.915 ;
        RECT 9.21 24.895 9.47 25.155 ;
        RECT 9.21 24.135 9.47 24.395 ;
        RECT 9.21 23.375 9.47 23.635 ;
        RECT 9.97 30.215 10.23 30.475 ;
        RECT 9.97 29.455 10.23 29.715 ;
        RECT 9.97 28.695 10.23 28.955 ;
        RECT 9.97 27.935 10.23 28.195 ;
        RECT 9.97 27.175 10.23 27.435 ;
        RECT 9.97 26.415 10.23 26.675 ;
        RECT 9.97 25.655 10.23 25.915 ;
        RECT 9.97 24.895 10.23 25.155 ;
        RECT 9.97 24.135 10.23 24.395 ;
        RECT 9.97 23.375 10.23 23.635 ;
        RECT 10.73 30.215 10.99 30.475 ;
        RECT 10.73 29.455 10.99 29.715 ;
        RECT 10.73 28.695 10.99 28.955 ;
        RECT 10.73 27.935 10.99 28.195 ;
        RECT 10.73 27.175 10.99 27.435 ;
        RECT 10.73 26.415 10.99 26.675 ;
        RECT 10.73 25.655 10.99 25.915 ;
        RECT 10.73 24.895 10.99 25.155 ;
        RECT 10.73 24.135 10.99 24.395 ;
        RECT 10.73 23.375 10.99 23.635 ;
        RECT 11.49 30.215 11.75 30.475 ;
        RECT 11.49 29.455 11.75 29.715 ;
        RECT 11.49 28.695 11.75 28.955 ;
        RECT 11.49 27.935 11.75 28.195 ;
        RECT 11.49 27.175 11.75 27.435 ;
        RECT 11.49 26.415 11.75 26.675 ;
        RECT 11.49 25.655 11.75 25.915 ;
        RECT 11.49 24.895 11.75 25.155 ;
        RECT 11.49 24.135 11.75 24.395 ;
        RECT 11.49 23.375 11.75 23.635 ;
        RECT 12.25 30.215 12.51 30.475 ;
        RECT 12.25 29.455 12.51 29.715 ;
        RECT 12.25 28.695 12.51 28.955 ;
        RECT 12.25 27.935 12.51 28.195 ;
        RECT 12.25 27.175 12.51 27.435 ;
        RECT 12.25 26.415 12.51 26.675 ;
        RECT 12.25 25.655 12.51 25.915 ;
        RECT 12.25 24.895 12.51 25.155 ;
        RECT 12.25 24.135 12.51 24.395 ;
        RECT 12.25 23.375 12.51 23.635 ;
        RECT 13.01 30.215 13.27 30.475 ;
        RECT 13.01 29.455 13.27 29.715 ;
        RECT 13.01 28.695 13.27 28.955 ;
        RECT 13.01 27.935 13.27 28.195 ;
        RECT 13.01 27.175 13.27 27.435 ;
        RECT 13.01 26.415 13.27 26.675 ;
        RECT 13.01 25.655 13.27 25.915 ;
        RECT 13.01 24.895 13.27 25.155 ;
        RECT 13.01 24.135 13.27 24.395 ;
        RECT 13.01 23.375 13.27 23.635 ;
        RECT 13.77 30.215 14.03 30.475 ;
        RECT 13.77 29.455 14.03 29.715 ;
        RECT 13.77 28.695 14.03 28.955 ;
        RECT 13.77 27.935 14.03 28.195 ;
        RECT 13.77 27.175 14.03 27.435 ;
        RECT 13.77 26.415 14.03 26.675 ;
        RECT 13.77 25.655 14.03 25.915 ;
        RECT 13.77 24.895 14.03 25.155 ;
        RECT 13.77 24.135 14.03 24.395 ;
        RECT 13.77 23.375 14.03 23.635 ;
        RECT 14.53 30.215 14.79 30.475 ;
        RECT 14.53 29.455 14.79 29.715 ;
        RECT 14.53 28.695 14.79 28.955 ;
        RECT 14.53 27.935 14.79 28.195 ;
        RECT 14.53 27.175 14.79 27.435 ;
        RECT 14.53 26.415 14.79 26.675 ;
        RECT 14.53 25.655 14.79 25.915 ;
        RECT 14.53 24.895 14.79 25.155 ;
        RECT 14.53 24.135 14.79 24.395 ;
        RECT 14.53 23.375 14.79 23.635 ;
        RECT 15.29 30.215 15.55 30.475 ;
        RECT 15.29 29.455 15.55 29.715 ;
        RECT 15.29 28.695 15.55 28.955 ;
        RECT 15.29 27.935 15.55 28.195 ;
        RECT 15.29 27.175 15.55 27.435 ;
        RECT 15.29 26.415 15.55 26.675 ;
        RECT 15.29 25.655 15.55 25.915 ;
        RECT 15.29 24.895 15.55 25.155 ;
        RECT 15.29 24.135 15.55 24.395 ;
        RECT 15.29 23.375 15.55 23.635 ;
        RECT 16.05 30.215 16.31 30.475 ;
        RECT 16.05 29.455 16.31 29.715 ;
        RECT 16.05 28.695 16.31 28.955 ;
        RECT 16.05 27.935 16.31 28.195 ;
        RECT 16.05 27.175 16.31 27.435 ;
        RECT 16.05 26.415 16.31 26.675 ;
        RECT 16.05 25.655 16.31 25.915 ;
        RECT 16.05 24.895 16.31 25.155 ;
        RECT 16.05 24.135 16.31 24.395 ;
        RECT 16.05 23.375 16.31 23.635 ;
        RECT 16.81 30.215 17.07 30.475 ;
        RECT 16.81 29.455 17.07 29.715 ;
        RECT 16.81 28.695 17.07 28.955 ;
        RECT 16.81 27.935 17.07 28.195 ;
        RECT 16.81 27.175 17.07 27.435 ;
        RECT 16.81 26.415 17.07 26.675 ;
        RECT 16.81 25.655 17.07 25.915 ;
        RECT 16.81 24.895 17.07 25.155 ;
        RECT 16.81 24.135 17.07 24.395 ;
        RECT 16.81 23.375 17.07 23.635 ;
        RECT 17.57 30.215 17.83 30.475 ;
        RECT 17.57 29.455 17.83 29.715 ;
        RECT 17.57 28.695 17.83 28.955 ;
        RECT 17.57 27.935 17.83 28.195 ;
        RECT 17.57 27.175 17.83 27.435 ;
        RECT 17.57 26.415 17.83 26.675 ;
        RECT 17.57 25.655 17.83 25.915 ;
        RECT 17.57 24.895 17.83 25.155 ;
        RECT 17.57 24.135 17.83 24.395 ;
        RECT 17.57 23.375 17.83 23.635 ;
        RECT 18.33 30.215 18.59 30.475 ;
        RECT 18.33 29.455 18.59 29.715 ;
        RECT 18.33 28.695 18.59 28.955 ;
        RECT 18.33 27.935 18.59 28.195 ;
        RECT 18.33 27.175 18.59 27.435 ;
        RECT 18.33 26.415 18.59 26.675 ;
        RECT 18.33 25.655 18.59 25.915 ;
        RECT 18.33 24.895 18.59 25.155 ;
        RECT 18.33 24.135 18.59 24.395 ;
        RECT 18.33 23.375 18.59 23.635 ;
        RECT 19.09 30.215 19.35 30.475 ;
        RECT 19.09 29.455 19.35 29.715 ;
        RECT 19.09 28.695 19.35 28.955 ;
        RECT 19.09 27.935 19.35 28.195 ;
        RECT 19.09 27.175 19.35 27.435 ;
        RECT 19.09 26.415 19.35 26.675 ;
        RECT 19.09 25.655 19.35 25.915 ;
        RECT 19.09 24.895 19.35 25.155 ;
        RECT 19.09 24.135 19.35 24.395 ;
        RECT 19.09 23.375 19.35 23.635 ;
        RECT 19.85 30.215 20.11 30.475 ;
        RECT 19.85 29.455 20.11 29.715 ;
        RECT 19.85 28.695 20.11 28.955 ;
        RECT 19.85 27.935 20.11 28.195 ;
        RECT 19.85 27.175 20.11 27.435 ;
        RECT 19.85 26.415 20.11 26.675 ;
        RECT 19.85 25.655 20.11 25.915 ;
        RECT 19.85 24.895 20.11 25.155 ;
        RECT 19.85 24.135 20.11 24.395 ;
        RECT 19.85 23.375 20.11 23.635 ;
        RECT 20.61 30.215 20.87 30.475 ;
        RECT 20.61 29.455 20.87 29.715 ;
        RECT 20.61 28.695 20.87 28.955 ;
        RECT 20.61 27.935 20.87 28.195 ;
        RECT 20.61 27.175 20.87 27.435 ;
        RECT 20.61 26.415 20.87 26.675 ;
        RECT 20.61 25.655 20.87 25.915 ;
        RECT 20.61 24.895 20.87 25.155 ;
        RECT 20.61 24.135 20.87 24.395 ;
        RECT 20.61 23.375 20.87 23.635 ;
        RECT 21.37 30.215 21.63 30.475 ;
        RECT 21.37 29.455 21.63 29.715 ;
        RECT 21.37 28.695 21.63 28.955 ;
        RECT 21.37 27.935 21.63 28.195 ;
        RECT 21.37 27.175 21.63 27.435 ;
        RECT 21.37 26.415 21.63 26.675 ;
        RECT 21.37 25.655 21.63 25.915 ;
        RECT 21.37 24.895 21.63 25.155 ;
        RECT 21.37 24.135 21.63 24.395 ;
        RECT 21.37 23.375 21.63 23.635 ;
        RECT 22.13 30.215 22.39 30.475 ;
        RECT 22.13 29.455 22.39 29.715 ;
        RECT 22.13 28.695 22.39 28.955 ;
        RECT 22.13 27.935 22.39 28.195 ;
        RECT 22.13 27.175 22.39 27.435 ;
        RECT 22.13 26.415 22.39 26.675 ;
        RECT 22.13 25.655 22.39 25.915 ;
        RECT 22.13 24.895 22.39 25.155 ;
        RECT 22.13 24.135 22.39 24.395 ;
        RECT 22.13 23.375 22.39 23.635 ;
        RECT 22.89 30.215 23.15 30.475 ;
        RECT 22.89 29.455 23.15 29.715 ;
        RECT 22.89 28.695 23.15 28.955 ;
        RECT 22.89 27.935 23.15 28.195 ;
        RECT 22.89 27.175 23.15 27.435 ;
        RECT 22.89 26.415 23.15 26.675 ;
        RECT 22.89 25.655 23.15 25.915 ;
        RECT 22.89 24.895 23.15 25.155 ;
        RECT 22.89 24.135 23.15 24.395 ;
        RECT 22.89 23.375 23.15 23.635 ;
        RECT 23.65 30.215 23.91 30.475 ;
        RECT 23.65 29.455 23.91 29.715 ;
        RECT 23.65 28.695 23.91 28.955 ;
        RECT 23.65 27.935 23.91 28.195 ;
        RECT 23.65 27.175 23.91 27.435 ;
        RECT 23.65 26.415 23.91 26.675 ;
        RECT 23.65 25.655 23.91 25.915 ;
        RECT 23.65 24.895 23.91 25.155 ;
        RECT 23.65 24.135 23.91 24.395 ;
        RECT 23.65 23.375 23.91 23.635 ;
        RECT 24.41 30.215 24.67 30.475 ;
        RECT 24.41 29.455 24.67 29.715 ;
        RECT 24.41 28.695 24.67 28.955 ;
        RECT 24.41 27.935 24.67 28.195 ;
        RECT 24.41 27.175 24.67 27.435 ;
        RECT 24.41 26.415 24.67 26.675 ;
        RECT 24.41 25.655 24.67 25.915 ;
        RECT 24.41 24.895 24.67 25.155 ;
        RECT 24.41 24.135 24.67 24.395 ;
        RECT 24.41 23.375 24.67 23.635 ;
        RECT 25.17 30.215 25.43 30.475 ;
        RECT 25.17 29.455 25.43 29.715 ;
        RECT 25.17 28.695 25.43 28.955 ;
        RECT 25.17 27.935 25.43 28.195 ;
        RECT 25.17 27.175 25.43 27.435 ;
        RECT 25.17 26.415 25.43 26.675 ;
        RECT 25.17 25.655 25.43 25.915 ;
        RECT 25.17 24.895 25.43 25.155 ;
        RECT 25.17 24.135 25.43 24.395 ;
        RECT 25.17 23.375 25.43 23.635 ;
        RECT 25.93 30.215 26.19 30.475 ;
        RECT 25.93 29.455 26.19 29.715 ;
        RECT 25.93 28.695 26.19 28.955 ;
        RECT 25.93 27.935 26.19 28.195 ;
        RECT 25.93 27.175 26.19 27.435 ;
        RECT 25.93 26.415 26.19 26.675 ;
        RECT 25.93 25.655 26.19 25.915 ;
        RECT 25.93 24.895 26.19 25.155 ;
        RECT 25.93 24.135 26.19 24.395 ;
        RECT 25.93 23.375 26.19 23.635 ;
        RECT 26.69 30.215 26.95 30.475 ;
        RECT 26.69 29.455 26.95 29.715 ;
        RECT 26.69 28.695 26.95 28.955 ;
        RECT 26.69 27.935 26.95 28.195 ;
        RECT 26.69 27.175 26.95 27.435 ;
        RECT 26.69 26.415 26.95 26.675 ;
        RECT 26.69 25.655 26.95 25.915 ;
        RECT 26.69 24.895 26.95 25.155 ;
        RECT 26.69 24.135 26.95 24.395 ;
        RECT 26.69 23.375 26.95 23.635 ;
        RECT 27.45 30.215 27.71 30.475 ;
        RECT 27.45 29.455 27.71 29.715 ;
        RECT 27.45 28.695 27.71 28.955 ;
        RECT 27.45 27.935 27.71 28.195 ;
        RECT 27.45 27.175 27.71 27.435 ;
        RECT 27.45 26.415 27.71 26.675 ;
        RECT 27.45 25.655 27.71 25.915 ;
        RECT 27.45 24.895 27.71 25.155 ;
        RECT 27.45 24.135 27.71 24.395 ;
        RECT 27.45 23.375 27.71 23.635 ;
        RECT 28.21 30.215 28.47 30.475 ;
        RECT 28.21 29.455 28.47 29.715 ;
        RECT 28.21 28.695 28.47 28.955 ;
        RECT 28.21 27.935 28.47 28.195 ;
        RECT 28.21 27.175 28.47 27.435 ;
        RECT 28.21 26.415 28.47 26.675 ;
        RECT 28.21 25.655 28.47 25.915 ;
        RECT 28.21 24.895 28.47 25.155 ;
        RECT 28.21 24.135 28.47 24.395 ;
        RECT 28.21 23.375 28.47 23.635 ;
        RECT 28.97 30.215 29.23 30.475 ;
        RECT 28.97 29.455 29.23 29.715 ;
        RECT 28.97 28.695 29.23 28.955 ;
        RECT 28.97 27.935 29.23 28.195 ;
        RECT 28.97 27.175 29.23 27.435 ;
        RECT 28.97 26.415 29.23 26.675 ;
        RECT 28.97 25.655 29.23 25.915 ;
        RECT 28.97 24.895 29.23 25.155 ;
        RECT 28.97 24.135 29.23 24.395 ;
        RECT 28.97 23.375 29.23 23.635 ;
        RECT 29.73 30.215 29.99 30.475 ;
        RECT 29.73 29.455 29.99 29.715 ;
        RECT 29.73 28.695 29.99 28.955 ;
        RECT 29.73 27.935 29.99 28.195 ;
        RECT 29.73 27.175 29.99 27.435 ;
        RECT 29.73 26.415 29.99 26.675 ;
        RECT 29.73 25.655 29.99 25.915 ;
        RECT 29.73 24.895 29.99 25.155 ;
        RECT 29.73 24.135 29.99 24.395 ;
        RECT 29.73 23.375 29.99 23.635 ;
        RECT 30.49 30.215 30.75 30.475 ;
        RECT 30.49 29.455 30.75 29.715 ;
        RECT 30.49 28.695 30.75 28.955 ;
        RECT 30.49 27.935 30.75 28.195 ;
        RECT 30.49 27.175 30.75 27.435 ;
        RECT 30.49 26.415 30.75 26.675 ;
        RECT 30.49 25.655 30.75 25.915 ;
        RECT 30.49 24.895 30.75 25.155 ;
        RECT 30.49 24.135 30.75 24.395 ;
        RECT 30.49 23.375 30.75 23.635 ;
        RECT 31.25 30.215 31.51 30.475 ;
        RECT 31.25 29.455 31.51 29.715 ;
        RECT 31.25 28.695 31.51 28.955 ;
        RECT 31.25 27.935 31.51 28.195 ;
        RECT 31.25 27.175 31.51 27.435 ;
        RECT 31.25 26.415 31.51 26.675 ;
        RECT 31.25 25.655 31.51 25.915 ;
        RECT 31.25 24.895 31.51 25.155 ;
        RECT 31.25 24.135 31.51 24.395 ;
        RECT 31.25 23.375 31.51 23.635 ;
        RECT 32.01 30.215 32.27 30.475 ;
        RECT 32.01 29.455 32.27 29.715 ;
        RECT 32.01 28.695 32.27 28.955 ;
        RECT 32.01 27.935 32.27 28.195 ;
        RECT 32.01 27.175 32.27 27.435 ;
        RECT 32.01 26.415 32.27 26.675 ;
        RECT 32.01 25.655 32.27 25.915 ;
        RECT 32.01 24.895 32.27 25.155 ;
        RECT 32.01 24.135 32.27 24.395 ;
        RECT 32.01 23.375 32.27 23.635 ;
        RECT 32.77 30.215 33.03 30.475 ;
        RECT 32.77 29.455 33.03 29.715 ;
        RECT 32.77 28.695 33.03 28.955 ;
        RECT 32.77 27.935 33.03 28.195 ;
        RECT 32.77 27.175 33.03 27.435 ;
        RECT 32.77 26.415 33.03 26.675 ;
        RECT 32.77 25.655 33.03 25.915 ;
        RECT 32.77 24.895 33.03 25.155 ;
        RECT 32.77 24.135 33.03 24.395 ;
        RECT 32.77 23.375 33.03 23.635 ;
        RECT 33.53 30.215 33.79 30.475 ;
        RECT 33.53 29.455 33.79 29.715 ;
        RECT 33.53 28.695 33.79 28.955 ;
        RECT 33.53 27.935 33.79 28.195 ;
        RECT 33.53 27.175 33.79 27.435 ;
        RECT 33.53 26.415 33.79 26.675 ;
        RECT 33.53 25.655 33.79 25.915 ;
        RECT 33.53 24.895 33.79 25.155 ;
        RECT 33.53 24.135 33.79 24.395 ;
        RECT 33.53 23.375 33.79 23.635 ;
        RECT 34.29 30.215 34.55 30.475 ;
        RECT 34.29 29.455 34.55 29.715 ;
        RECT 34.29 28.695 34.55 28.955 ;
        RECT 34.29 27.935 34.55 28.195 ;
        RECT 34.29 27.175 34.55 27.435 ;
        RECT 34.29 26.415 34.55 26.675 ;
        RECT 34.29 25.655 34.55 25.915 ;
        RECT 34.29 24.895 34.55 25.155 ;
        RECT 34.29 24.135 34.55 24.395 ;
        RECT 34.29 23.375 34.55 23.635 ;
        RECT 35.05 30.215 35.31 30.475 ;
        RECT 35.05 29.455 35.31 29.715 ;
        RECT 35.05 28.695 35.31 28.955 ;
        RECT 35.05 27.935 35.31 28.195 ;
        RECT 35.05 27.175 35.31 27.435 ;
        RECT 35.05 26.415 35.31 26.675 ;
        RECT 35.05 25.655 35.31 25.915 ;
        RECT 35.05 24.895 35.31 25.155 ;
        RECT 35.05 24.135 35.31 24.395 ;
        RECT 35.05 23.375 35.31 23.635 ;
        RECT 35.81 30.215 36.07 30.475 ;
        RECT 35.81 29.455 36.07 29.715 ;
        RECT 35.81 28.695 36.07 28.955 ;
        RECT 35.81 27.935 36.07 28.195 ;
        RECT 35.81 27.175 36.07 27.435 ;
        RECT 35.81 26.415 36.07 26.675 ;
        RECT 35.81 25.655 36.07 25.915 ;
        RECT 35.81 24.895 36.07 25.155 ;
        RECT 35.81 24.135 36.07 24.395 ;
        RECT 35.81 23.375 36.07 23.635 ;
        RECT 36.57 30.215 36.83 30.475 ;
        RECT 36.57 29.455 36.83 29.715 ;
        RECT 36.57 28.695 36.83 28.955 ;
        RECT 36.57 27.935 36.83 28.195 ;
        RECT 36.57 27.175 36.83 27.435 ;
        RECT 36.57 26.415 36.83 26.675 ;
        RECT 36.57 25.655 36.83 25.915 ;
        RECT 36.57 24.895 36.83 25.155 ;
        RECT 36.57 24.135 36.83 24.395 ;
        RECT 36.57 23.375 36.83 23.635 ;
        RECT 37.33 30.215 37.59 30.475 ;
        RECT 37.33 29.455 37.59 29.715 ;
        RECT 37.33 28.695 37.59 28.955 ;
        RECT 37.33 27.935 37.59 28.195 ;
        RECT 37.33 27.175 37.59 27.435 ;
        RECT 37.33 26.415 37.59 26.675 ;
        RECT 37.33 25.655 37.59 25.915 ;
        RECT 37.33 24.895 37.59 25.155 ;
        RECT 37.33 24.135 37.59 24.395 ;
        RECT 37.33 23.375 37.59 23.635 ;
        RECT 38.09 30.215 38.35 30.475 ;
        RECT 38.09 29.455 38.35 29.715 ;
        RECT 38.09 28.695 38.35 28.955 ;
        RECT 38.09 27.935 38.35 28.195 ;
        RECT 38.09 27.175 38.35 27.435 ;
        RECT 38.09 26.415 38.35 26.675 ;
        RECT 38.09 25.655 38.35 25.915 ;
        RECT 38.09 24.895 38.35 25.155 ;
        RECT 38.09 24.135 38.35 24.395 ;
        RECT 38.09 23.375 38.35 23.635 ;
        RECT 38.85 30.215 39.11 30.475 ;
        RECT 38.85 29.455 39.11 29.715 ;
        RECT 38.85 28.695 39.11 28.955 ;
        RECT 38.85 27.935 39.11 28.195 ;
        RECT 38.85 27.175 39.11 27.435 ;
        RECT 38.85 26.415 39.11 26.675 ;
        RECT 38.85 25.655 39.11 25.915 ;
        RECT 38.85 24.895 39.11 25.155 ;
        RECT 38.85 24.135 39.11 24.395 ;
        RECT 38.85 23.375 39.11 23.635 ;
        RECT 39.61 30.215 39.87 30.475 ;
        RECT 39.61 29.455 39.87 29.715 ;
        RECT 39.61 28.695 39.87 28.955 ;
        RECT 39.61 27.935 39.87 28.195 ;
        RECT 39.61 27.175 39.87 27.435 ;
        RECT 39.61 26.415 39.87 26.675 ;
        RECT 39.61 25.655 39.87 25.915 ;
        RECT 39.61 24.895 39.87 25.155 ;
        RECT 39.61 24.135 39.87 24.395 ;
        RECT 39.61 23.375 39.87 23.635 ;
        RECT 40.37 30.215 40.63 30.475 ;
        RECT 40.37 29.455 40.63 29.715 ;
        RECT 40.37 28.695 40.63 28.955 ;
        RECT 40.37 27.935 40.63 28.195 ;
        RECT 40.37 27.175 40.63 27.435 ;
        RECT 40.37 26.415 40.63 26.675 ;
        RECT 40.37 25.655 40.63 25.915 ;
        RECT 40.37 24.895 40.63 25.155 ;
        RECT 40.37 24.135 40.63 24.395 ;
        RECT 40.37 23.375 40.63 23.635 ;
        RECT 41.13 30.215 41.39 30.475 ;
        RECT 41.13 29.455 41.39 29.715 ;
        RECT 41.13 28.695 41.39 28.955 ;
        RECT 41.13 27.935 41.39 28.195 ;
        RECT 41.13 27.175 41.39 27.435 ;
        RECT 41.13 26.415 41.39 26.675 ;
        RECT 41.13 25.655 41.39 25.915 ;
        RECT 41.13 24.895 41.39 25.155 ;
        RECT 41.13 24.135 41.39 24.395 ;
        RECT 41.13 23.375 41.39 23.635 ;
        RECT 41.89 30.215 42.15 30.475 ;
        RECT 41.89 29.455 42.15 29.715 ;
        RECT 41.89 28.695 42.15 28.955 ;
        RECT 41.89 27.935 42.15 28.195 ;
        RECT 41.89 27.175 42.15 27.435 ;
        RECT 41.89 26.415 42.15 26.675 ;
        RECT 41.89 25.655 42.15 25.915 ;
        RECT 41.89 24.895 42.15 25.155 ;
        RECT 41.89 24.135 42.15 24.395 ;
        RECT 41.89 23.375 42.15 23.635 ;
        RECT 42.65 30.215 42.91 30.475 ;
        RECT 42.65 29.455 42.91 29.715 ;
        RECT 42.65 28.695 42.91 28.955 ;
        RECT 42.65 27.935 42.91 28.195 ;
        RECT 42.65 27.175 42.91 27.435 ;
        RECT 42.65 26.415 42.91 26.675 ;
        RECT 42.65 25.655 42.91 25.915 ;
        RECT 42.65 24.895 42.91 25.155 ;
        RECT 42.65 24.135 42.91 24.395 ;
        RECT 42.65 23.375 42.91 23.635 ;
        RECT 43.41 30.215 43.67 30.475 ;
        RECT 43.41 29.455 43.67 29.715 ;
        RECT 43.41 28.695 43.67 28.955 ;
        RECT 43.41 27.935 43.67 28.195 ;
        RECT 43.41 27.175 43.67 27.435 ;
        RECT 43.41 26.415 43.67 26.675 ;
        RECT 43.41 25.655 43.67 25.915 ;
        RECT 43.41 24.895 43.67 25.155 ;
        RECT 43.41 24.135 43.67 24.395 ;
        RECT 43.41 23.375 43.67 23.635 ;
        RECT 44.17 30.215 44.43 30.475 ;
        RECT 44.17 29.455 44.43 29.715 ;
        RECT 44.17 28.695 44.43 28.955 ;
        RECT 44.17 27.935 44.43 28.195 ;
        RECT 44.17 27.175 44.43 27.435 ;
        RECT 44.17 26.415 44.43 26.675 ;
        RECT 44.17 25.655 44.43 25.915 ;
        RECT 44.17 24.895 44.43 25.155 ;
        RECT 44.17 24.135 44.43 24.395 ;
        RECT 44.17 23.375 44.43 23.635 ;
        RECT 44.93 30.215 45.19 30.475 ;
        RECT 44.93 29.455 45.19 29.715 ;
        RECT 44.93 28.695 45.19 28.955 ;
        RECT 44.93 27.935 45.19 28.195 ;
        RECT 44.93 27.175 45.19 27.435 ;
        RECT 44.93 26.415 45.19 26.675 ;
        RECT 44.93 25.655 45.19 25.915 ;
        RECT 44.93 24.895 45.19 25.155 ;
        RECT 44.93 24.135 45.19 24.395 ;
        RECT 44.93 23.375 45.19 23.635 ;
        RECT 45.69 30.215 45.95 30.475 ;
        RECT 45.69 29.455 45.95 29.715 ;
        RECT 45.69 28.695 45.95 28.955 ;
        RECT 45.69 27.935 45.95 28.195 ;
        RECT 45.69 27.175 45.95 27.435 ;
        RECT 45.69 26.415 45.95 26.675 ;
        RECT 45.69 25.655 45.95 25.915 ;
        RECT 45.69 24.895 45.95 25.155 ;
        RECT 45.69 24.135 45.95 24.395 ;
        RECT 45.69 23.375 45.95 23.635 ;
        RECT 46.45 30.215 46.71 30.475 ;
        RECT 46.45 29.455 46.71 29.715 ;
        RECT 46.45 28.695 46.71 28.955 ;
        RECT 46.45 27.935 46.71 28.195 ;
        RECT 46.45 27.175 46.71 27.435 ;
        RECT 46.45 26.415 46.71 26.675 ;
        RECT 46.45 25.655 46.71 25.915 ;
        RECT 46.45 24.895 46.71 25.155 ;
        RECT 46.45 24.135 46.71 24.395 ;
        RECT 46.45 23.375 46.71 23.635 ;
        RECT 47.21 30.215 47.47 30.475 ;
        RECT 47.21 29.455 47.47 29.715 ;
        RECT 47.21 28.695 47.47 28.955 ;
        RECT 47.21 27.935 47.47 28.195 ;
        RECT 47.21 27.175 47.47 27.435 ;
        RECT 47.21 26.415 47.47 26.675 ;
        RECT 47.21 25.655 47.47 25.915 ;
        RECT 47.21 24.895 47.47 25.155 ;
        RECT 47.21 24.135 47.47 24.395 ;
        RECT 47.21 23.375 47.47 23.635 ;
        RECT 47.97 30.215 48.23 30.475 ;
        RECT 47.97 29.455 48.23 29.715 ;
        RECT 47.97 28.695 48.23 28.955 ;
        RECT 47.97 27.935 48.23 28.195 ;
        RECT 47.97 27.175 48.23 27.435 ;
        RECT 47.97 26.415 48.23 26.675 ;
        RECT 47.97 25.655 48.23 25.915 ;
        RECT 47.97 24.895 48.23 25.155 ;
        RECT 47.97 24.135 48.23 24.395 ;
        RECT 47.97 23.375 48.23 23.635 ;
        RECT 48.73 30.215 48.99 30.475 ;
        RECT 48.73 29.455 48.99 29.715 ;
        RECT 48.73 28.695 48.99 28.955 ;
        RECT 48.73 27.935 48.99 28.195 ;
        RECT 48.73 27.175 48.99 27.435 ;
        RECT 48.73 26.415 48.99 26.675 ;
        RECT 48.73 25.655 48.99 25.915 ;
        RECT 48.73 24.895 48.99 25.155 ;
        RECT 48.73 24.135 48.99 24.395 ;
        RECT 48.73 23.375 48.99 23.635 ;
        RECT 49.49 30.215 49.75 30.475 ;
        RECT 49.49 29.455 49.75 29.715 ;
        RECT 49.49 28.695 49.75 28.955 ;
        RECT 49.49 27.935 49.75 28.195 ;
        RECT 49.49 27.175 49.75 27.435 ;
        RECT 49.49 26.415 49.75 26.675 ;
        RECT 49.49 25.655 49.75 25.915 ;
        RECT 49.49 24.895 49.75 25.155 ;
        RECT 49.49 24.135 49.75 24.395 ;
        RECT 49.49 23.375 49.75 23.635 ;
        RECT 50.25 30.215 50.51 30.475 ;
        RECT 50.25 29.455 50.51 29.715 ;
        RECT 50.25 28.695 50.51 28.955 ;
        RECT 50.25 27.935 50.51 28.195 ;
        RECT 50.25 27.175 50.51 27.435 ;
        RECT 50.25 26.415 50.51 26.675 ;
        RECT 50.25 25.655 50.51 25.915 ;
        RECT 50.25 24.895 50.51 25.155 ;
        RECT 50.25 24.135 50.51 24.395 ;
        RECT 50.25 23.375 50.51 23.635 ;
        RECT 51.01 30.215 51.27 30.475 ;
        RECT 51.01 29.455 51.27 29.715 ;
        RECT 51.01 28.695 51.27 28.955 ;
        RECT 51.01 27.935 51.27 28.195 ;
        RECT 51.01 27.175 51.27 27.435 ;
        RECT 51.01 26.415 51.27 26.675 ;
        RECT 51.01 25.655 51.27 25.915 ;
        RECT 51.01 24.895 51.27 25.155 ;
        RECT 51.01 24.135 51.27 24.395 ;
        RECT 51.01 23.375 51.27 23.635 ;
        RECT 51.77 30.215 52.03 30.475 ;
        RECT 51.77 29.455 52.03 29.715 ;
        RECT 51.77 28.695 52.03 28.955 ;
        RECT 51.77 27.935 52.03 28.195 ;
        RECT 51.77 27.175 52.03 27.435 ;
        RECT 51.77 26.415 52.03 26.675 ;
        RECT 51.77 25.655 52.03 25.915 ;
        RECT 51.77 24.895 52.03 25.155 ;
        RECT 51.77 24.135 52.03 24.395 ;
        RECT 51.77 23.375 52.03 23.635 ;
        RECT 52.53 30.215 52.79 30.475 ;
        RECT 52.53 29.455 52.79 29.715 ;
        RECT 52.53 28.695 52.79 28.955 ;
        RECT 52.53 27.935 52.79 28.195 ;
        RECT 52.53 27.175 52.79 27.435 ;
        RECT 52.53 26.415 52.79 26.675 ;
        RECT 52.53 25.655 52.79 25.915 ;
        RECT 52.53 24.895 52.79 25.155 ;
        RECT 52.53 24.135 52.79 24.395 ;
        RECT 52.53 23.375 52.79 23.635 ;
        RECT 53.29 30.215 53.55 30.475 ;
        RECT 53.29 29.455 53.55 29.715 ;
        RECT 53.29 28.695 53.55 28.955 ;
        RECT 53.29 27.935 53.55 28.195 ;
        RECT 53.29 27.175 53.55 27.435 ;
        RECT 53.29 26.415 53.55 26.675 ;
        RECT 53.29 25.655 53.55 25.915 ;
        RECT 53.29 24.895 53.55 25.155 ;
        RECT 53.29 24.135 53.55 24.395 ;
        RECT 53.29 23.375 53.55 23.635 ;
        RECT 54.05 30.215 54.31 30.475 ;
        RECT 54.05 29.455 54.31 29.715 ;
        RECT 54.05 28.695 54.31 28.955 ;
        RECT 54.05 27.935 54.31 28.195 ;
        RECT 54.05 27.175 54.31 27.435 ;
        RECT 54.05 26.415 54.31 26.675 ;
        RECT 54.05 25.655 54.31 25.915 ;
        RECT 54.05 24.895 54.31 25.155 ;
        RECT 54.05 24.135 54.31 24.395 ;
        RECT 54.05 23.375 54.31 23.635 ;
        RECT 54.81 30.215 55.07 30.475 ;
        RECT 54.81 29.455 55.07 29.715 ;
        RECT 54.81 28.695 55.07 28.955 ;
        RECT 54.81 27.935 55.07 28.195 ;
        RECT 54.81 27.175 55.07 27.435 ;
        RECT 54.81 26.415 55.07 26.675 ;
        RECT 54.81 25.655 55.07 25.915 ;
        RECT 54.81 24.895 55.07 25.155 ;
        RECT 54.81 24.135 55.07 24.395 ;
        RECT 54.81 23.375 55.07 23.635 ;
        RECT 55.57 30.215 55.83 30.475 ;
        RECT 55.57 29.455 55.83 29.715 ;
        RECT 55.57 28.695 55.83 28.955 ;
        RECT 55.57 27.935 55.83 28.195 ;
        RECT 55.57 27.175 55.83 27.435 ;
        RECT 55.57 26.415 55.83 26.675 ;
        RECT 55.57 25.655 55.83 25.915 ;
        RECT 55.57 24.895 55.83 25.155 ;
        RECT 55.57 24.135 55.83 24.395 ;
        RECT 55.57 23.375 55.83 23.635 ;
        RECT 56.33 30.215 56.59 30.475 ;
        RECT 56.33 29.455 56.59 29.715 ;
        RECT 56.33 28.695 56.59 28.955 ;
        RECT 56.33 27.935 56.59 28.195 ;
        RECT 56.33 27.175 56.59 27.435 ;
        RECT 56.33 26.415 56.59 26.675 ;
        RECT 56.33 25.655 56.59 25.915 ;
        RECT 56.33 24.895 56.59 25.155 ;
        RECT 56.33 24.135 56.59 24.395 ;
        RECT 56.33 23.375 56.59 23.635 ;
        RECT 57.09 30.215 57.35 30.475 ;
        RECT 57.09 29.455 57.35 29.715 ;
        RECT 57.09 28.695 57.35 28.955 ;
        RECT 57.09 27.935 57.35 28.195 ;
        RECT 57.09 27.175 57.35 27.435 ;
        RECT 57.09 26.415 57.35 26.675 ;
        RECT 57.09 25.655 57.35 25.915 ;
        RECT 57.09 24.895 57.35 25.155 ;
        RECT 57.09 24.135 57.35 24.395 ;
        RECT 57.09 23.375 57.35 23.635 ;
        RECT 57.85 30.215 58.11 30.475 ;
        RECT 57.85 29.455 58.11 29.715 ;
        RECT 57.85 28.695 58.11 28.955 ;
        RECT 57.85 27.935 58.11 28.195 ;
        RECT 57.85 27.175 58.11 27.435 ;
        RECT 57.85 26.415 58.11 26.675 ;
        RECT 57.85 25.655 58.11 25.915 ;
        RECT 57.85 24.895 58.11 25.155 ;
        RECT 57.85 24.135 58.11 24.395 ;
        RECT 57.85 23.375 58.11 23.635 ;
        RECT 58.61 30.215 58.87 30.475 ;
        RECT 58.61 29.455 58.87 29.715 ;
        RECT 58.61 28.695 58.87 28.955 ;
        RECT 58.61 27.935 58.87 28.195 ;
        RECT 58.61 27.175 58.87 27.435 ;
        RECT 58.61 26.415 58.87 26.675 ;
        RECT 58.61 25.655 58.87 25.915 ;
        RECT 58.61 24.895 58.87 25.155 ;
        RECT 58.61 24.135 58.87 24.395 ;
        RECT 58.61 23.375 58.87 23.635 ;
        RECT 59.37 30.215 59.63 30.475 ;
        RECT 59.37 29.455 59.63 29.715 ;
        RECT 59.37 28.695 59.63 28.955 ;
        RECT 59.37 27.935 59.63 28.195 ;
        RECT 59.37 27.175 59.63 27.435 ;
        RECT 59.37 26.415 59.63 26.675 ;
        RECT 59.37 25.655 59.63 25.915 ;
        RECT 59.37 24.895 59.63 25.155 ;
        RECT 59.37 24.135 59.63 24.395 ;
        RECT 59.37 23.375 59.63 23.635 ;
        RECT 60.13 30.215 60.39 30.475 ;
        RECT 60.13 29.455 60.39 29.715 ;
        RECT 60.13 28.695 60.39 28.955 ;
        RECT 60.13 27.935 60.39 28.195 ;
        RECT 60.13 27.175 60.39 27.435 ;
        RECT 60.13 26.415 60.39 26.675 ;
        RECT 60.13 25.655 60.39 25.915 ;
        RECT 60.13 24.895 60.39 25.155 ;
        RECT 60.13 24.135 60.39 24.395 ;
        RECT 60.13 23.375 60.39 23.635 ;
        RECT 60.89 30.215 61.15 30.475 ;
        RECT 60.89 29.455 61.15 29.715 ;
        RECT 60.89 28.695 61.15 28.955 ;
        RECT 60.89 27.935 61.15 28.195 ;
        RECT 60.89 27.175 61.15 27.435 ;
        RECT 60.89 26.415 61.15 26.675 ;
        RECT 60.89 25.655 61.15 25.915 ;
        RECT 60.89 24.895 61.15 25.155 ;
        RECT 60.89 24.135 61.15 24.395 ;
        RECT 60.89 23.375 61.15 23.635 ;
        RECT 61.65 30.215 61.91 30.475 ;
        RECT 61.65 29.455 61.91 29.715 ;
        RECT 61.65 28.695 61.91 28.955 ;
        RECT 61.65 27.935 61.91 28.195 ;
        RECT 61.65 27.175 61.91 27.435 ;
        RECT 61.65 26.415 61.91 26.675 ;
        RECT 61.65 25.655 61.91 25.915 ;
        RECT 61.65 24.895 61.91 25.155 ;
        RECT 61.65 24.135 61.91 24.395 ;
        RECT 61.65 23.375 61.91 23.635 ;
        RECT 62.41 30.215 62.67 30.475 ;
        RECT 62.41 29.455 62.67 29.715 ;
        RECT 62.41 28.695 62.67 28.955 ;
        RECT 62.41 27.935 62.67 28.195 ;
        RECT 62.41 27.175 62.67 27.435 ;
        RECT 62.41 26.415 62.67 26.675 ;
        RECT 62.41 25.655 62.67 25.915 ;
        RECT 62.41 24.895 62.67 25.155 ;
        RECT 62.41 24.135 62.67 24.395 ;
        RECT 62.41 23.375 62.67 23.635 ;
        RECT 63.17 30.215 63.43 30.475 ;
        RECT 63.17 29.455 63.43 29.715 ;
        RECT 63.17 28.695 63.43 28.955 ;
        RECT 63.17 27.935 63.43 28.195 ;
        RECT 63.17 27.175 63.43 27.435 ;
        RECT 63.17 26.415 63.43 26.675 ;
        RECT 63.17 25.655 63.43 25.915 ;
        RECT 63.17 24.895 63.43 25.155 ;
        RECT 63.17 24.135 63.43 24.395 ;
        RECT 63.17 23.375 63.43 23.635 ;
        RECT 63.93 30.215 64.19 30.475 ;
        RECT 63.93 29.455 64.19 29.715 ;
        RECT 63.93 28.695 64.19 28.955 ;
        RECT 63.93 27.935 64.19 28.195 ;
        RECT 63.93 27.175 64.19 27.435 ;
        RECT 63.93 26.415 64.19 26.675 ;
        RECT 63.93 25.655 64.19 25.915 ;
        RECT 63.93 24.895 64.19 25.155 ;
        RECT 63.93 24.135 64.19 24.395 ;
        RECT 63.93 23.375 64.19 23.635 ;
        RECT 64.69 30.215 64.95 30.475 ;
        RECT 64.69 29.455 64.95 29.715 ;
        RECT 64.69 28.695 64.95 28.955 ;
        RECT 64.69 27.935 64.95 28.195 ;
        RECT 64.69 27.175 64.95 27.435 ;
        RECT 64.69 26.415 64.95 26.675 ;
        RECT 64.69 25.655 64.95 25.915 ;
        RECT 64.69 24.895 64.95 25.155 ;
        RECT 64.69 24.135 64.95 24.395 ;
        RECT 64.69 23.375 64.95 23.635 ;
        RECT 65.45 30.215 65.71 30.475 ;
        RECT 65.45 29.455 65.71 29.715 ;
        RECT 65.45 28.695 65.71 28.955 ;
        RECT 65.45 27.935 65.71 28.195 ;
        RECT 65.45 27.175 65.71 27.435 ;
        RECT 65.45 26.415 65.71 26.675 ;
        RECT 65.45 25.655 65.71 25.915 ;
        RECT 65.45 24.895 65.71 25.155 ;
        RECT 65.45 24.135 65.71 24.395 ;
        RECT 65.45 23.375 65.71 23.635 ;
        RECT 66.21 30.215 66.47 30.475 ;
        RECT 66.21 29.455 66.47 29.715 ;
        RECT 66.21 28.695 66.47 28.955 ;
        RECT 66.21 27.935 66.47 28.195 ;
        RECT 66.21 27.175 66.47 27.435 ;
        RECT 66.21 26.415 66.47 26.675 ;
        RECT 66.21 25.655 66.47 25.915 ;
        RECT 66.21 24.895 66.47 25.155 ;
        RECT 66.21 24.135 66.47 24.395 ;
        RECT 66.21 23.375 66.47 23.635 ;
        RECT 66.97 30.215 67.23 30.475 ;
        RECT 66.97 29.455 67.23 29.715 ;
        RECT 66.97 28.695 67.23 28.955 ;
        RECT 66.97 27.935 67.23 28.195 ;
        RECT 66.97 27.175 67.23 27.435 ;
        RECT 66.97 26.415 67.23 26.675 ;
        RECT 66.97 25.655 67.23 25.915 ;
        RECT 66.97 24.895 67.23 25.155 ;
        RECT 66.97 24.135 67.23 24.395 ;
        RECT 66.97 23.375 67.23 23.635 ;
        RECT 67.73 30.215 67.99 30.475 ;
        RECT 67.73 29.455 67.99 29.715 ;
        RECT 67.73 28.695 67.99 28.955 ;
        RECT 67.73 27.935 67.99 28.195 ;
        RECT 67.73 27.175 67.99 27.435 ;
        RECT 67.73 26.415 67.99 26.675 ;
        RECT 67.73 25.655 67.99 25.915 ;
        RECT 67.73 24.895 67.99 25.155 ;
        RECT 67.73 24.135 67.99 24.395 ;
        RECT 67.73 23.375 67.99 23.635 ;
        RECT 68.49 30.215 68.75 30.475 ;
        RECT 68.49 29.455 68.75 29.715 ;
        RECT 68.49 28.695 68.75 28.955 ;
        RECT 68.49 27.935 68.75 28.195 ;
        RECT 68.49 27.175 68.75 27.435 ;
        RECT 68.49 26.415 68.75 26.675 ;
        RECT 68.49 25.655 68.75 25.915 ;
        RECT 68.49 24.895 68.75 25.155 ;
        RECT 68.49 24.135 68.75 24.395 ;
        RECT 68.49 23.375 68.75 23.635 ;
        RECT 69.25 30.215 69.51 30.475 ;
        RECT 69.25 29.455 69.51 29.715 ;
        RECT 69.25 28.695 69.51 28.955 ;
        RECT 69.25 27.935 69.51 28.195 ;
        RECT 69.25 27.175 69.51 27.435 ;
        RECT 69.25 26.415 69.51 26.675 ;
        RECT 69.25 25.655 69.51 25.915 ;
        RECT 69.25 24.895 69.51 25.155 ;
        RECT 69.25 24.135 69.51 24.395 ;
        RECT 69.25 23.375 69.51 23.635 ;
        RECT 70.01 30.215 70.27 30.475 ;
        RECT 70.01 29.455 70.27 29.715 ;
        RECT 70.01 28.695 70.27 28.955 ;
        RECT 70.01 27.935 70.27 28.195 ;
        RECT 70.01 27.175 70.27 27.435 ;
        RECT 70.01 26.415 70.27 26.675 ;
        RECT 70.01 25.655 70.27 25.915 ;
        RECT 70.01 24.895 70.27 25.155 ;
        RECT 70.01 24.135 70.27 24.395 ;
        RECT 70.01 23.375 70.27 23.635 ;
        RECT 70.77 30.215 71.03 30.475 ;
        RECT 70.77 29.455 71.03 29.715 ;
        RECT 70.77 28.695 71.03 28.955 ;
        RECT 70.77 27.935 71.03 28.195 ;
        RECT 70.77 27.175 71.03 27.435 ;
        RECT 70.77 26.415 71.03 26.675 ;
        RECT 70.77 25.655 71.03 25.915 ;
        RECT 70.77 24.895 71.03 25.155 ;
        RECT 70.77 24.135 71.03 24.395 ;
        RECT 70.77 23.375 71.03 23.635 ;
        RECT 71.53 30.215 71.79 30.475 ;
        RECT 71.53 29.455 71.79 29.715 ;
        RECT 71.53 28.695 71.79 28.955 ;
        RECT 71.53 27.935 71.79 28.195 ;
        RECT 71.53 27.175 71.79 27.435 ;
        RECT 71.53 26.415 71.79 26.675 ;
        RECT 71.53 25.655 71.79 25.915 ;
        RECT 71.53 24.895 71.79 25.155 ;
        RECT 71.53 24.135 71.79 24.395 ;
        RECT 71.53 23.375 71.79 23.635 ;
        RECT 72.29 30.215 72.55 30.475 ;
        RECT 72.29 29.455 72.55 29.715 ;
        RECT 72.29 28.695 72.55 28.955 ;
        RECT 72.29 27.935 72.55 28.195 ;
        RECT 72.29 27.175 72.55 27.435 ;
        RECT 72.29 26.415 72.55 26.675 ;
        RECT 72.29 25.655 72.55 25.915 ;
        RECT 72.29 24.895 72.55 25.155 ;
        RECT 72.29 24.135 72.55 24.395 ;
        RECT 72.29 23.375 72.55 23.635 ;
        RECT 73.05 30.215 73.31 30.475 ;
        RECT 73.05 29.455 73.31 29.715 ;
        RECT 73.05 28.695 73.31 28.955 ;
        RECT 73.05 27.935 73.31 28.195 ;
        RECT 73.05 27.175 73.31 27.435 ;
        RECT 73.05 26.415 73.31 26.675 ;
        RECT 73.05 25.655 73.31 25.915 ;
        RECT 73.05 24.895 73.31 25.155 ;
        RECT 73.05 24.135 73.31 24.395 ;
        RECT 73.05 23.375 73.31 23.635 ;
        RECT 73.81 30.215 74.07 30.475 ;
        RECT 73.81 29.455 74.07 29.715 ;
        RECT 73.81 28.695 74.07 28.955 ;
        RECT 73.81 27.935 74.07 28.195 ;
        RECT 73.81 27.175 74.07 27.435 ;
        RECT 73.81 26.415 74.07 26.675 ;
        RECT 73.81 25.655 74.07 25.915 ;
        RECT 73.81 24.895 74.07 25.155 ;
        RECT 73.81 24.135 74.07 24.395 ;
        RECT 73.81 23.375 74.07 23.635 ;
        RECT 74.57 30.215 74.83 30.475 ;
        RECT 74.57 29.455 74.83 29.715 ;
        RECT 74.57 28.695 74.83 28.955 ;
        RECT 74.57 27.935 74.83 28.195 ;
        RECT 74.57 27.175 74.83 27.435 ;
        RECT 74.57 26.415 74.83 26.675 ;
        RECT 74.57 25.655 74.83 25.915 ;
        RECT 74.57 24.895 74.83 25.155 ;
        RECT 74.57 24.135 74.83 24.395 ;
        RECT 74.57 23.375 74.83 23.635 ;
        RECT 75.33 30.215 75.59 30.475 ;
        RECT 75.33 29.455 75.59 29.715 ;
        RECT 75.33 28.695 75.59 28.955 ;
        RECT 75.33 27.935 75.59 28.195 ;
        RECT 75.33 27.175 75.59 27.435 ;
        RECT 75.33 26.415 75.59 26.675 ;
        RECT 75.33 25.655 75.59 25.915 ;
        RECT 75.33 24.895 75.59 25.155 ;
        RECT 75.33 24.135 75.59 24.395 ;
        RECT 75.33 23.375 75.59 23.635 ;
        RECT 76.09 30.215 76.35 30.475 ;
        RECT 76.09 29.455 76.35 29.715 ;
        RECT 76.09 28.695 76.35 28.955 ;
        RECT 76.09 27.935 76.35 28.195 ;
        RECT 76.09 27.175 76.35 27.435 ;
        RECT 76.09 26.415 76.35 26.675 ;
        RECT 76.09 25.655 76.35 25.915 ;
        RECT 76.09 24.895 76.35 25.155 ;
        RECT 76.09 24.135 76.35 24.395 ;
        RECT 76.09 23.375 76.35 23.635 ;
        RECT 76.85 30.215 77.11 30.475 ;
        RECT 76.85 29.455 77.11 29.715 ;
        RECT 76.85 28.695 77.11 28.955 ;
        RECT 76.85 27.935 77.11 28.195 ;
        RECT 76.85 27.175 77.11 27.435 ;
        RECT 76.85 26.415 77.11 26.675 ;
        RECT 76.85 25.655 77.11 25.915 ;
        RECT 76.85 24.895 77.11 25.155 ;
        RECT 76.85 24.135 77.11 24.395 ;
        RECT 76.85 23.375 77.11 23.635 ;
        RECT 77.61 30.215 77.87 30.475 ;
        RECT 77.61 29.455 77.87 29.715 ;
        RECT 77.61 28.695 77.87 28.955 ;
        RECT 77.61 27.935 77.87 28.195 ;
        RECT 77.61 27.175 77.87 27.435 ;
        RECT 77.61 26.415 77.87 26.675 ;
        RECT 77.61 25.655 77.87 25.915 ;
        RECT 77.61 24.895 77.87 25.155 ;
        RECT 77.61 24.135 77.87 24.395 ;
        RECT 77.61 23.375 77.87 23.635 ;
        RECT 78.37 30.215 78.63 30.475 ;
        RECT 78.37 29.455 78.63 29.715 ;
        RECT 78.37 28.695 78.63 28.955 ;
        RECT 78.37 27.935 78.63 28.195 ;
        RECT 78.37 27.175 78.63 27.435 ;
        RECT 78.37 26.415 78.63 26.675 ;
        RECT 78.37 25.655 78.63 25.915 ;
        RECT 78.37 24.895 78.63 25.155 ;
        RECT 78.37 24.135 78.63 24.395 ;
        RECT 78.37 23.375 78.63 23.635 ;
        RECT 79.13 30.215 79.39 30.475 ;
        RECT 79.13 29.455 79.39 29.715 ;
        RECT 79.13 28.695 79.39 28.955 ;
        RECT 79.13 27.935 79.39 28.195 ;
        RECT 79.13 27.175 79.39 27.435 ;
        RECT 79.13 26.415 79.39 26.675 ;
        RECT 79.13 25.655 79.39 25.915 ;
        RECT 79.13 24.895 79.39 25.155 ;
        RECT 79.13 24.135 79.39 24.395 ;
        RECT 79.13 23.375 79.39 23.635 ;
        RECT 79.89 30.215 80.15 30.475 ;
        RECT 79.89 29.455 80.15 29.715 ;
        RECT 79.89 28.695 80.15 28.955 ;
        RECT 79.89 27.935 80.15 28.195 ;
        RECT 79.89 27.175 80.15 27.435 ;
        RECT 79.89 26.415 80.15 26.675 ;
        RECT 79.89 25.655 80.15 25.915 ;
        RECT 79.89 24.895 80.15 25.155 ;
        RECT 79.89 24.135 80.15 24.395 ;
        RECT 79.89 23.375 80.15 23.635 ;
    END
  END AVSS
  PIN AVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M3 ;
        RECT 0 10 100 20 ;
      LAYER M4 ;
        RECT 0 10 100 20 ;
      LAYER V4 ;
        RECT 80.65 18.24 80.91 18.5 ;
        RECT 80.65 17.48 80.91 17.74 ;
        RECT 80.65 16.72 80.91 16.98 ;
        RECT 80.65 15.96 80.91 16.22 ;
        RECT 80.65 15.2 80.91 15.46 ;
        RECT 80.65 14.44 80.91 14.7 ;
        RECT 80.65 13.68 80.91 13.94 ;
        RECT 80.65 12.92 80.91 13.18 ;
        RECT 80.65 12.16 80.91 12.42 ;
        RECT 80.65 11.4 80.91 11.66 ;
        RECT 81.41 18.24 81.67 18.5 ;
        RECT 81.41 17.48 81.67 17.74 ;
        RECT 81.41 16.72 81.67 16.98 ;
        RECT 81.41 15.96 81.67 16.22 ;
        RECT 81.41 15.2 81.67 15.46 ;
        RECT 81.41 14.44 81.67 14.7 ;
        RECT 81.41 13.68 81.67 13.94 ;
        RECT 81.41 12.92 81.67 13.18 ;
        RECT 81.41 12.16 81.67 12.42 ;
        RECT 81.41 11.4 81.67 11.66 ;
        RECT 82.17 18.24 82.43 18.5 ;
        RECT 82.17 17.48 82.43 17.74 ;
        RECT 82.17 16.72 82.43 16.98 ;
        RECT 82.17 15.96 82.43 16.22 ;
        RECT 82.17 15.2 82.43 15.46 ;
        RECT 82.17 14.44 82.43 14.7 ;
        RECT 82.17 13.68 82.43 13.94 ;
        RECT 82.17 12.92 82.43 13.18 ;
        RECT 82.17 12.16 82.43 12.42 ;
        RECT 82.17 11.4 82.43 11.66 ;
        RECT 82.93 18.24 83.19 18.5 ;
        RECT 82.93 17.48 83.19 17.74 ;
        RECT 82.93 16.72 83.19 16.98 ;
        RECT 82.93 15.96 83.19 16.22 ;
        RECT 82.93 15.2 83.19 15.46 ;
        RECT 82.93 14.44 83.19 14.7 ;
        RECT 82.93 13.68 83.19 13.94 ;
        RECT 82.93 12.92 83.19 13.18 ;
        RECT 82.93 12.16 83.19 12.42 ;
        RECT 82.93 11.4 83.19 11.66 ;
        RECT 83.69 18.24 83.95 18.5 ;
        RECT 83.69 17.48 83.95 17.74 ;
        RECT 83.69 16.72 83.95 16.98 ;
        RECT 83.69 15.96 83.95 16.22 ;
        RECT 83.69 15.2 83.95 15.46 ;
        RECT 83.69 14.44 83.95 14.7 ;
        RECT 83.69 13.68 83.95 13.94 ;
        RECT 83.69 12.92 83.95 13.18 ;
        RECT 83.69 12.16 83.95 12.42 ;
        RECT 83.69 11.4 83.95 11.66 ;
        RECT 84.45 18.24 84.71 18.5 ;
        RECT 84.45 17.48 84.71 17.74 ;
        RECT 84.45 16.72 84.71 16.98 ;
        RECT 84.45 15.96 84.71 16.22 ;
        RECT 84.45 15.2 84.71 15.46 ;
        RECT 84.45 14.44 84.71 14.7 ;
        RECT 84.45 13.68 84.71 13.94 ;
        RECT 84.45 12.92 84.71 13.18 ;
        RECT 84.45 12.16 84.71 12.42 ;
        RECT 84.45 11.4 84.71 11.66 ;
        RECT 85.21 18.24 85.47 18.5 ;
        RECT 85.21 17.48 85.47 17.74 ;
        RECT 85.21 16.72 85.47 16.98 ;
        RECT 85.21 15.96 85.47 16.22 ;
        RECT 85.21 15.2 85.47 15.46 ;
        RECT 85.21 14.44 85.47 14.7 ;
        RECT 85.21 13.68 85.47 13.94 ;
        RECT 85.21 12.92 85.47 13.18 ;
        RECT 85.21 12.16 85.47 12.42 ;
        RECT 85.21 11.4 85.47 11.66 ;
        RECT 85.97 18.24 86.23 18.5 ;
        RECT 85.97 17.48 86.23 17.74 ;
        RECT 85.97 16.72 86.23 16.98 ;
        RECT 85.97 15.96 86.23 16.22 ;
        RECT 85.97 15.2 86.23 15.46 ;
        RECT 85.97 14.44 86.23 14.7 ;
        RECT 85.97 13.68 86.23 13.94 ;
        RECT 85.97 12.92 86.23 13.18 ;
        RECT 85.97 12.16 86.23 12.42 ;
        RECT 85.97 11.4 86.23 11.66 ;
        RECT 86.73 18.24 86.99 18.5 ;
        RECT 86.73 17.48 86.99 17.74 ;
        RECT 86.73 16.72 86.99 16.98 ;
        RECT 86.73 15.96 86.99 16.22 ;
        RECT 86.73 15.2 86.99 15.46 ;
        RECT 86.73 14.44 86.99 14.7 ;
        RECT 86.73 13.68 86.99 13.94 ;
        RECT 86.73 12.92 86.99 13.18 ;
        RECT 86.73 12.16 86.99 12.42 ;
        RECT 86.73 11.4 86.99 11.66 ;
        RECT 87.49 18.24 87.75 18.5 ;
        RECT 87.49 17.48 87.75 17.74 ;
        RECT 87.49 16.72 87.75 16.98 ;
        RECT 87.49 15.96 87.75 16.22 ;
        RECT 87.49 15.2 87.75 15.46 ;
        RECT 87.49 14.44 87.75 14.7 ;
        RECT 87.49 13.68 87.75 13.94 ;
        RECT 87.49 12.92 87.75 13.18 ;
        RECT 87.49 12.16 87.75 12.42 ;
        RECT 87.49 11.4 87.75 11.66 ;
        RECT 88.25 18.24 88.51 18.5 ;
        RECT 88.25 17.48 88.51 17.74 ;
        RECT 88.25 16.72 88.51 16.98 ;
        RECT 88.25 15.96 88.51 16.22 ;
        RECT 88.25 15.2 88.51 15.46 ;
        RECT 88.25 14.44 88.51 14.7 ;
        RECT 88.25 13.68 88.51 13.94 ;
        RECT 88.25 12.92 88.51 13.18 ;
        RECT 88.25 12.16 88.51 12.42 ;
        RECT 88.25 11.4 88.51 11.66 ;
        RECT 89.01 18.24 89.27 18.5 ;
        RECT 89.01 17.48 89.27 17.74 ;
        RECT 89.01 16.72 89.27 16.98 ;
        RECT 89.01 15.96 89.27 16.22 ;
        RECT 89.01 15.2 89.27 15.46 ;
        RECT 89.01 14.44 89.27 14.7 ;
        RECT 89.01 13.68 89.27 13.94 ;
        RECT 89.01 12.92 89.27 13.18 ;
        RECT 89.01 12.16 89.27 12.42 ;
        RECT 89.01 11.4 89.27 11.66 ;
        RECT 89.77 18.24 90.03 18.5 ;
        RECT 89.77 17.48 90.03 17.74 ;
        RECT 89.77 16.72 90.03 16.98 ;
        RECT 89.77 15.96 90.03 16.22 ;
        RECT 89.77 15.2 90.03 15.46 ;
        RECT 89.77 14.44 90.03 14.7 ;
        RECT 89.77 13.68 90.03 13.94 ;
        RECT 89.77 12.92 90.03 13.18 ;
        RECT 89.77 12.16 90.03 12.42 ;
        RECT 89.77 11.4 90.03 11.66 ;
        RECT 90.53 18.24 90.79 18.5 ;
        RECT 90.53 17.48 90.79 17.74 ;
        RECT 90.53 16.72 90.79 16.98 ;
        RECT 90.53 15.96 90.79 16.22 ;
        RECT 90.53 15.2 90.79 15.46 ;
        RECT 90.53 14.44 90.79 14.7 ;
        RECT 90.53 13.68 90.79 13.94 ;
        RECT 90.53 12.92 90.79 13.18 ;
        RECT 90.53 12.16 90.79 12.42 ;
        RECT 90.53 11.4 90.79 11.66 ;
        RECT 91.29 18.24 91.55 18.5 ;
        RECT 91.29 17.48 91.55 17.74 ;
        RECT 91.29 16.72 91.55 16.98 ;
        RECT 91.29 15.96 91.55 16.22 ;
        RECT 91.29 15.2 91.55 15.46 ;
        RECT 91.29 14.44 91.55 14.7 ;
        RECT 91.29 13.68 91.55 13.94 ;
        RECT 91.29 12.92 91.55 13.18 ;
        RECT 91.29 12.16 91.55 12.42 ;
        RECT 91.29 11.4 91.55 11.66 ;
        RECT 92.05 18.24 92.31 18.5 ;
        RECT 92.05 17.48 92.31 17.74 ;
        RECT 92.05 16.72 92.31 16.98 ;
        RECT 92.05 15.96 92.31 16.22 ;
        RECT 92.05 15.2 92.31 15.46 ;
        RECT 92.05 14.44 92.31 14.7 ;
        RECT 92.05 13.68 92.31 13.94 ;
        RECT 92.05 12.92 92.31 13.18 ;
        RECT 92.05 12.16 92.31 12.42 ;
        RECT 92.05 11.4 92.31 11.66 ;
        RECT 92.81 18.24 93.07 18.5 ;
        RECT 92.81 17.48 93.07 17.74 ;
        RECT 92.81 16.72 93.07 16.98 ;
        RECT 92.81 15.96 93.07 16.22 ;
        RECT 92.81 15.2 93.07 15.46 ;
        RECT 92.81 14.44 93.07 14.7 ;
        RECT 92.81 13.68 93.07 13.94 ;
        RECT 92.81 12.92 93.07 13.18 ;
        RECT 92.81 12.16 93.07 12.42 ;
        RECT 92.81 11.4 93.07 11.66 ;
        RECT 93.57 18.24 93.83 18.5 ;
        RECT 93.57 17.48 93.83 17.74 ;
        RECT 93.57 16.72 93.83 16.98 ;
        RECT 93.57 15.96 93.83 16.22 ;
        RECT 93.57 15.2 93.83 15.46 ;
        RECT 93.57 14.44 93.83 14.7 ;
        RECT 93.57 13.68 93.83 13.94 ;
        RECT 93.57 12.92 93.83 13.18 ;
        RECT 93.57 12.16 93.83 12.42 ;
        RECT 93.57 11.4 93.83 11.66 ;
        RECT 94.33 18.24 94.59 18.5 ;
        RECT 94.33 17.48 94.59 17.74 ;
        RECT 94.33 16.72 94.59 16.98 ;
        RECT 94.33 15.96 94.59 16.22 ;
        RECT 94.33 15.2 94.59 15.46 ;
        RECT 94.33 14.44 94.59 14.7 ;
        RECT 94.33 13.68 94.59 13.94 ;
        RECT 94.33 12.92 94.59 13.18 ;
        RECT 94.33 12.16 94.59 12.42 ;
        RECT 94.33 11.4 94.59 11.66 ;
        RECT 95.09 18.24 95.35 18.5 ;
        RECT 95.09 17.48 95.35 17.74 ;
        RECT 95.09 16.72 95.35 16.98 ;
        RECT 95.09 15.96 95.35 16.22 ;
        RECT 95.09 15.2 95.35 15.46 ;
        RECT 95.09 14.44 95.35 14.7 ;
        RECT 95.09 13.68 95.35 13.94 ;
        RECT 95.09 12.92 95.35 13.18 ;
        RECT 95.09 12.16 95.35 12.42 ;
        RECT 95.09 11.4 95.35 11.66 ;
        RECT 4.65 18.24 4.91 18.5 ;
        RECT 4.65 17.48 4.91 17.74 ;
        RECT 4.65 16.72 4.91 16.98 ;
        RECT 4.65 15.96 4.91 16.22 ;
        RECT 4.65 15.2 4.91 15.46 ;
        RECT 4.65 14.44 4.91 14.7 ;
        RECT 4.65 13.68 4.91 13.94 ;
        RECT 4.65 12.92 4.91 13.18 ;
        RECT 4.65 12.16 4.91 12.42 ;
        RECT 4.65 11.4 4.91 11.66 ;
        RECT 5.41 18.24 5.67 18.5 ;
        RECT 5.41 17.48 5.67 17.74 ;
        RECT 5.41 16.72 5.67 16.98 ;
        RECT 5.41 15.96 5.67 16.22 ;
        RECT 5.41 15.2 5.67 15.46 ;
        RECT 5.41 14.44 5.67 14.7 ;
        RECT 5.41 13.68 5.67 13.94 ;
        RECT 5.41 12.92 5.67 13.18 ;
        RECT 5.41 12.16 5.67 12.42 ;
        RECT 5.41 11.4 5.67 11.66 ;
        RECT 6.17 18.24 6.43 18.5 ;
        RECT 6.17 17.48 6.43 17.74 ;
        RECT 6.17 16.72 6.43 16.98 ;
        RECT 6.17 15.96 6.43 16.22 ;
        RECT 6.17 15.2 6.43 15.46 ;
        RECT 6.17 14.44 6.43 14.7 ;
        RECT 6.17 13.68 6.43 13.94 ;
        RECT 6.17 12.92 6.43 13.18 ;
        RECT 6.17 12.16 6.43 12.42 ;
        RECT 6.17 11.4 6.43 11.66 ;
        RECT 6.93 18.24 7.19 18.5 ;
        RECT 6.93 17.48 7.19 17.74 ;
        RECT 6.93 16.72 7.19 16.98 ;
        RECT 6.93 15.96 7.19 16.22 ;
        RECT 6.93 15.2 7.19 15.46 ;
        RECT 6.93 14.44 7.19 14.7 ;
        RECT 6.93 13.68 7.19 13.94 ;
        RECT 6.93 12.92 7.19 13.18 ;
        RECT 6.93 12.16 7.19 12.42 ;
        RECT 6.93 11.4 7.19 11.66 ;
        RECT 7.69 18.24 7.95 18.5 ;
        RECT 7.69 17.48 7.95 17.74 ;
        RECT 7.69 16.72 7.95 16.98 ;
        RECT 7.69 15.96 7.95 16.22 ;
        RECT 7.69 15.2 7.95 15.46 ;
        RECT 7.69 14.44 7.95 14.7 ;
        RECT 7.69 13.68 7.95 13.94 ;
        RECT 7.69 12.92 7.95 13.18 ;
        RECT 7.69 12.16 7.95 12.42 ;
        RECT 7.69 11.4 7.95 11.66 ;
        RECT 8.45 18.24 8.71 18.5 ;
        RECT 8.45 17.48 8.71 17.74 ;
        RECT 8.45 16.72 8.71 16.98 ;
        RECT 8.45 15.96 8.71 16.22 ;
        RECT 8.45 15.2 8.71 15.46 ;
        RECT 8.45 14.44 8.71 14.7 ;
        RECT 8.45 13.68 8.71 13.94 ;
        RECT 8.45 12.92 8.71 13.18 ;
        RECT 8.45 12.16 8.71 12.42 ;
        RECT 8.45 11.4 8.71 11.66 ;
        RECT 9.21 18.24 9.47 18.5 ;
        RECT 9.21 17.48 9.47 17.74 ;
        RECT 9.21 16.72 9.47 16.98 ;
        RECT 9.21 15.96 9.47 16.22 ;
        RECT 9.21 15.2 9.47 15.46 ;
        RECT 9.21 14.44 9.47 14.7 ;
        RECT 9.21 13.68 9.47 13.94 ;
        RECT 9.21 12.92 9.47 13.18 ;
        RECT 9.21 12.16 9.47 12.42 ;
        RECT 9.21 11.4 9.47 11.66 ;
        RECT 9.97 18.24 10.23 18.5 ;
        RECT 9.97 17.48 10.23 17.74 ;
        RECT 9.97 16.72 10.23 16.98 ;
        RECT 9.97 15.96 10.23 16.22 ;
        RECT 9.97 15.2 10.23 15.46 ;
        RECT 9.97 14.44 10.23 14.7 ;
        RECT 9.97 13.68 10.23 13.94 ;
        RECT 9.97 12.92 10.23 13.18 ;
        RECT 9.97 12.16 10.23 12.42 ;
        RECT 9.97 11.4 10.23 11.66 ;
        RECT 10.73 18.24 10.99 18.5 ;
        RECT 10.73 17.48 10.99 17.74 ;
        RECT 10.73 16.72 10.99 16.98 ;
        RECT 10.73 15.96 10.99 16.22 ;
        RECT 10.73 15.2 10.99 15.46 ;
        RECT 10.73 14.44 10.99 14.7 ;
        RECT 10.73 13.68 10.99 13.94 ;
        RECT 10.73 12.92 10.99 13.18 ;
        RECT 10.73 12.16 10.99 12.42 ;
        RECT 10.73 11.4 10.99 11.66 ;
        RECT 11.49 18.24 11.75 18.5 ;
        RECT 11.49 17.48 11.75 17.74 ;
        RECT 11.49 16.72 11.75 16.98 ;
        RECT 11.49 15.96 11.75 16.22 ;
        RECT 11.49 15.2 11.75 15.46 ;
        RECT 11.49 14.44 11.75 14.7 ;
        RECT 11.49 13.68 11.75 13.94 ;
        RECT 11.49 12.92 11.75 13.18 ;
        RECT 11.49 12.16 11.75 12.42 ;
        RECT 11.49 11.4 11.75 11.66 ;
        RECT 12.25 18.24 12.51 18.5 ;
        RECT 12.25 17.48 12.51 17.74 ;
        RECT 12.25 16.72 12.51 16.98 ;
        RECT 12.25 15.96 12.51 16.22 ;
        RECT 12.25 15.2 12.51 15.46 ;
        RECT 12.25 14.44 12.51 14.7 ;
        RECT 12.25 13.68 12.51 13.94 ;
        RECT 12.25 12.92 12.51 13.18 ;
        RECT 12.25 12.16 12.51 12.42 ;
        RECT 12.25 11.4 12.51 11.66 ;
        RECT 13.01 18.24 13.27 18.5 ;
        RECT 13.01 17.48 13.27 17.74 ;
        RECT 13.01 16.72 13.27 16.98 ;
        RECT 13.01 15.96 13.27 16.22 ;
        RECT 13.01 15.2 13.27 15.46 ;
        RECT 13.01 14.44 13.27 14.7 ;
        RECT 13.01 13.68 13.27 13.94 ;
        RECT 13.01 12.92 13.27 13.18 ;
        RECT 13.01 12.16 13.27 12.42 ;
        RECT 13.01 11.4 13.27 11.66 ;
        RECT 13.77 18.24 14.03 18.5 ;
        RECT 13.77 17.48 14.03 17.74 ;
        RECT 13.77 16.72 14.03 16.98 ;
        RECT 13.77 15.96 14.03 16.22 ;
        RECT 13.77 15.2 14.03 15.46 ;
        RECT 13.77 14.44 14.03 14.7 ;
        RECT 13.77 13.68 14.03 13.94 ;
        RECT 13.77 12.92 14.03 13.18 ;
        RECT 13.77 12.16 14.03 12.42 ;
        RECT 13.77 11.4 14.03 11.66 ;
        RECT 14.53 18.24 14.79 18.5 ;
        RECT 14.53 17.48 14.79 17.74 ;
        RECT 14.53 16.72 14.79 16.98 ;
        RECT 14.53 15.96 14.79 16.22 ;
        RECT 14.53 15.2 14.79 15.46 ;
        RECT 14.53 14.44 14.79 14.7 ;
        RECT 14.53 13.68 14.79 13.94 ;
        RECT 14.53 12.92 14.79 13.18 ;
        RECT 14.53 12.16 14.79 12.42 ;
        RECT 14.53 11.4 14.79 11.66 ;
        RECT 15.29 18.24 15.55 18.5 ;
        RECT 15.29 17.48 15.55 17.74 ;
        RECT 15.29 16.72 15.55 16.98 ;
        RECT 15.29 15.96 15.55 16.22 ;
        RECT 15.29 15.2 15.55 15.46 ;
        RECT 15.29 14.44 15.55 14.7 ;
        RECT 15.29 13.68 15.55 13.94 ;
        RECT 15.29 12.92 15.55 13.18 ;
        RECT 15.29 12.16 15.55 12.42 ;
        RECT 15.29 11.4 15.55 11.66 ;
        RECT 16.05 18.24 16.31 18.5 ;
        RECT 16.05 17.48 16.31 17.74 ;
        RECT 16.05 16.72 16.31 16.98 ;
        RECT 16.05 15.96 16.31 16.22 ;
        RECT 16.05 15.2 16.31 15.46 ;
        RECT 16.05 14.44 16.31 14.7 ;
        RECT 16.05 13.68 16.31 13.94 ;
        RECT 16.05 12.92 16.31 13.18 ;
        RECT 16.05 12.16 16.31 12.42 ;
        RECT 16.05 11.4 16.31 11.66 ;
        RECT 16.81 18.24 17.07 18.5 ;
        RECT 16.81 17.48 17.07 17.74 ;
        RECT 16.81 16.72 17.07 16.98 ;
        RECT 16.81 15.96 17.07 16.22 ;
        RECT 16.81 15.2 17.07 15.46 ;
        RECT 16.81 14.44 17.07 14.7 ;
        RECT 16.81 13.68 17.07 13.94 ;
        RECT 16.81 12.92 17.07 13.18 ;
        RECT 16.81 12.16 17.07 12.42 ;
        RECT 16.81 11.4 17.07 11.66 ;
        RECT 17.57 18.24 17.83 18.5 ;
        RECT 17.57 17.48 17.83 17.74 ;
        RECT 17.57 16.72 17.83 16.98 ;
        RECT 17.57 15.96 17.83 16.22 ;
        RECT 17.57 15.2 17.83 15.46 ;
        RECT 17.57 14.44 17.83 14.7 ;
        RECT 17.57 13.68 17.83 13.94 ;
        RECT 17.57 12.92 17.83 13.18 ;
        RECT 17.57 12.16 17.83 12.42 ;
        RECT 17.57 11.4 17.83 11.66 ;
        RECT 18.33 18.24 18.59 18.5 ;
        RECT 18.33 17.48 18.59 17.74 ;
        RECT 18.33 16.72 18.59 16.98 ;
        RECT 18.33 15.96 18.59 16.22 ;
        RECT 18.33 15.2 18.59 15.46 ;
        RECT 18.33 14.44 18.59 14.7 ;
        RECT 18.33 13.68 18.59 13.94 ;
        RECT 18.33 12.92 18.59 13.18 ;
        RECT 18.33 12.16 18.59 12.42 ;
        RECT 18.33 11.4 18.59 11.66 ;
        RECT 19.09 18.24 19.35 18.5 ;
        RECT 19.09 17.48 19.35 17.74 ;
        RECT 19.09 16.72 19.35 16.98 ;
        RECT 19.09 15.96 19.35 16.22 ;
        RECT 19.09 15.2 19.35 15.46 ;
        RECT 19.09 14.44 19.35 14.7 ;
        RECT 19.09 13.68 19.35 13.94 ;
        RECT 19.09 12.92 19.35 13.18 ;
        RECT 19.09 12.16 19.35 12.42 ;
        RECT 19.09 11.4 19.35 11.66 ;
        RECT 19.85 18.24 20.11 18.5 ;
        RECT 19.85 17.48 20.11 17.74 ;
        RECT 19.85 16.72 20.11 16.98 ;
        RECT 19.85 15.96 20.11 16.22 ;
        RECT 19.85 15.2 20.11 15.46 ;
        RECT 19.85 14.44 20.11 14.7 ;
        RECT 19.85 13.68 20.11 13.94 ;
        RECT 19.85 12.92 20.11 13.18 ;
        RECT 19.85 12.16 20.11 12.42 ;
        RECT 19.85 11.4 20.11 11.66 ;
        RECT 20.61 18.24 20.87 18.5 ;
        RECT 20.61 17.48 20.87 17.74 ;
        RECT 20.61 16.72 20.87 16.98 ;
        RECT 20.61 15.96 20.87 16.22 ;
        RECT 20.61 15.2 20.87 15.46 ;
        RECT 20.61 14.44 20.87 14.7 ;
        RECT 20.61 13.68 20.87 13.94 ;
        RECT 20.61 12.92 20.87 13.18 ;
        RECT 20.61 12.16 20.87 12.42 ;
        RECT 20.61 11.4 20.87 11.66 ;
        RECT 21.37 18.24 21.63 18.5 ;
        RECT 21.37 17.48 21.63 17.74 ;
        RECT 21.37 16.72 21.63 16.98 ;
        RECT 21.37 15.96 21.63 16.22 ;
        RECT 21.37 15.2 21.63 15.46 ;
        RECT 21.37 14.44 21.63 14.7 ;
        RECT 21.37 13.68 21.63 13.94 ;
        RECT 21.37 12.92 21.63 13.18 ;
        RECT 21.37 12.16 21.63 12.42 ;
        RECT 21.37 11.4 21.63 11.66 ;
        RECT 22.13 18.24 22.39 18.5 ;
        RECT 22.13 17.48 22.39 17.74 ;
        RECT 22.13 16.72 22.39 16.98 ;
        RECT 22.13 15.96 22.39 16.22 ;
        RECT 22.13 15.2 22.39 15.46 ;
        RECT 22.13 14.44 22.39 14.7 ;
        RECT 22.13 13.68 22.39 13.94 ;
        RECT 22.13 12.92 22.39 13.18 ;
        RECT 22.13 12.16 22.39 12.42 ;
        RECT 22.13 11.4 22.39 11.66 ;
        RECT 22.89 18.24 23.15 18.5 ;
        RECT 22.89 17.48 23.15 17.74 ;
        RECT 22.89 16.72 23.15 16.98 ;
        RECT 22.89 15.96 23.15 16.22 ;
        RECT 22.89 15.2 23.15 15.46 ;
        RECT 22.89 14.44 23.15 14.7 ;
        RECT 22.89 13.68 23.15 13.94 ;
        RECT 22.89 12.92 23.15 13.18 ;
        RECT 22.89 12.16 23.15 12.42 ;
        RECT 22.89 11.4 23.15 11.66 ;
        RECT 23.65 18.24 23.91 18.5 ;
        RECT 23.65 17.48 23.91 17.74 ;
        RECT 23.65 16.72 23.91 16.98 ;
        RECT 23.65 15.96 23.91 16.22 ;
        RECT 23.65 15.2 23.91 15.46 ;
        RECT 23.65 14.44 23.91 14.7 ;
        RECT 23.65 13.68 23.91 13.94 ;
        RECT 23.65 12.92 23.91 13.18 ;
        RECT 23.65 12.16 23.91 12.42 ;
        RECT 23.65 11.4 23.91 11.66 ;
        RECT 24.41 18.24 24.67 18.5 ;
        RECT 24.41 17.48 24.67 17.74 ;
        RECT 24.41 16.72 24.67 16.98 ;
        RECT 24.41 15.96 24.67 16.22 ;
        RECT 24.41 15.2 24.67 15.46 ;
        RECT 24.41 14.44 24.67 14.7 ;
        RECT 24.41 13.68 24.67 13.94 ;
        RECT 24.41 12.92 24.67 13.18 ;
        RECT 24.41 12.16 24.67 12.42 ;
        RECT 24.41 11.4 24.67 11.66 ;
        RECT 25.17 18.24 25.43 18.5 ;
        RECT 25.17 17.48 25.43 17.74 ;
        RECT 25.17 16.72 25.43 16.98 ;
        RECT 25.17 15.96 25.43 16.22 ;
        RECT 25.17 15.2 25.43 15.46 ;
        RECT 25.17 14.44 25.43 14.7 ;
        RECT 25.17 13.68 25.43 13.94 ;
        RECT 25.17 12.92 25.43 13.18 ;
        RECT 25.17 12.16 25.43 12.42 ;
        RECT 25.17 11.4 25.43 11.66 ;
        RECT 25.93 18.24 26.19 18.5 ;
        RECT 25.93 17.48 26.19 17.74 ;
        RECT 25.93 16.72 26.19 16.98 ;
        RECT 25.93 15.96 26.19 16.22 ;
        RECT 25.93 15.2 26.19 15.46 ;
        RECT 25.93 14.44 26.19 14.7 ;
        RECT 25.93 13.68 26.19 13.94 ;
        RECT 25.93 12.92 26.19 13.18 ;
        RECT 25.93 12.16 26.19 12.42 ;
        RECT 25.93 11.4 26.19 11.66 ;
        RECT 26.69 18.24 26.95 18.5 ;
        RECT 26.69 17.48 26.95 17.74 ;
        RECT 26.69 16.72 26.95 16.98 ;
        RECT 26.69 15.96 26.95 16.22 ;
        RECT 26.69 15.2 26.95 15.46 ;
        RECT 26.69 14.44 26.95 14.7 ;
        RECT 26.69 13.68 26.95 13.94 ;
        RECT 26.69 12.92 26.95 13.18 ;
        RECT 26.69 12.16 26.95 12.42 ;
        RECT 26.69 11.4 26.95 11.66 ;
        RECT 27.45 18.24 27.71 18.5 ;
        RECT 27.45 17.48 27.71 17.74 ;
        RECT 27.45 16.72 27.71 16.98 ;
        RECT 27.45 15.96 27.71 16.22 ;
        RECT 27.45 15.2 27.71 15.46 ;
        RECT 27.45 14.44 27.71 14.7 ;
        RECT 27.45 13.68 27.71 13.94 ;
        RECT 27.45 12.92 27.71 13.18 ;
        RECT 27.45 12.16 27.71 12.42 ;
        RECT 27.45 11.4 27.71 11.66 ;
        RECT 28.21 18.24 28.47 18.5 ;
        RECT 28.21 17.48 28.47 17.74 ;
        RECT 28.21 16.72 28.47 16.98 ;
        RECT 28.21 15.96 28.47 16.22 ;
        RECT 28.21 15.2 28.47 15.46 ;
        RECT 28.21 14.44 28.47 14.7 ;
        RECT 28.21 13.68 28.47 13.94 ;
        RECT 28.21 12.92 28.47 13.18 ;
        RECT 28.21 12.16 28.47 12.42 ;
        RECT 28.21 11.4 28.47 11.66 ;
        RECT 28.97 18.24 29.23 18.5 ;
        RECT 28.97 17.48 29.23 17.74 ;
        RECT 28.97 16.72 29.23 16.98 ;
        RECT 28.97 15.96 29.23 16.22 ;
        RECT 28.97 15.2 29.23 15.46 ;
        RECT 28.97 14.44 29.23 14.7 ;
        RECT 28.97 13.68 29.23 13.94 ;
        RECT 28.97 12.92 29.23 13.18 ;
        RECT 28.97 12.16 29.23 12.42 ;
        RECT 28.97 11.4 29.23 11.66 ;
        RECT 29.73 18.24 29.99 18.5 ;
        RECT 29.73 17.48 29.99 17.74 ;
        RECT 29.73 16.72 29.99 16.98 ;
        RECT 29.73 15.96 29.99 16.22 ;
        RECT 29.73 15.2 29.99 15.46 ;
        RECT 29.73 14.44 29.99 14.7 ;
        RECT 29.73 13.68 29.99 13.94 ;
        RECT 29.73 12.92 29.99 13.18 ;
        RECT 29.73 12.16 29.99 12.42 ;
        RECT 29.73 11.4 29.99 11.66 ;
        RECT 30.49 18.24 30.75 18.5 ;
        RECT 30.49 17.48 30.75 17.74 ;
        RECT 30.49 16.72 30.75 16.98 ;
        RECT 30.49 15.96 30.75 16.22 ;
        RECT 30.49 15.2 30.75 15.46 ;
        RECT 30.49 14.44 30.75 14.7 ;
        RECT 30.49 13.68 30.75 13.94 ;
        RECT 30.49 12.92 30.75 13.18 ;
        RECT 30.49 12.16 30.75 12.42 ;
        RECT 30.49 11.4 30.75 11.66 ;
        RECT 31.25 18.24 31.51 18.5 ;
        RECT 31.25 17.48 31.51 17.74 ;
        RECT 31.25 16.72 31.51 16.98 ;
        RECT 31.25 15.96 31.51 16.22 ;
        RECT 31.25 15.2 31.51 15.46 ;
        RECT 31.25 14.44 31.51 14.7 ;
        RECT 31.25 13.68 31.51 13.94 ;
        RECT 31.25 12.92 31.51 13.18 ;
        RECT 31.25 12.16 31.51 12.42 ;
        RECT 31.25 11.4 31.51 11.66 ;
        RECT 32.01 18.24 32.27 18.5 ;
        RECT 32.01 17.48 32.27 17.74 ;
        RECT 32.01 16.72 32.27 16.98 ;
        RECT 32.01 15.96 32.27 16.22 ;
        RECT 32.01 15.2 32.27 15.46 ;
        RECT 32.01 14.44 32.27 14.7 ;
        RECT 32.01 13.68 32.27 13.94 ;
        RECT 32.01 12.92 32.27 13.18 ;
        RECT 32.01 12.16 32.27 12.42 ;
        RECT 32.01 11.4 32.27 11.66 ;
        RECT 32.77 18.24 33.03 18.5 ;
        RECT 32.77 17.48 33.03 17.74 ;
        RECT 32.77 16.72 33.03 16.98 ;
        RECT 32.77 15.96 33.03 16.22 ;
        RECT 32.77 15.2 33.03 15.46 ;
        RECT 32.77 14.44 33.03 14.7 ;
        RECT 32.77 13.68 33.03 13.94 ;
        RECT 32.77 12.92 33.03 13.18 ;
        RECT 32.77 12.16 33.03 12.42 ;
        RECT 32.77 11.4 33.03 11.66 ;
        RECT 33.53 18.24 33.79 18.5 ;
        RECT 33.53 17.48 33.79 17.74 ;
        RECT 33.53 16.72 33.79 16.98 ;
        RECT 33.53 15.96 33.79 16.22 ;
        RECT 33.53 15.2 33.79 15.46 ;
        RECT 33.53 14.44 33.79 14.7 ;
        RECT 33.53 13.68 33.79 13.94 ;
        RECT 33.53 12.92 33.79 13.18 ;
        RECT 33.53 12.16 33.79 12.42 ;
        RECT 33.53 11.4 33.79 11.66 ;
        RECT 34.29 18.24 34.55 18.5 ;
        RECT 34.29 17.48 34.55 17.74 ;
        RECT 34.29 16.72 34.55 16.98 ;
        RECT 34.29 15.96 34.55 16.22 ;
        RECT 34.29 15.2 34.55 15.46 ;
        RECT 34.29 14.44 34.55 14.7 ;
        RECT 34.29 13.68 34.55 13.94 ;
        RECT 34.29 12.92 34.55 13.18 ;
        RECT 34.29 12.16 34.55 12.42 ;
        RECT 34.29 11.4 34.55 11.66 ;
        RECT 35.05 18.24 35.31 18.5 ;
        RECT 35.05 17.48 35.31 17.74 ;
        RECT 35.05 16.72 35.31 16.98 ;
        RECT 35.05 15.96 35.31 16.22 ;
        RECT 35.05 15.2 35.31 15.46 ;
        RECT 35.05 14.44 35.31 14.7 ;
        RECT 35.05 13.68 35.31 13.94 ;
        RECT 35.05 12.92 35.31 13.18 ;
        RECT 35.05 12.16 35.31 12.42 ;
        RECT 35.05 11.4 35.31 11.66 ;
        RECT 35.81 18.24 36.07 18.5 ;
        RECT 35.81 17.48 36.07 17.74 ;
        RECT 35.81 16.72 36.07 16.98 ;
        RECT 35.81 15.96 36.07 16.22 ;
        RECT 35.81 15.2 36.07 15.46 ;
        RECT 35.81 14.44 36.07 14.7 ;
        RECT 35.81 13.68 36.07 13.94 ;
        RECT 35.81 12.92 36.07 13.18 ;
        RECT 35.81 12.16 36.07 12.42 ;
        RECT 35.81 11.4 36.07 11.66 ;
        RECT 36.57 18.24 36.83 18.5 ;
        RECT 36.57 17.48 36.83 17.74 ;
        RECT 36.57 16.72 36.83 16.98 ;
        RECT 36.57 15.96 36.83 16.22 ;
        RECT 36.57 15.2 36.83 15.46 ;
        RECT 36.57 14.44 36.83 14.7 ;
        RECT 36.57 13.68 36.83 13.94 ;
        RECT 36.57 12.92 36.83 13.18 ;
        RECT 36.57 12.16 36.83 12.42 ;
        RECT 36.57 11.4 36.83 11.66 ;
        RECT 37.33 18.24 37.59 18.5 ;
        RECT 37.33 17.48 37.59 17.74 ;
        RECT 37.33 16.72 37.59 16.98 ;
        RECT 37.33 15.96 37.59 16.22 ;
        RECT 37.33 15.2 37.59 15.46 ;
        RECT 37.33 14.44 37.59 14.7 ;
        RECT 37.33 13.68 37.59 13.94 ;
        RECT 37.33 12.92 37.59 13.18 ;
        RECT 37.33 12.16 37.59 12.42 ;
        RECT 37.33 11.4 37.59 11.66 ;
        RECT 38.09 18.24 38.35 18.5 ;
        RECT 38.09 17.48 38.35 17.74 ;
        RECT 38.09 16.72 38.35 16.98 ;
        RECT 38.09 15.96 38.35 16.22 ;
        RECT 38.09 15.2 38.35 15.46 ;
        RECT 38.09 14.44 38.35 14.7 ;
        RECT 38.09 13.68 38.35 13.94 ;
        RECT 38.09 12.92 38.35 13.18 ;
        RECT 38.09 12.16 38.35 12.42 ;
        RECT 38.09 11.4 38.35 11.66 ;
        RECT 38.85 18.24 39.11 18.5 ;
        RECT 38.85 17.48 39.11 17.74 ;
        RECT 38.85 16.72 39.11 16.98 ;
        RECT 38.85 15.96 39.11 16.22 ;
        RECT 38.85 15.2 39.11 15.46 ;
        RECT 38.85 14.44 39.11 14.7 ;
        RECT 38.85 13.68 39.11 13.94 ;
        RECT 38.85 12.92 39.11 13.18 ;
        RECT 38.85 12.16 39.11 12.42 ;
        RECT 38.85 11.4 39.11 11.66 ;
        RECT 39.61 18.24 39.87 18.5 ;
        RECT 39.61 17.48 39.87 17.74 ;
        RECT 39.61 16.72 39.87 16.98 ;
        RECT 39.61 15.96 39.87 16.22 ;
        RECT 39.61 15.2 39.87 15.46 ;
        RECT 39.61 14.44 39.87 14.7 ;
        RECT 39.61 13.68 39.87 13.94 ;
        RECT 39.61 12.92 39.87 13.18 ;
        RECT 39.61 12.16 39.87 12.42 ;
        RECT 39.61 11.4 39.87 11.66 ;
        RECT 40.37 18.24 40.63 18.5 ;
        RECT 40.37 17.48 40.63 17.74 ;
        RECT 40.37 16.72 40.63 16.98 ;
        RECT 40.37 15.96 40.63 16.22 ;
        RECT 40.37 15.2 40.63 15.46 ;
        RECT 40.37 14.44 40.63 14.7 ;
        RECT 40.37 13.68 40.63 13.94 ;
        RECT 40.37 12.92 40.63 13.18 ;
        RECT 40.37 12.16 40.63 12.42 ;
        RECT 40.37 11.4 40.63 11.66 ;
        RECT 41.13 18.24 41.39 18.5 ;
        RECT 41.13 17.48 41.39 17.74 ;
        RECT 41.13 16.72 41.39 16.98 ;
        RECT 41.13 15.96 41.39 16.22 ;
        RECT 41.13 15.2 41.39 15.46 ;
        RECT 41.13 14.44 41.39 14.7 ;
        RECT 41.13 13.68 41.39 13.94 ;
        RECT 41.13 12.92 41.39 13.18 ;
        RECT 41.13 12.16 41.39 12.42 ;
        RECT 41.13 11.4 41.39 11.66 ;
        RECT 41.89 18.24 42.15 18.5 ;
        RECT 41.89 17.48 42.15 17.74 ;
        RECT 41.89 16.72 42.15 16.98 ;
        RECT 41.89 15.96 42.15 16.22 ;
        RECT 41.89 15.2 42.15 15.46 ;
        RECT 41.89 14.44 42.15 14.7 ;
        RECT 41.89 13.68 42.15 13.94 ;
        RECT 41.89 12.92 42.15 13.18 ;
        RECT 41.89 12.16 42.15 12.42 ;
        RECT 41.89 11.4 42.15 11.66 ;
        RECT 42.65 18.24 42.91 18.5 ;
        RECT 42.65 17.48 42.91 17.74 ;
        RECT 42.65 16.72 42.91 16.98 ;
        RECT 42.65 15.96 42.91 16.22 ;
        RECT 42.65 15.2 42.91 15.46 ;
        RECT 42.65 14.44 42.91 14.7 ;
        RECT 42.65 13.68 42.91 13.94 ;
        RECT 42.65 12.92 42.91 13.18 ;
        RECT 42.65 12.16 42.91 12.42 ;
        RECT 42.65 11.4 42.91 11.66 ;
        RECT 43.41 18.24 43.67 18.5 ;
        RECT 43.41 17.48 43.67 17.74 ;
        RECT 43.41 16.72 43.67 16.98 ;
        RECT 43.41 15.96 43.67 16.22 ;
        RECT 43.41 15.2 43.67 15.46 ;
        RECT 43.41 14.44 43.67 14.7 ;
        RECT 43.41 13.68 43.67 13.94 ;
        RECT 43.41 12.92 43.67 13.18 ;
        RECT 43.41 12.16 43.67 12.42 ;
        RECT 43.41 11.4 43.67 11.66 ;
        RECT 44.17 18.24 44.43 18.5 ;
        RECT 44.17 17.48 44.43 17.74 ;
        RECT 44.17 16.72 44.43 16.98 ;
        RECT 44.17 15.96 44.43 16.22 ;
        RECT 44.17 15.2 44.43 15.46 ;
        RECT 44.17 14.44 44.43 14.7 ;
        RECT 44.17 13.68 44.43 13.94 ;
        RECT 44.17 12.92 44.43 13.18 ;
        RECT 44.17 12.16 44.43 12.42 ;
        RECT 44.17 11.4 44.43 11.66 ;
        RECT 44.93 18.24 45.19 18.5 ;
        RECT 44.93 17.48 45.19 17.74 ;
        RECT 44.93 16.72 45.19 16.98 ;
        RECT 44.93 15.96 45.19 16.22 ;
        RECT 44.93 15.2 45.19 15.46 ;
        RECT 44.93 14.44 45.19 14.7 ;
        RECT 44.93 13.68 45.19 13.94 ;
        RECT 44.93 12.92 45.19 13.18 ;
        RECT 44.93 12.16 45.19 12.42 ;
        RECT 44.93 11.4 45.19 11.66 ;
        RECT 45.69 18.24 45.95 18.5 ;
        RECT 45.69 17.48 45.95 17.74 ;
        RECT 45.69 16.72 45.95 16.98 ;
        RECT 45.69 15.96 45.95 16.22 ;
        RECT 45.69 15.2 45.95 15.46 ;
        RECT 45.69 14.44 45.95 14.7 ;
        RECT 45.69 13.68 45.95 13.94 ;
        RECT 45.69 12.92 45.95 13.18 ;
        RECT 45.69 12.16 45.95 12.42 ;
        RECT 45.69 11.4 45.95 11.66 ;
        RECT 46.45 18.24 46.71 18.5 ;
        RECT 46.45 17.48 46.71 17.74 ;
        RECT 46.45 16.72 46.71 16.98 ;
        RECT 46.45 15.96 46.71 16.22 ;
        RECT 46.45 15.2 46.71 15.46 ;
        RECT 46.45 14.44 46.71 14.7 ;
        RECT 46.45 13.68 46.71 13.94 ;
        RECT 46.45 12.92 46.71 13.18 ;
        RECT 46.45 12.16 46.71 12.42 ;
        RECT 46.45 11.4 46.71 11.66 ;
        RECT 47.21 18.24 47.47 18.5 ;
        RECT 47.21 17.48 47.47 17.74 ;
        RECT 47.21 16.72 47.47 16.98 ;
        RECT 47.21 15.96 47.47 16.22 ;
        RECT 47.21 15.2 47.47 15.46 ;
        RECT 47.21 14.44 47.47 14.7 ;
        RECT 47.21 13.68 47.47 13.94 ;
        RECT 47.21 12.92 47.47 13.18 ;
        RECT 47.21 12.16 47.47 12.42 ;
        RECT 47.21 11.4 47.47 11.66 ;
        RECT 47.97 18.24 48.23 18.5 ;
        RECT 47.97 17.48 48.23 17.74 ;
        RECT 47.97 16.72 48.23 16.98 ;
        RECT 47.97 15.96 48.23 16.22 ;
        RECT 47.97 15.2 48.23 15.46 ;
        RECT 47.97 14.44 48.23 14.7 ;
        RECT 47.97 13.68 48.23 13.94 ;
        RECT 47.97 12.92 48.23 13.18 ;
        RECT 47.97 12.16 48.23 12.42 ;
        RECT 47.97 11.4 48.23 11.66 ;
        RECT 48.73 18.24 48.99 18.5 ;
        RECT 48.73 17.48 48.99 17.74 ;
        RECT 48.73 16.72 48.99 16.98 ;
        RECT 48.73 15.96 48.99 16.22 ;
        RECT 48.73 15.2 48.99 15.46 ;
        RECT 48.73 14.44 48.99 14.7 ;
        RECT 48.73 13.68 48.99 13.94 ;
        RECT 48.73 12.92 48.99 13.18 ;
        RECT 48.73 12.16 48.99 12.42 ;
        RECT 48.73 11.4 48.99 11.66 ;
        RECT 49.49 18.24 49.75 18.5 ;
        RECT 49.49 17.48 49.75 17.74 ;
        RECT 49.49 16.72 49.75 16.98 ;
        RECT 49.49 15.96 49.75 16.22 ;
        RECT 49.49 15.2 49.75 15.46 ;
        RECT 49.49 14.44 49.75 14.7 ;
        RECT 49.49 13.68 49.75 13.94 ;
        RECT 49.49 12.92 49.75 13.18 ;
        RECT 49.49 12.16 49.75 12.42 ;
        RECT 49.49 11.4 49.75 11.66 ;
        RECT 50.25 18.24 50.51 18.5 ;
        RECT 50.25 17.48 50.51 17.74 ;
        RECT 50.25 16.72 50.51 16.98 ;
        RECT 50.25 15.96 50.51 16.22 ;
        RECT 50.25 15.2 50.51 15.46 ;
        RECT 50.25 14.44 50.51 14.7 ;
        RECT 50.25 13.68 50.51 13.94 ;
        RECT 50.25 12.92 50.51 13.18 ;
        RECT 50.25 12.16 50.51 12.42 ;
        RECT 50.25 11.4 50.51 11.66 ;
        RECT 51.01 18.24 51.27 18.5 ;
        RECT 51.01 17.48 51.27 17.74 ;
        RECT 51.01 16.72 51.27 16.98 ;
        RECT 51.01 15.96 51.27 16.22 ;
        RECT 51.01 15.2 51.27 15.46 ;
        RECT 51.01 14.44 51.27 14.7 ;
        RECT 51.01 13.68 51.27 13.94 ;
        RECT 51.01 12.92 51.27 13.18 ;
        RECT 51.01 12.16 51.27 12.42 ;
        RECT 51.01 11.4 51.27 11.66 ;
        RECT 51.77 18.24 52.03 18.5 ;
        RECT 51.77 17.48 52.03 17.74 ;
        RECT 51.77 16.72 52.03 16.98 ;
        RECT 51.77 15.96 52.03 16.22 ;
        RECT 51.77 15.2 52.03 15.46 ;
        RECT 51.77 14.44 52.03 14.7 ;
        RECT 51.77 13.68 52.03 13.94 ;
        RECT 51.77 12.92 52.03 13.18 ;
        RECT 51.77 12.16 52.03 12.42 ;
        RECT 51.77 11.4 52.03 11.66 ;
        RECT 52.53 18.24 52.79 18.5 ;
        RECT 52.53 17.48 52.79 17.74 ;
        RECT 52.53 16.72 52.79 16.98 ;
        RECT 52.53 15.96 52.79 16.22 ;
        RECT 52.53 15.2 52.79 15.46 ;
        RECT 52.53 14.44 52.79 14.7 ;
        RECT 52.53 13.68 52.79 13.94 ;
        RECT 52.53 12.92 52.79 13.18 ;
        RECT 52.53 12.16 52.79 12.42 ;
        RECT 52.53 11.4 52.79 11.66 ;
        RECT 53.29 18.24 53.55 18.5 ;
        RECT 53.29 17.48 53.55 17.74 ;
        RECT 53.29 16.72 53.55 16.98 ;
        RECT 53.29 15.96 53.55 16.22 ;
        RECT 53.29 15.2 53.55 15.46 ;
        RECT 53.29 14.44 53.55 14.7 ;
        RECT 53.29 13.68 53.55 13.94 ;
        RECT 53.29 12.92 53.55 13.18 ;
        RECT 53.29 12.16 53.55 12.42 ;
        RECT 53.29 11.4 53.55 11.66 ;
        RECT 54.05 18.24 54.31 18.5 ;
        RECT 54.05 17.48 54.31 17.74 ;
        RECT 54.05 16.72 54.31 16.98 ;
        RECT 54.05 15.96 54.31 16.22 ;
        RECT 54.05 15.2 54.31 15.46 ;
        RECT 54.05 14.44 54.31 14.7 ;
        RECT 54.05 13.68 54.31 13.94 ;
        RECT 54.05 12.92 54.31 13.18 ;
        RECT 54.05 12.16 54.31 12.42 ;
        RECT 54.05 11.4 54.31 11.66 ;
        RECT 54.81 18.24 55.07 18.5 ;
        RECT 54.81 17.48 55.07 17.74 ;
        RECT 54.81 16.72 55.07 16.98 ;
        RECT 54.81 15.96 55.07 16.22 ;
        RECT 54.81 15.2 55.07 15.46 ;
        RECT 54.81 14.44 55.07 14.7 ;
        RECT 54.81 13.68 55.07 13.94 ;
        RECT 54.81 12.92 55.07 13.18 ;
        RECT 54.81 12.16 55.07 12.42 ;
        RECT 54.81 11.4 55.07 11.66 ;
        RECT 55.57 18.24 55.83 18.5 ;
        RECT 55.57 17.48 55.83 17.74 ;
        RECT 55.57 16.72 55.83 16.98 ;
        RECT 55.57 15.96 55.83 16.22 ;
        RECT 55.57 15.2 55.83 15.46 ;
        RECT 55.57 14.44 55.83 14.7 ;
        RECT 55.57 13.68 55.83 13.94 ;
        RECT 55.57 12.92 55.83 13.18 ;
        RECT 55.57 12.16 55.83 12.42 ;
        RECT 55.57 11.4 55.83 11.66 ;
        RECT 56.33 18.24 56.59 18.5 ;
        RECT 56.33 17.48 56.59 17.74 ;
        RECT 56.33 16.72 56.59 16.98 ;
        RECT 56.33 15.96 56.59 16.22 ;
        RECT 56.33 15.2 56.59 15.46 ;
        RECT 56.33 14.44 56.59 14.7 ;
        RECT 56.33 13.68 56.59 13.94 ;
        RECT 56.33 12.92 56.59 13.18 ;
        RECT 56.33 12.16 56.59 12.42 ;
        RECT 56.33 11.4 56.59 11.66 ;
        RECT 57.09 18.24 57.35 18.5 ;
        RECT 57.09 17.48 57.35 17.74 ;
        RECT 57.09 16.72 57.35 16.98 ;
        RECT 57.09 15.96 57.35 16.22 ;
        RECT 57.09 15.2 57.35 15.46 ;
        RECT 57.09 14.44 57.35 14.7 ;
        RECT 57.09 13.68 57.35 13.94 ;
        RECT 57.09 12.92 57.35 13.18 ;
        RECT 57.09 12.16 57.35 12.42 ;
        RECT 57.09 11.4 57.35 11.66 ;
        RECT 57.85 18.24 58.11 18.5 ;
        RECT 57.85 17.48 58.11 17.74 ;
        RECT 57.85 16.72 58.11 16.98 ;
        RECT 57.85 15.96 58.11 16.22 ;
        RECT 57.85 15.2 58.11 15.46 ;
        RECT 57.85 14.44 58.11 14.7 ;
        RECT 57.85 13.68 58.11 13.94 ;
        RECT 57.85 12.92 58.11 13.18 ;
        RECT 57.85 12.16 58.11 12.42 ;
        RECT 57.85 11.4 58.11 11.66 ;
        RECT 58.61 18.24 58.87 18.5 ;
        RECT 58.61 17.48 58.87 17.74 ;
        RECT 58.61 16.72 58.87 16.98 ;
        RECT 58.61 15.96 58.87 16.22 ;
        RECT 58.61 15.2 58.87 15.46 ;
        RECT 58.61 14.44 58.87 14.7 ;
        RECT 58.61 13.68 58.87 13.94 ;
        RECT 58.61 12.92 58.87 13.18 ;
        RECT 58.61 12.16 58.87 12.42 ;
        RECT 58.61 11.4 58.87 11.66 ;
        RECT 59.37 18.24 59.63 18.5 ;
        RECT 59.37 17.48 59.63 17.74 ;
        RECT 59.37 16.72 59.63 16.98 ;
        RECT 59.37 15.96 59.63 16.22 ;
        RECT 59.37 15.2 59.63 15.46 ;
        RECT 59.37 14.44 59.63 14.7 ;
        RECT 59.37 13.68 59.63 13.94 ;
        RECT 59.37 12.92 59.63 13.18 ;
        RECT 59.37 12.16 59.63 12.42 ;
        RECT 59.37 11.4 59.63 11.66 ;
        RECT 60.13 18.24 60.39 18.5 ;
        RECT 60.13 17.48 60.39 17.74 ;
        RECT 60.13 16.72 60.39 16.98 ;
        RECT 60.13 15.96 60.39 16.22 ;
        RECT 60.13 15.2 60.39 15.46 ;
        RECT 60.13 14.44 60.39 14.7 ;
        RECT 60.13 13.68 60.39 13.94 ;
        RECT 60.13 12.92 60.39 13.18 ;
        RECT 60.13 12.16 60.39 12.42 ;
        RECT 60.13 11.4 60.39 11.66 ;
        RECT 60.89 18.24 61.15 18.5 ;
        RECT 60.89 17.48 61.15 17.74 ;
        RECT 60.89 16.72 61.15 16.98 ;
        RECT 60.89 15.96 61.15 16.22 ;
        RECT 60.89 15.2 61.15 15.46 ;
        RECT 60.89 14.44 61.15 14.7 ;
        RECT 60.89 13.68 61.15 13.94 ;
        RECT 60.89 12.92 61.15 13.18 ;
        RECT 60.89 12.16 61.15 12.42 ;
        RECT 60.89 11.4 61.15 11.66 ;
        RECT 61.65 18.24 61.91 18.5 ;
        RECT 61.65 17.48 61.91 17.74 ;
        RECT 61.65 16.72 61.91 16.98 ;
        RECT 61.65 15.96 61.91 16.22 ;
        RECT 61.65 15.2 61.91 15.46 ;
        RECT 61.65 14.44 61.91 14.7 ;
        RECT 61.65 13.68 61.91 13.94 ;
        RECT 61.65 12.92 61.91 13.18 ;
        RECT 61.65 12.16 61.91 12.42 ;
        RECT 61.65 11.4 61.91 11.66 ;
        RECT 62.41 18.24 62.67 18.5 ;
        RECT 62.41 17.48 62.67 17.74 ;
        RECT 62.41 16.72 62.67 16.98 ;
        RECT 62.41 15.96 62.67 16.22 ;
        RECT 62.41 15.2 62.67 15.46 ;
        RECT 62.41 14.44 62.67 14.7 ;
        RECT 62.41 13.68 62.67 13.94 ;
        RECT 62.41 12.92 62.67 13.18 ;
        RECT 62.41 12.16 62.67 12.42 ;
        RECT 62.41 11.4 62.67 11.66 ;
        RECT 63.17 18.24 63.43 18.5 ;
        RECT 63.17 17.48 63.43 17.74 ;
        RECT 63.17 16.72 63.43 16.98 ;
        RECT 63.17 15.96 63.43 16.22 ;
        RECT 63.17 15.2 63.43 15.46 ;
        RECT 63.17 14.44 63.43 14.7 ;
        RECT 63.17 13.68 63.43 13.94 ;
        RECT 63.17 12.92 63.43 13.18 ;
        RECT 63.17 12.16 63.43 12.42 ;
        RECT 63.17 11.4 63.43 11.66 ;
        RECT 63.93 18.24 64.19 18.5 ;
        RECT 63.93 17.48 64.19 17.74 ;
        RECT 63.93 16.72 64.19 16.98 ;
        RECT 63.93 15.96 64.19 16.22 ;
        RECT 63.93 15.2 64.19 15.46 ;
        RECT 63.93 14.44 64.19 14.7 ;
        RECT 63.93 13.68 64.19 13.94 ;
        RECT 63.93 12.92 64.19 13.18 ;
        RECT 63.93 12.16 64.19 12.42 ;
        RECT 63.93 11.4 64.19 11.66 ;
        RECT 64.69 18.24 64.95 18.5 ;
        RECT 64.69 17.48 64.95 17.74 ;
        RECT 64.69 16.72 64.95 16.98 ;
        RECT 64.69 15.96 64.95 16.22 ;
        RECT 64.69 15.2 64.95 15.46 ;
        RECT 64.69 14.44 64.95 14.7 ;
        RECT 64.69 13.68 64.95 13.94 ;
        RECT 64.69 12.92 64.95 13.18 ;
        RECT 64.69 12.16 64.95 12.42 ;
        RECT 64.69 11.4 64.95 11.66 ;
        RECT 65.45 18.24 65.71 18.5 ;
        RECT 65.45 17.48 65.71 17.74 ;
        RECT 65.45 16.72 65.71 16.98 ;
        RECT 65.45 15.96 65.71 16.22 ;
        RECT 65.45 15.2 65.71 15.46 ;
        RECT 65.45 14.44 65.71 14.7 ;
        RECT 65.45 13.68 65.71 13.94 ;
        RECT 65.45 12.92 65.71 13.18 ;
        RECT 65.45 12.16 65.71 12.42 ;
        RECT 65.45 11.4 65.71 11.66 ;
        RECT 66.21 18.24 66.47 18.5 ;
        RECT 66.21 17.48 66.47 17.74 ;
        RECT 66.21 16.72 66.47 16.98 ;
        RECT 66.21 15.96 66.47 16.22 ;
        RECT 66.21 15.2 66.47 15.46 ;
        RECT 66.21 14.44 66.47 14.7 ;
        RECT 66.21 13.68 66.47 13.94 ;
        RECT 66.21 12.92 66.47 13.18 ;
        RECT 66.21 12.16 66.47 12.42 ;
        RECT 66.21 11.4 66.47 11.66 ;
        RECT 66.97 18.24 67.23 18.5 ;
        RECT 66.97 17.48 67.23 17.74 ;
        RECT 66.97 16.72 67.23 16.98 ;
        RECT 66.97 15.96 67.23 16.22 ;
        RECT 66.97 15.2 67.23 15.46 ;
        RECT 66.97 14.44 67.23 14.7 ;
        RECT 66.97 13.68 67.23 13.94 ;
        RECT 66.97 12.92 67.23 13.18 ;
        RECT 66.97 12.16 67.23 12.42 ;
        RECT 66.97 11.4 67.23 11.66 ;
        RECT 67.73 18.24 67.99 18.5 ;
        RECT 67.73 17.48 67.99 17.74 ;
        RECT 67.73 16.72 67.99 16.98 ;
        RECT 67.73 15.96 67.99 16.22 ;
        RECT 67.73 15.2 67.99 15.46 ;
        RECT 67.73 14.44 67.99 14.7 ;
        RECT 67.73 13.68 67.99 13.94 ;
        RECT 67.73 12.92 67.99 13.18 ;
        RECT 67.73 12.16 67.99 12.42 ;
        RECT 67.73 11.4 67.99 11.66 ;
        RECT 68.49 18.24 68.75 18.5 ;
        RECT 68.49 17.48 68.75 17.74 ;
        RECT 68.49 16.72 68.75 16.98 ;
        RECT 68.49 15.96 68.75 16.22 ;
        RECT 68.49 15.2 68.75 15.46 ;
        RECT 68.49 14.44 68.75 14.7 ;
        RECT 68.49 13.68 68.75 13.94 ;
        RECT 68.49 12.92 68.75 13.18 ;
        RECT 68.49 12.16 68.75 12.42 ;
        RECT 68.49 11.4 68.75 11.66 ;
        RECT 69.25 18.24 69.51 18.5 ;
        RECT 69.25 17.48 69.51 17.74 ;
        RECT 69.25 16.72 69.51 16.98 ;
        RECT 69.25 15.96 69.51 16.22 ;
        RECT 69.25 15.2 69.51 15.46 ;
        RECT 69.25 14.44 69.51 14.7 ;
        RECT 69.25 13.68 69.51 13.94 ;
        RECT 69.25 12.92 69.51 13.18 ;
        RECT 69.25 12.16 69.51 12.42 ;
        RECT 69.25 11.4 69.51 11.66 ;
        RECT 70.01 18.24 70.27 18.5 ;
        RECT 70.01 17.48 70.27 17.74 ;
        RECT 70.01 16.72 70.27 16.98 ;
        RECT 70.01 15.96 70.27 16.22 ;
        RECT 70.01 15.2 70.27 15.46 ;
        RECT 70.01 14.44 70.27 14.7 ;
        RECT 70.01 13.68 70.27 13.94 ;
        RECT 70.01 12.92 70.27 13.18 ;
        RECT 70.01 12.16 70.27 12.42 ;
        RECT 70.01 11.4 70.27 11.66 ;
        RECT 70.77 18.24 71.03 18.5 ;
        RECT 70.77 17.48 71.03 17.74 ;
        RECT 70.77 16.72 71.03 16.98 ;
        RECT 70.77 15.96 71.03 16.22 ;
        RECT 70.77 15.2 71.03 15.46 ;
        RECT 70.77 14.44 71.03 14.7 ;
        RECT 70.77 13.68 71.03 13.94 ;
        RECT 70.77 12.92 71.03 13.18 ;
        RECT 70.77 12.16 71.03 12.42 ;
        RECT 70.77 11.4 71.03 11.66 ;
        RECT 71.53 18.24 71.79 18.5 ;
        RECT 71.53 17.48 71.79 17.74 ;
        RECT 71.53 16.72 71.79 16.98 ;
        RECT 71.53 15.96 71.79 16.22 ;
        RECT 71.53 15.2 71.79 15.46 ;
        RECT 71.53 14.44 71.79 14.7 ;
        RECT 71.53 13.68 71.79 13.94 ;
        RECT 71.53 12.92 71.79 13.18 ;
        RECT 71.53 12.16 71.79 12.42 ;
        RECT 71.53 11.4 71.79 11.66 ;
        RECT 72.29 18.24 72.55 18.5 ;
        RECT 72.29 17.48 72.55 17.74 ;
        RECT 72.29 16.72 72.55 16.98 ;
        RECT 72.29 15.96 72.55 16.22 ;
        RECT 72.29 15.2 72.55 15.46 ;
        RECT 72.29 14.44 72.55 14.7 ;
        RECT 72.29 13.68 72.55 13.94 ;
        RECT 72.29 12.92 72.55 13.18 ;
        RECT 72.29 12.16 72.55 12.42 ;
        RECT 72.29 11.4 72.55 11.66 ;
        RECT 73.05 18.24 73.31 18.5 ;
        RECT 73.05 17.48 73.31 17.74 ;
        RECT 73.05 16.72 73.31 16.98 ;
        RECT 73.05 15.96 73.31 16.22 ;
        RECT 73.05 15.2 73.31 15.46 ;
        RECT 73.05 14.44 73.31 14.7 ;
        RECT 73.05 13.68 73.31 13.94 ;
        RECT 73.05 12.92 73.31 13.18 ;
        RECT 73.05 12.16 73.31 12.42 ;
        RECT 73.05 11.4 73.31 11.66 ;
        RECT 73.81 18.24 74.07 18.5 ;
        RECT 73.81 17.48 74.07 17.74 ;
        RECT 73.81 16.72 74.07 16.98 ;
        RECT 73.81 15.96 74.07 16.22 ;
        RECT 73.81 15.2 74.07 15.46 ;
        RECT 73.81 14.44 74.07 14.7 ;
        RECT 73.81 13.68 74.07 13.94 ;
        RECT 73.81 12.92 74.07 13.18 ;
        RECT 73.81 12.16 74.07 12.42 ;
        RECT 73.81 11.4 74.07 11.66 ;
        RECT 74.57 18.24 74.83 18.5 ;
        RECT 74.57 17.48 74.83 17.74 ;
        RECT 74.57 16.72 74.83 16.98 ;
        RECT 74.57 15.96 74.83 16.22 ;
        RECT 74.57 15.2 74.83 15.46 ;
        RECT 74.57 14.44 74.83 14.7 ;
        RECT 74.57 13.68 74.83 13.94 ;
        RECT 74.57 12.92 74.83 13.18 ;
        RECT 74.57 12.16 74.83 12.42 ;
        RECT 74.57 11.4 74.83 11.66 ;
        RECT 75.33 18.24 75.59 18.5 ;
        RECT 75.33 17.48 75.59 17.74 ;
        RECT 75.33 16.72 75.59 16.98 ;
        RECT 75.33 15.96 75.59 16.22 ;
        RECT 75.33 15.2 75.59 15.46 ;
        RECT 75.33 14.44 75.59 14.7 ;
        RECT 75.33 13.68 75.59 13.94 ;
        RECT 75.33 12.92 75.59 13.18 ;
        RECT 75.33 12.16 75.59 12.42 ;
        RECT 75.33 11.4 75.59 11.66 ;
        RECT 76.09 18.24 76.35 18.5 ;
        RECT 76.09 17.48 76.35 17.74 ;
        RECT 76.09 16.72 76.35 16.98 ;
        RECT 76.09 15.96 76.35 16.22 ;
        RECT 76.09 15.2 76.35 15.46 ;
        RECT 76.09 14.44 76.35 14.7 ;
        RECT 76.09 13.68 76.35 13.94 ;
        RECT 76.09 12.92 76.35 13.18 ;
        RECT 76.09 12.16 76.35 12.42 ;
        RECT 76.09 11.4 76.35 11.66 ;
        RECT 76.85 18.24 77.11 18.5 ;
        RECT 76.85 17.48 77.11 17.74 ;
        RECT 76.85 16.72 77.11 16.98 ;
        RECT 76.85 15.96 77.11 16.22 ;
        RECT 76.85 15.2 77.11 15.46 ;
        RECT 76.85 14.44 77.11 14.7 ;
        RECT 76.85 13.68 77.11 13.94 ;
        RECT 76.85 12.92 77.11 13.18 ;
        RECT 76.85 12.16 77.11 12.42 ;
        RECT 76.85 11.4 77.11 11.66 ;
        RECT 77.61 18.24 77.87 18.5 ;
        RECT 77.61 17.48 77.87 17.74 ;
        RECT 77.61 16.72 77.87 16.98 ;
        RECT 77.61 15.96 77.87 16.22 ;
        RECT 77.61 15.2 77.87 15.46 ;
        RECT 77.61 14.44 77.87 14.7 ;
        RECT 77.61 13.68 77.87 13.94 ;
        RECT 77.61 12.92 77.87 13.18 ;
        RECT 77.61 12.16 77.87 12.42 ;
        RECT 77.61 11.4 77.87 11.66 ;
        RECT 78.37 18.24 78.63 18.5 ;
        RECT 78.37 17.48 78.63 17.74 ;
        RECT 78.37 16.72 78.63 16.98 ;
        RECT 78.37 15.96 78.63 16.22 ;
        RECT 78.37 15.2 78.63 15.46 ;
        RECT 78.37 14.44 78.63 14.7 ;
        RECT 78.37 13.68 78.63 13.94 ;
        RECT 78.37 12.92 78.63 13.18 ;
        RECT 78.37 12.16 78.63 12.42 ;
        RECT 78.37 11.4 78.63 11.66 ;
        RECT 79.13 18.24 79.39 18.5 ;
        RECT 79.13 17.48 79.39 17.74 ;
        RECT 79.13 16.72 79.39 16.98 ;
        RECT 79.13 15.96 79.39 16.22 ;
        RECT 79.13 15.2 79.39 15.46 ;
        RECT 79.13 14.44 79.39 14.7 ;
        RECT 79.13 13.68 79.39 13.94 ;
        RECT 79.13 12.92 79.39 13.18 ;
        RECT 79.13 12.16 79.39 12.42 ;
        RECT 79.13 11.4 79.39 11.66 ;
        RECT 79.89 18.24 80.15 18.5 ;
        RECT 79.89 17.48 80.15 17.74 ;
        RECT 79.89 16.72 80.15 16.98 ;
        RECT 79.89 15.96 80.15 16.22 ;
        RECT 79.89 15.2 80.15 15.46 ;
        RECT 79.89 14.44 80.15 14.7 ;
        RECT 79.89 13.68 80.15 13.94 ;
        RECT 79.89 12.92 80.15 13.18 ;
        RECT 79.89 12.16 80.15 12.42 ;
        RECT 79.89 11.4 80.15 11.66 ;
    END
  END AVDD
  PIN SUB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M3 ;
        RECT 0 4 100 8 ;
      LAYER M4 ;
        RECT 0 4 100 8 ;
      LAYER V4 ;
        RECT 4.65 6.59 4.91 6.85 ;
        RECT 4.65 5.83 4.91 6.09 ;
        RECT 4.65 5.07 4.91 5.33 ;
        RECT 5.41 6.59 5.67 6.85 ;
        RECT 5.41 5.83 5.67 6.09 ;
        RECT 5.41 5.07 5.67 5.33 ;
        RECT 6.17 6.59 6.43 6.85 ;
        RECT 6.17 5.83 6.43 6.09 ;
        RECT 6.17 5.07 6.43 5.33 ;
        RECT 6.93 6.59 7.19 6.85 ;
        RECT 6.93 5.83 7.19 6.09 ;
        RECT 6.93 5.07 7.19 5.33 ;
        RECT 7.69 6.59 7.95 6.85 ;
        RECT 7.69 5.83 7.95 6.09 ;
        RECT 7.69 5.07 7.95 5.33 ;
        RECT 8.45 6.59 8.71 6.85 ;
        RECT 8.45 5.83 8.71 6.09 ;
        RECT 8.45 5.07 8.71 5.33 ;
        RECT 9.21 6.59 9.47 6.85 ;
        RECT 9.21 5.83 9.47 6.09 ;
        RECT 9.21 5.07 9.47 5.33 ;
        RECT 9.97 6.59 10.23 6.85 ;
        RECT 9.97 5.83 10.23 6.09 ;
        RECT 9.97 5.07 10.23 5.33 ;
        RECT 10.73 6.59 10.99 6.85 ;
        RECT 10.73 5.83 10.99 6.09 ;
        RECT 10.73 5.07 10.99 5.33 ;
        RECT 11.49 6.59 11.75 6.85 ;
        RECT 11.49 5.83 11.75 6.09 ;
        RECT 11.49 5.07 11.75 5.33 ;
        RECT 12.25 6.59 12.51 6.85 ;
        RECT 12.25 5.83 12.51 6.09 ;
        RECT 12.25 5.07 12.51 5.33 ;
        RECT 13.01 6.59 13.27 6.85 ;
        RECT 13.01 5.83 13.27 6.09 ;
        RECT 13.01 5.07 13.27 5.33 ;
        RECT 13.77 6.59 14.03 6.85 ;
        RECT 13.77 5.83 14.03 6.09 ;
        RECT 13.77 5.07 14.03 5.33 ;
        RECT 14.53 6.59 14.79 6.85 ;
        RECT 14.53 5.83 14.79 6.09 ;
        RECT 14.53 5.07 14.79 5.33 ;
        RECT 15.29 6.59 15.55 6.85 ;
        RECT 15.29 5.83 15.55 6.09 ;
        RECT 15.29 5.07 15.55 5.33 ;
        RECT 16.05 6.59 16.31 6.85 ;
        RECT 16.05 5.83 16.31 6.09 ;
        RECT 16.05 5.07 16.31 5.33 ;
        RECT 16.81 6.59 17.07 6.85 ;
        RECT 16.81 5.83 17.07 6.09 ;
        RECT 16.81 5.07 17.07 5.33 ;
        RECT 17.57 6.59 17.83 6.85 ;
        RECT 17.57 5.83 17.83 6.09 ;
        RECT 17.57 5.07 17.83 5.33 ;
        RECT 18.33 6.59 18.59 6.85 ;
        RECT 18.33 5.83 18.59 6.09 ;
        RECT 18.33 5.07 18.59 5.33 ;
        RECT 19.09 6.59 19.35 6.85 ;
        RECT 19.09 5.83 19.35 6.09 ;
        RECT 19.09 5.07 19.35 5.33 ;
        RECT 19.85 6.59 20.11 6.85 ;
        RECT 19.85 5.83 20.11 6.09 ;
        RECT 19.85 5.07 20.11 5.33 ;
        RECT 20.61 6.59 20.87 6.85 ;
        RECT 20.61 5.83 20.87 6.09 ;
        RECT 20.61 5.07 20.87 5.33 ;
        RECT 21.37 6.59 21.63 6.85 ;
        RECT 21.37 5.83 21.63 6.09 ;
        RECT 21.37 5.07 21.63 5.33 ;
        RECT 22.13 6.59 22.39 6.85 ;
        RECT 22.13 5.83 22.39 6.09 ;
        RECT 22.13 5.07 22.39 5.33 ;
        RECT 22.89 6.59 23.15 6.85 ;
        RECT 22.89 5.83 23.15 6.09 ;
        RECT 22.89 5.07 23.15 5.33 ;
        RECT 23.65 6.59 23.91 6.85 ;
        RECT 23.65 5.83 23.91 6.09 ;
        RECT 23.65 5.07 23.91 5.33 ;
        RECT 24.41 6.59 24.67 6.85 ;
        RECT 24.41 5.83 24.67 6.09 ;
        RECT 24.41 5.07 24.67 5.33 ;
        RECT 25.17 6.59 25.43 6.85 ;
        RECT 25.17 5.83 25.43 6.09 ;
        RECT 25.17 5.07 25.43 5.33 ;
        RECT 25.93 6.59 26.19 6.85 ;
        RECT 25.93 5.83 26.19 6.09 ;
        RECT 25.93 5.07 26.19 5.33 ;
        RECT 26.69 6.59 26.95 6.85 ;
        RECT 26.69 5.83 26.95 6.09 ;
        RECT 26.69 5.07 26.95 5.33 ;
        RECT 27.45 6.59 27.71 6.85 ;
        RECT 27.45 5.83 27.71 6.09 ;
        RECT 27.45 5.07 27.71 5.33 ;
        RECT 28.21 6.59 28.47 6.85 ;
        RECT 28.21 5.83 28.47 6.09 ;
        RECT 28.21 5.07 28.47 5.33 ;
        RECT 28.97 6.59 29.23 6.85 ;
        RECT 28.97 5.83 29.23 6.09 ;
        RECT 28.97 5.07 29.23 5.33 ;
        RECT 29.73 6.59 29.99 6.85 ;
        RECT 29.73 5.83 29.99 6.09 ;
        RECT 29.73 5.07 29.99 5.33 ;
        RECT 30.49 6.59 30.75 6.85 ;
        RECT 30.49 5.83 30.75 6.09 ;
        RECT 30.49 5.07 30.75 5.33 ;
        RECT 31.25 6.59 31.51 6.85 ;
        RECT 31.25 5.83 31.51 6.09 ;
        RECT 31.25 5.07 31.51 5.33 ;
        RECT 32.01 6.59 32.27 6.85 ;
        RECT 32.01 5.83 32.27 6.09 ;
        RECT 32.01 5.07 32.27 5.33 ;
        RECT 32.77 6.59 33.03 6.85 ;
        RECT 32.77 5.83 33.03 6.09 ;
        RECT 32.77 5.07 33.03 5.33 ;
        RECT 33.53 6.59 33.79 6.85 ;
        RECT 33.53 5.83 33.79 6.09 ;
        RECT 33.53 5.07 33.79 5.33 ;
        RECT 34.29 6.59 34.55 6.85 ;
        RECT 34.29 5.83 34.55 6.09 ;
        RECT 34.29 5.07 34.55 5.33 ;
        RECT 35.05 6.59 35.31 6.85 ;
        RECT 35.05 5.83 35.31 6.09 ;
        RECT 35.05 5.07 35.31 5.33 ;
        RECT 35.81 6.59 36.07 6.85 ;
        RECT 35.81 5.83 36.07 6.09 ;
        RECT 35.81 5.07 36.07 5.33 ;
        RECT 36.57 6.59 36.83 6.85 ;
        RECT 36.57 5.83 36.83 6.09 ;
        RECT 36.57 5.07 36.83 5.33 ;
        RECT 37.33 6.59 37.59 6.85 ;
        RECT 37.33 5.83 37.59 6.09 ;
        RECT 37.33 5.07 37.59 5.33 ;
        RECT 38.09 6.59 38.35 6.85 ;
        RECT 38.09 5.83 38.35 6.09 ;
        RECT 38.09 5.07 38.35 5.33 ;
        RECT 38.85 6.59 39.11 6.85 ;
        RECT 38.85 5.83 39.11 6.09 ;
        RECT 38.85 5.07 39.11 5.33 ;
        RECT 39.61 6.59 39.87 6.85 ;
        RECT 39.61 5.83 39.87 6.09 ;
        RECT 39.61 5.07 39.87 5.33 ;
        RECT 40.37 6.59 40.63 6.85 ;
        RECT 40.37 5.83 40.63 6.09 ;
        RECT 40.37 5.07 40.63 5.33 ;
        RECT 41.13 6.59 41.39 6.85 ;
        RECT 41.13 5.83 41.39 6.09 ;
        RECT 41.13 5.07 41.39 5.33 ;
        RECT 41.89 6.59 42.15 6.85 ;
        RECT 41.89 5.83 42.15 6.09 ;
        RECT 41.89 5.07 42.15 5.33 ;
        RECT 42.65 6.59 42.91 6.85 ;
        RECT 42.65 5.83 42.91 6.09 ;
        RECT 42.65 5.07 42.91 5.33 ;
        RECT 43.41 6.59 43.67 6.85 ;
        RECT 43.41 5.83 43.67 6.09 ;
        RECT 43.41 5.07 43.67 5.33 ;
        RECT 44.17 6.59 44.43 6.85 ;
        RECT 44.17 5.83 44.43 6.09 ;
        RECT 44.17 5.07 44.43 5.33 ;
        RECT 44.93 6.59 45.19 6.85 ;
        RECT 44.93 5.83 45.19 6.09 ;
        RECT 44.93 5.07 45.19 5.33 ;
        RECT 45.69 6.59 45.95 6.85 ;
        RECT 45.69 5.83 45.95 6.09 ;
        RECT 45.69 5.07 45.95 5.33 ;
        RECT 46.45 6.59 46.71 6.85 ;
        RECT 46.45 5.83 46.71 6.09 ;
        RECT 46.45 5.07 46.71 5.33 ;
        RECT 47.21 6.59 47.47 6.85 ;
        RECT 47.21 5.83 47.47 6.09 ;
        RECT 47.21 5.07 47.47 5.33 ;
        RECT 47.97 6.59 48.23 6.85 ;
        RECT 47.97 5.83 48.23 6.09 ;
        RECT 47.97 5.07 48.23 5.33 ;
        RECT 48.73 6.59 48.99 6.85 ;
        RECT 48.73 5.83 48.99 6.09 ;
        RECT 48.73 5.07 48.99 5.33 ;
        RECT 49.49 6.59 49.75 6.85 ;
        RECT 49.49 5.83 49.75 6.09 ;
        RECT 49.49 5.07 49.75 5.33 ;
        RECT 50.25 6.59 50.51 6.85 ;
        RECT 50.25 5.83 50.51 6.09 ;
        RECT 50.25 5.07 50.51 5.33 ;
        RECT 51.01 6.59 51.27 6.85 ;
        RECT 51.01 5.83 51.27 6.09 ;
        RECT 51.01 5.07 51.27 5.33 ;
        RECT 51.77 6.59 52.03 6.85 ;
        RECT 51.77 5.83 52.03 6.09 ;
        RECT 51.77 5.07 52.03 5.33 ;
        RECT 52.53 6.59 52.79 6.85 ;
        RECT 52.53 5.83 52.79 6.09 ;
        RECT 52.53 5.07 52.79 5.33 ;
        RECT 53.29 6.59 53.55 6.85 ;
        RECT 53.29 5.83 53.55 6.09 ;
        RECT 53.29 5.07 53.55 5.33 ;
        RECT 54.05 6.59 54.31 6.85 ;
        RECT 54.05 5.83 54.31 6.09 ;
        RECT 54.05 5.07 54.31 5.33 ;
        RECT 54.81 6.59 55.07 6.85 ;
        RECT 54.81 5.83 55.07 6.09 ;
        RECT 54.81 5.07 55.07 5.33 ;
        RECT 55.57 6.59 55.83 6.85 ;
        RECT 55.57 5.83 55.83 6.09 ;
        RECT 55.57 5.07 55.83 5.33 ;
        RECT 56.33 6.59 56.59 6.85 ;
        RECT 56.33 5.83 56.59 6.09 ;
        RECT 56.33 5.07 56.59 5.33 ;
        RECT 57.09 6.59 57.35 6.85 ;
        RECT 57.09 5.83 57.35 6.09 ;
        RECT 57.09 5.07 57.35 5.33 ;
        RECT 57.85 6.59 58.11 6.85 ;
        RECT 57.85 5.83 58.11 6.09 ;
        RECT 57.85 5.07 58.11 5.33 ;
        RECT 58.61 6.59 58.87 6.85 ;
        RECT 58.61 5.83 58.87 6.09 ;
        RECT 58.61 5.07 58.87 5.33 ;
        RECT 59.37 6.59 59.63 6.85 ;
        RECT 59.37 5.83 59.63 6.09 ;
        RECT 59.37 5.07 59.63 5.33 ;
        RECT 60.13 6.59 60.39 6.85 ;
        RECT 60.13 5.83 60.39 6.09 ;
        RECT 60.13 5.07 60.39 5.33 ;
        RECT 60.89 6.59 61.15 6.85 ;
        RECT 60.89 5.83 61.15 6.09 ;
        RECT 60.89 5.07 61.15 5.33 ;
        RECT 61.65 6.59 61.91 6.85 ;
        RECT 61.65 5.83 61.91 6.09 ;
        RECT 61.65 5.07 61.91 5.33 ;
        RECT 62.41 6.59 62.67 6.85 ;
        RECT 62.41 5.83 62.67 6.09 ;
        RECT 62.41 5.07 62.67 5.33 ;
        RECT 63.17 6.59 63.43 6.85 ;
        RECT 63.17 5.83 63.43 6.09 ;
        RECT 63.17 5.07 63.43 5.33 ;
        RECT 63.93 6.59 64.19 6.85 ;
        RECT 63.93 5.83 64.19 6.09 ;
        RECT 63.93 5.07 64.19 5.33 ;
        RECT 64.69 6.59 64.95 6.85 ;
        RECT 64.69 5.83 64.95 6.09 ;
        RECT 64.69 5.07 64.95 5.33 ;
        RECT 65.45 6.59 65.71 6.85 ;
        RECT 65.45 5.83 65.71 6.09 ;
        RECT 65.45 5.07 65.71 5.33 ;
        RECT 66.21 6.59 66.47 6.85 ;
        RECT 66.21 5.83 66.47 6.09 ;
        RECT 66.21 5.07 66.47 5.33 ;
        RECT 66.97 6.59 67.23 6.85 ;
        RECT 66.97 5.83 67.23 6.09 ;
        RECT 66.97 5.07 67.23 5.33 ;
        RECT 67.73 6.59 67.99 6.85 ;
        RECT 67.73 5.83 67.99 6.09 ;
        RECT 67.73 5.07 67.99 5.33 ;
        RECT 68.49 6.59 68.75 6.85 ;
        RECT 68.49 5.83 68.75 6.09 ;
        RECT 68.49 5.07 68.75 5.33 ;
        RECT 69.25 6.59 69.51 6.85 ;
        RECT 69.25 5.83 69.51 6.09 ;
        RECT 69.25 5.07 69.51 5.33 ;
        RECT 70.01 6.59 70.27 6.85 ;
        RECT 70.01 5.83 70.27 6.09 ;
        RECT 70.01 5.07 70.27 5.33 ;
        RECT 70.77 6.59 71.03 6.85 ;
        RECT 70.77 5.83 71.03 6.09 ;
        RECT 70.77 5.07 71.03 5.33 ;
        RECT 71.53 6.59 71.79 6.85 ;
        RECT 71.53 5.83 71.79 6.09 ;
        RECT 71.53 5.07 71.79 5.33 ;
        RECT 72.29 6.59 72.55 6.85 ;
        RECT 72.29 5.83 72.55 6.09 ;
        RECT 72.29 5.07 72.55 5.33 ;
        RECT 73.05 6.59 73.31 6.85 ;
        RECT 73.05 5.83 73.31 6.09 ;
        RECT 73.05 5.07 73.31 5.33 ;
        RECT 73.81 6.59 74.07 6.85 ;
        RECT 73.81 5.83 74.07 6.09 ;
        RECT 73.81 5.07 74.07 5.33 ;
        RECT 74.57 6.59 74.83 6.85 ;
        RECT 74.57 5.83 74.83 6.09 ;
        RECT 74.57 5.07 74.83 5.33 ;
        RECT 75.33 6.59 75.59 6.85 ;
        RECT 75.33 5.83 75.59 6.09 ;
        RECT 75.33 5.07 75.59 5.33 ;
        RECT 76.09 6.59 76.35 6.85 ;
        RECT 76.09 5.83 76.35 6.09 ;
        RECT 76.09 5.07 76.35 5.33 ;
        RECT 76.85 6.59 77.11 6.85 ;
        RECT 76.85 5.83 77.11 6.09 ;
        RECT 76.85 5.07 77.11 5.33 ;
        RECT 77.61 6.59 77.87 6.85 ;
        RECT 77.61 5.83 77.87 6.09 ;
        RECT 77.61 5.07 77.87 5.33 ;
        RECT 78.37 6.59 78.63 6.85 ;
        RECT 78.37 5.83 78.63 6.09 ;
        RECT 78.37 5.07 78.63 5.33 ;
        RECT 79.13 6.59 79.39 6.85 ;
        RECT 79.13 5.83 79.39 6.09 ;
        RECT 79.13 5.07 79.39 5.33 ;
        RECT 79.89 6.59 80.15 6.85 ;
        RECT 79.89 5.83 80.15 6.09 ;
        RECT 79.89 5.07 80.15 5.33 ;
        RECT 80.65 6.59 80.91 6.85 ;
        RECT 80.65 5.83 80.91 6.09 ;
        RECT 80.65 5.07 80.91 5.33 ;
        RECT 81.41 6.59 81.67 6.85 ;
        RECT 81.41 5.83 81.67 6.09 ;
        RECT 81.41 5.07 81.67 5.33 ;
        RECT 82.17 6.59 82.43 6.85 ;
        RECT 82.17 5.83 82.43 6.09 ;
        RECT 82.17 5.07 82.43 5.33 ;
        RECT 82.93 6.59 83.19 6.85 ;
        RECT 82.93 5.83 83.19 6.09 ;
        RECT 82.93 5.07 83.19 5.33 ;
        RECT 83.69 6.59 83.95 6.85 ;
        RECT 83.69 5.83 83.95 6.09 ;
        RECT 83.69 5.07 83.95 5.33 ;
        RECT 84.45 6.59 84.71 6.85 ;
        RECT 84.45 5.83 84.71 6.09 ;
        RECT 84.45 5.07 84.71 5.33 ;
        RECT 85.21 6.59 85.47 6.85 ;
        RECT 85.21 5.83 85.47 6.09 ;
        RECT 85.21 5.07 85.47 5.33 ;
        RECT 85.97 6.59 86.23 6.85 ;
        RECT 85.97 5.83 86.23 6.09 ;
        RECT 85.97 5.07 86.23 5.33 ;
        RECT 86.73 6.59 86.99 6.85 ;
        RECT 86.73 5.83 86.99 6.09 ;
        RECT 86.73 5.07 86.99 5.33 ;
        RECT 87.49 6.59 87.75 6.85 ;
        RECT 87.49 5.83 87.75 6.09 ;
        RECT 87.49 5.07 87.75 5.33 ;
        RECT 88.25 6.59 88.51 6.85 ;
        RECT 88.25 5.83 88.51 6.09 ;
        RECT 88.25 5.07 88.51 5.33 ;
        RECT 89.01 6.59 89.27 6.85 ;
        RECT 89.01 5.83 89.27 6.09 ;
        RECT 89.01 5.07 89.27 5.33 ;
        RECT 89.77 6.59 90.03 6.85 ;
        RECT 89.77 5.83 90.03 6.09 ;
        RECT 89.77 5.07 90.03 5.33 ;
        RECT 90.53 6.59 90.79 6.85 ;
        RECT 90.53 5.83 90.79 6.09 ;
        RECT 90.53 5.07 90.79 5.33 ;
        RECT 91.29 6.59 91.55 6.85 ;
        RECT 91.29 5.83 91.55 6.09 ;
        RECT 91.29 5.07 91.55 5.33 ;
        RECT 92.05 6.59 92.31 6.85 ;
        RECT 92.05 5.83 92.31 6.09 ;
        RECT 92.05 5.07 92.31 5.33 ;
        RECT 92.81 6.59 93.07 6.85 ;
        RECT 92.81 5.83 93.07 6.09 ;
        RECT 92.81 5.07 93.07 5.33 ;
        RECT 93.57 6.59 93.83 6.85 ;
        RECT 93.57 5.83 93.83 6.09 ;
        RECT 93.57 5.07 93.83 5.33 ;
        RECT 94.33 6.59 94.59 6.85 ;
        RECT 94.33 5.83 94.59 6.09 ;
        RECT 94.33 5.07 94.59 5.33 ;
        RECT 95.09 6.59 95.35 6.85 ;
        RECT 95.09 5.83 95.35 6.09 ;
        RECT 95.09 5.07 95.35 5.33 ;
    END
  END SUB
  OBS
    LAYER M1 ;
      RECT 91.32 5.73 92.13 93.185 ;
      RECT 8.335 5.73 9.145 93.185 ;
      RECT 91.28 5.73 92.13 92.03 ;
      RECT 8.325 12.26 9.145 92.03 ;
      RECT 8.335 5.73 92.13 12.58 ;
      RECT 4.59 5.73 95.41 7.53 ;
      RECT 64.285 33.295 88.065 33.575 ;
      RECT 12.35 33.295 36.13 33.575 ;
      RECT 12.35 33.33 88.065 33.56 ;
      RECT 87.745 29.995 87.975 33.575 ;
      RECT 64.285 29.995 88.065 30.275 ;
      RECT 12.35 29.995 36.13 30.275 ;
      RECT 12.35 30.03 88.065 30.26 ;
      RECT 64.285 47.065 88.065 47.345 ;
      RECT 12.35 47.065 36.13 47.345 ;
      RECT 12.35 47.08 88.065 47.31 ;
      RECT 87.745 43.765 87.975 47.345 ;
      RECT 64.285 43.765 88.065 44.045 ;
      RECT 12.35 43.765 36.13 44.045 ;
      RECT 12.35 43.78 88.065 44.01 ;
      RECT 77.19 61.775 87.98 62.055 ;
      RECT 87.7 58.475 87.98 62.055 ;
      RECT 12.4 61.775 23.19 62.055 ;
      RECT 12.4 61.8 87.98 62.03 ;
      RECT 12.4 58.475 12.68 62.055 ;
      RECT 77.19 58.475 87.98 58.755 ;
      RECT 12.4 58.475 23.19 58.755 ;
      RECT 12.4 58.5 87.98 58.73 ;
      RECT 77.19 83.695 87.98 83.975 ;
      RECT 87.7 80.395 87.98 83.975 ;
      RECT 12.4 83.695 23.19 83.975 ;
      RECT 12.4 83.72 87.98 83.95 ;
      RECT 12.4 80.395 12.68 83.975 ;
      RECT 77.19 80.395 87.98 80.675 ;
      RECT 12.4 80.395 23.19 80.675 ;
      RECT 12.4 80.42 87.98 80.65 ;
      RECT 38.33 19.125 62.11 19.405 ;
      RECT 12.445 19.16 87.975 19.39 ;
      RECT 87.745 15.86 87.975 19.39 ;
      RECT 38.33 15.825 62.11 16.105 ;
      RECT 12.445 15.86 87.975 16.09 ;
      RECT 64.28 72.725 75.06 73.005 ;
      RECT 25.32 72.725 36.1 73.005 ;
      RECT 12.425 72.76 87.955 72.99 ;
      RECT 87.725 69.46 87.955 72.99 ;
      RECT 64.28 69.425 75.06 69.705 ;
      RECT 25.32 69.425 36.1 69.705 ;
      RECT 12.425 69.46 87.955 69.69 ;
      RECT 38.285 94.645 62.065 94.925 ;
      RECT 12.425 94.68 87.955 94.91 ;
      RECT 87.725 91.38 87.955 94.91 ;
      RECT 38.285 91.345 62.065 91.625 ;
      RECT 12.425 91.38 87.955 91.61 ;
      RECT 64.805 59.265 74.545 61.27 ;
      RECT 25.835 59.265 35.575 61.27 ;
      RECT 13.19 59.265 87.19 61.265 ;
      RECT 13.21 16.625 87.21 18.625 ;
      RECT 13.21 30.795 87.21 32.795 ;
      RECT 13.21 44.545 87.21 46.545 ;
      RECT 13.19 70.225 87.19 72.225 ;
      RECT 13.19 81.185 87.19 83.185 ;
      RECT 13.19 92.145 87.19 94.145 ;
    LAYER M2 ;
      RECT 4.64 5.68 95.36 7.58 ;
      RECT 4.59 5.73 95.41 7.53 ;
      RECT 64.21 29.46 88.21 33.835 ;
      RECT 64.19 14.67 88.19 30.49 ;
      RECT 64.19 15.29 88.21 19.665 ;
      RECT 64.19 39.18 75.19 61.84 ;
      RECT 64.19 39.18 88.19 56 ;
      RECT 64.19 43.505 88.21 47.88 ;
      RECT 77.19 58.475 88.19 73.185 ;
      RECT 77.19 58.455 88 73.185 ;
      RECT 38.19 15.09 62.19 95.105 ;
      RECT 38.19 43.545 62.21 47.98 ;
      RECT 38.19 29.36 62.21 33.795 ;
      RECT 38.19 15.19 62.21 19.625 ;
      RECT 12.21 29.46 36.21 33.835 ;
      RECT 12.19 14.67 36.19 30.49 ;
      RECT 12.19 15.29 36.21 19.665 ;
      RECT 25.19 39.18 36.19 61.84 ;
      RECT 12.19 39.18 36.19 56 ;
      RECT 12.19 43.505 36.21 47.88 ;
      RECT 12.19 58.475 23.19 73.185 ;
      RECT 12.38 58.455 23.19 73.185 ;
      RECT 77.19 79.745 88.19 95.105 ;
      RECT 64.19 69.375 75.19 84.045 ;
      RECT 25.19 69.375 36.19 84.045 ;
      RECT 12.19 79.745 23.19 95.105 ;
    LAYER TOP_M ;
      RECT 0 96 100 119.035 ;
  END
END PAD_DVDD

END LIBRARY
