// Library - TJ_Monopix_01, Cell - matrix_dac, View - schematic
// LAST TIME SAVED: May 19 19:21:00 2017
// NETLIST TIME: May 22 11:27:12 2017
`timescale 1ns / 1ns 

module matrix_dac ( DIG_MON_COMP, DIG_MON_HV, DIG_MON_PMOS,
     DIG_MON_PMOS_DPW, Data_COMP, Data_HV, Data_PMOS, Data_PMOS_DPW,
     OUTA_MON_L, OUTA_MON_R, nTOK_COMP, nTOK_HV, nTOK_PMOS,
     nTOK_PMOS_DPW, DACMON_IBIAS, DACMON_ICASN, DACMON_IDB,
     DACMON_IRESET, DACMON_ITHR, DACMON_VH, DACMON_VL, DACMON_VRESET_P,
     GNDA, GNDA_IDAC, GNDA_VDAC, GNDD, GND_Per, HV_DIODE, PSUB, PWELL,
     VDDA, VDDA_IDAC, VDDA_VDAC, VDDD, VDD_Per, BcidMtx, BiasSF,
     DIG_MON_SEL, FREEZE_COMP, FREEZE_HV, FREEZE_PMOS, FREEZE_PMOS_DPW,
     IBUFN_L_SET, IBUFN_R_SET, IBUFP_L_SET, IBUFP_R_SET, INJ_IN,
     INJ_IN_MON_L, INJ_IN_MON_R, INJ_ROW, MASKD, MASKH, MASKV,
     Read_COMP, Read_HV, Read_PMOS, Read_PMOS_DPW, SET_IBIAS,
     SET_ICASN, SET_IDB, SET_IRESET, SET_IRESET_BIT, SET_ITHR,
     SET_VCASN, SET_VCLIP, SET_VH, SET_VL, SET_VRESET_D, SET_VRESET_P,
     SWCNTL_DACMONI, SWCNTL_DACMONV, SWCNTL_IBIAS, SWCNTL_ICASN,
     SWCNTL_IDB, SWCNTL_IREF, SWCNTL_IRESET, SWCNTL_ITHR, SWCNTL_VCASN,
     SWCNTL_VCLIP, SWCNTL_VH, SWCNTL_VL, SWCNTL_VRESET_D,
     SWCNTL_VRESET_P, Vpc, nRST );

inout DACMON_IBIAS, DACMON_ICASN, DACMON_IDB, DACMON_IRESET,
     DACMON_ITHR, DACMON_VH, DACMON_VL, DACMON_VRESET_P, GNDA,
     GNDA_IDAC, GNDA_VDAC, GNDD, GND_Per, HV_DIODE, PSUB, PWELL, VDDA,
     VDDA_IDAC, VDDA_VDAC, VDDD, VDD_Per;

inout BiasSF, Vpc;
     
input INJ_IN_MON_L, INJ_IN_MON_R, SET_IRESET_BIT,
     SWCNTL_DACMONI, SWCNTL_DACMONV, SWCNTL_IBIAS, SWCNTL_ICASN,
     SWCNTL_IDB, SWCNTL_IREF, SWCNTL_IRESET, SWCNTL_ITHR, SWCNTL_VCASN,
     SWCNTL_VCLIP, SWCNTL_VH, SWCNTL_VL, SWCNTL_VRESET_D,
     SWCNTL_VRESET_P, nRST;

output [55:0]  nTOK_PMOS;
output [1175:0]  Data_COMP;
output [55:0]  nTOK_PMOS_DPW;
output [111:0]  DIG_MON_PMOS;
inout [3:0]  OUTA_MON_L;
output [1175:0]  Data_PMOS;
output [1175:0]  Data_HV;
output [1175:0]  Data_PMOS_DPW;
output [111:0]  DIG_MON_COMP;
output [111:0]  DIG_MON_PMOS_DPW;
inout [3:0]  OUTA_MON_R;
output [55:0]  nTOK_HV;
output [55:0]  nTOK_COMP;
output [111:0]  DIG_MON_HV;

input [127:0]  SET_ICASN;
input [127:0]  SET_VRESET_P;
input [447:0]  DIG_MON_SEL;
input [223:0]  INJ_ROW;
input [127:0]  SET_ITHR;
input [55:0]  FREEZE_COMP;
input [55:0]  Read_COMP;
input [55:0]  Read_HV;
input [127:0]  SET_VRESET_D;
input [55:0]  FREEZE_PMOS_DPW;
input [55:0]  Read_PMOS;
input [3:0]  IBUFN_R_SET;
input [127:0]  SET_VL;
input [127:0]  SET_IDB;
input [127:0]  SET_IBIAS;
input [223:0]  MASKH;
input [447:0]  INJ_IN;
input [55:0]  FREEZE_HV;
input [127:0]  SET_IRESET;
input [127:0]  SET_VCASN;
input [3:0]  IBUFP_R_SET;
input [447:0]  MASKV;
input [127:0]  SET_VCLIP;
input [55:0]  FREEZE_PMOS;
input [1343:0]  BcidMtx;
input [3:0]  IBUFP_L_SET;
input [3:0]  IBUFN_L_SET;
input [447:0]  MASKD;
input [127:0]  SET_VH;
input [55:0]  Read_PMOS_DPW;

//TODO: TB logic

endmodule
