VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO decoupling_cap_filler
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN decoupling_cap_filler 0 0 ;
  SIZE 20 BY 120 ;
  SYMMETRY X Y R90 ;
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER V4 ;
        RECT 3.005 91.14 3.265 91.4 ;
        RECT 3.005 90.38 3.265 90.64 ;
        RECT 3.005 89.62 3.265 89.88 ;
        RECT 3.005 88.86 3.265 89.12 ;
        RECT 3.005 88.1 3.265 88.36 ;
        RECT 3.005 87.34 3.265 87.6 ;
        RECT 3.005 86.58 3.265 86.84 ;
        RECT 3.005 85.82 3.265 86.08 ;
        RECT 3.005 85.06 3.265 85.32 ;
        RECT 3.005 84.3 3.265 84.56 ;
        RECT 3.005 83.54 3.265 83.8 ;
        RECT 3.005 82.78 3.265 83.04 ;
        RECT 3.005 82.02 3.265 82.28 ;
        RECT 3.005 81.26 3.265 81.52 ;
        RECT 3.005 80.5 3.265 80.76 ;
        RECT 3.005 79.74 3.265 80 ;
        RECT 3.005 78.98 3.265 79.24 ;
        RECT 3.005 78.22 3.265 78.48 ;
        RECT 3.005 77.46 3.265 77.72 ;
        RECT 3.005 76.7 3.265 76.96 ;
        RECT 3.005 75.94 3.265 76.2 ;
        RECT 3.005 75.18 3.265 75.44 ;
        RECT 3.005 74.42 3.265 74.68 ;
        RECT 3.005 73.66 3.265 73.92 ;
        RECT 3.005 72.9 3.265 73.16 ;
        RECT 3.005 72.14 3.265 72.4 ;
        RECT 3.005 71.38 3.265 71.64 ;
        RECT 3.005 70.62 3.265 70.88 ;
        RECT 3.005 69.86 3.265 70.12 ;
        RECT 3.005 69.1 3.265 69.36 ;
        RECT 3.765 91.14 4.025 91.4 ;
        RECT 3.765 90.38 4.025 90.64 ;
        RECT 3.765 89.62 4.025 89.88 ;
        RECT 3.765 88.86 4.025 89.12 ;
        RECT 3.765 88.1 4.025 88.36 ;
        RECT 3.765 87.34 4.025 87.6 ;
        RECT 3.765 86.58 4.025 86.84 ;
        RECT 3.765 85.82 4.025 86.08 ;
        RECT 3.765 85.06 4.025 85.32 ;
        RECT 3.765 84.3 4.025 84.56 ;
        RECT 3.765 83.54 4.025 83.8 ;
        RECT 3.765 82.78 4.025 83.04 ;
        RECT 3.765 82.02 4.025 82.28 ;
        RECT 3.765 81.26 4.025 81.52 ;
        RECT 3.765 80.5 4.025 80.76 ;
        RECT 3.765 79.74 4.025 80 ;
        RECT 3.765 78.98 4.025 79.24 ;
        RECT 3.765 78.22 4.025 78.48 ;
        RECT 3.765 77.46 4.025 77.72 ;
        RECT 3.765 76.7 4.025 76.96 ;
        RECT 3.765 75.94 4.025 76.2 ;
        RECT 3.765 75.18 4.025 75.44 ;
        RECT 3.765 74.42 4.025 74.68 ;
        RECT 3.765 73.66 4.025 73.92 ;
        RECT 3.765 72.9 4.025 73.16 ;
        RECT 3.765 72.14 4.025 72.4 ;
        RECT 3.765 71.38 4.025 71.64 ;
        RECT 3.765 70.62 4.025 70.88 ;
        RECT 3.765 69.86 4.025 70.12 ;
        RECT 3.765 69.1 4.025 69.36 ;
        RECT 4.525 91.14 4.785 91.4 ;
        RECT 4.525 90.38 4.785 90.64 ;
        RECT 4.525 89.62 4.785 89.88 ;
        RECT 4.525 88.86 4.785 89.12 ;
        RECT 4.525 88.1 4.785 88.36 ;
        RECT 4.525 87.34 4.785 87.6 ;
        RECT 4.525 86.58 4.785 86.84 ;
        RECT 4.525 85.82 4.785 86.08 ;
        RECT 4.525 85.06 4.785 85.32 ;
        RECT 4.525 84.3 4.785 84.56 ;
        RECT 4.525 83.54 4.785 83.8 ;
        RECT 4.525 82.78 4.785 83.04 ;
        RECT 4.525 82.02 4.785 82.28 ;
        RECT 4.525 81.26 4.785 81.52 ;
        RECT 4.525 80.5 4.785 80.76 ;
        RECT 4.525 79.74 4.785 80 ;
        RECT 4.525 78.98 4.785 79.24 ;
        RECT 4.525 78.22 4.785 78.48 ;
        RECT 4.525 77.46 4.785 77.72 ;
        RECT 4.525 76.7 4.785 76.96 ;
        RECT 4.525 75.94 4.785 76.2 ;
        RECT 4.525 75.18 4.785 75.44 ;
        RECT 4.525 74.42 4.785 74.68 ;
        RECT 4.525 73.66 4.785 73.92 ;
        RECT 4.525 72.9 4.785 73.16 ;
        RECT 4.525 72.14 4.785 72.4 ;
        RECT 4.525 71.38 4.785 71.64 ;
        RECT 4.525 70.62 4.785 70.88 ;
        RECT 4.525 69.86 4.785 70.12 ;
        RECT 4.525 69.1 4.785 69.36 ;
        RECT 5.285 91.14 5.545 91.4 ;
        RECT 5.285 90.38 5.545 90.64 ;
        RECT 5.285 89.62 5.545 89.88 ;
        RECT 5.285 88.86 5.545 89.12 ;
        RECT 5.285 88.1 5.545 88.36 ;
        RECT 5.285 87.34 5.545 87.6 ;
        RECT 5.285 86.58 5.545 86.84 ;
        RECT 5.285 85.82 5.545 86.08 ;
        RECT 5.285 85.06 5.545 85.32 ;
        RECT 5.285 84.3 5.545 84.56 ;
        RECT 5.285 83.54 5.545 83.8 ;
        RECT 5.285 82.78 5.545 83.04 ;
        RECT 5.285 82.02 5.545 82.28 ;
        RECT 5.285 81.26 5.545 81.52 ;
        RECT 5.285 80.5 5.545 80.76 ;
        RECT 5.285 79.74 5.545 80 ;
        RECT 5.285 78.98 5.545 79.24 ;
        RECT 5.285 78.22 5.545 78.48 ;
        RECT 5.285 77.46 5.545 77.72 ;
        RECT 5.285 76.7 5.545 76.96 ;
        RECT 5.285 75.94 5.545 76.2 ;
        RECT 5.285 75.18 5.545 75.44 ;
        RECT 5.285 74.42 5.545 74.68 ;
        RECT 5.285 73.66 5.545 73.92 ;
        RECT 5.285 72.9 5.545 73.16 ;
        RECT 5.285 72.14 5.545 72.4 ;
        RECT 5.285 71.38 5.545 71.64 ;
        RECT 5.285 70.62 5.545 70.88 ;
        RECT 5.285 69.86 5.545 70.12 ;
        RECT 5.285 69.1 5.545 69.36 ;
        RECT 6.045 91.14 6.305 91.4 ;
        RECT 6.045 90.38 6.305 90.64 ;
        RECT 6.045 89.62 6.305 89.88 ;
        RECT 6.045 88.86 6.305 89.12 ;
        RECT 6.045 88.1 6.305 88.36 ;
        RECT 6.045 87.34 6.305 87.6 ;
        RECT 6.045 86.58 6.305 86.84 ;
        RECT 6.045 85.82 6.305 86.08 ;
        RECT 6.045 85.06 6.305 85.32 ;
        RECT 6.045 84.3 6.305 84.56 ;
        RECT 6.045 83.54 6.305 83.8 ;
        RECT 6.045 82.78 6.305 83.04 ;
        RECT 6.045 82.02 6.305 82.28 ;
        RECT 6.045 81.26 6.305 81.52 ;
        RECT 6.045 80.5 6.305 80.76 ;
        RECT 6.045 79.74 6.305 80 ;
        RECT 6.045 78.98 6.305 79.24 ;
        RECT 6.045 78.22 6.305 78.48 ;
        RECT 6.045 77.46 6.305 77.72 ;
        RECT 6.045 76.7 6.305 76.96 ;
        RECT 6.045 75.94 6.305 76.2 ;
        RECT 6.045 75.18 6.305 75.44 ;
        RECT 6.045 74.42 6.305 74.68 ;
        RECT 6.045 73.66 6.305 73.92 ;
        RECT 6.045 72.9 6.305 73.16 ;
        RECT 6.045 72.14 6.305 72.4 ;
        RECT 6.045 71.38 6.305 71.64 ;
        RECT 6.045 70.62 6.305 70.88 ;
        RECT 6.045 69.86 6.305 70.12 ;
        RECT 6.045 69.1 6.305 69.36 ;
        RECT 6.805 91.14 7.065 91.4 ;
        RECT 6.805 90.38 7.065 90.64 ;
        RECT 6.805 89.62 7.065 89.88 ;
        RECT 6.805 88.86 7.065 89.12 ;
        RECT 6.805 88.1 7.065 88.36 ;
        RECT 6.805 87.34 7.065 87.6 ;
        RECT 6.805 86.58 7.065 86.84 ;
        RECT 6.805 85.82 7.065 86.08 ;
        RECT 6.805 85.06 7.065 85.32 ;
        RECT 6.805 84.3 7.065 84.56 ;
        RECT 6.805 83.54 7.065 83.8 ;
        RECT 6.805 82.78 7.065 83.04 ;
        RECT 6.805 82.02 7.065 82.28 ;
        RECT 6.805 81.26 7.065 81.52 ;
        RECT 6.805 80.5 7.065 80.76 ;
        RECT 6.805 79.74 7.065 80 ;
        RECT 6.805 78.98 7.065 79.24 ;
        RECT 6.805 78.22 7.065 78.48 ;
        RECT 6.805 77.46 7.065 77.72 ;
        RECT 6.805 76.7 7.065 76.96 ;
        RECT 6.805 75.94 7.065 76.2 ;
        RECT 6.805 75.18 7.065 75.44 ;
        RECT 6.805 74.42 7.065 74.68 ;
        RECT 6.805 73.66 7.065 73.92 ;
        RECT 6.805 72.9 7.065 73.16 ;
        RECT 6.805 72.14 7.065 72.4 ;
        RECT 6.805 71.38 7.065 71.64 ;
        RECT 6.805 70.62 7.065 70.88 ;
        RECT 6.805 69.86 7.065 70.12 ;
        RECT 6.805 69.1 7.065 69.36 ;
        RECT 7.565 91.14 7.825 91.4 ;
        RECT 7.565 90.38 7.825 90.64 ;
        RECT 7.565 89.62 7.825 89.88 ;
        RECT 7.565 88.86 7.825 89.12 ;
        RECT 7.565 88.1 7.825 88.36 ;
        RECT 7.565 87.34 7.825 87.6 ;
        RECT 7.565 86.58 7.825 86.84 ;
        RECT 7.565 85.82 7.825 86.08 ;
        RECT 7.565 85.06 7.825 85.32 ;
        RECT 7.565 84.3 7.825 84.56 ;
        RECT 7.565 83.54 7.825 83.8 ;
        RECT 7.565 82.78 7.825 83.04 ;
        RECT 7.565 82.02 7.825 82.28 ;
        RECT 7.565 81.26 7.825 81.52 ;
        RECT 7.565 80.5 7.825 80.76 ;
        RECT 7.565 79.74 7.825 80 ;
        RECT 7.565 78.98 7.825 79.24 ;
        RECT 7.565 78.22 7.825 78.48 ;
        RECT 7.565 77.46 7.825 77.72 ;
        RECT 7.565 76.7 7.825 76.96 ;
        RECT 7.565 75.94 7.825 76.2 ;
        RECT 7.565 75.18 7.825 75.44 ;
        RECT 7.565 74.42 7.825 74.68 ;
        RECT 7.565 73.66 7.825 73.92 ;
        RECT 7.565 72.9 7.825 73.16 ;
        RECT 7.565 72.14 7.825 72.4 ;
        RECT 7.565 71.38 7.825 71.64 ;
        RECT 7.565 70.62 7.825 70.88 ;
        RECT 7.565 69.86 7.825 70.12 ;
        RECT 7.565 69.1 7.825 69.36 ;
        RECT 8.325 91.14 8.585 91.4 ;
        RECT 8.325 90.38 8.585 90.64 ;
        RECT 8.325 89.62 8.585 89.88 ;
        RECT 8.325 88.86 8.585 89.12 ;
        RECT 8.325 88.1 8.585 88.36 ;
        RECT 8.325 87.34 8.585 87.6 ;
        RECT 8.325 86.58 8.585 86.84 ;
        RECT 8.325 85.82 8.585 86.08 ;
        RECT 8.325 85.06 8.585 85.32 ;
        RECT 8.325 84.3 8.585 84.56 ;
        RECT 8.325 83.54 8.585 83.8 ;
        RECT 8.325 82.78 8.585 83.04 ;
        RECT 8.325 82.02 8.585 82.28 ;
        RECT 8.325 81.26 8.585 81.52 ;
        RECT 8.325 80.5 8.585 80.76 ;
        RECT 8.325 79.74 8.585 80 ;
        RECT 8.325 78.98 8.585 79.24 ;
        RECT 8.325 78.22 8.585 78.48 ;
        RECT 8.325 77.46 8.585 77.72 ;
        RECT 8.325 76.7 8.585 76.96 ;
        RECT 8.325 75.94 8.585 76.2 ;
        RECT 8.325 75.18 8.585 75.44 ;
        RECT 8.325 74.42 8.585 74.68 ;
        RECT 8.325 73.66 8.585 73.92 ;
        RECT 8.325 72.9 8.585 73.16 ;
        RECT 8.325 72.14 8.585 72.4 ;
        RECT 8.325 71.38 8.585 71.64 ;
        RECT 8.325 70.62 8.585 70.88 ;
        RECT 8.325 69.86 8.585 70.12 ;
        RECT 8.325 69.1 8.585 69.36 ;
        RECT 9.085 91.14 9.345 91.4 ;
        RECT 9.085 90.38 9.345 90.64 ;
        RECT 9.085 89.62 9.345 89.88 ;
        RECT 9.085 88.86 9.345 89.12 ;
        RECT 9.085 88.1 9.345 88.36 ;
        RECT 9.085 87.34 9.345 87.6 ;
        RECT 9.085 86.58 9.345 86.84 ;
        RECT 9.085 85.82 9.345 86.08 ;
        RECT 9.085 85.06 9.345 85.32 ;
        RECT 9.085 84.3 9.345 84.56 ;
        RECT 9.085 83.54 9.345 83.8 ;
        RECT 9.085 82.78 9.345 83.04 ;
        RECT 9.085 82.02 9.345 82.28 ;
        RECT 9.085 81.26 9.345 81.52 ;
        RECT 9.085 80.5 9.345 80.76 ;
        RECT 9.085 79.74 9.345 80 ;
        RECT 9.085 78.98 9.345 79.24 ;
        RECT 9.085 78.22 9.345 78.48 ;
        RECT 9.085 77.46 9.345 77.72 ;
        RECT 9.085 76.7 9.345 76.96 ;
        RECT 9.085 75.94 9.345 76.2 ;
        RECT 9.085 75.18 9.345 75.44 ;
        RECT 9.085 74.42 9.345 74.68 ;
        RECT 9.085 73.66 9.345 73.92 ;
        RECT 9.085 72.9 9.345 73.16 ;
        RECT 9.085 72.14 9.345 72.4 ;
        RECT 9.085 71.38 9.345 71.64 ;
        RECT 9.085 70.62 9.345 70.88 ;
        RECT 9.085 69.86 9.345 70.12 ;
        RECT 9.085 69.1 9.345 69.36 ;
        RECT 9.845 91.14 10.105 91.4 ;
        RECT 9.845 90.38 10.105 90.64 ;
        RECT 9.845 89.62 10.105 89.88 ;
        RECT 9.845 88.86 10.105 89.12 ;
        RECT 9.845 88.1 10.105 88.36 ;
        RECT 9.845 87.34 10.105 87.6 ;
        RECT 9.845 86.58 10.105 86.84 ;
        RECT 9.845 85.82 10.105 86.08 ;
        RECT 9.845 85.06 10.105 85.32 ;
        RECT 9.845 84.3 10.105 84.56 ;
        RECT 9.845 83.54 10.105 83.8 ;
        RECT 9.845 82.78 10.105 83.04 ;
        RECT 9.845 82.02 10.105 82.28 ;
        RECT 9.845 81.26 10.105 81.52 ;
        RECT 9.845 80.5 10.105 80.76 ;
        RECT 9.845 79.74 10.105 80 ;
        RECT 9.845 78.98 10.105 79.24 ;
        RECT 9.845 78.22 10.105 78.48 ;
        RECT 9.845 77.46 10.105 77.72 ;
        RECT 9.845 76.7 10.105 76.96 ;
        RECT 9.845 75.94 10.105 76.2 ;
        RECT 9.845 75.18 10.105 75.44 ;
        RECT 9.845 74.42 10.105 74.68 ;
        RECT 9.845 73.66 10.105 73.92 ;
        RECT 9.845 72.9 10.105 73.16 ;
        RECT 9.845 72.14 10.105 72.4 ;
        RECT 9.845 71.38 10.105 71.64 ;
        RECT 9.845 70.62 10.105 70.88 ;
        RECT 9.845 69.86 10.105 70.12 ;
        RECT 9.845 69.1 10.105 69.36 ;
        RECT 10.605 91.14 10.865 91.4 ;
        RECT 10.605 90.38 10.865 90.64 ;
        RECT 10.605 89.62 10.865 89.88 ;
        RECT 10.605 88.86 10.865 89.12 ;
        RECT 10.605 88.1 10.865 88.36 ;
        RECT 10.605 87.34 10.865 87.6 ;
        RECT 10.605 86.58 10.865 86.84 ;
        RECT 10.605 85.82 10.865 86.08 ;
        RECT 10.605 85.06 10.865 85.32 ;
        RECT 10.605 84.3 10.865 84.56 ;
        RECT 10.605 83.54 10.865 83.8 ;
        RECT 10.605 82.78 10.865 83.04 ;
        RECT 10.605 82.02 10.865 82.28 ;
        RECT 10.605 81.26 10.865 81.52 ;
        RECT 10.605 80.5 10.865 80.76 ;
        RECT 10.605 79.74 10.865 80 ;
        RECT 10.605 78.98 10.865 79.24 ;
        RECT 10.605 78.22 10.865 78.48 ;
        RECT 10.605 77.46 10.865 77.72 ;
        RECT 10.605 76.7 10.865 76.96 ;
        RECT 10.605 75.94 10.865 76.2 ;
        RECT 10.605 75.18 10.865 75.44 ;
        RECT 10.605 74.42 10.865 74.68 ;
        RECT 10.605 73.66 10.865 73.92 ;
        RECT 10.605 72.9 10.865 73.16 ;
        RECT 10.605 72.14 10.865 72.4 ;
        RECT 10.605 71.38 10.865 71.64 ;
        RECT 10.605 70.62 10.865 70.88 ;
        RECT 10.605 69.86 10.865 70.12 ;
        RECT 10.605 69.1 10.865 69.36 ;
        RECT 11.365 91.14 11.625 91.4 ;
        RECT 11.365 90.38 11.625 90.64 ;
        RECT 11.365 89.62 11.625 89.88 ;
        RECT 11.365 88.86 11.625 89.12 ;
        RECT 11.365 88.1 11.625 88.36 ;
        RECT 11.365 87.34 11.625 87.6 ;
        RECT 11.365 86.58 11.625 86.84 ;
        RECT 11.365 85.82 11.625 86.08 ;
        RECT 11.365 85.06 11.625 85.32 ;
        RECT 11.365 84.3 11.625 84.56 ;
        RECT 11.365 83.54 11.625 83.8 ;
        RECT 11.365 82.78 11.625 83.04 ;
        RECT 11.365 82.02 11.625 82.28 ;
        RECT 11.365 81.26 11.625 81.52 ;
        RECT 11.365 80.5 11.625 80.76 ;
        RECT 11.365 79.74 11.625 80 ;
        RECT 11.365 78.98 11.625 79.24 ;
        RECT 11.365 78.22 11.625 78.48 ;
        RECT 11.365 77.46 11.625 77.72 ;
        RECT 11.365 76.7 11.625 76.96 ;
        RECT 11.365 75.94 11.625 76.2 ;
        RECT 11.365 75.18 11.625 75.44 ;
        RECT 11.365 74.42 11.625 74.68 ;
        RECT 11.365 73.66 11.625 73.92 ;
        RECT 11.365 72.9 11.625 73.16 ;
        RECT 11.365 72.14 11.625 72.4 ;
        RECT 11.365 71.38 11.625 71.64 ;
        RECT 11.365 70.62 11.625 70.88 ;
        RECT 11.365 69.86 11.625 70.12 ;
        RECT 11.365 69.1 11.625 69.36 ;
        RECT 12.125 91.14 12.385 91.4 ;
        RECT 12.125 90.38 12.385 90.64 ;
        RECT 12.125 89.62 12.385 89.88 ;
        RECT 12.125 88.86 12.385 89.12 ;
        RECT 12.125 88.1 12.385 88.36 ;
        RECT 12.125 87.34 12.385 87.6 ;
        RECT 12.125 86.58 12.385 86.84 ;
        RECT 12.125 85.82 12.385 86.08 ;
        RECT 12.125 85.06 12.385 85.32 ;
        RECT 12.125 84.3 12.385 84.56 ;
        RECT 12.125 83.54 12.385 83.8 ;
        RECT 12.125 82.78 12.385 83.04 ;
        RECT 12.125 82.02 12.385 82.28 ;
        RECT 12.125 81.26 12.385 81.52 ;
        RECT 12.125 80.5 12.385 80.76 ;
        RECT 12.125 79.74 12.385 80 ;
        RECT 12.125 78.98 12.385 79.24 ;
        RECT 12.125 78.22 12.385 78.48 ;
        RECT 12.125 77.46 12.385 77.72 ;
        RECT 12.125 76.7 12.385 76.96 ;
        RECT 12.125 75.94 12.385 76.2 ;
        RECT 12.125 75.18 12.385 75.44 ;
        RECT 12.125 74.42 12.385 74.68 ;
        RECT 12.125 73.66 12.385 73.92 ;
        RECT 12.125 72.9 12.385 73.16 ;
        RECT 12.125 72.14 12.385 72.4 ;
        RECT 12.125 71.38 12.385 71.64 ;
        RECT 12.125 70.62 12.385 70.88 ;
        RECT 12.125 69.86 12.385 70.12 ;
        RECT 12.125 69.1 12.385 69.36 ;
        RECT 12.885 91.14 13.145 91.4 ;
        RECT 12.885 90.38 13.145 90.64 ;
        RECT 12.885 89.62 13.145 89.88 ;
        RECT 12.885 88.86 13.145 89.12 ;
        RECT 12.885 88.1 13.145 88.36 ;
        RECT 12.885 87.34 13.145 87.6 ;
        RECT 12.885 86.58 13.145 86.84 ;
        RECT 12.885 85.82 13.145 86.08 ;
        RECT 12.885 85.06 13.145 85.32 ;
        RECT 12.885 84.3 13.145 84.56 ;
        RECT 12.885 83.54 13.145 83.8 ;
        RECT 12.885 82.78 13.145 83.04 ;
        RECT 12.885 82.02 13.145 82.28 ;
        RECT 12.885 81.26 13.145 81.52 ;
        RECT 12.885 80.5 13.145 80.76 ;
        RECT 12.885 79.74 13.145 80 ;
        RECT 12.885 78.98 13.145 79.24 ;
        RECT 12.885 78.22 13.145 78.48 ;
        RECT 12.885 77.46 13.145 77.72 ;
        RECT 12.885 76.7 13.145 76.96 ;
        RECT 12.885 75.94 13.145 76.2 ;
        RECT 12.885 75.18 13.145 75.44 ;
        RECT 12.885 74.42 13.145 74.68 ;
        RECT 12.885 73.66 13.145 73.92 ;
        RECT 12.885 72.9 13.145 73.16 ;
        RECT 12.885 72.14 13.145 72.4 ;
        RECT 12.885 71.38 13.145 71.64 ;
        RECT 12.885 70.62 13.145 70.88 ;
        RECT 12.885 69.86 13.145 70.12 ;
        RECT 12.885 69.1 13.145 69.36 ;
        RECT 13.645 91.14 13.905 91.4 ;
        RECT 13.645 90.38 13.905 90.64 ;
        RECT 13.645 89.62 13.905 89.88 ;
        RECT 13.645 88.86 13.905 89.12 ;
        RECT 13.645 88.1 13.905 88.36 ;
        RECT 13.645 87.34 13.905 87.6 ;
        RECT 13.645 86.58 13.905 86.84 ;
        RECT 13.645 85.82 13.905 86.08 ;
        RECT 13.645 85.06 13.905 85.32 ;
        RECT 13.645 84.3 13.905 84.56 ;
        RECT 13.645 83.54 13.905 83.8 ;
        RECT 13.645 82.78 13.905 83.04 ;
        RECT 13.645 82.02 13.905 82.28 ;
        RECT 13.645 81.26 13.905 81.52 ;
        RECT 13.645 80.5 13.905 80.76 ;
        RECT 13.645 79.74 13.905 80 ;
        RECT 13.645 78.98 13.905 79.24 ;
        RECT 13.645 78.22 13.905 78.48 ;
        RECT 13.645 77.46 13.905 77.72 ;
        RECT 13.645 76.7 13.905 76.96 ;
        RECT 13.645 75.94 13.905 76.2 ;
        RECT 13.645 75.18 13.905 75.44 ;
        RECT 13.645 74.42 13.905 74.68 ;
        RECT 13.645 73.66 13.905 73.92 ;
        RECT 13.645 72.9 13.905 73.16 ;
        RECT 13.645 72.14 13.905 72.4 ;
        RECT 13.645 71.38 13.905 71.64 ;
        RECT 13.645 70.62 13.905 70.88 ;
        RECT 13.645 69.86 13.905 70.12 ;
        RECT 13.645 69.1 13.905 69.36 ;
        RECT 14.405 91.14 14.665 91.4 ;
        RECT 14.405 90.38 14.665 90.64 ;
        RECT 14.405 89.62 14.665 89.88 ;
        RECT 14.405 88.86 14.665 89.12 ;
        RECT 14.405 88.1 14.665 88.36 ;
        RECT 14.405 87.34 14.665 87.6 ;
        RECT 14.405 86.58 14.665 86.84 ;
        RECT 14.405 85.82 14.665 86.08 ;
        RECT 14.405 85.06 14.665 85.32 ;
        RECT 14.405 84.3 14.665 84.56 ;
        RECT 14.405 83.54 14.665 83.8 ;
        RECT 14.405 82.78 14.665 83.04 ;
        RECT 14.405 82.02 14.665 82.28 ;
        RECT 14.405 81.26 14.665 81.52 ;
        RECT 14.405 80.5 14.665 80.76 ;
        RECT 14.405 79.74 14.665 80 ;
        RECT 14.405 78.98 14.665 79.24 ;
        RECT 14.405 78.22 14.665 78.48 ;
        RECT 14.405 77.46 14.665 77.72 ;
        RECT 14.405 76.7 14.665 76.96 ;
        RECT 14.405 75.94 14.665 76.2 ;
        RECT 14.405 75.18 14.665 75.44 ;
        RECT 14.405 74.42 14.665 74.68 ;
        RECT 14.405 73.66 14.665 73.92 ;
        RECT 14.405 72.9 14.665 73.16 ;
        RECT 14.405 72.14 14.665 72.4 ;
        RECT 14.405 71.38 14.665 71.64 ;
        RECT 14.405 70.62 14.665 70.88 ;
        RECT 14.405 69.86 14.665 70.12 ;
        RECT 14.405 69.1 14.665 69.36 ;
        RECT 15.165 91.14 15.425 91.4 ;
        RECT 15.165 90.38 15.425 90.64 ;
        RECT 15.165 89.62 15.425 89.88 ;
        RECT 15.165 88.86 15.425 89.12 ;
        RECT 15.165 88.1 15.425 88.36 ;
        RECT 15.165 87.34 15.425 87.6 ;
        RECT 15.165 86.58 15.425 86.84 ;
        RECT 15.165 85.82 15.425 86.08 ;
        RECT 15.165 85.06 15.425 85.32 ;
        RECT 15.165 84.3 15.425 84.56 ;
        RECT 15.165 83.54 15.425 83.8 ;
        RECT 15.165 82.78 15.425 83.04 ;
        RECT 15.165 82.02 15.425 82.28 ;
        RECT 15.165 81.26 15.425 81.52 ;
        RECT 15.165 80.5 15.425 80.76 ;
        RECT 15.165 79.74 15.425 80 ;
        RECT 15.165 78.98 15.425 79.24 ;
        RECT 15.165 78.22 15.425 78.48 ;
        RECT 15.165 77.46 15.425 77.72 ;
        RECT 15.165 76.7 15.425 76.96 ;
        RECT 15.165 75.94 15.425 76.2 ;
        RECT 15.165 75.18 15.425 75.44 ;
        RECT 15.165 74.42 15.425 74.68 ;
        RECT 15.165 73.66 15.425 73.92 ;
        RECT 15.165 72.9 15.425 73.16 ;
        RECT 15.165 72.14 15.425 72.4 ;
        RECT 15.165 71.38 15.425 71.64 ;
        RECT 15.165 70.62 15.425 70.88 ;
        RECT 15.165 69.86 15.425 70.12 ;
        RECT 15.165 69.1 15.425 69.36 ;
        RECT 15.925 91.14 16.185 91.4 ;
        RECT 15.925 90.38 16.185 90.64 ;
        RECT 15.925 89.62 16.185 89.88 ;
        RECT 15.925 88.86 16.185 89.12 ;
        RECT 15.925 88.1 16.185 88.36 ;
        RECT 15.925 87.34 16.185 87.6 ;
        RECT 15.925 86.58 16.185 86.84 ;
        RECT 15.925 85.82 16.185 86.08 ;
        RECT 15.925 85.06 16.185 85.32 ;
        RECT 15.925 84.3 16.185 84.56 ;
        RECT 15.925 83.54 16.185 83.8 ;
        RECT 15.925 82.78 16.185 83.04 ;
        RECT 15.925 82.02 16.185 82.28 ;
        RECT 15.925 81.26 16.185 81.52 ;
        RECT 15.925 80.5 16.185 80.76 ;
        RECT 15.925 79.74 16.185 80 ;
        RECT 15.925 78.98 16.185 79.24 ;
        RECT 15.925 78.22 16.185 78.48 ;
        RECT 15.925 77.46 16.185 77.72 ;
        RECT 15.925 76.7 16.185 76.96 ;
        RECT 15.925 75.94 16.185 76.2 ;
        RECT 15.925 75.18 16.185 75.44 ;
        RECT 15.925 74.42 16.185 74.68 ;
        RECT 15.925 73.66 16.185 73.92 ;
        RECT 15.925 72.9 16.185 73.16 ;
        RECT 15.925 72.14 16.185 72.4 ;
        RECT 15.925 71.38 16.185 71.64 ;
        RECT 15.925 70.62 16.185 70.88 ;
        RECT 15.925 69.86 16.185 70.12 ;
        RECT 15.925 69.1 16.185 69.36 ;
        RECT 16.685 91.14 16.945 91.4 ;
        RECT 16.685 90.38 16.945 90.64 ;
        RECT 16.685 89.62 16.945 89.88 ;
        RECT 16.685 88.86 16.945 89.12 ;
        RECT 16.685 88.1 16.945 88.36 ;
        RECT 16.685 87.34 16.945 87.6 ;
        RECT 16.685 86.58 16.945 86.84 ;
        RECT 16.685 85.82 16.945 86.08 ;
        RECT 16.685 85.06 16.945 85.32 ;
        RECT 16.685 84.3 16.945 84.56 ;
        RECT 16.685 83.54 16.945 83.8 ;
        RECT 16.685 82.78 16.945 83.04 ;
        RECT 16.685 82.02 16.945 82.28 ;
        RECT 16.685 81.26 16.945 81.52 ;
        RECT 16.685 80.5 16.945 80.76 ;
        RECT 16.685 79.74 16.945 80 ;
        RECT 16.685 78.98 16.945 79.24 ;
        RECT 16.685 78.22 16.945 78.48 ;
        RECT 16.685 77.46 16.945 77.72 ;
        RECT 16.685 76.7 16.945 76.96 ;
        RECT 16.685 75.94 16.945 76.2 ;
        RECT 16.685 75.18 16.945 75.44 ;
        RECT 16.685 74.42 16.945 74.68 ;
        RECT 16.685 73.66 16.945 73.92 ;
        RECT 16.685 72.9 16.945 73.16 ;
        RECT 16.685 72.14 16.945 72.4 ;
        RECT 16.685 71.38 16.945 71.64 ;
        RECT 16.685 70.62 16.945 70.88 ;
        RECT 16.685 69.86 16.945 70.12 ;
        RECT 16.685 69.1 16.945 69.36 ;
        RECT 17.445 91.14 17.705 91.4 ;
        RECT 17.445 90.38 17.705 90.64 ;
        RECT 17.445 89.62 17.705 89.88 ;
        RECT 17.445 88.86 17.705 89.12 ;
        RECT 17.445 88.1 17.705 88.36 ;
        RECT 17.445 87.34 17.705 87.6 ;
        RECT 17.445 86.58 17.705 86.84 ;
        RECT 17.445 85.82 17.705 86.08 ;
        RECT 17.445 85.06 17.705 85.32 ;
        RECT 17.445 84.3 17.705 84.56 ;
        RECT 17.445 83.54 17.705 83.8 ;
        RECT 17.445 82.78 17.705 83.04 ;
        RECT 17.445 82.02 17.705 82.28 ;
        RECT 17.445 81.26 17.705 81.52 ;
        RECT 17.445 80.5 17.705 80.76 ;
        RECT 17.445 79.74 17.705 80 ;
        RECT 17.445 78.98 17.705 79.24 ;
        RECT 17.445 78.22 17.705 78.48 ;
        RECT 17.445 77.46 17.705 77.72 ;
        RECT 17.445 76.7 17.705 76.96 ;
        RECT 17.445 75.94 17.705 76.2 ;
        RECT 17.445 75.18 17.705 75.44 ;
        RECT 17.445 74.42 17.705 74.68 ;
        RECT 17.445 73.66 17.705 73.92 ;
        RECT 17.445 72.9 17.705 73.16 ;
        RECT 17.445 72.14 17.705 72.4 ;
        RECT 17.445 71.38 17.705 71.64 ;
        RECT 17.445 70.62 17.705 70.88 ;
        RECT 17.445 69.86 17.705 70.12 ;
        RECT 17.445 69.1 17.705 69.36 ;
      LAYER V3 ;
        RECT 2.13 68.105 2.39 68.365 ;
        RECT 2.13 68.625 2.39 68.885 ;
        RECT 2.13 69.145 2.39 69.405 ;
        RECT 2.13 69.665 2.39 69.925 ;
        RECT 2.13 70.185 2.39 70.445 ;
        RECT 2.13 70.705 2.39 70.965 ;
        RECT 2.13 71.225 2.39 71.485 ;
        RECT 2.13 71.745 2.39 72.005 ;
        RECT 2.13 72.265 2.39 72.525 ;
        RECT 2.13 72.785 2.39 73.045 ;
        RECT 2.13 73.305 2.39 73.565 ;
        RECT 2.13 73.825 2.39 74.085 ;
        RECT 2.13 74.345 2.39 74.605 ;
        RECT 2.13 74.865 2.39 75.125 ;
        RECT 2.13 75.385 2.39 75.645 ;
        RECT 2.13 75.905 2.39 76.165 ;
        RECT 2.13 76.425 2.39 76.685 ;
        RECT 2.13 76.945 2.39 77.205 ;
        RECT 2.13 77.465 2.39 77.725 ;
        RECT 2.13 77.985 2.39 78.245 ;
        RECT 2.13 78.505 2.39 78.765 ;
        RECT 2.13 79.025 2.39 79.285 ;
        RECT 2.13 79.545 2.39 79.805 ;
        RECT 2.13 80.065 2.39 80.325 ;
        RECT 2.13 80.585 2.39 80.845 ;
        RECT 2.13 81.105 2.39 81.365 ;
        RECT 2.13 81.625 2.39 81.885 ;
        RECT 2.13 82.145 2.39 82.405 ;
        RECT 2.13 82.665 2.39 82.925 ;
        RECT 2.13 83.185 2.39 83.445 ;
        RECT 2.13 83.705 2.39 83.965 ;
        RECT 2.13 84.225 2.39 84.485 ;
        RECT 2.13 84.745 2.39 85.005 ;
        RECT 2.13 85.265 2.39 85.525 ;
        RECT 2.13 85.785 2.39 86.045 ;
        RECT 2.13 86.305 2.39 86.565 ;
        RECT 2.13 86.825 2.39 87.085 ;
        RECT 2.13 87.345 2.39 87.605 ;
        RECT 2.13 87.865 2.39 88.125 ;
        RECT 2.13 88.385 2.39 88.645 ;
        RECT 2.13 88.905 2.39 89.165 ;
        RECT 2.13 89.425 2.39 89.685 ;
        RECT 2.13 89.945 2.39 90.205 ;
        RECT 2.13 90.465 2.39 90.725 ;
        RECT 2.13 90.985 2.39 91.245 ;
        RECT 2.13 91.505 2.39 91.765 ;
        RECT 2.13 92.025 2.39 92.285 ;
        RECT 2.13 92.545 2.39 92.805 ;
        RECT 2.13 93.065 2.39 93.325 ;
        RECT 2.13 93.585 2.39 93.845 ;
        RECT 1.61 68.105 1.87 68.365 ;
        RECT 1.61 68.625 1.87 68.885 ;
        RECT 1.61 69.145 1.87 69.405 ;
        RECT 1.61 69.665 1.87 69.925 ;
        RECT 1.61 70.185 1.87 70.445 ;
        RECT 1.61 70.705 1.87 70.965 ;
        RECT 1.61 71.225 1.87 71.485 ;
        RECT 1.61 71.745 1.87 72.005 ;
        RECT 1.61 72.265 1.87 72.525 ;
        RECT 1.61 72.785 1.87 73.045 ;
        RECT 1.61 73.305 1.87 73.565 ;
        RECT 1.61 73.825 1.87 74.085 ;
        RECT 1.61 74.345 1.87 74.605 ;
        RECT 1.61 74.865 1.87 75.125 ;
        RECT 1.61 75.385 1.87 75.645 ;
        RECT 1.61 75.905 1.87 76.165 ;
        RECT 1.61 76.425 1.87 76.685 ;
        RECT 1.61 76.945 1.87 77.205 ;
        RECT 1.61 77.465 1.87 77.725 ;
        RECT 1.61 77.985 1.87 78.245 ;
        RECT 1.61 78.505 1.87 78.765 ;
        RECT 1.61 79.025 1.87 79.285 ;
        RECT 1.61 79.545 1.87 79.805 ;
        RECT 1.61 80.065 1.87 80.325 ;
        RECT 1.61 80.585 1.87 80.845 ;
        RECT 1.61 81.105 1.87 81.365 ;
        RECT 1.61 81.625 1.87 81.885 ;
        RECT 1.61 82.145 1.87 82.405 ;
        RECT 1.61 82.665 1.87 82.925 ;
        RECT 1.61 83.185 1.87 83.445 ;
        RECT 1.61 83.705 1.87 83.965 ;
        RECT 1.61 84.225 1.87 84.485 ;
        RECT 1.61 84.745 1.87 85.005 ;
        RECT 1.61 85.265 1.87 85.525 ;
        RECT 1.61 85.785 1.87 86.045 ;
        RECT 1.61 86.305 1.87 86.565 ;
        RECT 1.61 86.825 1.87 87.085 ;
        RECT 1.61 87.345 1.87 87.605 ;
        RECT 1.61 87.865 1.87 88.125 ;
        RECT 1.61 88.385 1.87 88.645 ;
        RECT 1.61 88.905 1.87 89.165 ;
        RECT 1.61 89.425 1.87 89.685 ;
        RECT 1.61 89.945 1.87 90.205 ;
        RECT 1.61 90.465 1.87 90.725 ;
        RECT 1.61 90.985 1.87 91.245 ;
        RECT 1.61 91.505 1.87 91.765 ;
        RECT 1.61 92.025 1.87 92.285 ;
        RECT 1.61 92.545 1.87 92.805 ;
        RECT 1.61 93.065 1.87 93.325 ;
        RECT 1.61 93.585 1.87 93.845 ;
      LAYER M4 ;
        RECT 0 66 20 96 ;
      LAYER M3 ;
        RECT 0 66 20 96 ;
    END
  END DVSS
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER V4 ;
        RECT 3.155 60.1 3.415 60.36 ;
        RECT 3.155 59.34 3.415 59.6 ;
        RECT 3.155 58.58 3.415 58.84 ;
        RECT 3.155 57.82 3.415 58.08 ;
        RECT 3.155 57.06 3.415 57.32 ;
        RECT 3.155 56.3 3.415 56.56 ;
        RECT 3.155 55.54 3.415 55.8 ;
        RECT 3.155 54.78 3.415 55.04 ;
        RECT 3.155 54.02 3.415 54.28 ;
        RECT 3.155 53.26 3.415 53.52 ;
        RECT 3.155 52.5 3.415 52.76 ;
        RECT 3.155 51.74 3.415 52 ;
        RECT 3.155 50.98 3.415 51.24 ;
        RECT 3.155 50.22 3.415 50.48 ;
        RECT 3.155 49.46 3.415 49.72 ;
        RECT 3.155 48.7 3.415 48.96 ;
        RECT 3.155 47.94 3.415 48.2 ;
        RECT 3.155 47.18 3.415 47.44 ;
        RECT 3.155 46.42 3.415 46.68 ;
        RECT 3.155 45.66 3.415 45.92 ;
        RECT 3.155 44.9 3.415 45.16 ;
        RECT 3.155 44.14 3.415 44.4 ;
        RECT 3.155 43.38 3.415 43.64 ;
        RECT 3.155 42.62 3.415 42.88 ;
        RECT 3.155 41.86 3.415 42.12 ;
        RECT 3.155 41.1 3.415 41.36 ;
        RECT 3.155 40.34 3.415 40.6 ;
        RECT 3.155 39.58 3.415 39.84 ;
        RECT 3.155 38.82 3.415 39.08 ;
        RECT 3.155 38.06 3.415 38.32 ;
        RECT 3.915 60.1 4.175 60.36 ;
        RECT 3.915 59.34 4.175 59.6 ;
        RECT 3.915 58.58 4.175 58.84 ;
        RECT 3.915 57.82 4.175 58.08 ;
        RECT 3.915 57.06 4.175 57.32 ;
        RECT 3.915 56.3 4.175 56.56 ;
        RECT 3.915 55.54 4.175 55.8 ;
        RECT 3.915 54.78 4.175 55.04 ;
        RECT 3.915 54.02 4.175 54.28 ;
        RECT 3.915 53.26 4.175 53.52 ;
        RECT 3.915 52.5 4.175 52.76 ;
        RECT 3.915 51.74 4.175 52 ;
        RECT 3.915 50.98 4.175 51.24 ;
        RECT 3.915 50.22 4.175 50.48 ;
        RECT 3.915 49.46 4.175 49.72 ;
        RECT 3.915 48.7 4.175 48.96 ;
        RECT 3.915 47.94 4.175 48.2 ;
        RECT 3.915 47.18 4.175 47.44 ;
        RECT 3.915 46.42 4.175 46.68 ;
        RECT 3.915 45.66 4.175 45.92 ;
        RECT 3.915 44.9 4.175 45.16 ;
        RECT 3.915 44.14 4.175 44.4 ;
        RECT 3.915 43.38 4.175 43.64 ;
        RECT 3.915 42.62 4.175 42.88 ;
        RECT 3.915 41.86 4.175 42.12 ;
        RECT 3.915 41.1 4.175 41.36 ;
        RECT 3.915 40.34 4.175 40.6 ;
        RECT 3.915 39.58 4.175 39.84 ;
        RECT 3.915 38.82 4.175 39.08 ;
        RECT 3.915 38.06 4.175 38.32 ;
        RECT 4.675 60.1 4.935 60.36 ;
        RECT 4.675 59.34 4.935 59.6 ;
        RECT 4.675 58.58 4.935 58.84 ;
        RECT 4.675 57.82 4.935 58.08 ;
        RECT 4.675 57.06 4.935 57.32 ;
        RECT 4.675 56.3 4.935 56.56 ;
        RECT 4.675 55.54 4.935 55.8 ;
        RECT 4.675 54.78 4.935 55.04 ;
        RECT 4.675 54.02 4.935 54.28 ;
        RECT 4.675 53.26 4.935 53.52 ;
        RECT 4.675 52.5 4.935 52.76 ;
        RECT 4.675 51.74 4.935 52 ;
        RECT 4.675 50.98 4.935 51.24 ;
        RECT 4.675 50.22 4.935 50.48 ;
        RECT 4.675 49.46 4.935 49.72 ;
        RECT 4.675 48.7 4.935 48.96 ;
        RECT 4.675 47.94 4.935 48.2 ;
        RECT 4.675 47.18 4.935 47.44 ;
        RECT 4.675 46.42 4.935 46.68 ;
        RECT 4.675 45.66 4.935 45.92 ;
        RECT 4.675 44.9 4.935 45.16 ;
        RECT 4.675 44.14 4.935 44.4 ;
        RECT 4.675 43.38 4.935 43.64 ;
        RECT 4.675 42.62 4.935 42.88 ;
        RECT 4.675 41.86 4.935 42.12 ;
        RECT 4.675 41.1 4.935 41.36 ;
        RECT 4.675 40.34 4.935 40.6 ;
        RECT 4.675 39.58 4.935 39.84 ;
        RECT 4.675 38.82 4.935 39.08 ;
        RECT 4.675 38.06 4.935 38.32 ;
        RECT 5.435 60.1 5.695 60.36 ;
        RECT 5.435 59.34 5.695 59.6 ;
        RECT 5.435 58.58 5.695 58.84 ;
        RECT 5.435 57.82 5.695 58.08 ;
        RECT 5.435 57.06 5.695 57.32 ;
        RECT 5.435 56.3 5.695 56.56 ;
        RECT 5.435 55.54 5.695 55.8 ;
        RECT 5.435 54.78 5.695 55.04 ;
        RECT 5.435 54.02 5.695 54.28 ;
        RECT 5.435 53.26 5.695 53.52 ;
        RECT 5.435 52.5 5.695 52.76 ;
        RECT 5.435 51.74 5.695 52 ;
        RECT 5.435 50.98 5.695 51.24 ;
        RECT 5.435 50.22 5.695 50.48 ;
        RECT 5.435 49.46 5.695 49.72 ;
        RECT 5.435 48.7 5.695 48.96 ;
        RECT 5.435 47.94 5.695 48.2 ;
        RECT 5.435 47.18 5.695 47.44 ;
        RECT 5.435 46.42 5.695 46.68 ;
        RECT 5.435 45.66 5.695 45.92 ;
        RECT 5.435 44.9 5.695 45.16 ;
        RECT 5.435 44.14 5.695 44.4 ;
        RECT 5.435 43.38 5.695 43.64 ;
        RECT 5.435 42.62 5.695 42.88 ;
        RECT 5.435 41.86 5.695 42.12 ;
        RECT 5.435 41.1 5.695 41.36 ;
        RECT 5.435 40.34 5.695 40.6 ;
        RECT 5.435 39.58 5.695 39.84 ;
        RECT 5.435 38.82 5.695 39.08 ;
        RECT 5.435 38.06 5.695 38.32 ;
        RECT 6.195 60.1 6.455 60.36 ;
        RECT 6.195 59.34 6.455 59.6 ;
        RECT 6.195 58.58 6.455 58.84 ;
        RECT 6.195 57.82 6.455 58.08 ;
        RECT 6.195 57.06 6.455 57.32 ;
        RECT 6.195 56.3 6.455 56.56 ;
        RECT 6.195 55.54 6.455 55.8 ;
        RECT 6.195 54.78 6.455 55.04 ;
        RECT 6.195 54.02 6.455 54.28 ;
        RECT 6.195 53.26 6.455 53.52 ;
        RECT 6.195 52.5 6.455 52.76 ;
        RECT 6.195 51.74 6.455 52 ;
        RECT 6.195 50.98 6.455 51.24 ;
        RECT 6.195 50.22 6.455 50.48 ;
        RECT 6.195 49.46 6.455 49.72 ;
        RECT 6.195 48.7 6.455 48.96 ;
        RECT 6.195 47.94 6.455 48.2 ;
        RECT 6.195 47.18 6.455 47.44 ;
        RECT 6.195 46.42 6.455 46.68 ;
        RECT 6.195 45.66 6.455 45.92 ;
        RECT 6.195 44.9 6.455 45.16 ;
        RECT 6.195 44.14 6.455 44.4 ;
        RECT 6.195 43.38 6.455 43.64 ;
        RECT 6.195 42.62 6.455 42.88 ;
        RECT 6.195 41.86 6.455 42.12 ;
        RECT 6.195 41.1 6.455 41.36 ;
        RECT 6.195 40.34 6.455 40.6 ;
        RECT 6.195 39.58 6.455 39.84 ;
        RECT 6.195 38.82 6.455 39.08 ;
        RECT 6.195 38.06 6.455 38.32 ;
        RECT 6.955 60.1 7.215 60.36 ;
        RECT 6.955 59.34 7.215 59.6 ;
        RECT 6.955 58.58 7.215 58.84 ;
        RECT 6.955 57.82 7.215 58.08 ;
        RECT 6.955 57.06 7.215 57.32 ;
        RECT 6.955 56.3 7.215 56.56 ;
        RECT 6.955 55.54 7.215 55.8 ;
        RECT 6.955 54.78 7.215 55.04 ;
        RECT 6.955 54.02 7.215 54.28 ;
        RECT 6.955 53.26 7.215 53.52 ;
        RECT 6.955 52.5 7.215 52.76 ;
        RECT 6.955 51.74 7.215 52 ;
        RECT 6.955 50.98 7.215 51.24 ;
        RECT 6.955 50.22 7.215 50.48 ;
        RECT 6.955 49.46 7.215 49.72 ;
        RECT 6.955 48.7 7.215 48.96 ;
        RECT 6.955 47.94 7.215 48.2 ;
        RECT 6.955 47.18 7.215 47.44 ;
        RECT 6.955 46.42 7.215 46.68 ;
        RECT 6.955 45.66 7.215 45.92 ;
        RECT 6.955 44.9 7.215 45.16 ;
        RECT 6.955 44.14 7.215 44.4 ;
        RECT 6.955 43.38 7.215 43.64 ;
        RECT 6.955 42.62 7.215 42.88 ;
        RECT 6.955 41.86 7.215 42.12 ;
        RECT 6.955 41.1 7.215 41.36 ;
        RECT 6.955 40.34 7.215 40.6 ;
        RECT 6.955 39.58 7.215 39.84 ;
        RECT 6.955 38.82 7.215 39.08 ;
        RECT 6.955 38.06 7.215 38.32 ;
        RECT 7.715 60.1 7.975 60.36 ;
        RECT 7.715 59.34 7.975 59.6 ;
        RECT 7.715 58.58 7.975 58.84 ;
        RECT 7.715 57.82 7.975 58.08 ;
        RECT 7.715 57.06 7.975 57.32 ;
        RECT 7.715 56.3 7.975 56.56 ;
        RECT 7.715 55.54 7.975 55.8 ;
        RECT 7.715 54.78 7.975 55.04 ;
        RECT 7.715 54.02 7.975 54.28 ;
        RECT 7.715 53.26 7.975 53.52 ;
        RECT 7.715 52.5 7.975 52.76 ;
        RECT 7.715 51.74 7.975 52 ;
        RECT 7.715 50.98 7.975 51.24 ;
        RECT 7.715 50.22 7.975 50.48 ;
        RECT 7.715 49.46 7.975 49.72 ;
        RECT 7.715 48.7 7.975 48.96 ;
        RECT 7.715 47.94 7.975 48.2 ;
        RECT 7.715 47.18 7.975 47.44 ;
        RECT 7.715 46.42 7.975 46.68 ;
        RECT 7.715 45.66 7.975 45.92 ;
        RECT 7.715 44.9 7.975 45.16 ;
        RECT 7.715 44.14 7.975 44.4 ;
        RECT 7.715 43.38 7.975 43.64 ;
        RECT 7.715 42.62 7.975 42.88 ;
        RECT 7.715 41.86 7.975 42.12 ;
        RECT 7.715 41.1 7.975 41.36 ;
        RECT 7.715 40.34 7.975 40.6 ;
        RECT 7.715 39.58 7.975 39.84 ;
        RECT 7.715 38.82 7.975 39.08 ;
        RECT 7.715 38.06 7.975 38.32 ;
        RECT 8.475 60.1 8.735 60.36 ;
        RECT 8.475 59.34 8.735 59.6 ;
        RECT 8.475 58.58 8.735 58.84 ;
        RECT 8.475 57.82 8.735 58.08 ;
        RECT 8.475 57.06 8.735 57.32 ;
        RECT 8.475 56.3 8.735 56.56 ;
        RECT 8.475 55.54 8.735 55.8 ;
        RECT 8.475 54.78 8.735 55.04 ;
        RECT 8.475 54.02 8.735 54.28 ;
        RECT 8.475 53.26 8.735 53.52 ;
        RECT 8.475 52.5 8.735 52.76 ;
        RECT 8.475 51.74 8.735 52 ;
        RECT 8.475 50.98 8.735 51.24 ;
        RECT 8.475 50.22 8.735 50.48 ;
        RECT 8.475 49.46 8.735 49.72 ;
        RECT 8.475 48.7 8.735 48.96 ;
        RECT 8.475 47.94 8.735 48.2 ;
        RECT 8.475 47.18 8.735 47.44 ;
        RECT 8.475 46.42 8.735 46.68 ;
        RECT 8.475 45.66 8.735 45.92 ;
        RECT 8.475 44.9 8.735 45.16 ;
        RECT 8.475 44.14 8.735 44.4 ;
        RECT 8.475 43.38 8.735 43.64 ;
        RECT 8.475 42.62 8.735 42.88 ;
        RECT 8.475 41.86 8.735 42.12 ;
        RECT 8.475 41.1 8.735 41.36 ;
        RECT 8.475 40.34 8.735 40.6 ;
        RECT 8.475 39.58 8.735 39.84 ;
        RECT 8.475 38.82 8.735 39.08 ;
        RECT 8.475 38.06 8.735 38.32 ;
        RECT 9.235 60.1 9.495 60.36 ;
        RECT 9.235 59.34 9.495 59.6 ;
        RECT 9.235 58.58 9.495 58.84 ;
        RECT 9.235 57.82 9.495 58.08 ;
        RECT 9.235 57.06 9.495 57.32 ;
        RECT 9.235 56.3 9.495 56.56 ;
        RECT 9.235 55.54 9.495 55.8 ;
        RECT 9.235 54.78 9.495 55.04 ;
        RECT 9.235 54.02 9.495 54.28 ;
        RECT 9.235 53.26 9.495 53.52 ;
        RECT 9.235 52.5 9.495 52.76 ;
        RECT 9.235 51.74 9.495 52 ;
        RECT 9.235 50.98 9.495 51.24 ;
        RECT 9.235 50.22 9.495 50.48 ;
        RECT 9.235 49.46 9.495 49.72 ;
        RECT 9.235 48.7 9.495 48.96 ;
        RECT 9.235 47.94 9.495 48.2 ;
        RECT 9.235 47.18 9.495 47.44 ;
        RECT 9.235 46.42 9.495 46.68 ;
        RECT 9.235 45.66 9.495 45.92 ;
        RECT 9.235 44.9 9.495 45.16 ;
        RECT 9.235 44.14 9.495 44.4 ;
        RECT 9.235 43.38 9.495 43.64 ;
        RECT 9.235 42.62 9.495 42.88 ;
        RECT 9.235 41.86 9.495 42.12 ;
        RECT 9.235 41.1 9.495 41.36 ;
        RECT 9.235 40.34 9.495 40.6 ;
        RECT 9.235 39.58 9.495 39.84 ;
        RECT 9.235 38.82 9.495 39.08 ;
        RECT 9.235 38.06 9.495 38.32 ;
        RECT 9.995 60.1 10.255 60.36 ;
        RECT 9.995 59.34 10.255 59.6 ;
        RECT 9.995 58.58 10.255 58.84 ;
        RECT 9.995 57.82 10.255 58.08 ;
        RECT 9.995 57.06 10.255 57.32 ;
        RECT 9.995 56.3 10.255 56.56 ;
        RECT 9.995 55.54 10.255 55.8 ;
        RECT 9.995 54.78 10.255 55.04 ;
        RECT 9.995 54.02 10.255 54.28 ;
        RECT 9.995 53.26 10.255 53.52 ;
        RECT 9.995 52.5 10.255 52.76 ;
        RECT 9.995 51.74 10.255 52 ;
        RECT 9.995 50.98 10.255 51.24 ;
        RECT 9.995 50.22 10.255 50.48 ;
        RECT 9.995 49.46 10.255 49.72 ;
        RECT 9.995 48.7 10.255 48.96 ;
        RECT 9.995 47.94 10.255 48.2 ;
        RECT 9.995 47.18 10.255 47.44 ;
        RECT 9.995 46.42 10.255 46.68 ;
        RECT 9.995 45.66 10.255 45.92 ;
        RECT 9.995 44.9 10.255 45.16 ;
        RECT 9.995 44.14 10.255 44.4 ;
        RECT 9.995 43.38 10.255 43.64 ;
        RECT 9.995 42.62 10.255 42.88 ;
        RECT 9.995 41.86 10.255 42.12 ;
        RECT 9.995 41.1 10.255 41.36 ;
        RECT 9.995 40.34 10.255 40.6 ;
        RECT 9.995 39.58 10.255 39.84 ;
        RECT 9.995 38.82 10.255 39.08 ;
        RECT 9.995 38.06 10.255 38.32 ;
        RECT 10.755 60.1 11.015 60.36 ;
        RECT 10.755 59.34 11.015 59.6 ;
        RECT 10.755 58.58 11.015 58.84 ;
        RECT 10.755 57.82 11.015 58.08 ;
        RECT 10.755 57.06 11.015 57.32 ;
        RECT 10.755 56.3 11.015 56.56 ;
        RECT 10.755 55.54 11.015 55.8 ;
        RECT 10.755 54.78 11.015 55.04 ;
        RECT 10.755 54.02 11.015 54.28 ;
        RECT 10.755 53.26 11.015 53.52 ;
        RECT 10.755 52.5 11.015 52.76 ;
        RECT 10.755 51.74 11.015 52 ;
        RECT 10.755 50.98 11.015 51.24 ;
        RECT 10.755 50.22 11.015 50.48 ;
        RECT 10.755 49.46 11.015 49.72 ;
        RECT 10.755 48.7 11.015 48.96 ;
        RECT 10.755 47.94 11.015 48.2 ;
        RECT 10.755 47.18 11.015 47.44 ;
        RECT 10.755 46.42 11.015 46.68 ;
        RECT 10.755 45.66 11.015 45.92 ;
        RECT 10.755 44.9 11.015 45.16 ;
        RECT 10.755 44.14 11.015 44.4 ;
        RECT 10.755 43.38 11.015 43.64 ;
        RECT 10.755 42.62 11.015 42.88 ;
        RECT 10.755 41.86 11.015 42.12 ;
        RECT 10.755 41.1 11.015 41.36 ;
        RECT 10.755 40.34 11.015 40.6 ;
        RECT 10.755 39.58 11.015 39.84 ;
        RECT 10.755 38.82 11.015 39.08 ;
        RECT 10.755 38.06 11.015 38.32 ;
        RECT 11.515 60.1 11.775 60.36 ;
        RECT 11.515 59.34 11.775 59.6 ;
        RECT 11.515 58.58 11.775 58.84 ;
        RECT 11.515 57.82 11.775 58.08 ;
        RECT 11.515 57.06 11.775 57.32 ;
        RECT 11.515 56.3 11.775 56.56 ;
        RECT 11.515 55.54 11.775 55.8 ;
        RECT 11.515 54.78 11.775 55.04 ;
        RECT 11.515 54.02 11.775 54.28 ;
        RECT 11.515 53.26 11.775 53.52 ;
        RECT 11.515 52.5 11.775 52.76 ;
        RECT 11.515 51.74 11.775 52 ;
        RECT 11.515 50.98 11.775 51.24 ;
        RECT 11.515 50.22 11.775 50.48 ;
        RECT 11.515 49.46 11.775 49.72 ;
        RECT 11.515 48.7 11.775 48.96 ;
        RECT 11.515 47.94 11.775 48.2 ;
        RECT 11.515 47.18 11.775 47.44 ;
        RECT 11.515 46.42 11.775 46.68 ;
        RECT 11.515 45.66 11.775 45.92 ;
        RECT 11.515 44.9 11.775 45.16 ;
        RECT 11.515 44.14 11.775 44.4 ;
        RECT 11.515 43.38 11.775 43.64 ;
        RECT 11.515 42.62 11.775 42.88 ;
        RECT 11.515 41.86 11.775 42.12 ;
        RECT 11.515 41.1 11.775 41.36 ;
        RECT 11.515 40.34 11.775 40.6 ;
        RECT 11.515 39.58 11.775 39.84 ;
        RECT 11.515 38.82 11.775 39.08 ;
        RECT 11.515 38.06 11.775 38.32 ;
        RECT 12.275 60.1 12.535 60.36 ;
        RECT 12.275 59.34 12.535 59.6 ;
        RECT 12.275 58.58 12.535 58.84 ;
        RECT 12.275 57.82 12.535 58.08 ;
        RECT 12.275 57.06 12.535 57.32 ;
        RECT 12.275 56.3 12.535 56.56 ;
        RECT 12.275 55.54 12.535 55.8 ;
        RECT 12.275 54.78 12.535 55.04 ;
        RECT 12.275 54.02 12.535 54.28 ;
        RECT 12.275 53.26 12.535 53.52 ;
        RECT 12.275 52.5 12.535 52.76 ;
        RECT 12.275 51.74 12.535 52 ;
        RECT 12.275 50.98 12.535 51.24 ;
        RECT 12.275 50.22 12.535 50.48 ;
        RECT 12.275 49.46 12.535 49.72 ;
        RECT 12.275 48.7 12.535 48.96 ;
        RECT 12.275 47.94 12.535 48.2 ;
        RECT 12.275 47.18 12.535 47.44 ;
        RECT 12.275 46.42 12.535 46.68 ;
        RECT 12.275 45.66 12.535 45.92 ;
        RECT 12.275 44.9 12.535 45.16 ;
        RECT 12.275 44.14 12.535 44.4 ;
        RECT 12.275 43.38 12.535 43.64 ;
        RECT 12.275 42.62 12.535 42.88 ;
        RECT 12.275 41.86 12.535 42.12 ;
        RECT 12.275 41.1 12.535 41.36 ;
        RECT 12.275 40.34 12.535 40.6 ;
        RECT 12.275 39.58 12.535 39.84 ;
        RECT 12.275 38.82 12.535 39.08 ;
        RECT 12.275 38.06 12.535 38.32 ;
        RECT 13.035 60.1 13.295 60.36 ;
        RECT 13.035 59.34 13.295 59.6 ;
        RECT 13.035 58.58 13.295 58.84 ;
        RECT 13.035 57.82 13.295 58.08 ;
        RECT 13.035 57.06 13.295 57.32 ;
        RECT 13.035 56.3 13.295 56.56 ;
        RECT 13.035 55.54 13.295 55.8 ;
        RECT 13.035 54.78 13.295 55.04 ;
        RECT 13.035 54.02 13.295 54.28 ;
        RECT 13.035 53.26 13.295 53.52 ;
        RECT 13.035 52.5 13.295 52.76 ;
        RECT 13.035 51.74 13.295 52 ;
        RECT 13.035 50.98 13.295 51.24 ;
        RECT 13.035 50.22 13.295 50.48 ;
        RECT 13.035 49.46 13.295 49.72 ;
        RECT 13.035 48.7 13.295 48.96 ;
        RECT 13.035 47.94 13.295 48.2 ;
        RECT 13.035 47.18 13.295 47.44 ;
        RECT 13.035 46.42 13.295 46.68 ;
        RECT 13.035 45.66 13.295 45.92 ;
        RECT 13.035 44.9 13.295 45.16 ;
        RECT 13.035 44.14 13.295 44.4 ;
        RECT 13.035 43.38 13.295 43.64 ;
        RECT 13.035 42.62 13.295 42.88 ;
        RECT 13.035 41.86 13.295 42.12 ;
        RECT 13.035 41.1 13.295 41.36 ;
        RECT 13.035 40.34 13.295 40.6 ;
        RECT 13.035 39.58 13.295 39.84 ;
        RECT 13.035 38.82 13.295 39.08 ;
        RECT 13.035 38.06 13.295 38.32 ;
        RECT 13.795 60.1 14.055 60.36 ;
        RECT 13.795 59.34 14.055 59.6 ;
        RECT 13.795 58.58 14.055 58.84 ;
        RECT 13.795 57.82 14.055 58.08 ;
        RECT 13.795 57.06 14.055 57.32 ;
        RECT 13.795 56.3 14.055 56.56 ;
        RECT 13.795 55.54 14.055 55.8 ;
        RECT 13.795 54.78 14.055 55.04 ;
        RECT 13.795 54.02 14.055 54.28 ;
        RECT 13.795 53.26 14.055 53.52 ;
        RECT 13.795 52.5 14.055 52.76 ;
        RECT 13.795 51.74 14.055 52 ;
        RECT 13.795 50.98 14.055 51.24 ;
        RECT 13.795 50.22 14.055 50.48 ;
        RECT 13.795 49.46 14.055 49.72 ;
        RECT 13.795 48.7 14.055 48.96 ;
        RECT 13.795 47.94 14.055 48.2 ;
        RECT 13.795 47.18 14.055 47.44 ;
        RECT 13.795 46.42 14.055 46.68 ;
        RECT 13.795 45.66 14.055 45.92 ;
        RECT 13.795 44.9 14.055 45.16 ;
        RECT 13.795 44.14 14.055 44.4 ;
        RECT 13.795 43.38 14.055 43.64 ;
        RECT 13.795 42.62 14.055 42.88 ;
        RECT 13.795 41.86 14.055 42.12 ;
        RECT 13.795 41.1 14.055 41.36 ;
        RECT 13.795 40.34 14.055 40.6 ;
        RECT 13.795 39.58 14.055 39.84 ;
        RECT 13.795 38.82 14.055 39.08 ;
        RECT 13.795 38.06 14.055 38.32 ;
        RECT 14.555 60.1 14.815 60.36 ;
        RECT 14.555 59.34 14.815 59.6 ;
        RECT 14.555 58.58 14.815 58.84 ;
        RECT 14.555 57.82 14.815 58.08 ;
        RECT 14.555 57.06 14.815 57.32 ;
        RECT 14.555 56.3 14.815 56.56 ;
        RECT 14.555 55.54 14.815 55.8 ;
        RECT 14.555 54.78 14.815 55.04 ;
        RECT 14.555 54.02 14.815 54.28 ;
        RECT 14.555 53.26 14.815 53.52 ;
        RECT 14.555 52.5 14.815 52.76 ;
        RECT 14.555 51.74 14.815 52 ;
        RECT 14.555 50.98 14.815 51.24 ;
        RECT 14.555 50.22 14.815 50.48 ;
        RECT 14.555 49.46 14.815 49.72 ;
        RECT 14.555 48.7 14.815 48.96 ;
        RECT 14.555 47.94 14.815 48.2 ;
        RECT 14.555 47.18 14.815 47.44 ;
        RECT 14.555 46.42 14.815 46.68 ;
        RECT 14.555 45.66 14.815 45.92 ;
        RECT 14.555 44.9 14.815 45.16 ;
        RECT 14.555 44.14 14.815 44.4 ;
        RECT 14.555 43.38 14.815 43.64 ;
        RECT 14.555 42.62 14.815 42.88 ;
        RECT 14.555 41.86 14.815 42.12 ;
        RECT 14.555 41.1 14.815 41.36 ;
        RECT 14.555 40.34 14.815 40.6 ;
        RECT 14.555 39.58 14.815 39.84 ;
        RECT 14.555 38.82 14.815 39.08 ;
        RECT 14.555 38.06 14.815 38.32 ;
        RECT 15.315 60.1 15.575 60.36 ;
        RECT 15.315 59.34 15.575 59.6 ;
        RECT 15.315 58.58 15.575 58.84 ;
        RECT 15.315 57.82 15.575 58.08 ;
        RECT 15.315 57.06 15.575 57.32 ;
        RECT 15.315 56.3 15.575 56.56 ;
        RECT 15.315 55.54 15.575 55.8 ;
        RECT 15.315 54.78 15.575 55.04 ;
        RECT 15.315 54.02 15.575 54.28 ;
        RECT 15.315 53.26 15.575 53.52 ;
        RECT 15.315 52.5 15.575 52.76 ;
        RECT 15.315 51.74 15.575 52 ;
        RECT 15.315 50.98 15.575 51.24 ;
        RECT 15.315 50.22 15.575 50.48 ;
        RECT 15.315 49.46 15.575 49.72 ;
        RECT 15.315 48.7 15.575 48.96 ;
        RECT 15.315 47.94 15.575 48.2 ;
        RECT 15.315 47.18 15.575 47.44 ;
        RECT 15.315 46.42 15.575 46.68 ;
        RECT 15.315 45.66 15.575 45.92 ;
        RECT 15.315 44.9 15.575 45.16 ;
        RECT 15.315 44.14 15.575 44.4 ;
        RECT 15.315 43.38 15.575 43.64 ;
        RECT 15.315 42.62 15.575 42.88 ;
        RECT 15.315 41.86 15.575 42.12 ;
        RECT 15.315 41.1 15.575 41.36 ;
        RECT 15.315 40.34 15.575 40.6 ;
        RECT 15.315 39.58 15.575 39.84 ;
        RECT 15.315 38.82 15.575 39.08 ;
        RECT 15.315 38.06 15.575 38.32 ;
        RECT 16.075 60.1 16.335 60.36 ;
        RECT 16.075 59.34 16.335 59.6 ;
        RECT 16.075 58.58 16.335 58.84 ;
        RECT 16.075 57.82 16.335 58.08 ;
        RECT 16.075 57.06 16.335 57.32 ;
        RECT 16.075 56.3 16.335 56.56 ;
        RECT 16.075 55.54 16.335 55.8 ;
        RECT 16.075 54.78 16.335 55.04 ;
        RECT 16.075 54.02 16.335 54.28 ;
        RECT 16.075 53.26 16.335 53.52 ;
        RECT 16.075 52.5 16.335 52.76 ;
        RECT 16.075 51.74 16.335 52 ;
        RECT 16.075 50.98 16.335 51.24 ;
        RECT 16.075 50.22 16.335 50.48 ;
        RECT 16.075 49.46 16.335 49.72 ;
        RECT 16.075 48.7 16.335 48.96 ;
        RECT 16.075 47.94 16.335 48.2 ;
        RECT 16.075 47.18 16.335 47.44 ;
        RECT 16.075 46.42 16.335 46.68 ;
        RECT 16.075 45.66 16.335 45.92 ;
        RECT 16.075 44.9 16.335 45.16 ;
        RECT 16.075 44.14 16.335 44.4 ;
        RECT 16.075 43.38 16.335 43.64 ;
        RECT 16.075 42.62 16.335 42.88 ;
        RECT 16.075 41.86 16.335 42.12 ;
        RECT 16.075 41.1 16.335 41.36 ;
        RECT 16.075 40.34 16.335 40.6 ;
        RECT 16.075 39.58 16.335 39.84 ;
        RECT 16.075 38.82 16.335 39.08 ;
        RECT 16.075 38.06 16.335 38.32 ;
        RECT 16.835 60.1 17.095 60.36 ;
        RECT 16.835 59.34 17.095 59.6 ;
        RECT 16.835 58.58 17.095 58.84 ;
        RECT 16.835 57.82 17.095 58.08 ;
        RECT 16.835 57.06 17.095 57.32 ;
        RECT 16.835 56.3 17.095 56.56 ;
        RECT 16.835 55.54 17.095 55.8 ;
        RECT 16.835 54.78 17.095 55.04 ;
        RECT 16.835 54.02 17.095 54.28 ;
        RECT 16.835 53.26 17.095 53.52 ;
        RECT 16.835 52.5 17.095 52.76 ;
        RECT 16.835 51.74 17.095 52 ;
        RECT 16.835 50.98 17.095 51.24 ;
        RECT 16.835 50.22 17.095 50.48 ;
        RECT 16.835 49.46 17.095 49.72 ;
        RECT 16.835 48.7 17.095 48.96 ;
        RECT 16.835 47.94 17.095 48.2 ;
        RECT 16.835 47.18 17.095 47.44 ;
        RECT 16.835 46.42 17.095 46.68 ;
        RECT 16.835 45.66 17.095 45.92 ;
        RECT 16.835 44.9 17.095 45.16 ;
        RECT 16.835 44.14 17.095 44.4 ;
        RECT 16.835 43.38 17.095 43.64 ;
        RECT 16.835 42.62 17.095 42.88 ;
        RECT 16.835 41.86 17.095 42.12 ;
        RECT 16.835 41.1 17.095 41.36 ;
        RECT 16.835 40.34 17.095 40.6 ;
        RECT 16.835 39.58 17.095 39.84 ;
        RECT 16.835 38.82 17.095 39.08 ;
        RECT 16.835 38.06 17.095 38.32 ;
        RECT 17.595 60.1 17.855 60.36 ;
        RECT 17.595 59.34 17.855 59.6 ;
        RECT 17.595 58.58 17.855 58.84 ;
        RECT 17.595 57.82 17.855 58.08 ;
        RECT 17.595 57.06 17.855 57.32 ;
        RECT 17.595 56.3 17.855 56.56 ;
        RECT 17.595 55.54 17.855 55.8 ;
        RECT 17.595 54.78 17.855 55.04 ;
        RECT 17.595 54.02 17.855 54.28 ;
        RECT 17.595 53.26 17.855 53.52 ;
        RECT 17.595 52.5 17.855 52.76 ;
        RECT 17.595 51.74 17.855 52 ;
        RECT 17.595 50.98 17.855 51.24 ;
        RECT 17.595 50.22 17.855 50.48 ;
        RECT 17.595 49.46 17.855 49.72 ;
        RECT 17.595 48.7 17.855 48.96 ;
        RECT 17.595 47.94 17.855 48.2 ;
        RECT 17.595 47.18 17.855 47.44 ;
        RECT 17.595 46.42 17.855 46.68 ;
        RECT 17.595 45.66 17.855 45.92 ;
        RECT 17.595 44.9 17.855 45.16 ;
        RECT 17.595 44.14 17.855 44.4 ;
        RECT 17.595 43.38 17.855 43.64 ;
        RECT 17.595 42.62 17.855 42.88 ;
        RECT 17.595 41.86 17.855 42.12 ;
        RECT 17.595 41.1 17.855 41.36 ;
        RECT 17.595 40.34 17.855 40.6 ;
        RECT 17.595 39.58 17.855 39.84 ;
        RECT 17.595 38.82 17.855 39.08 ;
        RECT 17.595 38.06 17.855 38.32 ;
      LAYER V3 ;
        RECT 18.13 35.705 18.39 35.965 ;
        RECT 18.13 36.225 18.39 36.485 ;
        RECT 18.13 36.745 18.39 37.005 ;
        RECT 18.13 37.265 18.39 37.525 ;
        RECT 18.13 37.785 18.39 38.045 ;
        RECT 18.13 38.305 18.39 38.565 ;
        RECT 18.13 38.825 18.39 39.085 ;
        RECT 18.13 39.345 18.39 39.605 ;
        RECT 18.13 39.865 18.39 40.125 ;
        RECT 18.13 40.385 18.39 40.645 ;
        RECT 18.13 40.905 18.39 41.165 ;
        RECT 18.13 41.425 18.39 41.685 ;
        RECT 18.13 41.945 18.39 42.205 ;
        RECT 18.13 42.465 18.39 42.725 ;
        RECT 18.13 42.985 18.39 43.245 ;
        RECT 18.13 43.505 18.39 43.765 ;
        RECT 18.13 44.025 18.39 44.285 ;
        RECT 18.13 44.545 18.39 44.805 ;
        RECT 18.13 45.065 18.39 45.325 ;
        RECT 18.13 45.585 18.39 45.845 ;
        RECT 18.13 46.105 18.39 46.365 ;
        RECT 18.13 46.625 18.39 46.885 ;
        RECT 18.13 47.145 18.39 47.405 ;
        RECT 18.13 47.665 18.39 47.925 ;
        RECT 18.13 48.185 18.39 48.445 ;
        RECT 18.13 48.705 18.39 48.965 ;
        RECT 18.13 49.225 18.39 49.485 ;
        RECT 18.13 49.745 18.39 50.005 ;
        RECT 18.13 50.265 18.39 50.525 ;
        RECT 18.13 50.785 18.39 51.045 ;
        RECT 18.13 51.305 18.39 51.565 ;
        RECT 18.13 51.825 18.39 52.085 ;
        RECT 18.13 52.345 18.39 52.605 ;
        RECT 18.13 52.865 18.39 53.125 ;
        RECT 18.13 53.385 18.39 53.645 ;
        RECT 18.13 53.905 18.39 54.165 ;
        RECT 18.13 54.425 18.39 54.685 ;
        RECT 18.13 54.945 18.39 55.205 ;
        RECT 18.13 55.465 18.39 55.725 ;
        RECT 18.13 55.985 18.39 56.245 ;
        RECT 18.13 56.505 18.39 56.765 ;
        RECT 18.13 57.025 18.39 57.285 ;
        RECT 18.13 57.545 18.39 57.805 ;
        RECT 18.13 58.065 18.39 58.325 ;
        RECT 18.13 58.585 18.39 58.845 ;
        RECT 18.13 59.105 18.39 59.365 ;
        RECT 18.13 59.625 18.39 59.885 ;
        RECT 18.13 60.145 18.39 60.405 ;
        RECT 18.13 60.665 18.39 60.925 ;
        RECT 18.13 61.185 18.39 61.445 ;
        RECT 17.61 35.705 17.87 35.965 ;
        RECT 17.61 36.225 17.87 36.485 ;
        RECT 17.61 36.745 17.87 37.005 ;
        RECT 17.61 37.265 17.87 37.525 ;
        RECT 17.61 37.785 17.87 38.045 ;
        RECT 17.61 38.305 17.87 38.565 ;
        RECT 17.61 38.825 17.87 39.085 ;
        RECT 17.61 39.345 17.87 39.605 ;
        RECT 17.61 39.865 17.87 40.125 ;
        RECT 17.61 40.385 17.87 40.645 ;
        RECT 17.61 40.905 17.87 41.165 ;
        RECT 17.61 41.425 17.87 41.685 ;
        RECT 17.61 41.945 17.87 42.205 ;
        RECT 17.61 42.465 17.87 42.725 ;
        RECT 17.61 42.985 17.87 43.245 ;
        RECT 17.61 43.505 17.87 43.765 ;
        RECT 17.61 44.025 17.87 44.285 ;
        RECT 17.61 44.545 17.87 44.805 ;
        RECT 17.61 45.065 17.87 45.325 ;
        RECT 17.61 45.585 17.87 45.845 ;
        RECT 17.61 46.105 17.87 46.365 ;
        RECT 17.61 46.625 17.87 46.885 ;
        RECT 17.61 47.145 17.87 47.405 ;
        RECT 17.61 47.665 17.87 47.925 ;
        RECT 17.61 48.185 17.87 48.445 ;
        RECT 17.61 48.705 17.87 48.965 ;
        RECT 17.61 49.225 17.87 49.485 ;
        RECT 17.61 49.745 17.87 50.005 ;
        RECT 17.61 50.265 17.87 50.525 ;
        RECT 17.61 50.785 17.87 51.045 ;
        RECT 17.61 51.305 17.87 51.565 ;
        RECT 17.61 51.825 17.87 52.085 ;
        RECT 17.61 52.345 17.87 52.605 ;
        RECT 17.61 52.865 17.87 53.125 ;
        RECT 17.61 53.385 17.87 53.645 ;
        RECT 17.61 53.905 17.87 54.165 ;
        RECT 17.61 54.425 17.87 54.685 ;
        RECT 17.61 54.945 17.87 55.205 ;
        RECT 17.61 55.465 17.87 55.725 ;
        RECT 17.61 55.985 17.87 56.245 ;
        RECT 17.61 56.505 17.87 56.765 ;
        RECT 17.61 57.025 17.87 57.285 ;
        RECT 17.61 57.545 17.87 57.805 ;
        RECT 17.61 58.065 17.87 58.325 ;
        RECT 17.61 58.585 17.87 58.845 ;
        RECT 17.61 59.105 17.87 59.365 ;
        RECT 17.61 59.625 17.87 59.885 ;
        RECT 17.61 60.145 17.87 60.405 ;
        RECT 17.61 60.665 17.87 60.925 ;
        RECT 17.61 61.185 17.87 61.445 ;
      LAYER M4 ;
        RECT 0 34 20 64 ;
      LAYER M3 ;
        RECT 0 34 20 64 ;
    END
  END DVDD
  PIN AVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER V4 ;
        RECT 2.56 30.03 2.82 30.29 ;
        RECT 2.56 29.27 2.82 29.53 ;
        RECT 2.56 28.51 2.82 28.77 ;
        RECT 2.56 27.75 2.82 28.01 ;
        RECT 2.56 26.99 2.82 27.25 ;
        RECT 2.56 26.23 2.82 26.49 ;
        RECT 2.56 25.47 2.82 25.73 ;
        RECT 2.56 24.71 2.82 24.97 ;
        RECT 2.56 23.95 2.82 24.21 ;
        RECT 2.56 23.19 2.82 23.45 ;
        RECT 3.32 30.03 3.58 30.29 ;
        RECT 3.32 29.27 3.58 29.53 ;
        RECT 3.32 28.51 3.58 28.77 ;
        RECT 3.32 27.75 3.58 28.01 ;
        RECT 3.32 26.99 3.58 27.25 ;
        RECT 3.32 26.23 3.58 26.49 ;
        RECT 3.32 25.47 3.58 25.73 ;
        RECT 3.32 24.71 3.58 24.97 ;
        RECT 3.32 23.95 3.58 24.21 ;
        RECT 3.32 23.19 3.58 23.45 ;
        RECT 4.08 30.03 4.34 30.29 ;
        RECT 4.08 29.27 4.34 29.53 ;
        RECT 4.08 28.51 4.34 28.77 ;
        RECT 4.08 27.75 4.34 28.01 ;
        RECT 4.08 26.99 4.34 27.25 ;
        RECT 4.08 26.23 4.34 26.49 ;
        RECT 4.08 25.47 4.34 25.73 ;
        RECT 4.08 24.71 4.34 24.97 ;
        RECT 4.08 23.95 4.34 24.21 ;
        RECT 4.08 23.19 4.34 23.45 ;
        RECT 4.84 30.03 5.1 30.29 ;
        RECT 4.84 29.27 5.1 29.53 ;
        RECT 4.84 28.51 5.1 28.77 ;
        RECT 4.84 27.75 5.1 28.01 ;
        RECT 4.84 26.99 5.1 27.25 ;
        RECT 4.84 26.23 5.1 26.49 ;
        RECT 4.84 25.47 5.1 25.73 ;
        RECT 4.84 24.71 5.1 24.97 ;
        RECT 4.84 23.95 5.1 24.21 ;
        RECT 4.84 23.19 5.1 23.45 ;
        RECT 5.6 30.03 5.86 30.29 ;
        RECT 5.6 29.27 5.86 29.53 ;
        RECT 5.6 28.51 5.86 28.77 ;
        RECT 5.6 27.75 5.86 28.01 ;
        RECT 5.6 26.99 5.86 27.25 ;
        RECT 5.6 26.23 5.86 26.49 ;
        RECT 5.6 25.47 5.86 25.73 ;
        RECT 5.6 24.71 5.86 24.97 ;
        RECT 5.6 23.95 5.86 24.21 ;
        RECT 5.6 23.19 5.86 23.45 ;
        RECT 6.36 30.03 6.62 30.29 ;
        RECT 6.36 29.27 6.62 29.53 ;
        RECT 6.36 28.51 6.62 28.77 ;
        RECT 6.36 27.75 6.62 28.01 ;
        RECT 6.36 26.99 6.62 27.25 ;
        RECT 6.36 26.23 6.62 26.49 ;
        RECT 6.36 25.47 6.62 25.73 ;
        RECT 6.36 24.71 6.62 24.97 ;
        RECT 6.36 23.95 6.62 24.21 ;
        RECT 6.36 23.19 6.62 23.45 ;
        RECT 7.12 30.03 7.38 30.29 ;
        RECT 7.12 29.27 7.38 29.53 ;
        RECT 7.12 28.51 7.38 28.77 ;
        RECT 7.12 27.75 7.38 28.01 ;
        RECT 7.12 26.99 7.38 27.25 ;
        RECT 7.12 26.23 7.38 26.49 ;
        RECT 7.12 25.47 7.38 25.73 ;
        RECT 7.12 24.71 7.38 24.97 ;
        RECT 7.12 23.95 7.38 24.21 ;
        RECT 7.12 23.19 7.38 23.45 ;
        RECT 7.88 30.03 8.14 30.29 ;
        RECT 7.88 29.27 8.14 29.53 ;
        RECT 7.88 28.51 8.14 28.77 ;
        RECT 7.88 27.75 8.14 28.01 ;
        RECT 7.88 26.99 8.14 27.25 ;
        RECT 7.88 26.23 8.14 26.49 ;
        RECT 7.88 25.47 8.14 25.73 ;
        RECT 7.88 24.71 8.14 24.97 ;
        RECT 7.88 23.95 8.14 24.21 ;
        RECT 7.88 23.19 8.14 23.45 ;
        RECT 8.64 30.03 8.9 30.29 ;
        RECT 8.64 29.27 8.9 29.53 ;
        RECT 8.64 28.51 8.9 28.77 ;
        RECT 8.64 27.75 8.9 28.01 ;
        RECT 8.64 26.99 8.9 27.25 ;
        RECT 8.64 26.23 8.9 26.49 ;
        RECT 8.64 25.47 8.9 25.73 ;
        RECT 8.64 24.71 8.9 24.97 ;
        RECT 8.64 23.95 8.9 24.21 ;
        RECT 8.64 23.19 8.9 23.45 ;
        RECT 9.4 30.03 9.66 30.29 ;
        RECT 9.4 29.27 9.66 29.53 ;
        RECT 9.4 28.51 9.66 28.77 ;
        RECT 9.4 27.75 9.66 28.01 ;
        RECT 9.4 26.99 9.66 27.25 ;
        RECT 9.4 26.23 9.66 26.49 ;
        RECT 9.4 25.47 9.66 25.73 ;
        RECT 9.4 24.71 9.66 24.97 ;
        RECT 9.4 23.95 9.66 24.21 ;
        RECT 9.4 23.19 9.66 23.45 ;
        RECT 10.16 30.03 10.42 30.29 ;
        RECT 10.16 29.27 10.42 29.53 ;
        RECT 10.16 28.51 10.42 28.77 ;
        RECT 10.16 27.75 10.42 28.01 ;
        RECT 10.16 26.99 10.42 27.25 ;
        RECT 10.16 26.23 10.42 26.49 ;
        RECT 10.16 25.47 10.42 25.73 ;
        RECT 10.16 24.71 10.42 24.97 ;
        RECT 10.16 23.95 10.42 24.21 ;
        RECT 10.16 23.19 10.42 23.45 ;
        RECT 10.92 30.03 11.18 30.29 ;
        RECT 10.92 29.27 11.18 29.53 ;
        RECT 10.92 28.51 11.18 28.77 ;
        RECT 10.92 27.75 11.18 28.01 ;
        RECT 10.92 26.99 11.18 27.25 ;
        RECT 10.92 26.23 11.18 26.49 ;
        RECT 10.92 25.47 11.18 25.73 ;
        RECT 10.92 24.71 11.18 24.97 ;
        RECT 10.92 23.95 11.18 24.21 ;
        RECT 10.92 23.19 11.18 23.45 ;
        RECT 11.68 30.03 11.94 30.29 ;
        RECT 11.68 29.27 11.94 29.53 ;
        RECT 11.68 28.51 11.94 28.77 ;
        RECT 11.68 27.75 11.94 28.01 ;
        RECT 11.68 26.99 11.94 27.25 ;
        RECT 11.68 26.23 11.94 26.49 ;
        RECT 11.68 25.47 11.94 25.73 ;
        RECT 11.68 24.71 11.94 24.97 ;
        RECT 11.68 23.95 11.94 24.21 ;
        RECT 11.68 23.19 11.94 23.45 ;
        RECT 12.44 30.03 12.7 30.29 ;
        RECT 12.44 29.27 12.7 29.53 ;
        RECT 12.44 28.51 12.7 28.77 ;
        RECT 12.44 27.75 12.7 28.01 ;
        RECT 12.44 26.99 12.7 27.25 ;
        RECT 12.44 26.23 12.7 26.49 ;
        RECT 12.44 25.47 12.7 25.73 ;
        RECT 12.44 24.71 12.7 24.97 ;
        RECT 12.44 23.95 12.7 24.21 ;
        RECT 12.44 23.19 12.7 23.45 ;
        RECT 13.2 30.03 13.46 30.29 ;
        RECT 13.2 29.27 13.46 29.53 ;
        RECT 13.2 28.51 13.46 28.77 ;
        RECT 13.2 27.75 13.46 28.01 ;
        RECT 13.2 26.99 13.46 27.25 ;
        RECT 13.2 26.23 13.46 26.49 ;
        RECT 13.2 25.47 13.46 25.73 ;
        RECT 13.2 24.71 13.46 24.97 ;
        RECT 13.2 23.95 13.46 24.21 ;
        RECT 13.2 23.19 13.46 23.45 ;
        RECT 13.96 30.03 14.22 30.29 ;
        RECT 13.96 29.27 14.22 29.53 ;
        RECT 13.96 28.51 14.22 28.77 ;
        RECT 13.96 27.75 14.22 28.01 ;
        RECT 13.96 26.99 14.22 27.25 ;
        RECT 13.96 26.23 14.22 26.49 ;
        RECT 13.96 25.47 14.22 25.73 ;
        RECT 13.96 24.71 14.22 24.97 ;
        RECT 13.96 23.95 14.22 24.21 ;
        RECT 13.96 23.19 14.22 23.45 ;
        RECT 14.72 30.03 14.98 30.29 ;
        RECT 14.72 29.27 14.98 29.53 ;
        RECT 14.72 28.51 14.98 28.77 ;
        RECT 14.72 27.75 14.98 28.01 ;
        RECT 14.72 26.99 14.98 27.25 ;
        RECT 14.72 26.23 14.98 26.49 ;
        RECT 14.72 25.47 14.98 25.73 ;
        RECT 14.72 24.71 14.98 24.97 ;
        RECT 14.72 23.95 14.98 24.21 ;
        RECT 14.72 23.19 14.98 23.45 ;
        RECT 15.48 30.03 15.74 30.29 ;
        RECT 15.48 29.27 15.74 29.53 ;
        RECT 15.48 28.51 15.74 28.77 ;
        RECT 15.48 27.75 15.74 28.01 ;
        RECT 15.48 26.99 15.74 27.25 ;
        RECT 15.48 26.23 15.74 26.49 ;
        RECT 15.48 25.47 15.74 25.73 ;
        RECT 15.48 24.71 15.74 24.97 ;
        RECT 15.48 23.95 15.74 24.21 ;
        RECT 15.48 23.19 15.74 23.45 ;
        RECT 16.24 30.03 16.5 30.29 ;
        RECT 16.24 29.27 16.5 29.53 ;
        RECT 16.24 28.51 16.5 28.77 ;
        RECT 16.24 27.75 16.5 28.01 ;
        RECT 16.24 26.99 16.5 27.25 ;
        RECT 16.24 26.23 16.5 26.49 ;
        RECT 16.24 25.47 16.5 25.73 ;
        RECT 16.24 24.71 16.5 24.97 ;
        RECT 16.24 23.95 16.5 24.21 ;
        RECT 16.24 23.19 16.5 23.45 ;
        RECT 17 30.03 17.26 30.29 ;
        RECT 17 29.27 17.26 29.53 ;
        RECT 17 28.51 17.26 28.77 ;
        RECT 17 27.75 17.26 28.01 ;
        RECT 17 26.99 17.26 27.25 ;
        RECT 17 26.23 17.26 26.49 ;
        RECT 17 25.47 17.26 25.73 ;
        RECT 17 24.71 17.26 24.97 ;
        RECT 17 23.95 17.26 24.21 ;
        RECT 17 23.19 17.26 23.45 ;
      LAYER M4 ;
        RECT 0 22 20 32 ;
      LAYER M3 ;
        RECT 0 22 20 32 ;
    END
  END AVSS
  PIN AVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER V4 ;
        RECT 2.71 17.91 2.97 18.17 ;
        RECT 2.71 17.15 2.97 17.41 ;
        RECT 2.71 16.39 2.97 16.65 ;
        RECT 2.71 15.63 2.97 15.89 ;
        RECT 2.71 14.87 2.97 15.13 ;
        RECT 2.71 14.11 2.97 14.37 ;
        RECT 2.71 13.35 2.97 13.61 ;
        RECT 2.71 12.59 2.97 12.85 ;
        RECT 2.71 11.83 2.97 12.09 ;
        RECT 2.71 11.07 2.97 11.33 ;
        RECT 3.47 17.91 3.73 18.17 ;
        RECT 3.47 17.15 3.73 17.41 ;
        RECT 3.47 16.39 3.73 16.65 ;
        RECT 3.47 15.63 3.73 15.89 ;
        RECT 3.47 14.87 3.73 15.13 ;
        RECT 3.47 14.11 3.73 14.37 ;
        RECT 3.47 13.35 3.73 13.61 ;
        RECT 3.47 12.59 3.73 12.85 ;
        RECT 3.47 11.83 3.73 12.09 ;
        RECT 3.47 11.07 3.73 11.33 ;
        RECT 4.23 17.91 4.49 18.17 ;
        RECT 4.23 17.15 4.49 17.41 ;
        RECT 4.23 16.39 4.49 16.65 ;
        RECT 4.23 15.63 4.49 15.89 ;
        RECT 4.23 14.87 4.49 15.13 ;
        RECT 4.23 14.11 4.49 14.37 ;
        RECT 4.23 13.35 4.49 13.61 ;
        RECT 4.23 12.59 4.49 12.85 ;
        RECT 4.23 11.83 4.49 12.09 ;
        RECT 4.23 11.07 4.49 11.33 ;
        RECT 4.99 17.91 5.25 18.17 ;
        RECT 4.99 17.15 5.25 17.41 ;
        RECT 4.99 16.39 5.25 16.65 ;
        RECT 4.99 15.63 5.25 15.89 ;
        RECT 4.99 14.87 5.25 15.13 ;
        RECT 4.99 14.11 5.25 14.37 ;
        RECT 4.99 13.35 5.25 13.61 ;
        RECT 4.99 12.59 5.25 12.85 ;
        RECT 4.99 11.83 5.25 12.09 ;
        RECT 4.99 11.07 5.25 11.33 ;
        RECT 5.75 17.91 6.01 18.17 ;
        RECT 5.75 17.15 6.01 17.41 ;
        RECT 5.75 16.39 6.01 16.65 ;
        RECT 5.75 15.63 6.01 15.89 ;
        RECT 5.75 14.87 6.01 15.13 ;
        RECT 5.75 14.11 6.01 14.37 ;
        RECT 5.75 13.35 6.01 13.61 ;
        RECT 5.75 12.59 6.01 12.85 ;
        RECT 5.75 11.83 6.01 12.09 ;
        RECT 5.75 11.07 6.01 11.33 ;
        RECT 6.51 17.91 6.77 18.17 ;
        RECT 6.51 17.15 6.77 17.41 ;
        RECT 6.51 16.39 6.77 16.65 ;
        RECT 6.51 15.63 6.77 15.89 ;
        RECT 6.51 14.87 6.77 15.13 ;
        RECT 6.51 14.11 6.77 14.37 ;
        RECT 6.51 13.35 6.77 13.61 ;
        RECT 6.51 12.59 6.77 12.85 ;
        RECT 6.51 11.83 6.77 12.09 ;
        RECT 6.51 11.07 6.77 11.33 ;
        RECT 7.27 17.91 7.53 18.17 ;
        RECT 7.27 17.15 7.53 17.41 ;
        RECT 7.27 16.39 7.53 16.65 ;
        RECT 7.27 15.63 7.53 15.89 ;
        RECT 7.27 14.87 7.53 15.13 ;
        RECT 7.27 14.11 7.53 14.37 ;
        RECT 7.27 13.35 7.53 13.61 ;
        RECT 7.27 12.59 7.53 12.85 ;
        RECT 7.27 11.83 7.53 12.09 ;
        RECT 7.27 11.07 7.53 11.33 ;
        RECT 8.03 17.91 8.29 18.17 ;
        RECT 8.03 17.15 8.29 17.41 ;
        RECT 8.03 16.39 8.29 16.65 ;
        RECT 8.03 15.63 8.29 15.89 ;
        RECT 8.03 14.87 8.29 15.13 ;
        RECT 8.03 14.11 8.29 14.37 ;
        RECT 8.03 13.35 8.29 13.61 ;
        RECT 8.03 12.59 8.29 12.85 ;
        RECT 8.03 11.83 8.29 12.09 ;
        RECT 8.03 11.07 8.29 11.33 ;
        RECT 8.79 17.91 9.05 18.17 ;
        RECT 8.79 17.15 9.05 17.41 ;
        RECT 8.79 16.39 9.05 16.65 ;
        RECT 8.79 15.63 9.05 15.89 ;
        RECT 8.79 14.87 9.05 15.13 ;
        RECT 8.79 14.11 9.05 14.37 ;
        RECT 8.79 13.35 9.05 13.61 ;
        RECT 8.79 12.59 9.05 12.85 ;
        RECT 8.79 11.83 9.05 12.09 ;
        RECT 8.79 11.07 9.05 11.33 ;
        RECT 9.55 17.91 9.81 18.17 ;
        RECT 9.55 17.15 9.81 17.41 ;
        RECT 9.55 16.39 9.81 16.65 ;
        RECT 9.55 15.63 9.81 15.89 ;
        RECT 9.55 14.87 9.81 15.13 ;
        RECT 9.55 14.11 9.81 14.37 ;
        RECT 9.55 13.35 9.81 13.61 ;
        RECT 9.55 12.59 9.81 12.85 ;
        RECT 9.55 11.83 9.81 12.09 ;
        RECT 9.55 11.07 9.81 11.33 ;
        RECT 10.31 17.91 10.57 18.17 ;
        RECT 10.31 17.15 10.57 17.41 ;
        RECT 10.31 16.39 10.57 16.65 ;
        RECT 10.31 15.63 10.57 15.89 ;
        RECT 10.31 14.87 10.57 15.13 ;
        RECT 10.31 14.11 10.57 14.37 ;
        RECT 10.31 13.35 10.57 13.61 ;
        RECT 10.31 12.59 10.57 12.85 ;
        RECT 10.31 11.83 10.57 12.09 ;
        RECT 10.31 11.07 10.57 11.33 ;
        RECT 11.07 17.91 11.33 18.17 ;
        RECT 11.07 17.15 11.33 17.41 ;
        RECT 11.07 16.39 11.33 16.65 ;
        RECT 11.07 15.63 11.33 15.89 ;
        RECT 11.07 14.87 11.33 15.13 ;
        RECT 11.07 14.11 11.33 14.37 ;
        RECT 11.07 13.35 11.33 13.61 ;
        RECT 11.07 12.59 11.33 12.85 ;
        RECT 11.07 11.83 11.33 12.09 ;
        RECT 11.07 11.07 11.33 11.33 ;
        RECT 11.83 17.91 12.09 18.17 ;
        RECT 11.83 17.15 12.09 17.41 ;
        RECT 11.83 16.39 12.09 16.65 ;
        RECT 11.83 15.63 12.09 15.89 ;
        RECT 11.83 14.87 12.09 15.13 ;
        RECT 11.83 14.11 12.09 14.37 ;
        RECT 11.83 13.35 12.09 13.61 ;
        RECT 11.83 12.59 12.09 12.85 ;
        RECT 11.83 11.83 12.09 12.09 ;
        RECT 11.83 11.07 12.09 11.33 ;
        RECT 12.59 17.91 12.85 18.17 ;
        RECT 12.59 17.15 12.85 17.41 ;
        RECT 12.59 16.39 12.85 16.65 ;
        RECT 12.59 15.63 12.85 15.89 ;
        RECT 12.59 14.87 12.85 15.13 ;
        RECT 12.59 14.11 12.85 14.37 ;
        RECT 12.59 13.35 12.85 13.61 ;
        RECT 12.59 12.59 12.85 12.85 ;
        RECT 12.59 11.83 12.85 12.09 ;
        RECT 12.59 11.07 12.85 11.33 ;
        RECT 13.35 17.91 13.61 18.17 ;
        RECT 13.35 17.15 13.61 17.41 ;
        RECT 13.35 16.39 13.61 16.65 ;
        RECT 13.35 15.63 13.61 15.89 ;
        RECT 13.35 14.87 13.61 15.13 ;
        RECT 13.35 14.11 13.61 14.37 ;
        RECT 13.35 13.35 13.61 13.61 ;
        RECT 13.35 12.59 13.61 12.85 ;
        RECT 13.35 11.83 13.61 12.09 ;
        RECT 13.35 11.07 13.61 11.33 ;
        RECT 14.11 17.91 14.37 18.17 ;
        RECT 14.11 17.15 14.37 17.41 ;
        RECT 14.11 16.39 14.37 16.65 ;
        RECT 14.11 15.63 14.37 15.89 ;
        RECT 14.11 14.87 14.37 15.13 ;
        RECT 14.11 14.11 14.37 14.37 ;
        RECT 14.11 13.35 14.37 13.61 ;
        RECT 14.11 12.59 14.37 12.85 ;
        RECT 14.11 11.83 14.37 12.09 ;
        RECT 14.11 11.07 14.37 11.33 ;
        RECT 14.87 17.91 15.13 18.17 ;
        RECT 14.87 17.15 15.13 17.41 ;
        RECT 14.87 16.39 15.13 16.65 ;
        RECT 14.87 15.63 15.13 15.89 ;
        RECT 14.87 14.87 15.13 15.13 ;
        RECT 14.87 14.11 15.13 14.37 ;
        RECT 14.87 13.35 15.13 13.61 ;
        RECT 14.87 12.59 15.13 12.85 ;
        RECT 14.87 11.83 15.13 12.09 ;
        RECT 14.87 11.07 15.13 11.33 ;
        RECT 15.63 17.91 15.89 18.17 ;
        RECT 15.63 17.15 15.89 17.41 ;
        RECT 15.63 16.39 15.89 16.65 ;
        RECT 15.63 15.63 15.89 15.89 ;
        RECT 15.63 14.87 15.89 15.13 ;
        RECT 15.63 14.11 15.89 14.37 ;
        RECT 15.63 13.35 15.89 13.61 ;
        RECT 15.63 12.59 15.89 12.85 ;
        RECT 15.63 11.83 15.89 12.09 ;
        RECT 15.63 11.07 15.89 11.33 ;
        RECT 16.39 17.91 16.65 18.17 ;
        RECT 16.39 17.15 16.65 17.41 ;
        RECT 16.39 16.39 16.65 16.65 ;
        RECT 16.39 15.63 16.65 15.89 ;
        RECT 16.39 14.87 16.65 15.13 ;
        RECT 16.39 14.11 16.65 14.37 ;
        RECT 16.39 13.35 16.65 13.61 ;
        RECT 16.39 12.59 16.65 12.85 ;
        RECT 16.39 11.83 16.65 12.09 ;
        RECT 16.39 11.07 16.65 11.33 ;
        RECT 17.15 17.91 17.41 18.17 ;
        RECT 17.15 17.15 17.41 17.41 ;
        RECT 17.15 16.39 17.41 16.65 ;
        RECT 17.15 15.63 17.41 15.89 ;
        RECT 17.15 14.87 17.41 15.13 ;
        RECT 17.15 14.11 17.41 14.37 ;
        RECT 17.15 13.35 17.41 13.61 ;
        RECT 17.15 12.59 17.41 12.85 ;
        RECT 17.15 11.83 17.41 12.09 ;
        RECT 17.15 11.07 17.41 11.33 ;
      LAYER M4 ;
        RECT 0 10 20 20 ;
      LAYER M3 ;
        RECT 0 10 20 20 ;
    END
  END AVDD
  PIN SUB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER V4 ;
        RECT 2.855 6.76 3.115 7.02 ;
        RECT 2.855 6 3.115 6.26 ;
        RECT 2.855 5.24 3.115 5.5 ;
        RECT 2.855 4.48 3.115 4.74 ;
        RECT 3.615 6.76 3.875 7.02 ;
        RECT 3.615 6 3.875 6.26 ;
        RECT 3.615 5.24 3.875 5.5 ;
        RECT 3.615 4.48 3.875 4.74 ;
        RECT 4.375 6.76 4.635 7.02 ;
        RECT 4.375 6 4.635 6.26 ;
        RECT 4.375 5.24 4.635 5.5 ;
        RECT 4.375 4.48 4.635 4.74 ;
        RECT 5.135 6.76 5.395 7.02 ;
        RECT 5.135 6 5.395 6.26 ;
        RECT 5.135 5.24 5.395 5.5 ;
        RECT 5.135 4.48 5.395 4.74 ;
        RECT 5.895 6.76 6.155 7.02 ;
        RECT 5.895 6 6.155 6.26 ;
        RECT 5.895 5.24 6.155 5.5 ;
        RECT 5.895 4.48 6.155 4.74 ;
        RECT 6.655 6.76 6.915 7.02 ;
        RECT 6.655 6 6.915 6.26 ;
        RECT 6.655 5.24 6.915 5.5 ;
        RECT 6.655 4.48 6.915 4.74 ;
        RECT 7.415 6.76 7.675 7.02 ;
        RECT 7.415 6 7.675 6.26 ;
        RECT 7.415 5.24 7.675 5.5 ;
        RECT 7.415 4.48 7.675 4.74 ;
        RECT 8.175 6.76 8.435 7.02 ;
        RECT 8.175 6 8.435 6.26 ;
        RECT 8.175 5.24 8.435 5.5 ;
        RECT 8.175 4.48 8.435 4.74 ;
        RECT 8.935 6.76 9.195 7.02 ;
        RECT 8.935 6 9.195 6.26 ;
        RECT 8.935 5.24 9.195 5.5 ;
        RECT 8.935 4.48 9.195 4.74 ;
        RECT 9.695 6.76 9.955 7.02 ;
        RECT 9.695 6 9.955 6.26 ;
        RECT 9.695 5.24 9.955 5.5 ;
        RECT 9.695 4.48 9.955 4.74 ;
        RECT 10.455 6.76 10.715 7.02 ;
        RECT 10.455 6 10.715 6.26 ;
        RECT 10.455 5.24 10.715 5.5 ;
        RECT 10.455 4.48 10.715 4.74 ;
        RECT 11.215 6.76 11.475 7.02 ;
        RECT 11.215 6 11.475 6.26 ;
        RECT 11.215 5.24 11.475 5.5 ;
        RECT 11.215 4.48 11.475 4.74 ;
        RECT 11.975 6.76 12.235 7.02 ;
        RECT 11.975 6 12.235 6.26 ;
        RECT 11.975 5.24 12.235 5.5 ;
        RECT 11.975 4.48 12.235 4.74 ;
        RECT 12.735 6.76 12.995 7.02 ;
        RECT 12.735 6 12.995 6.26 ;
        RECT 12.735 5.24 12.995 5.5 ;
        RECT 12.735 4.48 12.995 4.74 ;
        RECT 13.495 6.76 13.755 7.02 ;
        RECT 13.495 6 13.755 6.26 ;
        RECT 13.495 5.24 13.755 5.5 ;
        RECT 13.495 4.48 13.755 4.74 ;
        RECT 14.255 6.76 14.515 7.02 ;
        RECT 14.255 6 14.515 6.26 ;
        RECT 14.255 5.24 14.515 5.5 ;
        RECT 14.255 4.48 14.515 4.74 ;
        RECT 15.015 6.76 15.275 7.02 ;
        RECT 15.015 6 15.275 6.26 ;
        RECT 15.015 5.24 15.275 5.5 ;
        RECT 15.015 4.48 15.275 4.74 ;
        RECT 15.775 6.76 16.035 7.02 ;
        RECT 15.775 6 16.035 6.26 ;
        RECT 15.775 5.24 16.035 5.5 ;
        RECT 15.775 4.48 16.035 4.74 ;
        RECT 16.535 6.76 16.795 7.02 ;
        RECT 16.535 6 16.795 6.26 ;
        RECT 16.535 5.24 16.795 5.5 ;
        RECT 16.535 4.48 16.795 4.74 ;
        RECT 17.295 6.76 17.555 7.02 ;
        RECT 17.295 6 17.555 6.26 ;
        RECT 17.295 5.24 17.555 5.5 ;
        RECT 17.295 4.48 17.555 4.74 ;
      LAYER V3 ;
        RECT 19.28 4.26 19.54 4.52 ;
        RECT 19.28 4.78 19.54 5.04 ;
        RECT 19.28 5.3 19.54 5.56 ;
        RECT 19.28 5.82 19.54 6.08 ;
        RECT 19.28 6.34 19.54 6.6 ;
        RECT 19.28 6.86 19.54 7.12 ;
        RECT 19.28 7.38 19.54 7.64 ;
        RECT 0.46 4.26 0.72 4.52 ;
        RECT 0.46 4.78 0.72 5.04 ;
        RECT 0.46 5.3 0.72 5.56 ;
        RECT 0.46 5.82 0.72 6.08 ;
        RECT 0.46 6.34 0.72 6.6 ;
        RECT 0.46 6.86 0.72 7.12 ;
        RECT 0.46 7.38 0.72 7.64 ;
      LAYER M4 ;
        RECT 0 4 20 8 ;
      LAYER M3 ;
        RECT 0 4 20 8 ;
    END
  END SUB
  OBS
    LAYER M1 ;
      RECT 6.36 5.65 7.17 5.99 ;
      RECT 8.99 5.65 9.8 5.99 ;
      RECT 11.62 5.65 12.43 5.99 ;
      RECT 6.36 5.65 6.66 6.91 ;
      RECT 5.9 6.61 6.66 6.91 ;
      RECT 8.99 5.65 9.29 6.91 ;
      RECT 8.53 6.61 9.29 6.91 ;
      RECT 11.62 5.65 11.92 6.91 ;
      RECT 11.16 6.61 11.92 6.91 ;
      RECT 1.5 8.245 14.965 9.245 ;
      RECT 5.9 6.61 6.2 10.88 ;
      RECT 8.53 6.61 8.91 10.88 ;
      RECT 11.16 6.61 11.54 10.88 ;
      RECT 5.9 10.58 6.66 10.88 ;
      RECT 8.53 10.58 9.29 10.88 ;
      RECT 11.16 10.58 11.92 10.88 ;
      RECT 13.825 6.61 14.17 10.88 ;
      RECT 6.36 10.58 6.66 11.84 ;
      RECT 8.99 10.58 9.29 11.84 ;
      RECT 11.62 10.58 11.92 11.84 ;
      RECT 6.36 11.5 7.17 11.84 ;
      RECT 8.99 11.5 9.8 11.84 ;
      RECT 11.62 11.5 12.43 11.84 ;
      RECT 6.36 17.03 7.17 17.37 ;
      RECT 8.99 17.03 9.8 17.37 ;
      RECT 11.62 17.03 12.43 17.37 ;
      RECT 6.36 17.03 6.66 18.29 ;
      RECT 5.9 17.99 6.66 18.29 ;
      RECT 8.99 17.03 9.29 18.29 ;
      RECT 8.53 17.99 9.29 18.29 ;
      RECT 11.62 17.03 11.92 18.29 ;
      RECT 11.16 17.99 11.92 18.29 ;
      RECT 1.5 19.625 14.965 20.625 ;
      RECT 5.9 17.99 6.2 22.26 ;
      RECT 8.53 17.99 8.91 22.26 ;
      RECT 11.16 17.99 11.54 22.26 ;
      RECT 5.9 21.96 6.66 22.26 ;
      RECT 8.53 21.96 9.29 22.26 ;
      RECT 11.16 21.96 11.92 22.26 ;
      RECT 13.825 17.99 14.17 22.26 ;
      RECT 6.36 21.96 6.66 23.22 ;
      RECT 8.99 21.96 9.29 23.22 ;
      RECT 11.62 21.96 11.92 23.22 ;
      RECT 6.36 22.88 7.17 23.22 ;
      RECT 8.99 22.88 9.8 23.22 ;
      RECT 11.62 22.88 12.43 23.22 ;
      RECT 6.36 28.41 7.17 28.75 ;
      RECT 8.99 28.41 9.8 28.75 ;
      RECT 11.62 28.41 12.43 28.75 ;
      RECT 6.36 28.41 6.66 29.67 ;
      RECT 5.9 29.37 6.66 29.67 ;
      RECT 8.99 28.41 9.29 29.67 ;
      RECT 8.53 29.37 9.29 29.67 ;
      RECT 11.62 28.41 11.92 29.67 ;
      RECT 11.16 29.37 11.92 29.67 ;
      RECT 1.5 31.005 14.965 32.005 ;
      RECT 5.9 29.37 6.2 33.64 ;
      RECT 8.53 29.37 8.91 33.64 ;
      RECT 11.16 29.37 11.54 33.64 ;
      RECT 5.9 33.34 6.66 33.64 ;
      RECT 8.53 33.34 9.29 33.64 ;
      RECT 11.16 33.34 11.92 33.64 ;
      RECT 13.825 29.37 14.17 33.64 ;
      RECT 6.36 33.34 6.66 34.6 ;
      RECT 8.99 33.34 9.29 34.6 ;
      RECT 11.62 33.34 11.92 34.6 ;
      RECT 6.36 34.26 7.17 34.6 ;
      RECT 8.99 34.26 9.8 34.6 ;
      RECT 11.62 34.26 12.43 34.6 ;
      RECT 6.36 39.79 7.17 40.13 ;
      RECT 8.99 39.79 9.8 40.13 ;
      RECT 11.62 39.79 12.43 40.13 ;
      RECT 6.36 39.79 6.66 41.05 ;
      RECT 5.9 40.75 6.66 41.05 ;
      RECT 8.99 39.79 9.29 41.05 ;
      RECT 8.53 40.75 9.29 41.05 ;
      RECT 11.62 39.79 11.92 41.05 ;
      RECT 11.16 40.75 11.92 41.05 ;
      RECT 1.5 42.385 14.965 43.385 ;
      RECT 5.9 40.75 6.2 45.02 ;
      RECT 8.53 40.75 8.91 45.02 ;
      RECT 11.16 40.75 11.54 45.02 ;
      RECT 5.9 44.72 6.66 45.02 ;
      RECT 8.53 44.72 9.29 45.02 ;
      RECT 11.16 44.72 11.92 45.02 ;
      RECT 13.825 40.75 14.17 45.02 ;
      RECT 6.36 44.72 6.66 45.98 ;
      RECT 8.99 44.72 9.29 45.98 ;
      RECT 11.62 44.72 11.92 45.98 ;
      RECT 6.36 45.64 7.17 45.98 ;
      RECT 8.99 45.64 9.8 45.98 ;
      RECT 11.62 45.64 12.43 45.98 ;
      RECT 6.36 51.17 7.17 51.51 ;
      RECT 8.99 51.17 9.8 51.51 ;
      RECT 11.62 51.17 12.43 51.51 ;
      RECT 6.36 51.17 6.66 52.43 ;
      RECT 5.9 52.13 6.66 52.43 ;
      RECT 8.99 51.17 9.29 52.43 ;
      RECT 8.53 52.13 9.29 52.43 ;
      RECT 11.62 51.17 11.92 52.43 ;
      RECT 11.16 52.13 11.92 52.43 ;
      RECT 1.5 53.765 14.965 54.765 ;
      RECT 5.9 52.13 6.2 56.4 ;
      RECT 8.53 52.13 8.91 56.4 ;
      RECT 11.16 52.13 11.54 56.4 ;
      RECT 5.9 56.1 6.66 56.4 ;
      RECT 8.53 56.1 9.29 56.4 ;
      RECT 11.16 56.1 11.92 56.4 ;
      RECT 13.825 52.13 14.17 56.4 ;
      RECT 6.36 56.1 6.66 57.36 ;
      RECT 8.99 56.1 9.29 57.36 ;
      RECT 11.62 56.1 11.92 57.36 ;
      RECT 6.36 57.02 7.17 57.36 ;
      RECT 8.99 57.02 9.8 57.36 ;
      RECT 11.62 57.02 12.43 57.36 ;
      RECT 6.36 62.55 7.17 62.89 ;
      RECT 8.99 62.55 9.8 62.89 ;
      RECT 11.62 62.55 12.43 62.89 ;
      RECT 6.36 62.55 6.66 63.81 ;
      RECT 5.9 63.51 6.66 63.81 ;
      RECT 8.99 62.55 9.29 63.81 ;
      RECT 8.53 63.51 9.29 63.81 ;
      RECT 11.62 62.55 11.92 63.81 ;
      RECT 11.16 63.51 11.92 63.81 ;
      RECT 1.5 65.145 14.965 66.145 ;
      RECT 5.9 63.51 6.2 67.78 ;
      RECT 8.53 63.51 8.91 67.78 ;
      RECT 11.16 63.51 11.54 67.78 ;
      RECT 5.9 67.48 6.66 67.78 ;
      RECT 8.53 67.48 9.29 67.78 ;
      RECT 11.16 67.48 11.92 67.78 ;
      RECT 13.825 63.51 14.17 67.78 ;
      RECT 6.36 67.48 6.66 68.74 ;
      RECT 8.99 67.48 9.29 68.74 ;
      RECT 11.62 67.48 11.92 68.74 ;
      RECT 6.36 68.4 7.17 68.74 ;
      RECT 8.99 68.4 9.8 68.74 ;
      RECT 11.62 68.4 12.43 68.74 ;
      RECT 6.36 73.93 7.17 74.27 ;
      RECT 8.99 73.93 9.8 74.27 ;
      RECT 11.62 73.93 12.43 74.27 ;
      RECT 6.36 73.93 6.66 75.19 ;
      RECT 5.9 74.89 6.66 75.19 ;
      RECT 8.99 73.93 9.29 75.19 ;
      RECT 8.53 74.89 9.29 75.19 ;
      RECT 11.62 73.93 11.92 75.19 ;
      RECT 11.16 74.89 11.92 75.19 ;
      RECT 1.5 76.525 14.965 77.525 ;
      RECT 5.9 74.89 6.2 79.16 ;
      RECT 8.53 74.89 8.91 79.16 ;
      RECT 11.16 74.89 11.54 79.16 ;
      RECT 5.9 78.86 6.66 79.16 ;
      RECT 8.53 78.86 9.29 79.16 ;
      RECT 11.16 78.86 11.92 79.16 ;
      RECT 13.825 74.89 14.17 79.16 ;
      RECT 6.36 78.86 6.66 80.12 ;
      RECT 8.99 78.86 9.29 80.12 ;
      RECT 11.62 78.86 11.92 80.12 ;
      RECT 6.36 79.78 7.17 80.12 ;
      RECT 8.99 79.78 9.8 80.12 ;
      RECT 11.62 79.78 12.43 80.12 ;
      RECT 6.36 85.31 7.17 85.65 ;
      RECT 8.99 85.31 9.8 85.65 ;
      RECT 11.62 85.31 12.43 85.65 ;
      RECT 6.36 85.31 6.66 86.57 ;
      RECT 5.9 86.27 6.66 86.57 ;
      RECT 8.99 85.31 9.29 86.57 ;
      RECT 8.53 86.27 9.29 86.57 ;
      RECT 11.62 85.31 11.92 86.57 ;
      RECT 11.16 86.27 11.92 86.57 ;
      RECT 1.5 87.905 14.965 88.905 ;
      RECT 5.9 86.27 6.2 90.54 ;
      RECT 8.53 86.27 8.91 90.54 ;
      RECT 11.16 86.27 11.54 90.54 ;
      RECT 5.9 90.24 6.66 90.54 ;
      RECT 8.53 90.24 9.29 90.54 ;
      RECT 11.16 90.24 11.92 90.54 ;
      RECT 13.825 86.27 14.17 90.54 ;
      RECT 6.36 90.24 6.66 91.5 ;
      RECT 8.99 90.24 9.29 91.5 ;
      RECT 11.62 90.24 11.92 91.5 ;
      RECT 6.36 91.16 7.17 91.5 ;
      RECT 8.99 91.16 9.8 91.5 ;
      RECT 11.62 91.16 12.43 91.5 ;
      RECT 6.36 96.69 7.17 97.03 ;
      RECT 8.99 96.69 9.8 97.03 ;
      RECT 11.62 96.69 12.43 97.03 ;
      RECT 6.36 96.69 6.66 97.95 ;
      RECT 5.9 97.65 6.66 97.95 ;
      RECT 8.99 96.69 9.29 97.95 ;
      RECT 8.53 97.65 9.29 97.95 ;
      RECT 11.62 96.69 11.92 97.95 ;
      RECT 11.16 97.65 11.92 97.95 ;
      RECT 1.5 99.285 14.965 100.285 ;
      RECT 5.9 97.65 6.2 101.92 ;
      RECT 8.53 97.65 8.91 101.92 ;
      RECT 11.16 97.65 11.54 101.92 ;
      RECT 5.9 101.62 6.66 101.92 ;
      RECT 8.53 101.62 9.29 101.92 ;
      RECT 11.16 101.62 11.92 101.92 ;
      RECT 13.825 97.65 14.17 101.92 ;
      RECT 6.36 101.62 6.66 102.88 ;
      RECT 8.99 101.62 9.29 102.88 ;
      RECT 11.62 101.62 11.92 102.88 ;
      RECT 6.36 102.54 7.17 102.88 ;
      RECT 8.99 102.54 9.8 102.88 ;
      RECT 11.62 102.54 12.43 102.88 ;
      RECT 6.36 108.07 7.17 108.41 ;
      RECT 8.99 108.07 9.8 108.41 ;
      RECT 11.62 108.07 12.43 108.41 ;
      RECT 6.36 108.07 6.66 109.33 ;
      RECT 5.9 109.03 6.66 109.33 ;
      RECT 8.99 108.07 9.29 109.33 ;
      RECT 8.53 109.03 9.29 109.33 ;
      RECT 11.62 108.07 11.92 109.33 ;
      RECT 11.16 109.03 11.92 109.33 ;
      RECT 1.5 8.245 2.5 111.665 ;
      RECT 1.5 110.665 14.965 111.665 ;
      RECT 5.9 109.03 6.2 113.3 ;
      RECT 8.53 109.03 8.91 113.3 ;
      RECT 11.16 109.03 11.54 113.3 ;
      RECT 5.9 113 6.66 113.3 ;
      RECT 8.53 113 9.29 113.3 ;
      RECT 11.16 113 11.92 113.3 ;
      RECT 13.825 109.03 14.17 113.3 ;
      RECT 6.36 113 6.66 114.26 ;
      RECT 8.99 113 9.29 114.26 ;
      RECT 11.62 113 11.92 114.26 ;
      RECT 6.36 113.92 7.17 114.26 ;
      RECT 8.99 113.92 9.8 114.26 ;
      RECT 11.62 113.92 12.43 114.26 ;
      RECT 5.035 2.555 18.5 3.555 ;
      RECT 5.9 2.555 6.2 5.35 ;
      RECT 8.53 2.555 8.83 5.35 ;
      RECT 8.07 5.05 8.83 5.35 ;
      RECT 11.16 2.555 11.46 5.35 ;
      RECT 10.7 5.05 11.46 5.35 ;
      RECT 13.79 2.555 14.09 5.35 ;
      RECT 13.33 5.05 14.09 5.35 ;
      RECT 8.07 5.05 8.37 6.31 ;
      RECT 7.56 5.97 8.37 6.31 ;
      RECT 10.7 5.05 11 6.31 ;
      RECT 10.19 5.97 11 6.31 ;
      RECT 13.33 5.05 13.63 6.31 ;
      RECT 12.82 5.97 13.63 6.31 ;
      RECT 7.56 11.18 8.37 11.52 ;
      RECT 10.19 11.18 11 11.52 ;
      RECT 12.82 11.18 13.63 11.52 ;
      RECT 8.07 11.18 8.37 12.44 ;
      RECT 10.7 11.18 11 12.44 ;
      RECT 13.33 11.18 13.63 12.44 ;
      RECT 8.07 12.14 8.83 12.44 ;
      RECT 10.7 12.14 11.46 12.44 ;
      RECT 13.33 12.14 14.09 12.44 ;
      RECT 5.035 13.935 18.5 14.935 ;
      RECT 5.9 12.14 6.2 16.73 ;
      RECT 8.53 12.14 8.83 16.73 ;
      RECT 8.07 16.43 8.83 16.73 ;
      RECT 11.16 12.14 11.46 16.73 ;
      RECT 10.7 16.43 11.46 16.73 ;
      RECT 13.79 12.14 14.09 16.73 ;
      RECT 13.33 16.43 14.09 16.73 ;
      RECT 8.07 16.43 8.37 17.69 ;
      RECT 7.56 17.35 8.37 17.69 ;
      RECT 10.7 16.43 11 17.69 ;
      RECT 10.19 17.35 11 17.69 ;
      RECT 13.33 16.43 13.63 17.69 ;
      RECT 12.82 17.35 13.63 17.69 ;
      RECT 7.56 22.56 8.37 22.9 ;
      RECT 10.19 22.56 11 22.9 ;
      RECT 12.82 22.56 13.63 22.9 ;
      RECT 8.07 22.56 8.37 23.82 ;
      RECT 10.7 22.56 11 23.82 ;
      RECT 13.33 22.56 13.63 23.82 ;
      RECT 8.07 23.52 8.83 23.82 ;
      RECT 10.7 23.52 11.46 23.82 ;
      RECT 13.33 23.52 14.09 23.82 ;
      RECT 5.035 25.315 18.5 26.315 ;
      RECT 5.9 23.52 6.2 28.11 ;
      RECT 8.53 23.52 8.83 28.11 ;
      RECT 8.07 27.81 8.83 28.11 ;
      RECT 11.16 23.52 11.46 28.11 ;
      RECT 10.7 27.81 11.46 28.11 ;
      RECT 13.79 23.52 14.09 28.11 ;
      RECT 13.33 27.81 14.09 28.11 ;
      RECT 8.07 27.81 8.37 29.07 ;
      RECT 7.56 28.73 8.37 29.07 ;
      RECT 10.7 27.81 11 29.07 ;
      RECT 10.19 28.73 11 29.07 ;
      RECT 13.33 27.81 13.63 29.07 ;
      RECT 12.82 28.73 13.63 29.07 ;
      RECT 7.56 33.94 8.37 34.28 ;
      RECT 10.19 33.94 11 34.28 ;
      RECT 12.82 33.94 13.63 34.28 ;
      RECT 8.07 33.94 8.37 35.2 ;
      RECT 10.7 33.94 11 35.2 ;
      RECT 13.33 33.94 13.63 35.2 ;
      RECT 8.07 34.9 8.83 35.2 ;
      RECT 10.7 34.9 11.46 35.2 ;
      RECT 13.33 34.9 14.09 35.2 ;
      RECT 5.035 36.695 18.5 37.695 ;
      RECT 5.9 34.9 6.2 39.49 ;
      RECT 8.53 34.9 8.83 39.49 ;
      RECT 8.07 39.19 8.83 39.49 ;
      RECT 11.16 34.9 11.46 39.49 ;
      RECT 10.7 39.19 11.46 39.49 ;
      RECT 13.79 34.9 14.09 39.49 ;
      RECT 13.33 39.19 14.09 39.49 ;
      RECT 8.07 39.19 8.37 40.45 ;
      RECT 7.56 40.11 8.37 40.45 ;
      RECT 10.7 39.19 11 40.45 ;
      RECT 10.19 40.11 11 40.45 ;
      RECT 13.33 39.19 13.63 40.45 ;
      RECT 12.82 40.11 13.63 40.45 ;
      RECT 7.56 45.32 8.37 45.66 ;
      RECT 10.19 45.32 11 45.66 ;
      RECT 12.82 45.32 13.63 45.66 ;
      RECT 8.07 45.32 8.37 46.58 ;
      RECT 10.7 45.32 11 46.58 ;
      RECT 13.33 45.32 13.63 46.58 ;
      RECT 8.07 46.28 8.83 46.58 ;
      RECT 10.7 46.28 11.46 46.58 ;
      RECT 13.33 46.28 14.09 46.58 ;
      RECT 5.035 48.075 18.5 49.075 ;
      RECT 5.9 46.28 6.2 50.87 ;
      RECT 8.53 46.28 8.83 50.87 ;
      RECT 8.07 50.57 8.83 50.87 ;
      RECT 11.16 46.28 11.46 50.87 ;
      RECT 10.7 50.57 11.46 50.87 ;
      RECT 13.79 46.28 14.09 50.87 ;
      RECT 13.33 50.57 14.09 50.87 ;
      RECT 8.07 50.57 8.37 51.83 ;
      RECT 7.56 51.49 8.37 51.83 ;
      RECT 10.7 50.57 11 51.83 ;
      RECT 10.19 51.49 11 51.83 ;
      RECT 13.33 50.57 13.63 51.83 ;
      RECT 12.82 51.49 13.63 51.83 ;
      RECT 7.56 56.7 8.37 57.04 ;
      RECT 10.19 56.7 11 57.04 ;
      RECT 12.82 56.7 13.63 57.04 ;
      RECT 8.07 56.7 8.37 57.96 ;
      RECT 10.7 56.7 11 57.96 ;
      RECT 13.33 56.7 13.63 57.96 ;
      RECT 8.07 57.66 8.83 57.96 ;
      RECT 10.7 57.66 11.46 57.96 ;
      RECT 13.33 57.66 14.09 57.96 ;
      RECT 5.035 59.455 18.5 60.455 ;
      RECT 5.9 57.66 6.2 62.25 ;
      RECT 8.53 57.66 8.83 62.25 ;
      RECT 8.07 61.95 8.83 62.25 ;
      RECT 11.16 57.66 11.46 62.25 ;
      RECT 10.7 61.95 11.46 62.25 ;
      RECT 13.79 57.66 14.09 62.25 ;
      RECT 13.33 61.95 14.09 62.25 ;
      RECT 8.07 61.95 8.37 63.21 ;
      RECT 7.56 62.87 8.37 63.21 ;
      RECT 10.7 61.95 11 63.21 ;
      RECT 10.19 62.87 11 63.21 ;
      RECT 13.33 61.95 13.63 63.21 ;
      RECT 12.82 62.87 13.63 63.21 ;
      RECT 7.56 68.08 8.37 68.42 ;
      RECT 10.19 68.08 11 68.42 ;
      RECT 12.82 68.08 13.63 68.42 ;
      RECT 8.07 68.08 8.37 69.34 ;
      RECT 10.7 68.08 11 69.34 ;
      RECT 13.33 68.08 13.63 69.34 ;
      RECT 8.07 69.04 8.83 69.34 ;
      RECT 10.7 69.04 11.46 69.34 ;
      RECT 13.33 69.04 14.09 69.34 ;
      RECT 5.035 70.835 18.5 71.835 ;
      RECT 5.9 69.04 6.2 73.63 ;
      RECT 8.53 69.04 8.83 73.63 ;
      RECT 8.07 73.33 8.83 73.63 ;
      RECT 11.16 69.04 11.46 73.63 ;
      RECT 10.7 73.33 11.46 73.63 ;
      RECT 13.79 69.04 14.09 73.63 ;
      RECT 13.33 73.33 14.09 73.63 ;
      RECT 8.07 73.33 8.37 74.59 ;
      RECT 7.56 74.25 8.37 74.59 ;
      RECT 10.7 73.33 11 74.59 ;
      RECT 10.19 74.25 11 74.59 ;
      RECT 13.33 73.33 13.63 74.59 ;
      RECT 12.82 74.25 13.63 74.59 ;
      RECT 7.56 79.46 8.37 79.8 ;
      RECT 10.19 79.46 11 79.8 ;
      RECT 12.82 79.46 13.63 79.8 ;
      RECT 8.07 79.46 8.37 80.72 ;
      RECT 10.7 79.46 11 80.72 ;
      RECT 13.33 79.46 13.63 80.72 ;
      RECT 8.07 80.42 8.83 80.72 ;
      RECT 10.7 80.42 11.46 80.72 ;
      RECT 13.33 80.42 14.09 80.72 ;
      RECT 5.035 82.215 18.5 83.215 ;
      RECT 5.9 80.42 6.2 85.01 ;
      RECT 8.53 80.42 8.83 85.01 ;
      RECT 8.07 84.71 8.83 85.01 ;
      RECT 11.16 80.42 11.46 85.01 ;
      RECT 10.7 84.71 11.46 85.01 ;
      RECT 13.79 80.42 14.09 85.01 ;
      RECT 13.33 84.71 14.09 85.01 ;
      RECT 8.07 84.71 8.37 85.97 ;
      RECT 7.56 85.63 8.37 85.97 ;
      RECT 10.7 84.71 11 85.97 ;
      RECT 10.19 85.63 11 85.97 ;
      RECT 13.33 84.71 13.63 85.97 ;
      RECT 12.82 85.63 13.63 85.97 ;
      RECT 7.56 90.84 8.37 91.18 ;
      RECT 10.19 90.84 11 91.18 ;
      RECT 12.82 90.84 13.63 91.18 ;
      RECT 8.07 90.84 8.37 92.1 ;
      RECT 10.7 90.84 11 92.1 ;
      RECT 13.33 90.84 13.63 92.1 ;
      RECT 8.07 91.8 8.83 92.1 ;
      RECT 10.7 91.8 11.46 92.1 ;
      RECT 13.33 91.8 14.09 92.1 ;
      RECT 5.035 93.595 18.5 94.595 ;
      RECT 5.9 91.8 6.2 96.39 ;
      RECT 8.53 91.8 8.83 96.39 ;
      RECT 8.07 96.09 8.83 96.39 ;
      RECT 11.16 91.8 11.46 96.39 ;
      RECT 10.7 96.09 11.46 96.39 ;
      RECT 13.79 91.8 14.09 96.39 ;
      RECT 13.33 96.09 14.09 96.39 ;
      RECT 8.07 96.09 8.37 97.35 ;
      RECT 7.56 97.01 8.37 97.35 ;
      RECT 10.7 96.09 11 97.35 ;
      RECT 10.19 97.01 11 97.35 ;
      RECT 13.33 96.09 13.63 97.35 ;
      RECT 12.82 97.01 13.63 97.35 ;
      RECT 7.56 102.22 8.37 102.56 ;
      RECT 10.19 102.22 11 102.56 ;
      RECT 12.82 102.22 13.63 102.56 ;
      RECT 8.07 102.22 8.37 103.48 ;
      RECT 10.7 102.22 11 103.48 ;
      RECT 13.33 102.22 13.63 103.48 ;
      RECT 8.07 103.18 8.83 103.48 ;
      RECT 10.7 103.18 11.46 103.48 ;
      RECT 13.33 103.18 14.09 103.48 ;
      RECT 5.035 104.975 18.5 105.975 ;
      RECT 5.9 103.18 6.2 107.77 ;
      RECT 8.53 103.18 8.83 107.77 ;
      RECT 8.07 107.47 8.83 107.77 ;
      RECT 11.16 103.18 11.46 107.77 ;
      RECT 10.7 107.47 11.46 107.77 ;
      RECT 13.79 103.18 14.09 107.77 ;
      RECT 13.33 107.47 14.09 107.77 ;
      RECT 8.07 107.47 8.37 108.73 ;
      RECT 7.56 108.39 8.37 108.73 ;
      RECT 10.7 107.47 11 108.73 ;
      RECT 10.19 108.39 11 108.73 ;
      RECT 13.33 107.47 13.63 108.73 ;
      RECT 12.82 108.39 13.63 108.73 ;
      RECT 7.56 113.6 8.37 113.94 ;
      RECT 10.19 113.6 11 113.94 ;
      RECT 12.82 113.6 13.63 113.94 ;
      RECT 8.07 113.6 8.37 114.86 ;
      RECT 10.7 113.6 11 114.86 ;
      RECT 13.33 113.6 13.63 114.86 ;
      RECT 8.07 114.56 8.83 114.86 ;
      RECT 10.7 114.56 11.46 114.86 ;
      RECT 13.33 114.56 14.09 114.86 ;
      RECT 5.9 114.56 6.2 117.355 ;
      RECT 8.53 114.56 8.83 117.355 ;
      RECT 11.16 114.56 11.46 117.355 ;
      RECT 13.79 114.56 14.09 117.355 ;
      RECT 17.5 2.555 18.5 117.355 ;
      RECT 5.035 116.355 18.5 117.355 ;
      RECT 0.42 0.42 19.58 0.76 ;
      RECT 0.42 0.42 0.76 119.58 ;
      RECT 19.24 0.42 19.58 119.58 ;
      RECT 0.42 119.24 19.58 119.58 ;
    LAYER M2 ;
      RECT 0.45 4.2 0.73 7.7 ;
      RECT 1.55 68.095 2.45 93.855 ;
      RECT 17.55 35.695 18.45 61.455 ;
      RECT 19.27 4.2 19.55 7.7 ;
  END
END decoupling_cap_filler

END LIBRARY
