VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO digital_ring
  CLASS BLOCK ;
  ORIGIN -13.415 -16.245 ;
  FOREIGN digital_ring 13.415 16.245 ;
  SIZE 18162.76 BY 402.9 ;
  SYMMETRY X Y R90 ;
  PIN PSUB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 18171.195 20.725 18172.195 419.145 ;
        RECT 17.395 20.725 18172.195 21.725 ;
        RECT 17.395 20.725 18.395 419.145 ;
    END
  END PSUB
  PIN VDDP
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 26.67 404.43 18162.92 405.93 ;
        RECT 18161.42 30 18162.92 405.93 ;
        RECT 26.67 30 18162.92 31.5 ;
        RECT 26.67 30 28.17 405.93 ;
    END
  END VDDP
END digital_ring

END LIBRARY
