VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  MACRO CatenaDesignType STRING ;
END PROPERTYDEFINITIONS

MACRO matrix_dac
  CLASS BLOCK ;
  ORIGIN -326.66 -187.44 ;
  FOREIGN matrix_dac 326.66 187.44 ;
  SIZE 18163.8 BY 8426.125 ;
  SYMMETRY X Y R90 ;
  PIN BcidMtx[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 493.705 187.44 493.985 188.44 ;
    END
  END BcidMtx[5]
  PIN BcidMtx[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 493.145 187.44 493.425 188.44 ;
    END
  END BcidMtx[4]
  PIN BcidMtx[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 492.585 187.44 492.865 188.44 ;
    END
  END BcidMtx[3]
  PIN BcidMtx[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 490.905 187.44 491.185 188.44 ;
    END
  END BcidMtx[2]
  PIN BcidMtx[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 490.345 187.44 490.625 188.44 ;
    END
  END BcidMtx[1]
  PIN BcidMtx[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 489.785 187.44 490.065 188.44 ;
    END
  END BcidMtx[0]
  PIN Data_PMOS[1175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9392.665 187.44 9392.945 188.44 ;
    END
  END Data_PMOS[1175]
  PIN Data_PMOS[1174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9394.345 187.44 9394.625 188.44 ;
    END
  END Data_PMOS[1174]
  PIN Data_PMOS[1173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9396.025 187.44 9396.305 188.44 ;
    END
  END Data_PMOS[1173]
  PIN Data_PMOS[1172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9362.425 187.44 9362.705 188.44 ;
    END
  END Data_PMOS[1172]
  PIN Data_PMOS[1171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9364.665 187.44 9364.945 188.44 ;
    END
  END Data_PMOS[1171]
  PIN Data_PMOS[1170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9366.345 187.44 9366.625 188.44 ;
    END
  END Data_PMOS[1170]
  PIN Data_PMOS[1169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9392.105 187.44 9392.385 188.44 ;
    END
  END Data_PMOS[1169]
  PIN Data_PMOS[1168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9393.225 187.44 9393.505 188.44 ;
    END
  END Data_PMOS[1168]
  PIN Data_PMOS[1167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9394.905 187.44 9395.185 188.44 ;
    END
  END Data_PMOS[1167]
  PIN Data_PMOS[1166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9364.105 187.44 9364.385 188.44 ;
    END
  END Data_PMOS[1166]
  PIN Data_PMOS[1165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9365.785 187.44 9366.065 188.44 ;
    END
  END Data_PMOS[1165]
  PIN Data_PMOS[1164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9366.905 187.44 9367.185 188.44 ;
    END
  END Data_PMOS[1164]
  PIN Data_PMOS[1163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9395.465 187.44 9395.745 188.44 ;
    END
  END Data_PMOS[1163]
  PIN Data_PMOS[1162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9391.545 187.44 9391.825 188.44 ;
    END
  END Data_PMOS[1162]
  PIN Data_PMOS[1161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9390.985 187.44 9391.265 188.44 ;
    END
  END Data_PMOS[1161]
  PIN Data_PMOS[1160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9393.785 187.44 9394.065 188.44 ;
    END
  END Data_PMOS[1160]
  PIN Data_PMOS[1159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9365.225 187.44 9365.505 188.44 ;
    END
  END Data_PMOS[1159]
  PIN Data_PMOS[1158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9368.025 187.44 9368.305 188.44 ;
    END
  END Data_PMOS[1158]
  PIN Data_PMOS[1157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9367.465 187.44 9367.745 188.44 ;
    END
  END Data_PMOS[1157]
  PIN Data_PMOS[1156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9363.545 187.44 9363.825 188.44 ;
    END
  END Data_PMOS[1156]
  PIN Data_PMOS[1155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9362.985 187.44 9363.265 188.44 ;
    END
  END Data_PMOS[1155]
  PIN Data_PMOS[1154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9310.905 187.44 9311.185 188.44 ;
    END
  END Data_PMOS[1154]
  PIN Data_PMOS[1153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9312.585 187.44 9312.865 188.44 ;
    END
  END Data_PMOS[1153]
  PIN Data_PMOS[1152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9314.265 187.44 9314.545 188.44 ;
    END
  END Data_PMOS[1152]
  PIN Data_PMOS[1151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9258.265 187.44 9258.545 188.44 ;
    END
  END Data_PMOS[1151]
  PIN Data_PMOS[1150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9260.505 187.44 9260.785 188.44 ;
    END
  END Data_PMOS[1150]
  PIN Data_PMOS[1149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9287.665 187.44 9287.945 188.44 ;
    END
  END Data_PMOS[1149]
  PIN Data_PMOS[1148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9310.345 187.44 9310.625 188.44 ;
    END
  END Data_PMOS[1148]
  PIN Data_PMOS[1147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9311.465 187.44 9311.745 188.44 ;
    END
  END Data_PMOS[1147]
  PIN Data_PMOS[1146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9313.145 187.44 9313.425 188.44 ;
    END
  END Data_PMOS[1146]
  PIN Data_PMOS[1145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9259.945 187.44 9260.225 188.44 ;
    END
  END Data_PMOS[1145]
  PIN Data_PMOS[1144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9287.105 187.44 9287.385 188.44 ;
    END
  END Data_PMOS[1144]
  PIN Data_PMOS[1143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9288.225 187.44 9288.505 188.44 ;
    END
  END Data_PMOS[1143]
  PIN Data_PMOS[1142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9313.705 187.44 9313.985 188.44 ;
    END
  END Data_PMOS[1142]
  PIN Data_PMOS[1141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9309.785 187.44 9310.065 188.44 ;
    END
  END Data_PMOS[1141]
  PIN Data_PMOS[1140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9300.825 187.44 9301.105 188.44 ;
    END
  END Data_PMOS[1140]
  PIN Data_PMOS[1139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9312.025 187.44 9312.305 188.44 ;
    END
  END Data_PMOS[1139]
  PIN Data_PMOS[1138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9261.065 187.44 9261.345 188.44 ;
    END
  END Data_PMOS[1138]
  PIN Data_PMOS[1137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9289.345 187.44 9289.625 188.44 ;
    END
  END Data_PMOS[1137]
  PIN Data_PMOS[1136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9288.785 187.44 9289.065 188.44 ;
    END
  END Data_PMOS[1136]
  PIN Data_PMOS[1135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9259.385 187.44 9259.665 188.44 ;
    END
  END Data_PMOS[1135]
  PIN Data_PMOS[1134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9258.825 187.44 9259.105 188.44 ;
    END
  END Data_PMOS[1134]
  PIN Data_PMOS[1133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9232.505 187.44 9232.785 188.44 ;
    END
  END Data_PMOS[1133]
  PIN Data_PMOS[1132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9234.185 187.44 9234.465 188.44 ;
    END
  END Data_PMOS[1132]
  PIN Data_PMOS[1131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9248.745 187.44 9249.025 188.44 ;
    END
  END Data_PMOS[1131]
  PIN Data_PMOS[1130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9177.065 187.44 9177.345 188.44 ;
    END
  END Data_PMOS[1130]
  PIN Data_PMOS[1129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9179.305 187.44 9179.585 188.44 ;
    END
  END Data_PMOS[1129]
  PIN Data_PMOS[1128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9180.985 187.44 9181.265 188.44 ;
    END
  END Data_PMOS[1128]
  PIN Data_PMOS[1127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9231.945 187.44 9232.225 188.44 ;
    END
  END Data_PMOS[1127]
  PIN Data_PMOS[1126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9233.065 187.44 9233.345 188.44 ;
    END
  END Data_PMOS[1126]
  PIN Data_PMOS[1125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9234.745 187.44 9235.025 188.44 ;
    END
  END Data_PMOS[1125]
  PIN Data_PMOS[1124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9178.745 187.44 9179.025 188.44 ;
    END
  END Data_PMOS[1124]
  PIN Data_PMOS[1123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9180.425 187.44 9180.705 188.44 ;
    END
  END Data_PMOS[1123]
  PIN Data_PMOS[1122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9181.545 187.44 9181.825 188.44 ;
    END
  END Data_PMOS[1122]
  PIN Data_PMOS[1121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9248.185 187.44 9248.465 188.44 ;
    END
  END Data_PMOS[1121]
  PIN Data_PMOS[1120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9231.385 187.44 9231.665 188.44 ;
    END
  END Data_PMOS[1120]
  PIN Data_PMOS[1119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9230.825 187.44 9231.105 188.44 ;
    END
  END Data_PMOS[1119]
  PIN Data_PMOS[1118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9233.625 187.44 9233.905 188.44 ;
    END
  END Data_PMOS[1118]
  PIN Data_PMOS[1117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9179.865 187.44 9180.145 188.44 ;
    END
  END Data_PMOS[1117]
  PIN Data_PMOS[1116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9182.665 187.44 9182.945 188.44 ;
    END
  END Data_PMOS[1116]
  PIN Data_PMOS[1115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9182.105 187.44 9182.385 188.44 ;
    END
  END Data_PMOS[1115]
  PIN Data_PMOS[1114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9178.185 187.44 9178.465 188.44 ;
    END
  END Data_PMOS[1114]
  PIN Data_PMOS[1113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9177.625 187.44 9177.905 188.44 ;
    END
  END Data_PMOS[1113]
  PIN Data_PMOS[1112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9155.785 187.44 9156.065 188.44 ;
    END
  END Data_PMOS[1112]
  PIN Data_PMOS[1111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9157.465 187.44 9157.745 188.44 ;
    END
  END Data_PMOS[1111]
  PIN Data_PMOS[1110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9159.145 187.44 9159.425 188.44 ;
    END
  END Data_PMOS[1110]
  PIN Data_PMOS[1109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9111.545 187.44 9111.825 188.44 ;
    END
  END Data_PMOS[1109]
  PIN Data_PMOS[1108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9113.785 187.44 9114.065 188.44 ;
    END
  END Data_PMOS[1108]
  PIN Data_PMOS[1107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9115.465 187.44 9115.745 188.44 ;
    END
  END Data_PMOS[1107]
  PIN Data_PMOS[1106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9155.225 187.44 9155.505 188.44 ;
    END
  END Data_PMOS[1106]
  PIN Data_PMOS[1105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9156.345 187.44 9156.625 188.44 ;
    END
  END Data_PMOS[1105]
  PIN Data_PMOS[1104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9158.025 187.44 9158.305 188.44 ;
    END
  END Data_PMOS[1104]
  PIN Data_PMOS[1103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9113.225 187.44 9113.505 188.44 ;
    END
  END Data_PMOS[1103]
  PIN Data_PMOS[1102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9114.905 187.44 9115.185 188.44 ;
    END
  END Data_PMOS[1102]
  PIN Data_PMOS[1101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9116.025 187.44 9116.305 188.44 ;
    END
  END Data_PMOS[1101]
  PIN Data_PMOS[1100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9158.585 187.44 9158.865 188.44 ;
    END
  END Data_PMOS[1100]
  PIN Data_PMOS[1099]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9154.665 187.44 9154.945 188.44 ;
    END
  END Data_PMOS[1099]
  PIN Data_PMOS[1098]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9154.105 187.44 9154.385 188.44 ;
    END
  END Data_PMOS[1098]
  PIN Data_PMOS[1097]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9156.905 187.44 9157.185 188.44 ;
    END
  END Data_PMOS[1097]
  PIN Data_PMOS[1096]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9114.345 187.44 9114.625 188.44 ;
    END
  END Data_PMOS[1096]
  PIN Data_PMOS[1095]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9117.145 187.44 9117.425 188.44 ;
    END
  END Data_PMOS[1095]
  PIN Data_PMOS[1094]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9116.585 187.44 9116.865 188.44 ;
    END
  END Data_PMOS[1094]
  PIN Data_PMOS[1093]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9112.665 187.44 9112.945 188.44 ;
    END
  END Data_PMOS[1093]
  PIN Data_PMOS[1092]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9112.105 187.44 9112.385 188.44 ;
    END
  END Data_PMOS[1092]
  PIN Data_PMOS[1091]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9085.785 187.44 9086.065 188.44 ;
    END
  END Data_PMOS[1091]
  PIN Data_PMOS[1090]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9087.465 187.44 9087.745 188.44 ;
    END
  END Data_PMOS[1090]
  PIN Data_PMOS[1089]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9089.145 187.44 9089.425 188.44 ;
    END
  END Data_PMOS[1089]
  PIN Data_PMOS[1088]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9029.785 187.44 9030.065 188.44 ;
    END
  END Data_PMOS[1088]
  PIN Data_PMOS[1087]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9032.025 187.44 9032.305 188.44 ;
    END
  END Data_PMOS[1087]
  PIN Data_PMOS[1086]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9033.705 187.44 9033.985 188.44 ;
    END
  END Data_PMOS[1086]
  PIN Data_PMOS[1085]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9085.225 187.44 9085.505 188.44 ;
    END
  END Data_PMOS[1085]
  PIN Data_PMOS[1084]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9086.345 187.44 9086.625 188.44 ;
    END
  END Data_PMOS[1084]
  PIN Data_PMOS[1083]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9088.025 187.44 9088.305 188.44 ;
    END
  END Data_PMOS[1083]
  PIN Data_PMOS[1082]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9031.465 187.44 9031.745 188.44 ;
    END
  END Data_PMOS[1082]
  PIN Data_PMOS[1081]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9033.145 187.44 9033.425 188.44 ;
    END
  END Data_PMOS[1081]
  PIN Data_PMOS[1080]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9034.265 187.44 9034.545 188.44 ;
    END
  END Data_PMOS[1080]
  PIN Data_PMOS[1079]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9088.585 187.44 9088.865 188.44 ;
    END
  END Data_PMOS[1079]
  PIN Data_PMOS[1078]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9084.665 187.44 9084.945 188.44 ;
    END
  END Data_PMOS[1078]
  PIN Data_PMOS[1077]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9084.105 187.44 9084.385 188.44 ;
    END
  END Data_PMOS[1077]
  PIN Data_PMOS[1076]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9086.905 187.44 9087.185 188.44 ;
    END
  END Data_PMOS[1076]
  PIN Data_PMOS[1075]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9032.585 187.44 9032.865 188.44 ;
    END
  END Data_PMOS[1075]
  PIN Data_PMOS[1074]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9035.385 187.44 9035.665 188.44 ;
    END
  END Data_PMOS[1074]
  PIN Data_PMOS[1073]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9034.825 187.44 9035.105 188.44 ;
    END
  END Data_PMOS[1073]
  PIN Data_PMOS[1072]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9030.905 187.44 9031.185 188.44 ;
    END
  END Data_PMOS[1072]
  PIN Data_PMOS[1071]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9030.345 187.44 9030.625 188.44 ;
    END
  END Data_PMOS[1071]
  PIN Data_PMOS[1070]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8981.065 187.44 8981.345 188.44 ;
    END
  END Data_PMOS[1070]
  PIN Data_PMOS[1069]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9008.225 187.44 9008.505 188.44 ;
    END
  END Data_PMOS[1069]
  PIN Data_PMOS[1068]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9009.905 187.44 9010.185 188.44 ;
    END
  END Data_PMOS[1068]
  PIN Data_PMOS[1067]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8951.385 187.44 8951.665 188.44 ;
    END
  END Data_PMOS[1067]
  PIN Data_PMOS[1066]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8953.625 187.44 8953.905 188.44 ;
    END
  END Data_PMOS[1066]
  PIN Data_PMOS[1065]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8955.305 187.44 8955.585 188.44 ;
    END
  END Data_PMOS[1065]
  PIN Data_PMOS[1064]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8980.505 187.44 8980.785 188.44 ;
    END
  END Data_PMOS[1064]
  PIN Data_PMOS[1063]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8981.625 187.44 8981.905 188.44 ;
    END
  END Data_PMOS[1063]
  PIN Data_PMOS[1062]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9008.785 187.44 9009.065 188.44 ;
    END
  END Data_PMOS[1062]
  PIN Data_PMOS[1061]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8953.065 187.44 8953.345 188.44 ;
    END
  END Data_PMOS[1061]
  PIN Data_PMOS[1060]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8954.745 187.44 8955.025 188.44 ;
    END
  END Data_PMOS[1060]
  PIN Data_PMOS[1059]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8968.745 187.44 8969.025 188.44 ;
    END
  END Data_PMOS[1059]
  PIN Data_PMOS[1058]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9009.345 187.44 9009.625 188.44 ;
    END
  END Data_PMOS[1058]
  PIN Data_PMOS[1057]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8979.945 187.44 8980.225 188.44 ;
    END
  END Data_PMOS[1057]
  PIN Data_PMOS[1056]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8979.385 187.44 8979.665 188.44 ;
    END
  END Data_PMOS[1056]
  PIN Data_PMOS[1055]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9007.665 187.44 9007.945 188.44 ;
    END
  END Data_PMOS[1055]
  PIN Data_PMOS[1054]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8954.185 187.44 8954.465 188.44 ;
    END
  END Data_PMOS[1054]
  PIN Data_PMOS[1053]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8969.865 187.44 8970.145 188.44 ;
    END
  END Data_PMOS[1053]
  PIN Data_PMOS[1052]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8969.305 187.44 8969.585 188.44 ;
    END
  END Data_PMOS[1052]
  PIN Data_PMOS[1051]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8952.505 187.44 8952.785 188.44 ;
    END
  END Data_PMOS[1051]
  PIN Data_PMOS[1050]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8951.945 187.44 8952.225 188.44 ;
    END
  END Data_PMOS[1050]
  PIN Data_PMOS[1049]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8898.745 187.44 8899.025 188.44 ;
    END
  END Data_PMOS[1049]
  PIN Data_PMOS[1048]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8900.425 187.44 8900.705 188.44 ;
    END
  END Data_PMOS[1048]
  PIN Data_PMOS[1047]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8902.105 187.44 8902.385 188.44 ;
    END
  END Data_PMOS[1047]
  PIN Data_PMOS[1046]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8873.545 187.44 8873.825 188.44 ;
    END
  END Data_PMOS[1046]
  PIN Data_PMOS[1045]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8875.785 187.44 8876.065 188.44 ;
    END
  END Data_PMOS[1045]
  PIN Data_PMOS[1044]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8877.465 187.44 8877.745 188.44 ;
    END
  END Data_PMOS[1044]
  PIN Data_PMOS[1043]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8898.185 187.44 8898.465 188.44 ;
    END
  END Data_PMOS[1043]
  PIN Data_PMOS[1042]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8899.305 187.44 8899.585 188.44 ;
    END
  END Data_PMOS[1042]
  PIN Data_PMOS[1041]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8900.985 187.44 8901.265 188.44 ;
    END
  END Data_PMOS[1041]
  PIN Data_PMOS[1040]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8875.225 187.44 8875.505 188.44 ;
    END
  END Data_PMOS[1040]
  PIN Data_PMOS[1039]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8876.905 187.44 8877.185 188.44 ;
    END
  END Data_PMOS[1039]
  PIN Data_PMOS[1038]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8878.025 187.44 8878.305 188.44 ;
    END
  END Data_PMOS[1038]
  PIN Data_PMOS[1037]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8901.545 187.44 8901.825 188.44 ;
    END
  END Data_PMOS[1037]
  PIN Data_PMOS[1036]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8897.625 187.44 8897.905 188.44 ;
    END
  END Data_PMOS[1036]
  PIN Data_PMOS[1035]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8897.065 187.44 8897.345 188.44 ;
    END
  END Data_PMOS[1035]
  PIN Data_PMOS[1034]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8899.865 187.44 8900.145 188.44 ;
    END
  END Data_PMOS[1034]
  PIN Data_PMOS[1033]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8876.345 187.44 8876.625 188.44 ;
    END
  END Data_PMOS[1033]
  PIN Data_PMOS[1032]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8879.145 187.44 8879.425 188.44 ;
    END
  END Data_PMOS[1032]
  PIN Data_PMOS[1031]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8878.585 187.44 8878.865 188.44 ;
    END
  END Data_PMOS[1031]
  PIN Data_PMOS[1030]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8874.665 187.44 8874.945 188.44 ;
    END
  END Data_PMOS[1030]
  PIN Data_PMOS[1029]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8874.105 187.44 8874.385 188.44 ;
    END
  END Data_PMOS[1029]
  PIN Data_PMOS[1028]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8832.665 187.44 8832.945 188.44 ;
    END
  END Data_PMOS[1028]
  PIN Data_PMOS[1027]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8834.345 187.44 8834.625 188.44 ;
    END
  END Data_PMOS[1027]
  PIN Data_PMOS[1026]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8836.025 187.44 8836.305 188.44 ;
    END
  END Data_PMOS[1026]
  PIN Data_PMOS[1025]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8802.425 187.44 8802.705 188.44 ;
    END
  END Data_PMOS[1025]
  PIN Data_PMOS[1024]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8804.665 187.44 8804.945 188.44 ;
    END
  END Data_PMOS[1024]
  PIN Data_PMOS[1023]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8806.345 187.44 8806.625 188.44 ;
    END
  END Data_PMOS[1023]
  PIN Data_PMOS[1022]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8832.105 187.44 8832.385 188.44 ;
    END
  END Data_PMOS[1022]
  PIN Data_PMOS[1021]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8833.225 187.44 8833.505 188.44 ;
    END
  END Data_PMOS[1021]
  PIN Data_PMOS[1020]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8834.905 187.44 8835.185 188.44 ;
    END
  END Data_PMOS[1020]
  PIN Data_PMOS[1019]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8804.105 187.44 8804.385 188.44 ;
    END
  END Data_PMOS[1019]
  PIN Data_PMOS[1018]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8805.785 187.44 8806.065 188.44 ;
    END
  END Data_PMOS[1018]
  PIN Data_PMOS[1017]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8806.905 187.44 8807.185 188.44 ;
    END
  END Data_PMOS[1017]
  PIN Data_PMOS[1016]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8835.465 187.44 8835.745 188.44 ;
    END
  END Data_PMOS[1016]
  PIN Data_PMOS[1015]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8831.545 187.44 8831.825 188.44 ;
    END
  END Data_PMOS[1015]
  PIN Data_PMOS[1014]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8830.985 187.44 8831.265 188.44 ;
    END
  END Data_PMOS[1014]
  PIN Data_PMOS[1013]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8833.785 187.44 8834.065 188.44 ;
    END
  END Data_PMOS[1013]
  PIN Data_PMOS[1012]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8805.225 187.44 8805.505 188.44 ;
    END
  END Data_PMOS[1012]
  PIN Data_PMOS[1011]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8808.025 187.44 8808.305 188.44 ;
    END
  END Data_PMOS[1011]
  PIN Data_PMOS[1010]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8807.465 187.44 8807.745 188.44 ;
    END
  END Data_PMOS[1010]
  PIN Data_PMOS[1009]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8803.545 187.44 8803.825 188.44 ;
    END
  END Data_PMOS[1009]
  PIN Data_PMOS[1008]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8802.985 187.44 8803.265 188.44 ;
    END
  END Data_PMOS[1008]
  PIN Data_PMOS[1007]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8750.905 187.44 8751.185 188.44 ;
    END
  END Data_PMOS[1007]
  PIN Data_PMOS[1006]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8752.585 187.44 8752.865 188.44 ;
    END
  END Data_PMOS[1006]
  PIN Data_PMOS[1005]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8754.265 187.44 8754.545 188.44 ;
    END
  END Data_PMOS[1005]
  PIN Data_PMOS[1004]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8698.265 187.44 8698.545 188.44 ;
    END
  END Data_PMOS[1004]
  PIN Data_PMOS[1003]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8700.505 187.44 8700.785 188.44 ;
    END
  END Data_PMOS[1003]
  PIN Data_PMOS[1002]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8727.665 187.44 8727.945 188.44 ;
    END
  END Data_PMOS[1002]
  PIN Data_PMOS[1001]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8750.345 187.44 8750.625 188.44 ;
    END
  END Data_PMOS[1001]
  PIN Data_PMOS[1000]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8751.465 187.44 8751.745 188.44 ;
    END
  END Data_PMOS[1000]
  PIN Data_PMOS[999]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8753.145 187.44 8753.425 188.44 ;
    END
  END Data_PMOS[999]
  PIN Data_PMOS[998]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8699.945 187.44 8700.225 188.44 ;
    END
  END Data_PMOS[998]
  PIN Data_PMOS[997]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8727.105 187.44 8727.385 188.44 ;
    END
  END Data_PMOS[997]
  PIN Data_PMOS[996]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8728.225 187.44 8728.505 188.44 ;
    END
  END Data_PMOS[996]
  PIN Data_PMOS[995]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8753.705 187.44 8753.985 188.44 ;
    END
  END Data_PMOS[995]
  PIN Data_PMOS[994]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8749.785 187.44 8750.065 188.44 ;
    END
  END Data_PMOS[994]
  PIN Data_PMOS[993]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8740.825 187.44 8741.105 188.44 ;
    END
  END Data_PMOS[993]
  PIN Data_PMOS[992]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8752.025 187.44 8752.305 188.44 ;
    END
  END Data_PMOS[992]
  PIN Data_PMOS[991]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8701.065 187.44 8701.345 188.44 ;
    END
  END Data_PMOS[991]
  PIN Data_PMOS[990]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8729.345 187.44 8729.625 188.44 ;
    END
  END Data_PMOS[990]
  PIN Data_PMOS[989]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8728.785 187.44 8729.065 188.44 ;
    END
  END Data_PMOS[989]
  PIN Data_PMOS[988]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8699.385 187.44 8699.665 188.44 ;
    END
  END Data_PMOS[988]
  PIN Data_PMOS[987]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8698.825 187.44 8699.105 188.44 ;
    END
  END Data_PMOS[987]
  PIN Data_PMOS[986]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8672.505 187.44 8672.785 188.44 ;
    END
  END Data_PMOS[986]
  PIN Data_PMOS[985]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8674.185 187.44 8674.465 188.44 ;
    END
  END Data_PMOS[985]
  PIN Data_PMOS[984]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8688.745 187.44 8689.025 188.44 ;
    END
  END Data_PMOS[984]
  PIN Data_PMOS[983]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8617.065 187.44 8617.345 188.44 ;
    END
  END Data_PMOS[983]
  PIN Data_PMOS[982]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8619.305 187.44 8619.585 188.44 ;
    END
  END Data_PMOS[982]
  PIN Data_PMOS[981]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8620.985 187.44 8621.265 188.44 ;
    END
  END Data_PMOS[981]
  PIN Data_PMOS[980]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8671.945 187.44 8672.225 188.44 ;
    END
  END Data_PMOS[980]
  PIN Data_PMOS[979]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8673.065 187.44 8673.345 188.44 ;
    END
  END Data_PMOS[979]
  PIN Data_PMOS[978]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8674.745 187.44 8675.025 188.44 ;
    END
  END Data_PMOS[978]
  PIN Data_PMOS[977]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8618.745 187.44 8619.025 188.44 ;
    END
  END Data_PMOS[977]
  PIN Data_PMOS[976]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8620.425 187.44 8620.705 188.44 ;
    END
  END Data_PMOS[976]
  PIN Data_PMOS[975]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8621.545 187.44 8621.825 188.44 ;
    END
  END Data_PMOS[975]
  PIN Data_PMOS[974]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8688.185 187.44 8688.465 188.44 ;
    END
  END Data_PMOS[974]
  PIN Data_PMOS[973]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8671.385 187.44 8671.665 188.44 ;
    END
  END Data_PMOS[973]
  PIN Data_PMOS[972]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8670.825 187.44 8671.105 188.44 ;
    END
  END Data_PMOS[972]
  PIN Data_PMOS[971]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8673.625 187.44 8673.905 188.44 ;
    END
  END Data_PMOS[971]
  PIN Data_PMOS[970]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8619.865 187.44 8620.145 188.44 ;
    END
  END Data_PMOS[970]
  PIN Data_PMOS[969]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8622.665 187.44 8622.945 188.44 ;
    END
  END Data_PMOS[969]
  PIN Data_PMOS[968]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8622.105 187.44 8622.385 188.44 ;
    END
  END Data_PMOS[968]
  PIN Data_PMOS[967]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8618.185 187.44 8618.465 188.44 ;
    END
  END Data_PMOS[967]
  PIN Data_PMOS[966]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8617.625 187.44 8617.905 188.44 ;
    END
  END Data_PMOS[966]
  PIN Data_PMOS[965]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8595.785 187.44 8596.065 188.44 ;
    END
  END Data_PMOS[965]
  PIN Data_PMOS[964]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8597.465 187.44 8597.745 188.44 ;
    END
  END Data_PMOS[964]
  PIN Data_PMOS[963]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8599.145 187.44 8599.425 188.44 ;
    END
  END Data_PMOS[963]
  PIN Data_PMOS[962]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8551.545 187.44 8551.825 188.44 ;
    END
  END Data_PMOS[962]
  PIN Data_PMOS[961]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8553.785 187.44 8554.065 188.44 ;
    END
  END Data_PMOS[961]
  PIN Data_PMOS[960]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8555.465 187.44 8555.745 188.44 ;
    END
  END Data_PMOS[960]
  PIN Data_PMOS[959]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8595.225 187.44 8595.505 188.44 ;
    END
  END Data_PMOS[959]
  PIN Data_PMOS[958]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8596.345 187.44 8596.625 188.44 ;
    END
  END Data_PMOS[958]
  PIN Data_PMOS[957]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8598.025 187.44 8598.305 188.44 ;
    END
  END Data_PMOS[957]
  PIN Data_PMOS[956]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8553.225 187.44 8553.505 188.44 ;
    END
  END Data_PMOS[956]
  PIN Data_PMOS[955]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8554.905 187.44 8555.185 188.44 ;
    END
  END Data_PMOS[955]
  PIN Data_PMOS[954]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8556.025 187.44 8556.305 188.44 ;
    END
  END Data_PMOS[954]
  PIN Data_PMOS[953]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8598.585 187.44 8598.865 188.44 ;
    END
  END Data_PMOS[953]
  PIN Data_PMOS[952]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8594.665 187.44 8594.945 188.44 ;
    END
  END Data_PMOS[952]
  PIN Data_PMOS[951]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8594.105 187.44 8594.385 188.44 ;
    END
  END Data_PMOS[951]
  PIN Data_PMOS[950]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8596.905 187.44 8597.185 188.44 ;
    END
  END Data_PMOS[950]
  PIN Data_PMOS[949]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8554.345 187.44 8554.625 188.44 ;
    END
  END Data_PMOS[949]
  PIN Data_PMOS[948]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8557.145 187.44 8557.425 188.44 ;
    END
  END Data_PMOS[948]
  PIN Data_PMOS[947]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8556.585 187.44 8556.865 188.44 ;
    END
  END Data_PMOS[947]
  PIN Data_PMOS[946]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8552.665 187.44 8552.945 188.44 ;
    END
  END Data_PMOS[946]
  PIN Data_PMOS[945]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8552.105 187.44 8552.385 188.44 ;
    END
  END Data_PMOS[945]
  PIN Data_PMOS[944]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8525.785 187.44 8526.065 188.44 ;
    END
  END Data_PMOS[944]
  PIN Data_PMOS[943]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8527.465 187.44 8527.745 188.44 ;
    END
  END Data_PMOS[943]
  PIN Data_PMOS[942]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8529.145 187.44 8529.425 188.44 ;
    END
  END Data_PMOS[942]
  PIN Data_PMOS[941]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8469.785 187.44 8470.065 188.44 ;
    END
  END Data_PMOS[941]
  PIN Data_PMOS[940]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8472.025 187.44 8472.305 188.44 ;
    END
  END Data_PMOS[940]
  PIN Data_PMOS[939]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8473.705 187.44 8473.985 188.44 ;
    END
  END Data_PMOS[939]
  PIN Data_PMOS[938]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8525.225 187.44 8525.505 188.44 ;
    END
  END Data_PMOS[938]
  PIN Data_PMOS[937]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8526.345 187.44 8526.625 188.44 ;
    END
  END Data_PMOS[937]
  PIN Data_PMOS[936]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8528.025 187.44 8528.305 188.44 ;
    END
  END Data_PMOS[936]
  PIN Data_PMOS[935]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8471.465 187.44 8471.745 188.44 ;
    END
  END Data_PMOS[935]
  PIN Data_PMOS[934]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8473.145 187.44 8473.425 188.44 ;
    END
  END Data_PMOS[934]
  PIN Data_PMOS[933]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8474.265 187.44 8474.545 188.44 ;
    END
  END Data_PMOS[933]
  PIN Data_PMOS[932]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8528.585 187.44 8528.865 188.44 ;
    END
  END Data_PMOS[932]
  PIN Data_PMOS[931]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8524.665 187.44 8524.945 188.44 ;
    END
  END Data_PMOS[931]
  PIN Data_PMOS[930]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8524.105 187.44 8524.385 188.44 ;
    END
  END Data_PMOS[930]
  PIN Data_PMOS[929]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8526.905 187.44 8527.185 188.44 ;
    END
  END Data_PMOS[929]
  PIN Data_PMOS[928]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8472.585 187.44 8472.865 188.44 ;
    END
  END Data_PMOS[928]
  PIN Data_PMOS[927]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8475.385 187.44 8475.665 188.44 ;
    END
  END Data_PMOS[927]
  PIN Data_PMOS[926]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8474.825 187.44 8475.105 188.44 ;
    END
  END Data_PMOS[926]
  PIN Data_PMOS[925]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8470.905 187.44 8471.185 188.44 ;
    END
  END Data_PMOS[925]
  PIN Data_PMOS[924]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8470.345 187.44 8470.625 188.44 ;
    END
  END Data_PMOS[924]
  PIN Data_PMOS[923]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8421.065 187.44 8421.345 188.44 ;
    END
  END Data_PMOS[923]
  PIN Data_PMOS[922]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8448.225 187.44 8448.505 188.44 ;
    END
  END Data_PMOS[922]
  PIN Data_PMOS[921]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8449.905 187.44 8450.185 188.44 ;
    END
  END Data_PMOS[921]
  PIN Data_PMOS[920]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8391.385 187.44 8391.665 188.44 ;
    END
  END Data_PMOS[920]
  PIN Data_PMOS[919]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8393.625 187.44 8393.905 188.44 ;
    END
  END Data_PMOS[919]
  PIN Data_PMOS[918]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8395.305 187.44 8395.585 188.44 ;
    END
  END Data_PMOS[918]
  PIN Data_PMOS[917]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8420.505 187.44 8420.785 188.44 ;
    END
  END Data_PMOS[917]
  PIN Data_PMOS[916]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8421.625 187.44 8421.905 188.44 ;
    END
  END Data_PMOS[916]
  PIN Data_PMOS[915]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8448.785 187.44 8449.065 188.44 ;
    END
  END Data_PMOS[915]
  PIN Data_PMOS[914]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8393.065 187.44 8393.345 188.44 ;
    END
  END Data_PMOS[914]
  PIN Data_PMOS[913]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8394.745 187.44 8395.025 188.44 ;
    END
  END Data_PMOS[913]
  PIN Data_PMOS[912]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8408.745 187.44 8409.025 188.44 ;
    END
  END Data_PMOS[912]
  PIN Data_PMOS[911]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8449.345 187.44 8449.625 188.44 ;
    END
  END Data_PMOS[911]
  PIN Data_PMOS[910]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8419.945 187.44 8420.225 188.44 ;
    END
  END Data_PMOS[910]
  PIN Data_PMOS[909]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8419.385 187.44 8419.665 188.44 ;
    END
  END Data_PMOS[909]
  PIN Data_PMOS[908]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8447.665 187.44 8447.945 188.44 ;
    END
  END Data_PMOS[908]
  PIN Data_PMOS[907]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8394.185 187.44 8394.465 188.44 ;
    END
  END Data_PMOS[907]
  PIN Data_PMOS[906]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8409.865 187.44 8410.145 188.44 ;
    END
  END Data_PMOS[906]
  PIN Data_PMOS[905]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8409.305 187.44 8409.585 188.44 ;
    END
  END Data_PMOS[905]
  PIN Data_PMOS[904]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8392.505 187.44 8392.785 188.44 ;
    END
  END Data_PMOS[904]
  PIN Data_PMOS[903]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8391.945 187.44 8392.225 188.44 ;
    END
  END Data_PMOS[903]
  PIN Data_PMOS[902]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8338.745 187.44 8339.025 188.44 ;
    END
  END Data_PMOS[902]
  PIN Data_PMOS[901]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8340.425 187.44 8340.705 188.44 ;
    END
  END Data_PMOS[901]
  PIN Data_PMOS[900]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8342.105 187.44 8342.385 188.44 ;
    END
  END Data_PMOS[900]
  PIN Data_PMOS[899]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8313.545 187.44 8313.825 188.44 ;
    END
  END Data_PMOS[899]
  PIN Data_PMOS[898]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8315.785 187.44 8316.065 188.44 ;
    END
  END Data_PMOS[898]
  PIN Data_PMOS[897]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8317.465 187.44 8317.745 188.44 ;
    END
  END Data_PMOS[897]
  PIN Data_PMOS[896]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8338.185 187.44 8338.465 188.44 ;
    END
  END Data_PMOS[896]
  PIN Data_PMOS[895]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8339.305 187.44 8339.585 188.44 ;
    END
  END Data_PMOS[895]
  PIN Data_PMOS[894]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8340.985 187.44 8341.265 188.44 ;
    END
  END Data_PMOS[894]
  PIN Data_PMOS[893]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8315.225 187.44 8315.505 188.44 ;
    END
  END Data_PMOS[893]
  PIN Data_PMOS[892]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8316.905 187.44 8317.185 188.44 ;
    END
  END Data_PMOS[892]
  PIN Data_PMOS[891]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8318.025 187.44 8318.305 188.44 ;
    END
  END Data_PMOS[891]
  PIN Data_PMOS[890]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8341.545 187.44 8341.825 188.44 ;
    END
  END Data_PMOS[890]
  PIN Data_PMOS[889]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8337.625 187.44 8337.905 188.44 ;
    END
  END Data_PMOS[889]
  PIN Data_PMOS[888]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8337.065 187.44 8337.345 188.44 ;
    END
  END Data_PMOS[888]
  PIN Data_PMOS[887]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8339.865 187.44 8340.145 188.44 ;
    END
  END Data_PMOS[887]
  PIN Data_PMOS[886]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8316.345 187.44 8316.625 188.44 ;
    END
  END Data_PMOS[886]
  PIN Data_PMOS[885]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8319.145 187.44 8319.425 188.44 ;
    END
  END Data_PMOS[885]
  PIN Data_PMOS[884]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8318.585 187.44 8318.865 188.44 ;
    END
  END Data_PMOS[884]
  PIN Data_PMOS[883]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8314.665 187.44 8314.945 188.44 ;
    END
  END Data_PMOS[883]
  PIN Data_PMOS[882]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8314.105 187.44 8314.385 188.44 ;
    END
  END Data_PMOS[882]
  PIN Data_PMOS[881]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8272.665 187.44 8272.945 188.44 ;
    END
  END Data_PMOS[881]
  PIN Data_PMOS[880]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8274.345 187.44 8274.625 188.44 ;
    END
  END Data_PMOS[880]
  PIN Data_PMOS[879]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8276.025 187.44 8276.305 188.44 ;
    END
  END Data_PMOS[879]
  PIN Data_PMOS[878]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8242.425 187.44 8242.705 188.44 ;
    END
  END Data_PMOS[878]
  PIN Data_PMOS[877]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8244.665 187.44 8244.945 188.44 ;
    END
  END Data_PMOS[877]
  PIN Data_PMOS[876]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8246.345 187.44 8246.625 188.44 ;
    END
  END Data_PMOS[876]
  PIN Data_PMOS[875]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8272.105 187.44 8272.385 188.44 ;
    END
  END Data_PMOS[875]
  PIN Data_PMOS[874]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8273.225 187.44 8273.505 188.44 ;
    END
  END Data_PMOS[874]
  PIN Data_PMOS[873]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8274.905 187.44 8275.185 188.44 ;
    END
  END Data_PMOS[873]
  PIN Data_PMOS[872]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8244.105 187.44 8244.385 188.44 ;
    END
  END Data_PMOS[872]
  PIN Data_PMOS[871]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8245.785 187.44 8246.065 188.44 ;
    END
  END Data_PMOS[871]
  PIN Data_PMOS[870]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8246.905 187.44 8247.185 188.44 ;
    END
  END Data_PMOS[870]
  PIN Data_PMOS[869]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8275.465 187.44 8275.745 188.44 ;
    END
  END Data_PMOS[869]
  PIN Data_PMOS[868]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8271.545 187.44 8271.825 188.44 ;
    END
  END Data_PMOS[868]
  PIN Data_PMOS[867]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8270.985 187.44 8271.265 188.44 ;
    END
  END Data_PMOS[867]
  PIN Data_PMOS[866]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8273.785 187.44 8274.065 188.44 ;
    END
  END Data_PMOS[866]
  PIN Data_PMOS[865]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8245.225 187.44 8245.505 188.44 ;
    END
  END Data_PMOS[865]
  PIN Data_PMOS[864]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8248.025 187.44 8248.305 188.44 ;
    END
  END Data_PMOS[864]
  PIN Data_PMOS[863]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8247.465 187.44 8247.745 188.44 ;
    END
  END Data_PMOS[863]
  PIN Data_PMOS[862]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8243.545 187.44 8243.825 188.44 ;
    END
  END Data_PMOS[862]
  PIN Data_PMOS[861]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8242.985 187.44 8243.265 188.44 ;
    END
  END Data_PMOS[861]
  PIN Data_PMOS[860]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8190.905 187.44 8191.185 188.44 ;
    END
  END Data_PMOS[860]
  PIN Data_PMOS[859]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8192.585 187.44 8192.865 188.44 ;
    END
  END Data_PMOS[859]
  PIN Data_PMOS[858]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8194.265 187.44 8194.545 188.44 ;
    END
  END Data_PMOS[858]
  PIN Data_PMOS[857]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8138.265 187.44 8138.545 188.44 ;
    END
  END Data_PMOS[857]
  PIN Data_PMOS[856]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8140.505 187.44 8140.785 188.44 ;
    END
  END Data_PMOS[856]
  PIN Data_PMOS[855]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8167.665 187.44 8167.945 188.44 ;
    END
  END Data_PMOS[855]
  PIN Data_PMOS[854]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8190.345 187.44 8190.625 188.44 ;
    END
  END Data_PMOS[854]
  PIN Data_PMOS[853]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8191.465 187.44 8191.745 188.44 ;
    END
  END Data_PMOS[853]
  PIN Data_PMOS[852]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8193.145 187.44 8193.425 188.44 ;
    END
  END Data_PMOS[852]
  PIN Data_PMOS[851]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8139.945 187.44 8140.225 188.44 ;
    END
  END Data_PMOS[851]
  PIN Data_PMOS[850]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8167.105 187.44 8167.385 188.44 ;
    END
  END Data_PMOS[850]
  PIN Data_PMOS[849]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8168.225 187.44 8168.505 188.44 ;
    END
  END Data_PMOS[849]
  PIN Data_PMOS[848]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8193.705 187.44 8193.985 188.44 ;
    END
  END Data_PMOS[848]
  PIN Data_PMOS[847]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8189.785 187.44 8190.065 188.44 ;
    END
  END Data_PMOS[847]
  PIN Data_PMOS[846]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8180.825 187.44 8181.105 188.44 ;
    END
  END Data_PMOS[846]
  PIN Data_PMOS[845]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8192.025 187.44 8192.305 188.44 ;
    END
  END Data_PMOS[845]
  PIN Data_PMOS[844]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8141.065 187.44 8141.345 188.44 ;
    END
  END Data_PMOS[844]
  PIN Data_PMOS[843]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8169.345 187.44 8169.625 188.44 ;
    END
  END Data_PMOS[843]
  PIN Data_PMOS[842]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8168.785 187.44 8169.065 188.44 ;
    END
  END Data_PMOS[842]
  PIN Data_PMOS[841]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8139.385 187.44 8139.665 188.44 ;
    END
  END Data_PMOS[841]
  PIN Data_PMOS[840]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8138.825 187.44 8139.105 188.44 ;
    END
  END Data_PMOS[840]
  PIN Data_PMOS[839]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8112.505 187.44 8112.785 188.44 ;
    END
  END Data_PMOS[839]
  PIN Data_PMOS[838]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8114.185 187.44 8114.465 188.44 ;
    END
  END Data_PMOS[838]
  PIN Data_PMOS[837]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8128.745 187.44 8129.025 188.44 ;
    END
  END Data_PMOS[837]
  PIN Data_PMOS[836]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8057.065 187.44 8057.345 188.44 ;
    END
  END Data_PMOS[836]
  PIN Data_PMOS[835]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8059.305 187.44 8059.585 188.44 ;
    END
  END Data_PMOS[835]
  PIN Data_PMOS[834]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8060.985 187.44 8061.265 188.44 ;
    END
  END Data_PMOS[834]
  PIN Data_PMOS[833]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8111.945 187.44 8112.225 188.44 ;
    END
  END Data_PMOS[833]
  PIN Data_PMOS[832]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8113.065 187.44 8113.345 188.44 ;
    END
  END Data_PMOS[832]
  PIN Data_PMOS[831]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8114.745 187.44 8115.025 188.44 ;
    END
  END Data_PMOS[831]
  PIN Data_PMOS[830]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8058.745 187.44 8059.025 188.44 ;
    END
  END Data_PMOS[830]
  PIN Data_PMOS[829]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8060.425 187.44 8060.705 188.44 ;
    END
  END Data_PMOS[829]
  PIN Data_PMOS[828]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8061.545 187.44 8061.825 188.44 ;
    END
  END Data_PMOS[828]
  PIN Data_PMOS[827]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8128.185 187.44 8128.465 188.44 ;
    END
  END Data_PMOS[827]
  PIN Data_PMOS[826]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8111.385 187.44 8111.665 188.44 ;
    END
  END Data_PMOS[826]
  PIN Data_PMOS[825]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8110.825 187.44 8111.105 188.44 ;
    END
  END Data_PMOS[825]
  PIN Data_PMOS[824]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8113.625 187.44 8113.905 188.44 ;
    END
  END Data_PMOS[824]
  PIN Data_PMOS[823]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8059.865 187.44 8060.145 188.44 ;
    END
  END Data_PMOS[823]
  PIN Data_PMOS[822]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8062.665 187.44 8062.945 188.44 ;
    END
  END Data_PMOS[822]
  PIN Data_PMOS[821]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8062.105 187.44 8062.385 188.44 ;
    END
  END Data_PMOS[821]
  PIN Data_PMOS[820]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8058.185 187.44 8058.465 188.44 ;
    END
  END Data_PMOS[820]
  PIN Data_PMOS[819]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8057.625 187.44 8057.905 188.44 ;
    END
  END Data_PMOS[819]
  PIN Data_PMOS[818]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8035.785 187.44 8036.065 188.44 ;
    END
  END Data_PMOS[818]
  PIN Data_PMOS[817]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8037.465 187.44 8037.745 188.44 ;
    END
  END Data_PMOS[817]
  PIN Data_PMOS[816]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8039.145 187.44 8039.425 188.44 ;
    END
  END Data_PMOS[816]
  PIN Data_PMOS[815]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7991.545 187.44 7991.825 188.44 ;
    END
  END Data_PMOS[815]
  PIN Data_PMOS[814]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7993.785 187.44 7994.065 188.44 ;
    END
  END Data_PMOS[814]
  PIN Data_PMOS[813]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7995.465 187.44 7995.745 188.44 ;
    END
  END Data_PMOS[813]
  PIN Data_PMOS[812]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8035.225 187.44 8035.505 188.44 ;
    END
  END Data_PMOS[812]
  PIN Data_PMOS[811]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8036.345 187.44 8036.625 188.44 ;
    END
  END Data_PMOS[811]
  PIN Data_PMOS[810]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8038.025 187.44 8038.305 188.44 ;
    END
  END Data_PMOS[810]
  PIN Data_PMOS[809]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7993.225 187.44 7993.505 188.44 ;
    END
  END Data_PMOS[809]
  PIN Data_PMOS[808]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7994.905 187.44 7995.185 188.44 ;
    END
  END Data_PMOS[808]
  PIN Data_PMOS[807]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7996.025 187.44 7996.305 188.44 ;
    END
  END Data_PMOS[807]
  PIN Data_PMOS[806]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8038.585 187.44 8038.865 188.44 ;
    END
  END Data_PMOS[806]
  PIN Data_PMOS[805]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8034.665 187.44 8034.945 188.44 ;
    END
  END Data_PMOS[805]
  PIN Data_PMOS[804]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8034.105 187.44 8034.385 188.44 ;
    END
  END Data_PMOS[804]
  PIN Data_PMOS[803]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8036.905 187.44 8037.185 188.44 ;
    END
  END Data_PMOS[803]
  PIN Data_PMOS[802]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7994.345 187.44 7994.625 188.44 ;
    END
  END Data_PMOS[802]
  PIN Data_PMOS[801]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7997.145 187.44 7997.425 188.44 ;
    END
  END Data_PMOS[801]
  PIN Data_PMOS[800]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7996.585 187.44 7996.865 188.44 ;
    END
  END Data_PMOS[800]
  PIN Data_PMOS[799]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7992.665 187.44 7992.945 188.44 ;
    END
  END Data_PMOS[799]
  PIN Data_PMOS[798]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7992.105 187.44 7992.385 188.44 ;
    END
  END Data_PMOS[798]
  PIN Data_PMOS[797]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7965.785 187.44 7966.065 188.44 ;
    END
  END Data_PMOS[797]
  PIN Data_PMOS[796]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7967.465 187.44 7967.745 188.44 ;
    END
  END Data_PMOS[796]
  PIN Data_PMOS[795]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7969.145 187.44 7969.425 188.44 ;
    END
  END Data_PMOS[795]
  PIN Data_PMOS[794]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7909.785 187.44 7910.065 188.44 ;
    END
  END Data_PMOS[794]
  PIN Data_PMOS[793]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7912.025 187.44 7912.305 188.44 ;
    END
  END Data_PMOS[793]
  PIN Data_PMOS[792]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7913.705 187.44 7913.985 188.44 ;
    END
  END Data_PMOS[792]
  PIN Data_PMOS[791]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7965.225 187.44 7965.505 188.44 ;
    END
  END Data_PMOS[791]
  PIN Data_PMOS[790]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7966.345 187.44 7966.625 188.44 ;
    END
  END Data_PMOS[790]
  PIN Data_PMOS[789]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7968.025 187.44 7968.305 188.44 ;
    END
  END Data_PMOS[789]
  PIN Data_PMOS[788]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7911.465 187.44 7911.745 188.44 ;
    END
  END Data_PMOS[788]
  PIN Data_PMOS[787]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7913.145 187.44 7913.425 188.44 ;
    END
  END Data_PMOS[787]
  PIN Data_PMOS[786]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7914.265 187.44 7914.545 188.44 ;
    END
  END Data_PMOS[786]
  PIN Data_PMOS[785]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7968.585 187.44 7968.865 188.44 ;
    END
  END Data_PMOS[785]
  PIN Data_PMOS[784]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7964.665 187.44 7964.945 188.44 ;
    END
  END Data_PMOS[784]
  PIN Data_PMOS[783]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7964.105 187.44 7964.385 188.44 ;
    END
  END Data_PMOS[783]
  PIN Data_PMOS[782]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7966.905 187.44 7967.185 188.44 ;
    END
  END Data_PMOS[782]
  PIN Data_PMOS[781]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7912.585 187.44 7912.865 188.44 ;
    END
  END Data_PMOS[781]
  PIN Data_PMOS[780]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7915.385 187.44 7915.665 188.44 ;
    END
  END Data_PMOS[780]
  PIN Data_PMOS[779]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7914.825 187.44 7915.105 188.44 ;
    END
  END Data_PMOS[779]
  PIN Data_PMOS[778]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7910.905 187.44 7911.185 188.44 ;
    END
  END Data_PMOS[778]
  PIN Data_PMOS[777]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7910.345 187.44 7910.625 188.44 ;
    END
  END Data_PMOS[777]
  PIN Data_PMOS[776]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7861.065 187.44 7861.345 188.44 ;
    END
  END Data_PMOS[776]
  PIN Data_PMOS[775]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7888.225 187.44 7888.505 188.44 ;
    END
  END Data_PMOS[775]
  PIN Data_PMOS[774]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7889.905 187.44 7890.185 188.44 ;
    END
  END Data_PMOS[774]
  PIN Data_PMOS[773]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7831.385 187.44 7831.665 188.44 ;
    END
  END Data_PMOS[773]
  PIN Data_PMOS[772]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7833.625 187.44 7833.905 188.44 ;
    END
  END Data_PMOS[772]
  PIN Data_PMOS[771]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7835.305 187.44 7835.585 188.44 ;
    END
  END Data_PMOS[771]
  PIN Data_PMOS[770]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7860.505 187.44 7860.785 188.44 ;
    END
  END Data_PMOS[770]
  PIN Data_PMOS[769]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7861.625 187.44 7861.905 188.44 ;
    END
  END Data_PMOS[769]
  PIN Data_PMOS[768]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7888.785 187.44 7889.065 188.44 ;
    END
  END Data_PMOS[768]
  PIN Data_PMOS[767]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7833.065 187.44 7833.345 188.44 ;
    END
  END Data_PMOS[767]
  PIN Data_PMOS[766]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7834.745 187.44 7835.025 188.44 ;
    END
  END Data_PMOS[766]
  PIN Data_PMOS[765]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7848.745 187.44 7849.025 188.44 ;
    END
  END Data_PMOS[765]
  PIN Data_PMOS[764]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7889.345 187.44 7889.625 188.44 ;
    END
  END Data_PMOS[764]
  PIN Data_PMOS[763]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7859.945 187.44 7860.225 188.44 ;
    END
  END Data_PMOS[763]
  PIN Data_PMOS[762]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7859.385 187.44 7859.665 188.44 ;
    END
  END Data_PMOS[762]
  PIN Data_PMOS[761]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7887.665 187.44 7887.945 188.44 ;
    END
  END Data_PMOS[761]
  PIN Data_PMOS[760]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7834.185 187.44 7834.465 188.44 ;
    END
  END Data_PMOS[760]
  PIN Data_PMOS[759]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7849.865 187.44 7850.145 188.44 ;
    END
  END Data_PMOS[759]
  PIN Data_PMOS[758]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7849.305 187.44 7849.585 188.44 ;
    END
  END Data_PMOS[758]
  PIN Data_PMOS[757]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7832.505 187.44 7832.785 188.44 ;
    END
  END Data_PMOS[757]
  PIN Data_PMOS[756]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7831.945 187.44 7832.225 188.44 ;
    END
  END Data_PMOS[756]
  PIN Data_PMOS[755]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7778.745 187.44 7779.025 188.44 ;
    END
  END Data_PMOS[755]
  PIN Data_PMOS[754]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7780.425 187.44 7780.705 188.44 ;
    END
  END Data_PMOS[754]
  PIN Data_PMOS[753]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7782.105 187.44 7782.385 188.44 ;
    END
  END Data_PMOS[753]
  PIN Data_PMOS[752]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7753.545 187.44 7753.825 188.44 ;
    END
  END Data_PMOS[752]
  PIN Data_PMOS[751]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7755.785 187.44 7756.065 188.44 ;
    END
  END Data_PMOS[751]
  PIN Data_PMOS[750]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7757.465 187.44 7757.745 188.44 ;
    END
  END Data_PMOS[750]
  PIN Data_PMOS[749]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7778.185 187.44 7778.465 188.44 ;
    END
  END Data_PMOS[749]
  PIN Data_PMOS[748]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7779.305 187.44 7779.585 188.44 ;
    END
  END Data_PMOS[748]
  PIN Data_PMOS[747]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7780.985 187.44 7781.265 188.44 ;
    END
  END Data_PMOS[747]
  PIN Data_PMOS[746]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7755.225 187.44 7755.505 188.44 ;
    END
  END Data_PMOS[746]
  PIN Data_PMOS[745]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7756.905 187.44 7757.185 188.44 ;
    END
  END Data_PMOS[745]
  PIN Data_PMOS[744]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7758.025 187.44 7758.305 188.44 ;
    END
  END Data_PMOS[744]
  PIN Data_PMOS[743]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7781.545 187.44 7781.825 188.44 ;
    END
  END Data_PMOS[743]
  PIN Data_PMOS[742]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7777.625 187.44 7777.905 188.44 ;
    END
  END Data_PMOS[742]
  PIN Data_PMOS[741]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7777.065 187.44 7777.345 188.44 ;
    END
  END Data_PMOS[741]
  PIN Data_PMOS[740]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7779.865 187.44 7780.145 188.44 ;
    END
  END Data_PMOS[740]
  PIN Data_PMOS[739]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7756.345 187.44 7756.625 188.44 ;
    END
  END Data_PMOS[739]
  PIN Data_PMOS[738]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7759.145 187.44 7759.425 188.44 ;
    END
  END Data_PMOS[738]
  PIN Data_PMOS[737]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7758.585 187.44 7758.865 188.44 ;
    END
  END Data_PMOS[737]
  PIN Data_PMOS[736]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7754.665 187.44 7754.945 188.44 ;
    END
  END Data_PMOS[736]
  PIN Data_PMOS[735]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7754.105 187.44 7754.385 188.44 ;
    END
  END Data_PMOS[735]
  PIN Data_PMOS[734]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7712.665 187.44 7712.945 188.44 ;
    END
  END Data_PMOS[734]
  PIN Data_PMOS[733]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7714.345 187.44 7714.625 188.44 ;
    END
  END Data_PMOS[733]
  PIN Data_PMOS[732]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7716.025 187.44 7716.305 188.44 ;
    END
  END Data_PMOS[732]
  PIN Data_PMOS[731]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7682.425 187.44 7682.705 188.44 ;
    END
  END Data_PMOS[731]
  PIN Data_PMOS[730]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7684.665 187.44 7684.945 188.44 ;
    END
  END Data_PMOS[730]
  PIN Data_PMOS[729]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7686.345 187.44 7686.625 188.44 ;
    END
  END Data_PMOS[729]
  PIN Data_PMOS[728]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7712.105 187.44 7712.385 188.44 ;
    END
  END Data_PMOS[728]
  PIN Data_PMOS[727]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7713.225 187.44 7713.505 188.44 ;
    END
  END Data_PMOS[727]
  PIN Data_PMOS[726]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7714.905 187.44 7715.185 188.44 ;
    END
  END Data_PMOS[726]
  PIN Data_PMOS[725]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7684.105 187.44 7684.385 188.44 ;
    END
  END Data_PMOS[725]
  PIN Data_PMOS[724]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7685.785 187.44 7686.065 188.44 ;
    END
  END Data_PMOS[724]
  PIN Data_PMOS[723]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7686.905 187.44 7687.185 188.44 ;
    END
  END Data_PMOS[723]
  PIN Data_PMOS[722]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7715.465 187.44 7715.745 188.44 ;
    END
  END Data_PMOS[722]
  PIN Data_PMOS[721]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7711.545 187.44 7711.825 188.44 ;
    END
  END Data_PMOS[721]
  PIN Data_PMOS[720]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7710.985 187.44 7711.265 188.44 ;
    END
  END Data_PMOS[720]
  PIN Data_PMOS[719]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7713.785 187.44 7714.065 188.44 ;
    END
  END Data_PMOS[719]
  PIN Data_PMOS[718]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7685.225 187.44 7685.505 188.44 ;
    END
  END Data_PMOS[718]
  PIN Data_PMOS[717]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7688.025 187.44 7688.305 188.44 ;
    END
  END Data_PMOS[717]
  PIN Data_PMOS[716]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7687.465 187.44 7687.745 188.44 ;
    END
  END Data_PMOS[716]
  PIN Data_PMOS[715]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7683.545 187.44 7683.825 188.44 ;
    END
  END Data_PMOS[715]
  PIN Data_PMOS[714]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7682.985 187.44 7683.265 188.44 ;
    END
  END Data_PMOS[714]
  PIN Data_PMOS[713]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7630.905 187.44 7631.185 188.44 ;
    END
  END Data_PMOS[713]
  PIN Data_PMOS[712]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7632.585 187.44 7632.865 188.44 ;
    END
  END Data_PMOS[712]
  PIN Data_PMOS[711]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7634.265 187.44 7634.545 188.44 ;
    END
  END Data_PMOS[711]
  PIN Data_PMOS[710]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7578.265 187.44 7578.545 188.44 ;
    END
  END Data_PMOS[710]
  PIN Data_PMOS[709]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7580.505 187.44 7580.785 188.44 ;
    END
  END Data_PMOS[709]
  PIN Data_PMOS[708]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7607.665 187.44 7607.945 188.44 ;
    END
  END Data_PMOS[708]
  PIN Data_PMOS[707]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7630.345 187.44 7630.625 188.44 ;
    END
  END Data_PMOS[707]
  PIN Data_PMOS[706]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7631.465 187.44 7631.745 188.44 ;
    END
  END Data_PMOS[706]
  PIN Data_PMOS[705]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7633.145 187.44 7633.425 188.44 ;
    END
  END Data_PMOS[705]
  PIN Data_PMOS[704]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7579.945 187.44 7580.225 188.44 ;
    END
  END Data_PMOS[704]
  PIN Data_PMOS[703]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7607.105 187.44 7607.385 188.44 ;
    END
  END Data_PMOS[703]
  PIN Data_PMOS[702]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7608.225 187.44 7608.505 188.44 ;
    END
  END Data_PMOS[702]
  PIN Data_PMOS[701]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7633.705 187.44 7633.985 188.44 ;
    END
  END Data_PMOS[701]
  PIN Data_PMOS[700]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7629.785 187.44 7630.065 188.44 ;
    END
  END Data_PMOS[700]
  PIN Data_PMOS[699]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7620.825 187.44 7621.105 188.44 ;
    END
  END Data_PMOS[699]
  PIN Data_PMOS[698]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7632.025 187.44 7632.305 188.44 ;
    END
  END Data_PMOS[698]
  PIN Data_PMOS[697]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7581.065 187.44 7581.345 188.44 ;
    END
  END Data_PMOS[697]
  PIN Data_PMOS[696]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7609.345 187.44 7609.625 188.44 ;
    END
  END Data_PMOS[696]
  PIN Data_PMOS[695]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7608.785 187.44 7609.065 188.44 ;
    END
  END Data_PMOS[695]
  PIN Data_PMOS[694]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7579.385 187.44 7579.665 188.44 ;
    END
  END Data_PMOS[694]
  PIN Data_PMOS[693]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7578.825 187.44 7579.105 188.44 ;
    END
  END Data_PMOS[693]
  PIN Data_PMOS[692]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7552.505 187.44 7552.785 188.44 ;
    END
  END Data_PMOS[692]
  PIN Data_PMOS[691]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7554.185 187.44 7554.465 188.44 ;
    END
  END Data_PMOS[691]
  PIN Data_PMOS[690]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7568.745 187.44 7569.025 188.44 ;
    END
  END Data_PMOS[690]
  PIN Data_PMOS[689]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7497.065 187.44 7497.345 188.44 ;
    END
  END Data_PMOS[689]
  PIN Data_PMOS[688]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7499.305 187.44 7499.585 188.44 ;
    END
  END Data_PMOS[688]
  PIN Data_PMOS[687]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7500.985 187.44 7501.265 188.44 ;
    END
  END Data_PMOS[687]
  PIN Data_PMOS[686]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7551.945 187.44 7552.225 188.44 ;
    END
  END Data_PMOS[686]
  PIN Data_PMOS[685]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7553.065 187.44 7553.345 188.44 ;
    END
  END Data_PMOS[685]
  PIN Data_PMOS[684]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7554.745 187.44 7555.025 188.44 ;
    END
  END Data_PMOS[684]
  PIN Data_PMOS[683]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7498.745 187.44 7499.025 188.44 ;
    END
  END Data_PMOS[683]
  PIN Data_PMOS[682]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7500.425 187.44 7500.705 188.44 ;
    END
  END Data_PMOS[682]
  PIN Data_PMOS[681]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7501.545 187.44 7501.825 188.44 ;
    END
  END Data_PMOS[681]
  PIN Data_PMOS[680]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7568.185 187.44 7568.465 188.44 ;
    END
  END Data_PMOS[680]
  PIN Data_PMOS[679]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7551.385 187.44 7551.665 188.44 ;
    END
  END Data_PMOS[679]
  PIN Data_PMOS[678]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7550.825 187.44 7551.105 188.44 ;
    END
  END Data_PMOS[678]
  PIN Data_PMOS[677]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7553.625 187.44 7553.905 188.44 ;
    END
  END Data_PMOS[677]
  PIN Data_PMOS[676]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7499.865 187.44 7500.145 188.44 ;
    END
  END Data_PMOS[676]
  PIN Data_PMOS[675]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7502.665 187.44 7502.945 188.44 ;
    END
  END Data_PMOS[675]
  PIN Data_PMOS[674]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7502.105 187.44 7502.385 188.44 ;
    END
  END Data_PMOS[674]
  PIN Data_PMOS[673]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7498.185 187.44 7498.465 188.44 ;
    END
  END Data_PMOS[673]
  PIN Data_PMOS[672]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7497.625 187.44 7497.905 188.44 ;
    END
  END Data_PMOS[672]
  PIN Data_PMOS[671]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7475.785 187.44 7476.065 188.44 ;
    END
  END Data_PMOS[671]
  PIN Data_PMOS[670]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7477.465 187.44 7477.745 188.44 ;
    END
  END Data_PMOS[670]
  PIN Data_PMOS[669]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7479.145 187.44 7479.425 188.44 ;
    END
  END Data_PMOS[669]
  PIN Data_PMOS[668]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7431.545 187.44 7431.825 188.44 ;
    END
  END Data_PMOS[668]
  PIN Data_PMOS[667]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7433.785 187.44 7434.065 188.44 ;
    END
  END Data_PMOS[667]
  PIN Data_PMOS[666]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7435.465 187.44 7435.745 188.44 ;
    END
  END Data_PMOS[666]
  PIN Data_PMOS[665]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7475.225 187.44 7475.505 188.44 ;
    END
  END Data_PMOS[665]
  PIN Data_PMOS[664]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7476.345 187.44 7476.625 188.44 ;
    END
  END Data_PMOS[664]
  PIN Data_PMOS[663]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7478.025 187.44 7478.305 188.44 ;
    END
  END Data_PMOS[663]
  PIN Data_PMOS[662]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7433.225 187.44 7433.505 188.44 ;
    END
  END Data_PMOS[662]
  PIN Data_PMOS[661]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7434.905 187.44 7435.185 188.44 ;
    END
  END Data_PMOS[661]
  PIN Data_PMOS[660]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7436.025 187.44 7436.305 188.44 ;
    END
  END Data_PMOS[660]
  PIN Data_PMOS[659]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7478.585 187.44 7478.865 188.44 ;
    END
  END Data_PMOS[659]
  PIN Data_PMOS[658]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7474.665 187.44 7474.945 188.44 ;
    END
  END Data_PMOS[658]
  PIN Data_PMOS[657]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7474.105 187.44 7474.385 188.44 ;
    END
  END Data_PMOS[657]
  PIN Data_PMOS[656]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7476.905 187.44 7477.185 188.44 ;
    END
  END Data_PMOS[656]
  PIN Data_PMOS[655]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7434.345 187.44 7434.625 188.44 ;
    END
  END Data_PMOS[655]
  PIN Data_PMOS[654]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7437.145 187.44 7437.425 188.44 ;
    END
  END Data_PMOS[654]
  PIN Data_PMOS[653]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7436.585 187.44 7436.865 188.44 ;
    END
  END Data_PMOS[653]
  PIN Data_PMOS[652]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7432.665 187.44 7432.945 188.44 ;
    END
  END Data_PMOS[652]
  PIN Data_PMOS[651]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7432.105 187.44 7432.385 188.44 ;
    END
  END Data_PMOS[651]
  PIN Data_PMOS[650]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7405.785 187.44 7406.065 188.44 ;
    END
  END Data_PMOS[650]
  PIN Data_PMOS[649]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7407.465 187.44 7407.745 188.44 ;
    END
  END Data_PMOS[649]
  PIN Data_PMOS[648]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7409.145 187.44 7409.425 188.44 ;
    END
  END Data_PMOS[648]
  PIN Data_PMOS[647]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7349.785 187.44 7350.065 188.44 ;
    END
  END Data_PMOS[647]
  PIN Data_PMOS[646]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7352.025 187.44 7352.305 188.44 ;
    END
  END Data_PMOS[646]
  PIN Data_PMOS[645]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7353.705 187.44 7353.985 188.44 ;
    END
  END Data_PMOS[645]
  PIN Data_PMOS[644]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7405.225 187.44 7405.505 188.44 ;
    END
  END Data_PMOS[644]
  PIN Data_PMOS[643]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7406.345 187.44 7406.625 188.44 ;
    END
  END Data_PMOS[643]
  PIN Data_PMOS[642]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7408.025 187.44 7408.305 188.44 ;
    END
  END Data_PMOS[642]
  PIN Data_PMOS[641]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7351.465 187.44 7351.745 188.44 ;
    END
  END Data_PMOS[641]
  PIN Data_PMOS[640]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7353.145 187.44 7353.425 188.44 ;
    END
  END Data_PMOS[640]
  PIN Data_PMOS[639]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7354.265 187.44 7354.545 188.44 ;
    END
  END Data_PMOS[639]
  PIN Data_PMOS[638]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7408.585 187.44 7408.865 188.44 ;
    END
  END Data_PMOS[638]
  PIN Data_PMOS[637]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7404.665 187.44 7404.945 188.44 ;
    END
  END Data_PMOS[637]
  PIN Data_PMOS[636]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7404.105 187.44 7404.385 188.44 ;
    END
  END Data_PMOS[636]
  PIN Data_PMOS[635]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7406.905 187.44 7407.185 188.44 ;
    END
  END Data_PMOS[635]
  PIN Data_PMOS[634]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7352.585 187.44 7352.865 188.44 ;
    END
  END Data_PMOS[634]
  PIN Data_PMOS[633]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7355.385 187.44 7355.665 188.44 ;
    END
  END Data_PMOS[633]
  PIN Data_PMOS[632]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7354.825 187.44 7355.105 188.44 ;
    END
  END Data_PMOS[632]
  PIN Data_PMOS[631]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7350.905 187.44 7351.185 188.44 ;
    END
  END Data_PMOS[631]
  PIN Data_PMOS[630]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7350.345 187.44 7350.625 188.44 ;
    END
  END Data_PMOS[630]
  PIN Data_PMOS[629]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7301.065 187.44 7301.345 188.44 ;
    END
  END Data_PMOS[629]
  PIN Data_PMOS[628]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7328.225 187.44 7328.505 188.44 ;
    END
  END Data_PMOS[628]
  PIN Data_PMOS[627]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7329.905 187.44 7330.185 188.44 ;
    END
  END Data_PMOS[627]
  PIN Data_PMOS[626]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7271.385 187.44 7271.665 188.44 ;
    END
  END Data_PMOS[626]
  PIN Data_PMOS[625]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7273.625 187.44 7273.905 188.44 ;
    END
  END Data_PMOS[625]
  PIN Data_PMOS[624]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7275.305 187.44 7275.585 188.44 ;
    END
  END Data_PMOS[624]
  PIN Data_PMOS[623]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7300.505 187.44 7300.785 188.44 ;
    END
  END Data_PMOS[623]
  PIN Data_PMOS[622]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7301.625 187.44 7301.905 188.44 ;
    END
  END Data_PMOS[622]
  PIN Data_PMOS[621]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7328.785 187.44 7329.065 188.44 ;
    END
  END Data_PMOS[621]
  PIN Data_PMOS[620]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7273.065 187.44 7273.345 188.44 ;
    END
  END Data_PMOS[620]
  PIN Data_PMOS[619]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7274.745 187.44 7275.025 188.44 ;
    END
  END Data_PMOS[619]
  PIN Data_PMOS[618]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7288.745 187.44 7289.025 188.44 ;
    END
  END Data_PMOS[618]
  PIN Data_PMOS[617]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7329.345 187.44 7329.625 188.44 ;
    END
  END Data_PMOS[617]
  PIN Data_PMOS[616]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7299.945 187.44 7300.225 188.44 ;
    END
  END Data_PMOS[616]
  PIN Data_PMOS[615]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7299.385 187.44 7299.665 188.44 ;
    END
  END Data_PMOS[615]
  PIN Data_PMOS[614]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7327.665 187.44 7327.945 188.44 ;
    END
  END Data_PMOS[614]
  PIN Data_PMOS[613]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7274.185 187.44 7274.465 188.44 ;
    END
  END Data_PMOS[613]
  PIN Data_PMOS[612]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7289.865 187.44 7290.145 188.44 ;
    END
  END Data_PMOS[612]
  PIN Data_PMOS[611]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7289.305 187.44 7289.585 188.44 ;
    END
  END Data_PMOS[611]
  PIN Data_PMOS[610]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7272.505 187.44 7272.785 188.44 ;
    END
  END Data_PMOS[610]
  PIN Data_PMOS[609]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7271.945 187.44 7272.225 188.44 ;
    END
  END Data_PMOS[609]
  PIN Data_PMOS[608]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7218.745 187.44 7219.025 188.44 ;
    END
  END Data_PMOS[608]
  PIN Data_PMOS[607]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7220.425 187.44 7220.705 188.44 ;
    END
  END Data_PMOS[607]
  PIN Data_PMOS[606]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7222.105 187.44 7222.385 188.44 ;
    END
  END Data_PMOS[606]
  PIN Data_PMOS[605]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7193.545 187.44 7193.825 188.44 ;
    END
  END Data_PMOS[605]
  PIN Data_PMOS[604]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7195.785 187.44 7196.065 188.44 ;
    END
  END Data_PMOS[604]
  PIN Data_PMOS[603]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7197.465 187.44 7197.745 188.44 ;
    END
  END Data_PMOS[603]
  PIN Data_PMOS[602]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7218.185 187.44 7218.465 188.44 ;
    END
  END Data_PMOS[602]
  PIN Data_PMOS[601]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7219.305 187.44 7219.585 188.44 ;
    END
  END Data_PMOS[601]
  PIN Data_PMOS[600]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7220.985 187.44 7221.265 188.44 ;
    END
  END Data_PMOS[600]
  PIN Data_PMOS[599]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7195.225 187.44 7195.505 188.44 ;
    END
  END Data_PMOS[599]
  PIN Data_PMOS[598]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7196.905 187.44 7197.185 188.44 ;
    END
  END Data_PMOS[598]
  PIN Data_PMOS[597]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7198.025 187.44 7198.305 188.44 ;
    END
  END Data_PMOS[597]
  PIN Data_PMOS[596]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7221.545 187.44 7221.825 188.44 ;
    END
  END Data_PMOS[596]
  PIN Data_PMOS[595]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7217.625 187.44 7217.905 188.44 ;
    END
  END Data_PMOS[595]
  PIN Data_PMOS[594]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7217.065 187.44 7217.345 188.44 ;
    END
  END Data_PMOS[594]
  PIN Data_PMOS[593]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7219.865 187.44 7220.145 188.44 ;
    END
  END Data_PMOS[593]
  PIN Data_PMOS[592]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7196.345 187.44 7196.625 188.44 ;
    END
  END Data_PMOS[592]
  PIN Data_PMOS[591]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7199.145 187.44 7199.425 188.44 ;
    END
  END Data_PMOS[591]
  PIN Data_PMOS[590]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7198.585 187.44 7198.865 188.44 ;
    END
  END Data_PMOS[590]
  PIN Data_PMOS[589]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7194.665 187.44 7194.945 188.44 ;
    END
  END Data_PMOS[589]
  PIN Data_PMOS[588]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7194.105 187.44 7194.385 188.44 ;
    END
  END Data_PMOS[588]
  PIN Data_PMOS[587]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7152.665 187.44 7152.945 188.44 ;
    END
  END Data_PMOS[587]
  PIN Data_PMOS[586]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7154.345 187.44 7154.625 188.44 ;
    END
  END Data_PMOS[586]
  PIN Data_PMOS[585]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7156.025 187.44 7156.305 188.44 ;
    END
  END Data_PMOS[585]
  PIN Data_PMOS[584]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7122.425 187.44 7122.705 188.44 ;
    END
  END Data_PMOS[584]
  PIN Data_PMOS[583]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7124.665 187.44 7124.945 188.44 ;
    END
  END Data_PMOS[583]
  PIN Data_PMOS[582]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7126.345 187.44 7126.625 188.44 ;
    END
  END Data_PMOS[582]
  PIN Data_PMOS[581]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7152.105 187.44 7152.385 188.44 ;
    END
  END Data_PMOS[581]
  PIN Data_PMOS[580]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7153.225 187.44 7153.505 188.44 ;
    END
  END Data_PMOS[580]
  PIN Data_PMOS[579]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7154.905 187.44 7155.185 188.44 ;
    END
  END Data_PMOS[579]
  PIN Data_PMOS[578]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7124.105 187.44 7124.385 188.44 ;
    END
  END Data_PMOS[578]
  PIN Data_PMOS[577]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7125.785 187.44 7126.065 188.44 ;
    END
  END Data_PMOS[577]
  PIN Data_PMOS[576]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7126.905 187.44 7127.185 188.44 ;
    END
  END Data_PMOS[576]
  PIN Data_PMOS[575]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7155.465 187.44 7155.745 188.44 ;
    END
  END Data_PMOS[575]
  PIN Data_PMOS[574]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7151.545 187.44 7151.825 188.44 ;
    END
  END Data_PMOS[574]
  PIN Data_PMOS[573]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7150.985 187.44 7151.265 188.44 ;
    END
  END Data_PMOS[573]
  PIN Data_PMOS[572]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7153.785 187.44 7154.065 188.44 ;
    END
  END Data_PMOS[572]
  PIN Data_PMOS[571]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7125.225 187.44 7125.505 188.44 ;
    END
  END Data_PMOS[571]
  PIN Data_PMOS[570]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7128.025 187.44 7128.305 188.44 ;
    END
  END Data_PMOS[570]
  PIN Data_PMOS[569]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7127.465 187.44 7127.745 188.44 ;
    END
  END Data_PMOS[569]
  PIN Data_PMOS[568]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7123.545 187.44 7123.825 188.44 ;
    END
  END Data_PMOS[568]
  PIN Data_PMOS[567]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7122.985 187.44 7123.265 188.44 ;
    END
  END Data_PMOS[567]
  PIN Data_PMOS[566]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7070.905 187.44 7071.185 188.44 ;
    END
  END Data_PMOS[566]
  PIN Data_PMOS[565]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7072.585 187.44 7072.865 188.44 ;
    END
  END Data_PMOS[565]
  PIN Data_PMOS[564]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7074.265 187.44 7074.545 188.44 ;
    END
  END Data_PMOS[564]
  PIN Data_PMOS[563]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7018.265 187.44 7018.545 188.44 ;
    END
  END Data_PMOS[563]
  PIN Data_PMOS[562]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7020.505 187.44 7020.785 188.44 ;
    END
  END Data_PMOS[562]
  PIN Data_PMOS[561]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7047.665 187.44 7047.945 188.44 ;
    END
  END Data_PMOS[561]
  PIN Data_PMOS[560]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7070.345 187.44 7070.625 188.44 ;
    END
  END Data_PMOS[560]
  PIN Data_PMOS[559]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7071.465 187.44 7071.745 188.44 ;
    END
  END Data_PMOS[559]
  PIN Data_PMOS[558]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7073.145 187.44 7073.425 188.44 ;
    END
  END Data_PMOS[558]
  PIN Data_PMOS[557]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7019.945 187.44 7020.225 188.44 ;
    END
  END Data_PMOS[557]
  PIN Data_PMOS[556]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7047.105 187.44 7047.385 188.44 ;
    END
  END Data_PMOS[556]
  PIN Data_PMOS[555]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7048.225 187.44 7048.505 188.44 ;
    END
  END Data_PMOS[555]
  PIN Data_PMOS[554]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7073.705 187.44 7073.985 188.44 ;
    END
  END Data_PMOS[554]
  PIN Data_PMOS[553]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7069.785 187.44 7070.065 188.44 ;
    END
  END Data_PMOS[553]
  PIN Data_PMOS[552]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7060.825 187.44 7061.105 188.44 ;
    END
  END Data_PMOS[552]
  PIN Data_PMOS[551]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7072.025 187.44 7072.305 188.44 ;
    END
  END Data_PMOS[551]
  PIN Data_PMOS[550]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7021.065 187.44 7021.345 188.44 ;
    END
  END Data_PMOS[550]
  PIN Data_PMOS[549]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7049.345 187.44 7049.625 188.44 ;
    END
  END Data_PMOS[549]
  PIN Data_PMOS[548]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7048.785 187.44 7049.065 188.44 ;
    END
  END Data_PMOS[548]
  PIN Data_PMOS[547]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7019.385 187.44 7019.665 188.44 ;
    END
  END Data_PMOS[547]
  PIN Data_PMOS[546]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7018.825 187.44 7019.105 188.44 ;
    END
  END Data_PMOS[546]
  PIN Data_PMOS[545]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6992.505 187.44 6992.785 188.44 ;
    END
  END Data_PMOS[545]
  PIN Data_PMOS[544]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6994.185 187.44 6994.465 188.44 ;
    END
  END Data_PMOS[544]
  PIN Data_PMOS[543]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7008.745 187.44 7009.025 188.44 ;
    END
  END Data_PMOS[543]
  PIN Data_PMOS[542]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6937.065 187.44 6937.345 188.44 ;
    END
  END Data_PMOS[542]
  PIN Data_PMOS[541]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6939.305 187.44 6939.585 188.44 ;
    END
  END Data_PMOS[541]
  PIN Data_PMOS[540]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6940.985 187.44 6941.265 188.44 ;
    END
  END Data_PMOS[540]
  PIN Data_PMOS[539]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6991.945 187.44 6992.225 188.44 ;
    END
  END Data_PMOS[539]
  PIN Data_PMOS[538]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6993.065 187.44 6993.345 188.44 ;
    END
  END Data_PMOS[538]
  PIN Data_PMOS[537]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6994.745 187.44 6995.025 188.44 ;
    END
  END Data_PMOS[537]
  PIN Data_PMOS[536]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6938.745 187.44 6939.025 188.44 ;
    END
  END Data_PMOS[536]
  PIN Data_PMOS[535]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6940.425 187.44 6940.705 188.44 ;
    END
  END Data_PMOS[535]
  PIN Data_PMOS[534]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6941.545 187.44 6941.825 188.44 ;
    END
  END Data_PMOS[534]
  PIN Data_PMOS[533]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7008.185 187.44 7008.465 188.44 ;
    END
  END Data_PMOS[533]
  PIN Data_PMOS[532]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6991.385 187.44 6991.665 188.44 ;
    END
  END Data_PMOS[532]
  PIN Data_PMOS[531]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6990.825 187.44 6991.105 188.44 ;
    END
  END Data_PMOS[531]
  PIN Data_PMOS[530]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6993.625 187.44 6993.905 188.44 ;
    END
  END Data_PMOS[530]
  PIN Data_PMOS[529]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6939.865 187.44 6940.145 188.44 ;
    END
  END Data_PMOS[529]
  PIN Data_PMOS[528]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6942.665 187.44 6942.945 188.44 ;
    END
  END Data_PMOS[528]
  PIN Data_PMOS[527]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6942.105 187.44 6942.385 188.44 ;
    END
  END Data_PMOS[527]
  PIN Data_PMOS[526]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6938.185 187.44 6938.465 188.44 ;
    END
  END Data_PMOS[526]
  PIN Data_PMOS[525]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6937.625 187.44 6937.905 188.44 ;
    END
  END Data_PMOS[525]
  PIN Data_PMOS[524]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6915.785 187.44 6916.065 188.44 ;
    END
  END Data_PMOS[524]
  PIN Data_PMOS[523]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6917.465 187.44 6917.745 188.44 ;
    END
  END Data_PMOS[523]
  PIN Data_PMOS[522]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6919.145 187.44 6919.425 188.44 ;
    END
  END Data_PMOS[522]
  PIN Data_PMOS[521]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6871.545 187.44 6871.825 188.44 ;
    END
  END Data_PMOS[521]
  PIN Data_PMOS[520]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6873.785 187.44 6874.065 188.44 ;
    END
  END Data_PMOS[520]
  PIN Data_PMOS[519]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6875.465 187.44 6875.745 188.44 ;
    END
  END Data_PMOS[519]
  PIN Data_PMOS[518]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6915.225 187.44 6915.505 188.44 ;
    END
  END Data_PMOS[518]
  PIN Data_PMOS[517]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6916.345 187.44 6916.625 188.44 ;
    END
  END Data_PMOS[517]
  PIN Data_PMOS[516]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6918.025 187.44 6918.305 188.44 ;
    END
  END Data_PMOS[516]
  PIN Data_PMOS[515]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6873.225 187.44 6873.505 188.44 ;
    END
  END Data_PMOS[515]
  PIN Data_PMOS[514]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6874.905 187.44 6875.185 188.44 ;
    END
  END Data_PMOS[514]
  PIN Data_PMOS[513]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6876.025 187.44 6876.305 188.44 ;
    END
  END Data_PMOS[513]
  PIN Data_PMOS[512]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6918.585 187.44 6918.865 188.44 ;
    END
  END Data_PMOS[512]
  PIN Data_PMOS[511]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6914.665 187.44 6914.945 188.44 ;
    END
  END Data_PMOS[511]
  PIN Data_PMOS[510]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6914.105 187.44 6914.385 188.44 ;
    END
  END Data_PMOS[510]
  PIN Data_PMOS[509]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6916.905 187.44 6917.185 188.44 ;
    END
  END Data_PMOS[509]
  PIN Data_PMOS[508]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6874.345 187.44 6874.625 188.44 ;
    END
  END Data_PMOS[508]
  PIN Data_PMOS[507]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6877.145 187.44 6877.425 188.44 ;
    END
  END Data_PMOS[507]
  PIN Data_PMOS[506]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6876.585 187.44 6876.865 188.44 ;
    END
  END Data_PMOS[506]
  PIN Data_PMOS[505]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6872.665 187.44 6872.945 188.44 ;
    END
  END Data_PMOS[505]
  PIN Data_PMOS[504]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6872.105 187.44 6872.385 188.44 ;
    END
  END Data_PMOS[504]
  PIN Data_PMOS[503]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6845.785 187.44 6846.065 188.44 ;
    END
  END Data_PMOS[503]
  PIN Data_PMOS[502]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6847.465 187.44 6847.745 188.44 ;
    END
  END Data_PMOS[502]
  PIN Data_PMOS[501]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6849.145 187.44 6849.425 188.44 ;
    END
  END Data_PMOS[501]
  PIN Data_PMOS[500]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6789.785 187.44 6790.065 188.44 ;
    END
  END Data_PMOS[500]
  PIN Data_PMOS[499]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6792.025 187.44 6792.305 188.44 ;
    END
  END Data_PMOS[499]
  PIN Data_PMOS[498]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6793.705 187.44 6793.985 188.44 ;
    END
  END Data_PMOS[498]
  PIN Data_PMOS[497]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6845.225 187.44 6845.505 188.44 ;
    END
  END Data_PMOS[497]
  PIN Data_PMOS[496]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6846.345 187.44 6846.625 188.44 ;
    END
  END Data_PMOS[496]
  PIN Data_PMOS[495]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6848.025 187.44 6848.305 188.44 ;
    END
  END Data_PMOS[495]
  PIN Data_PMOS[494]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6791.465 187.44 6791.745 188.44 ;
    END
  END Data_PMOS[494]
  PIN Data_PMOS[493]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6793.145 187.44 6793.425 188.44 ;
    END
  END Data_PMOS[493]
  PIN Data_PMOS[492]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6794.265 187.44 6794.545 188.44 ;
    END
  END Data_PMOS[492]
  PIN Data_PMOS[491]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6848.585 187.44 6848.865 188.44 ;
    END
  END Data_PMOS[491]
  PIN Data_PMOS[490]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6844.665 187.44 6844.945 188.44 ;
    END
  END Data_PMOS[490]
  PIN Data_PMOS[489]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6844.105 187.44 6844.385 188.44 ;
    END
  END Data_PMOS[489]
  PIN Data_PMOS[488]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6846.905 187.44 6847.185 188.44 ;
    END
  END Data_PMOS[488]
  PIN Data_PMOS[487]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6792.585 187.44 6792.865 188.44 ;
    END
  END Data_PMOS[487]
  PIN Data_PMOS[486]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6795.385 187.44 6795.665 188.44 ;
    END
  END Data_PMOS[486]
  PIN Data_PMOS[485]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6794.825 187.44 6795.105 188.44 ;
    END
  END Data_PMOS[485]
  PIN Data_PMOS[484]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6790.905 187.44 6791.185 188.44 ;
    END
  END Data_PMOS[484]
  PIN Data_PMOS[483]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6790.345 187.44 6790.625 188.44 ;
    END
  END Data_PMOS[483]
  PIN Data_PMOS[482]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6741.065 187.44 6741.345 188.44 ;
    END
  END Data_PMOS[482]
  PIN Data_PMOS[481]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6768.225 187.44 6768.505 188.44 ;
    END
  END Data_PMOS[481]
  PIN Data_PMOS[480]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6769.905 187.44 6770.185 188.44 ;
    END
  END Data_PMOS[480]
  PIN Data_PMOS[479]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6711.385 187.44 6711.665 188.44 ;
    END
  END Data_PMOS[479]
  PIN Data_PMOS[478]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6713.625 187.44 6713.905 188.44 ;
    END
  END Data_PMOS[478]
  PIN Data_PMOS[477]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6715.305 187.44 6715.585 188.44 ;
    END
  END Data_PMOS[477]
  PIN Data_PMOS[476]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6740.505 187.44 6740.785 188.44 ;
    END
  END Data_PMOS[476]
  PIN Data_PMOS[475]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6741.625 187.44 6741.905 188.44 ;
    END
  END Data_PMOS[475]
  PIN Data_PMOS[474]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6768.785 187.44 6769.065 188.44 ;
    END
  END Data_PMOS[474]
  PIN Data_PMOS[473]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6713.065 187.44 6713.345 188.44 ;
    END
  END Data_PMOS[473]
  PIN Data_PMOS[472]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6714.745 187.44 6715.025 188.44 ;
    END
  END Data_PMOS[472]
  PIN Data_PMOS[471]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6728.745 187.44 6729.025 188.44 ;
    END
  END Data_PMOS[471]
  PIN Data_PMOS[470]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6769.345 187.44 6769.625 188.44 ;
    END
  END Data_PMOS[470]
  PIN Data_PMOS[469]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6739.945 187.44 6740.225 188.44 ;
    END
  END Data_PMOS[469]
  PIN Data_PMOS[468]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6739.385 187.44 6739.665 188.44 ;
    END
  END Data_PMOS[468]
  PIN Data_PMOS[467]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6767.665 187.44 6767.945 188.44 ;
    END
  END Data_PMOS[467]
  PIN Data_PMOS[466]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6714.185 187.44 6714.465 188.44 ;
    END
  END Data_PMOS[466]
  PIN Data_PMOS[465]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6729.865 187.44 6730.145 188.44 ;
    END
  END Data_PMOS[465]
  PIN Data_PMOS[464]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6729.305 187.44 6729.585 188.44 ;
    END
  END Data_PMOS[464]
  PIN Data_PMOS[463]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6712.505 187.44 6712.785 188.44 ;
    END
  END Data_PMOS[463]
  PIN Data_PMOS[462]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6711.945 187.44 6712.225 188.44 ;
    END
  END Data_PMOS[462]
  PIN Data_PMOS[461]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6658.745 187.44 6659.025 188.44 ;
    END
  END Data_PMOS[461]
  PIN Data_PMOS[460]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6660.425 187.44 6660.705 188.44 ;
    END
  END Data_PMOS[460]
  PIN Data_PMOS[459]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6662.105 187.44 6662.385 188.44 ;
    END
  END Data_PMOS[459]
  PIN Data_PMOS[458]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6633.545 187.44 6633.825 188.44 ;
    END
  END Data_PMOS[458]
  PIN Data_PMOS[457]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6635.785 187.44 6636.065 188.44 ;
    END
  END Data_PMOS[457]
  PIN Data_PMOS[456]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6637.465 187.44 6637.745 188.44 ;
    END
  END Data_PMOS[456]
  PIN Data_PMOS[455]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6658.185 187.44 6658.465 188.44 ;
    END
  END Data_PMOS[455]
  PIN Data_PMOS[454]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6659.305 187.44 6659.585 188.44 ;
    END
  END Data_PMOS[454]
  PIN Data_PMOS[453]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6660.985 187.44 6661.265 188.44 ;
    END
  END Data_PMOS[453]
  PIN Data_PMOS[452]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6635.225 187.44 6635.505 188.44 ;
    END
  END Data_PMOS[452]
  PIN Data_PMOS[451]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6636.905 187.44 6637.185 188.44 ;
    END
  END Data_PMOS[451]
  PIN Data_PMOS[450]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6638.025 187.44 6638.305 188.44 ;
    END
  END Data_PMOS[450]
  PIN Data_PMOS[449]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6661.545 187.44 6661.825 188.44 ;
    END
  END Data_PMOS[449]
  PIN Data_PMOS[448]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6657.625 187.44 6657.905 188.44 ;
    END
  END Data_PMOS[448]
  PIN Data_PMOS[447]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6657.065 187.44 6657.345 188.44 ;
    END
  END Data_PMOS[447]
  PIN Data_PMOS[446]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6659.865 187.44 6660.145 188.44 ;
    END
  END Data_PMOS[446]
  PIN Data_PMOS[445]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6636.345 187.44 6636.625 188.44 ;
    END
  END Data_PMOS[445]
  PIN Data_PMOS[444]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6639.145 187.44 6639.425 188.44 ;
    END
  END Data_PMOS[444]
  PIN Data_PMOS[443]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6638.585 187.44 6638.865 188.44 ;
    END
  END Data_PMOS[443]
  PIN Data_PMOS[442]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6634.665 187.44 6634.945 188.44 ;
    END
  END Data_PMOS[442]
  PIN Data_PMOS[441]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6634.105 187.44 6634.385 188.44 ;
    END
  END Data_PMOS[441]
  PIN Data_PMOS[440]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6592.665 187.44 6592.945 188.44 ;
    END
  END Data_PMOS[440]
  PIN Data_PMOS[439]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6594.345 187.44 6594.625 188.44 ;
    END
  END Data_PMOS[439]
  PIN Data_PMOS[438]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6596.025 187.44 6596.305 188.44 ;
    END
  END Data_PMOS[438]
  PIN Data_PMOS[437]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6562.425 187.44 6562.705 188.44 ;
    END
  END Data_PMOS[437]
  PIN Data_PMOS[436]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6564.665 187.44 6564.945 188.44 ;
    END
  END Data_PMOS[436]
  PIN Data_PMOS[435]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6566.345 187.44 6566.625 188.44 ;
    END
  END Data_PMOS[435]
  PIN Data_PMOS[434]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6592.105 187.44 6592.385 188.44 ;
    END
  END Data_PMOS[434]
  PIN Data_PMOS[433]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6593.225 187.44 6593.505 188.44 ;
    END
  END Data_PMOS[433]
  PIN Data_PMOS[432]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6594.905 187.44 6595.185 188.44 ;
    END
  END Data_PMOS[432]
  PIN Data_PMOS[431]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6564.105 187.44 6564.385 188.44 ;
    END
  END Data_PMOS[431]
  PIN Data_PMOS[430]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6565.785 187.44 6566.065 188.44 ;
    END
  END Data_PMOS[430]
  PIN Data_PMOS[429]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6566.905 187.44 6567.185 188.44 ;
    END
  END Data_PMOS[429]
  PIN Data_PMOS[428]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6595.465 187.44 6595.745 188.44 ;
    END
  END Data_PMOS[428]
  PIN Data_PMOS[427]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6591.545 187.44 6591.825 188.44 ;
    END
  END Data_PMOS[427]
  PIN Data_PMOS[426]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6590.985 187.44 6591.265 188.44 ;
    END
  END Data_PMOS[426]
  PIN Data_PMOS[425]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6593.785 187.44 6594.065 188.44 ;
    END
  END Data_PMOS[425]
  PIN Data_PMOS[424]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6565.225 187.44 6565.505 188.44 ;
    END
  END Data_PMOS[424]
  PIN Data_PMOS[423]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6568.025 187.44 6568.305 188.44 ;
    END
  END Data_PMOS[423]
  PIN Data_PMOS[422]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6567.465 187.44 6567.745 188.44 ;
    END
  END Data_PMOS[422]
  PIN Data_PMOS[421]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6563.545 187.44 6563.825 188.44 ;
    END
  END Data_PMOS[421]
  PIN Data_PMOS[420]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6562.985 187.44 6563.265 188.44 ;
    END
  END Data_PMOS[420]
  PIN Data_PMOS[419]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6510.905 187.44 6511.185 188.44 ;
    END
  END Data_PMOS[419]
  PIN Data_PMOS[418]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6512.585 187.44 6512.865 188.44 ;
    END
  END Data_PMOS[418]
  PIN Data_PMOS[417]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6514.265 187.44 6514.545 188.44 ;
    END
  END Data_PMOS[417]
  PIN Data_PMOS[416]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6458.265 187.44 6458.545 188.44 ;
    END
  END Data_PMOS[416]
  PIN Data_PMOS[415]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6460.505 187.44 6460.785 188.44 ;
    END
  END Data_PMOS[415]
  PIN Data_PMOS[414]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6487.665 187.44 6487.945 188.44 ;
    END
  END Data_PMOS[414]
  PIN Data_PMOS[413]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6510.345 187.44 6510.625 188.44 ;
    END
  END Data_PMOS[413]
  PIN Data_PMOS[412]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6511.465 187.44 6511.745 188.44 ;
    END
  END Data_PMOS[412]
  PIN Data_PMOS[411]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6513.145 187.44 6513.425 188.44 ;
    END
  END Data_PMOS[411]
  PIN Data_PMOS[410]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6459.945 187.44 6460.225 188.44 ;
    END
  END Data_PMOS[410]
  PIN Data_PMOS[409]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6487.105 187.44 6487.385 188.44 ;
    END
  END Data_PMOS[409]
  PIN Data_PMOS[408]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6488.225 187.44 6488.505 188.44 ;
    END
  END Data_PMOS[408]
  PIN Data_PMOS[407]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6513.705 187.44 6513.985 188.44 ;
    END
  END Data_PMOS[407]
  PIN Data_PMOS[406]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6509.785 187.44 6510.065 188.44 ;
    END
  END Data_PMOS[406]
  PIN Data_PMOS[405]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6500.825 187.44 6501.105 188.44 ;
    END
  END Data_PMOS[405]
  PIN Data_PMOS[404]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6512.025 187.44 6512.305 188.44 ;
    END
  END Data_PMOS[404]
  PIN Data_PMOS[403]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6461.065 187.44 6461.345 188.44 ;
    END
  END Data_PMOS[403]
  PIN Data_PMOS[402]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6489.345 187.44 6489.625 188.44 ;
    END
  END Data_PMOS[402]
  PIN Data_PMOS[401]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6488.785 187.44 6489.065 188.44 ;
    END
  END Data_PMOS[401]
  PIN Data_PMOS[400]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6459.385 187.44 6459.665 188.44 ;
    END
  END Data_PMOS[400]
  PIN Data_PMOS[399]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6458.825 187.44 6459.105 188.44 ;
    END
  END Data_PMOS[399]
  PIN Data_PMOS[398]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6432.505 187.44 6432.785 188.44 ;
    END
  END Data_PMOS[398]
  PIN Data_PMOS[397]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6434.185 187.44 6434.465 188.44 ;
    END
  END Data_PMOS[397]
  PIN Data_PMOS[396]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6448.745 187.44 6449.025 188.44 ;
    END
  END Data_PMOS[396]
  PIN Data_PMOS[395]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6377.065 187.44 6377.345 188.44 ;
    END
  END Data_PMOS[395]
  PIN Data_PMOS[394]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6379.305 187.44 6379.585 188.44 ;
    END
  END Data_PMOS[394]
  PIN Data_PMOS[393]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6380.985 187.44 6381.265 188.44 ;
    END
  END Data_PMOS[393]
  PIN Data_PMOS[392]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6431.945 187.44 6432.225 188.44 ;
    END
  END Data_PMOS[392]
  PIN Data_PMOS[391]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6433.065 187.44 6433.345 188.44 ;
    END
  END Data_PMOS[391]
  PIN Data_PMOS[390]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6434.745 187.44 6435.025 188.44 ;
    END
  END Data_PMOS[390]
  PIN Data_PMOS[389]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6378.745 187.44 6379.025 188.44 ;
    END
  END Data_PMOS[389]
  PIN Data_PMOS[388]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6380.425 187.44 6380.705 188.44 ;
    END
  END Data_PMOS[388]
  PIN Data_PMOS[387]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6381.545 187.44 6381.825 188.44 ;
    END
  END Data_PMOS[387]
  PIN Data_PMOS[386]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6448.185 187.44 6448.465 188.44 ;
    END
  END Data_PMOS[386]
  PIN Data_PMOS[385]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6431.385 187.44 6431.665 188.44 ;
    END
  END Data_PMOS[385]
  PIN Data_PMOS[384]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6430.825 187.44 6431.105 188.44 ;
    END
  END Data_PMOS[384]
  PIN Data_PMOS[383]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6433.625 187.44 6433.905 188.44 ;
    END
  END Data_PMOS[383]
  PIN Data_PMOS[382]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6379.865 187.44 6380.145 188.44 ;
    END
  END Data_PMOS[382]
  PIN Data_PMOS[381]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6382.665 187.44 6382.945 188.44 ;
    END
  END Data_PMOS[381]
  PIN Data_PMOS[380]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6382.105 187.44 6382.385 188.44 ;
    END
  END Data_PMOS[380]
  PIN Data_PMOS[379]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6378.185 187.44 6378.465 188.44 ;
    END
  END Data_PMOS[379]
  PIN Data_PMOS[378]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6377.625 187.44 6377.905 188.44 ;
    END
  END Data_PMOS[378]
  PIN Data_PMOS[377]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6355.785 187.44 6356.065 188.44 ;
    END
  END Data_PMOS[377]
  PIN Data_PMOS[376]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6357.465 187.44 6357.745 188.44 ;
    END
  END Data_PMOS[376]
  PIN Data_PMOS[375]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6359.145 187.44 6359.425 188.44 ;
    END
  END Data_PMOS[375]
  PIN Data_PMOS[374]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6311.545 187.44 6311.825 188.44 ;
    END
  END Data_PMOS[374]
  PIN Data_PMOS[373]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6313.785 187.44 6314.065 188.44 ;
    END
  END Data_PMOS[373]
  PIN Data_PMOS[372]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6315.465 187.44 6315.745 188.44 ;
    END
  END Data_PMOS[372]
  PIN Data_PMOS[371]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6355.225 187.44 6355.505 188.44 ;
    END
  END Data_PMOS[371]
  PIN Data_PMOS[370]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6356.345 187.44 6356.625 188.44 ;
    END
  END Data_PMOS[370]
  PIN Data_PMOS[369]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6358.025 187.44 6358.305 188.44 ;
    END
  END Data_PMOS[369]
  PIN Data_PMOS[368]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6313.225 187.44 6313.505 188.44 ;
    END
  END Data_PMOS[368]
  PIN Data_PMOS[367]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6314.905 187.44 6315.185 188.44 ;
    END
  END Data_PMOS[367]
  PIN Data_PMOS[366]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6316.025 187.44 6316.305 188.44 ;
    END
  END Data_PMOS[366]
  PIN Data_PMOS[365]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6358.585 187.44 6358.865 188.44 ;
    END
  END Data_PMOS[365]
  PIN Data_PMOS[364]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6354.665 187.44 6354.945 188.44 ;
    END
  END Data_PMOS[364]
  PIN Data_PMOS[363]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6354.105 187.44 6354.385 188.44 ;
    END
  END Data_PMOS[363]
  PIN Data_PMOS[362]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6356.905 187.44 6357.185 188.44 ;
    END
  END Data_PMOS[362]
  PIN Data_PMOS[361]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6314.345 187.44 6314.625 188.44 ;
    END
  END Data_PMOS[361]
  PIN Data_PMOS[360]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6317.145 187.44 6317.425 188.44 ;
    END
  END Data_PMOS[360]
  PIN Data_PMOS[359]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6316.585 187.44 6316.865 188.44 ;
    END
  END Data_PMOS[359]
  PIN Data_PMOS[358]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6312.665 187.44 6312.945 188.44 ;
    END
  END Data_PMOS[358]
  PIN Data_PMOS[357]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6312.105 187.44 6312.385 188.44 ;
    END
  END Data_PMOS[357]
  PIN Data_PMOS[356]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6285.785 187.44 6286.065 188.44 ;
    END
  END Data_PMOS[356]
  PIN Data_PMOS[355]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6287.465 187.44 6287.745 188.44 ;
    END
  END Data_PMOS[355]
  PIN Data_PMOS[354]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6289.145 187.44 6289.425 188.44 ;
    END
  END Data_PMOS[354]
  PIN Data_PMOS[353]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6229.785 187.44 6230.065 188.44 ;
    END
  END Data_PMOS[353]
  PIN Data_PMOS[352]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6232.025 187.44 6232.305 188.44 ;
    END
  END Data_PMOS[352]
  PIN Data_PMOS[351]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6233.705 187.44 6233.985 188.44 ;
    END
  END Data_PMOS[351]
  PIN Data_PMOS[350]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6285.225 187.44 6285.505 188.44 ;
    END
  END Data_PMOS[350]
  PIN Data_PMOS[349]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6286.345 187.44 6286.625 188.44 ;
    END
  END Data_PMOS[349]
  PIN Data_PMOS[348]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6288.025 187.44 6288.305 188.44 ;
    END
  END Data_PMOS[348]
  PIN Data_PMOS[347]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6231.465 187.44 6231.745 188.44 ;
    END
  END Data_PMOS[347]
  PIN Data_PMOS[346]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6233.145 187.44 6233.425 188.44 ;
    END
  END Data_PMOS[346]
  PIN Data_PMOS[345]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6234.265 187.44 6234.545 188.44 ;
    END
  END Data_PMOS[345]
  PIN Data_PMOS[344]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6288.585 187.44 6288.865 188.44 ;
    END
  END Data_PMOS[344]
  PIN Data_PMOS[343]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6284.665 187.44 6284.945 188.44 ;
    END
  END Data_PMOS[343]
  PIN Data_PMOS[342]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6284.105 187.44 6284.385 188.44 ;
    END
  END Data_PMOS[342]
  PIN Data_PMOS[341]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6286.905 187.44 6287.185 188.44 ;
    END
  END Data_PMOS[341]
  PIN Data_PMOS[340]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6232.585 187.44 6232.865 188.44 ;
    END
  END Data_PMOS[340]
  PIN Data_PMOS[339]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6235.385 187.44 6235.665 188.44 ;
    END
  END Data_PMOS[339]
  PIN Data_PMOS[338]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6234.825 187.44 6235.105 188.44 ;
    END
  END Data_PMOS[338]
  PIN Data_PMOS[337]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6230.905 187.44 6231.185 188.44 ;
    END
  END Data_PMOS[337]
  PIN Data_PMOS[336]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6230.345 187.44 6230.625 188.44 ;
    END
  END Data_PMOS[336]
  PIN Data_PMOS[335]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6181.065 187.44 6181.345 188.44 ;
    END
  END Data_PMOS[335]
  PIN Data_PMOS[334]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6208.225 187.44 6208.505 188.44 ;
    END
  END Data_PMOS[334]
  PIN Data_PMOS[333]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6209.905 187.44 6210.185 188.44 ;
    END
  END Data_PMOS[333]
  PIN Data_PMOS[332]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6151.385 187.44 6151.665 188.44 ;
    END
  END Data_PMOS[332]
  PIN Data_PMOS[331]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6153.625 187.44 6153.905 188.44 ;
    END
  END Data_PMOS[331]
  PIN Data_PMOS[330]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6155.305 187.44 6155.585 188.44 ;
    END
  END Data_PMOS[330]
  PIN Data_PMOS[329]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6180.505 187.44 6180.785 188.44 ;
    END
  END Data_PMOS[329]
  PIN Data_PMOS[328]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6181.625 187.44 6181.905 188.44 ;
    END
  END Data_PMOS[328]
  PIN Data_PMOS[327]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6208.785 187.44 6209.065 188.44 ;
    END
  END Data_PMOS[327]
  PIN Data_PMOS[326]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6153.065 187.44 6153.345 188.44 ;
    END
  END Data_PMOS[326]
  PIN Data_PMOS[325]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6154.745 187.44 6155.025 188.44 ;
    END
  END Data_PMOS[325]
  PIN Data_PMOS[324]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6168.745 187.44 6169.025 188.44 ;
    END
  END Data_PMOS[324]
  PIN Data_PMOS[323]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6209.345 187.44 6209.625 188.44 ;
    END
  END Data_PMOS[323]
  PIN Data_PMOS[322]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6179.945 187.44 6180.225 188.44 ;
    END
  END Data_PMOS[322]
  PIN Data_PMOS[321]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6179.385 187.44 6179.665 188.44 ;
    END
  END Data_PMOS[321]
  PIN Data_PMOS[320]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6207.665 187.44 6207.945 188.44 ;
    END
  END Data_PMOS[320]
  PIN Data_PMOS[319]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6154.185 187.44 6154.465 188.44 ;
    END
  END Data_PMOS[319]
  PIN Data_PMOS[318]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6169.865 187.44 6170.145 188.44 ;
    END
  END Data_PMOS[318]
  PIN Data_PMOS[317]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6169.305 187.44 6169.585 188.44 ;
    END
  END Data_PMOS[317]
  PIN Data_PMOS[316]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6152.505 187.44 6152.785 188.44 ;
    END
  END Data_PMOS[316]
  PIN Data_PMOS[315]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6151.945 187.44 6152.225 188.44 ;
    END
  END Data_PMOS[315]
  PIN Data_PMOS[314]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6098.745 187.44 6099.025 188.44 ;
    END
  END Data_PMOS[314]
  PIN Data_PMOS[313]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6100.425 187.44 6100.705 188.44 ;
    END
  END Data_PMOS[313]
  PIN Data_PMOS[312]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6102.105 187.44 6102.385 188.44 ;
    END
  END Data_PMOS[312]
  PIN Data_PMOS[311]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6073.545 187.44 6073.825 188.44 ;
    END
  END Data_PMOS[311]
  PIN Data_PMOS[310]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6075.785 187.44 6076.065 188.44 ;
    END
  END Data_PMOS[310]
  PIN Data_PMOS[309]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6077.465 187.44 6077.745 188.44 ;
    END
  END Data_PMOS[309]
  PIN Data_PMOS[308]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6098.185 187.44 6098.465 188.44 ;
    END
  END Data_PMOS[308]
  PIN Data_PMOS[307]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6099.305 187.44 6099.585 188.44 ;
    END
  END Data_PMOS[307]
  PIN Data_PMOS[306]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6100.985 187.44 6101.265 188.44 ;
    END
  END Data_PMOS[306]
  PIN Data_PMOS[305]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6075.225 187.44 6075.505 188.44 ;
    END
  END Data_PMOS[305]
  PIN Data_PMOS[304]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6076.905 187.44 6077.185 188.44 ;
    END
  END Data_PMOS[304]
  PIN Data_PMOS[303]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6078.025 187.44 6078.305 188.44 ;
    END
  END Data_PMOS[303]
  PIN Data_PMOS[302]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6101.545 187.44 6101.825 188.44 ;
    END
  END Data_PMOS[302]
  PIN Data_PMOS[301]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6097.625 187.44 6097.905 188.44 ;
    END
  END Data_PMOS[301]
  PIN Data_PMOS[300]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6097.065 187.44 6097.345 188.44 ;
    END
  END Data_PMOS[300]
  PIN Data_PMOS[299]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6099.865 187.44 6100.145 188.44 ;
    END
  END Data_PMOS[299]
  PIN Data_PMOS[298]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6076.345 187.44 6076.625 188.44 ;
    END
  END Data_PMOS[298]
  PIN Data_PMOS[297]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6079.145 187.44 6079.425 188.44 ;
    END
  END Data_PMOS[297]
  PIN Data_PMOS[296]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6078.585 187.44 6078.865 188.44 ;
    END
  END Data_PMOS[296]
  PIN Data_PMOS[295]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6074.665 187.44 6074.945 188.44 ;
    END
  END Data_PMOS[295]
  PIN Data_PMOS[294]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6074.105 187.44 6074.385 188.44 ;
    END
  END Data_PMOS[294]
  PIN Data_PMOS[293]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6032.665 187.44 6032.945 188.44 ;
    END
  END Data_PMOS[293]
  PIN Data_PMOS[292]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6034.345 187.44 6034.625 188.44 ;
    END
  END Data_PMOS[292]
  PIN Data_PMOS[291]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6036.025 187.44 6036.305 188.44 ;
    END
  END Data_PMOS[291]
  PIN Data_PMOS[290]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6002.425 187.44 6002.705 188.44 ;
    END
  END Data_PMOS[290]
  PIN Data_PMOS[289]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6004.665 187.44 6004.945 188.44 ;
    END
  END Data_PMOS[289]
  PIN Data_PMOS[288]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6006.345 187.44 6006.625 188.44 ;
    END
  END Data_PMOS[288]
  PIN Data_PMOS[287]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6032.105 187.44 6032.385 188.44 ;
    END
  END Data_PMOS[287]
  PIN Data_PMOS[286]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6033.225 187.44 6033.505 188.44 ;
    END
  END Data_PMOS[286]
  PIN Data_PMOS[285]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6034.905 187.44 6035.185 188.44 ;
    END
  END Data_PMOS[285]
  PIN Data_PMOS[284]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6004.105 187.44 6004.385 188.44 ;
    END
  END Data_PMOS[284]
  PIN Data_PMOS[283]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6005.785 187.44 6006.065 188.44 ;
    END
  END Data_PMOS[283]
  PIN Data_PMOS[282]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6006.905 187.44 6007.185 188.44 ;
    END
  END Data_PMOS[282]
  PIN Data_PMOS[281]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6035.465 187.44 6035.745 188.44 ;
    END
  END Data_PMOS[281]
  PIN Data_PMOS[280]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6031.545 187.44 6031.825 188.44 ;
    END
  END Data_PMOS[280]
  PIN Data_PMOS[279]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6030.985 187.44 6031.265 188.44 ;
    END
  END Data_PMOS[279]
  PIN Data_PMOS[278]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6033.785 187.44 6034.065 188.44 ;
    END
  END Data_PMOS[278]
  PIN Data_PMOS[277]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6005.225 187.44 6005.505 188.44 ;
    END
  END Data_PMOS[277]
  PIN Data_PMOS[276]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6008.025 187.44 6008.305 188.44 ;
    END
  END Data_PMOS[276]
  PIN Data_PMOS[275]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6007.465 187.44 6007.745 188.44 ;
    END
  END Data_PMOS[275]
  PIN Data_PMOS[274]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6003.545 187.44 6003.825 188.44 ;
    END
  END Data_PMOS[274]
  PIN Data_PMOS[273]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6002.985 187.44 6003.265 188.44 ;
    END
  END Data_PMOS[273]
  PIN Data_PMOS[272]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5950.905 187.44 5951.185 188.44 ;
    END
  END Data_PMOS[272]
  PIN Data_PMOS[271]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5952.585 187.44 5952.865 188.44 ;
    END
  END Data_PMOS[271]
  PIN Data_PMOS[270]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5954.265 187.44 5954.545 188.44 ;
    END
  END Data_PMOS[270]
  PIN Data_PMOS[269]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5898.265 187.44 5898.545 188.44 ;
    END
  END Data_PMOS[269]
  PIN Data_PMOS[268]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5900.505 187.44 5900.785 188.44 ;
    END
  END Data_PMOS[268]
  PIN Data_PMOS[267]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5927.665 187.44 5927.945 188.44 ;
    END
  END Data_PMOS[267]
  PIN Data_PMOS[266]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5950.345 187.44 5950.625 188.44 ;
    END
  END Data_PMOS[266]
  PIN Data_PMOS[265]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5951.465 187.44 5951.745 188.44 ;
    END
  END Data_PMOS[265]
  PIN Data_PMOS[264]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5953.145 187.44 5953.425 188.44 ;
    END
  END Data_PMOS[264]
  PIN Data_PMOS[263]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5899.945 187.44 5900.225 188.44 ;
    END
  END Data_PMOS[263]
  PIN Data_PMOS[262]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5927.105 187.44 5927.385 188.44 ;
    END
  END Data_PMOS[262]
  PIN Data_PMOS[261]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5928.225 187.44 5928.505 188.44 ;
    END
  END Data_PMOS[261]
  PIN Data_PMOS[260]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5953.705 187.44 5953.985 188.44 ;
    END
  END Data_PMOS[260]
  PIN Data_PMOS[259]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5949.785 187.44 5950.065 188.44 ;
    END
  END Data_PMOS[259]
  PIN Data_PMOS[258]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5940.825 187.44 5941.105 188.44 ;
    END
  END Data_PMOS[258]
  PIN Data_PMOS[257]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5952.025 187.44 5952.305 188.44 ;
    END
  END Data_PMOS[257]
  PIN Data_PMOS[256]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5901.065 187.44 5901.345 188.44 ;
    END
  END Data_PMOS[256]
  PIN Data_PMOS[255]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5929.345 187.44 5929.625 188.44 ;
    END
  END Data_PMOS[255]
  PIN Data_PMOS[254]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5928.785 187.44 5929.065 188.44 ;
    END
  END Data_PMOS[254]
  PIN Data_PMOS[253]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5899.385 187.44 5899.665 188.44 ;
    END
  END Data_PMOS[253]
  PIN Data_PMOS[252]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5898.825 187.44 5899.105 188.44 ;
    END
  END Data_PMOS[252]
  PIN Data_PMOS[251]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5872.505 187.44 5872.785 188.44 ;
    END
  END Data_PMOS[251]
  PIN Data_PMOS[250]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5874.185 187.44 5874.465 188.44 ;
    END
  END Data_PMOS[250]
  PIN Data_PMOS[249]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5888.745 187.44 5889.025 188.44 ;
    END
  END Data_PMOS[249]
  PIN Data_PMOS[248]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5817.065 187.44 5817.345 188.44 ;
    END
  END Data_PMOS[248]
  PIN Data_PMOS[247]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5819.305 187.44 5819.585 188.44 ;
    END
  END Data_PMOS[247]
  PIN Data_PMOS[246]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5820.985 187.44 5821.265 188.44 ;
    END
  END Data_PMOS[246]
  PIN Data_PMOS[245]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5871.945 187.44 5872.225 188.44 ;
    END
  END Data_PMOS[245]
  PIN Data_PMOS[244]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5873.065 187.44 5873.345 188.44 ;
    END
  END Data_PMOS[244]
  PIN Data_PMOS[243]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5874.745 187.44 5875.025 188.44 ;
    END
  END Data_PMOS[243]
  PIN Data_PMOS[242]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5818.745 187.44 5819.025 188.44 ;
    END
  END Data_PMOS[242]
  PIN Data_PMOS[241]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5820.425 187.44 5820.705 188.44 ;
    END
  END Data_PMOS[241]
  PIN Data_PMOS[240]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5821.545 187.44 5821.825 188.44 ;
    END
  END Data_PMOS[240]
  PIN Data_PMOS[239]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5888.185 187.44 5888.465 188.44 ;
    END
  END Data_PMOS[239]
  PIN Data_PMOS[238]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5871.385 187.44 5871.665 188.44 ;
    END
  END Data_PMOS[238]
  PIN Data_PMOS[237]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5870.825 187.44 5871.105 188.44 ;
    END
  END Data_PMOS[237]
  PIN Data_PMOS[236]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5873.625 187.44 5873.905 188.44 ;
    END
  END Data_PMOS[236]
  PIN Data_PMOS[235]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5819.865 187.44 5820.145 188.44 ;
    END
  END Data_PMOS[235]
  PIN Data_PMOS[234]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5822.665 187.44 5822.945 188.44 ;
    END
  END Data_PMOS[234]
  PIN Data_PMOS[233]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5822.105 187.44 5822.385 188.44 ;
    END
  END Data_PMOS[233]
  PIN Data_PMOS[232]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5818.185 187.44 5818.465 188.44 ;
    END
  END Data_PMOS[232]
  PIN Data_PMOS[231]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5817.625 187.44 5817.905 188.44 ;
    END
  END Data_PMOS[231]
  PIN Data_PMOS[230]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5795.785 187.44 5796.065 188.44 ;
    END
  END Data_PMOS[230]
  PIN Data_PMOS[229]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5797.465 187.44 5797.745 188.44 ;
    END
  END Data_PMOS[229]
  PIN Data_PMOS[228]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5799.145 187.44 5799.425 188.44 ;
    END
  END Data_PMOS[228]
  PIN Data_PMOS[227]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5751.545 187.44 5751.825 188.44 ;
    END
  END Data_PMOS[227]
  PIN Data_PMOS[226]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5753.785 187.44 5754.065 188.44 ;
    END
  END Data_PMOS[226]
  PIN Data_PMOS[225]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5755.465 187.44 5755.745 188.44 ;
    END
  END Data_PMOS[225]
  PIN Data_PMOS[224]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5795.225 187.44 5795.505 188.44 ;
    END
  END Data_PMOS[224]
  PIN Data_PMOS[223]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5796.345 187.44 5796.625 188.44 ;
    END
  END Data_PMOS[223]
  PIN Data_PMOS[222]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5798.025 187.44 5798.305 188.44 ;
    END
  END Data_PMOS[222]
  PIN Data_PMOS[221]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5753.225 187.44 5753.505 188.44 ;
    END
  END Data_PMOS[221]
  PIN Data_PMOS[220]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5754.905 187.44 5755.185 188.44 ;
    END
  END Data_PMOS[220]
  PIN Data_PMOS[219]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5756.025 187.44 5756.305 188.44 ;
    END
  END Data_PMOS[219]
  PIN Data_PMOS[218]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5798.585 187.44 5798.865 188.44 ;
    END
  END Data_PMOS[218]
  PIN Data_PMOS[217]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5794.665 187.44 5794.945 188.44 ;
    END
  END Data_PMOS[217]
  PIN Data_PMOS[216]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5794.105 187.44 5794.385 188.44 ;
    END
  END Data_PMOS[216]
  PIN Data_PMOS[215]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5796.905 187.44 5797.185 188.44 ;
    END
  END Data_PMOS[215]
  PIN Data_PMOS[214]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5754.345 187.44 5754.625 188.44 ;
    END
  END Data_PMOS[214]
  PIN Data_PMOS[213]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5757.145 187.44 5757.425 188.44 ;
    END
  END Data_PMOS[213]
  PIN Data_PMOS[212]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5756.585 187.44 5756.865 188.44 ;
    END
  END Data_PMOS[212]
  PIN Data_PMOS[211]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5752.665 187.44 5752.945 188.44 ;
    END
  END Data_PMOS[211]
  PIN Data_PMOS[210]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5752.105 187.44 5752.385 188.44 ;
    END
  END Data_PMOS[210]
  PIN Data_PMOS[209]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5725.785 187.44 5726.065 188.44 ;
    END
  END Data_PMOS[209]
  PIN Data_PMOS[208]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5727.465 187.44 5727.745 188.44 ;
    END
  END Data_PMOS[208]
  PIN Data_PMOS[207]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5729.145 187.44 5729.425 188.44 ;
    END
  END Data_PMOS[207]
  PIN Data_PMOS[206]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5669.785 187.44 5670.065 188.44 ;
    END
  END Data_PMOS[206]
  PIN Data_PMOS[205]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5672.025 187.44 5672.305 188.44 ;
    END
  END Data_PMOS[205]
  PIN Data_PMOS[204]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5673.705 187.44 5673.985 188.44 ;
    END
  END Data_PMOS[204]
  PIN Data_PMOS[203]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5725.225 187.44 5725.505 188.44 ;
    END
  END Data_PMOS[203]
  PIN Data_PMOS[202]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5726.345 187.44 5726.625 188.44 ;
    END
  END Data_PMOS[202]
  PIN Data_PMOS[201]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5728.025 187.44 5728.305 188.44 ;
    END
  END Data_PMOS[201]
  PIN Data_PMOS[200]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5671.465 187.44 5671.745 188.44 ;
    END
  END Data_PMOS[200]
  PIN Data_PMOS[199]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5673.145 187.44 5673.425 188.44 ;
    END
  END Data_PMOS[199]
  PIN Data_PMOS[198]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5674.265 187.44 5674.545 188.44 ;
    END
  END Data_PMOS[198]
  PIN Data_PMOS[197]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5728.585 187.44 5728.865 188.44 ;
    END
  END Data_PMOS[197]
  PIN Data_PMOS[196]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5724.665 187.44 5724.945 188.44 ;
    END
  END Data_PMOS[196]
  PIN Data_PMOS[195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5724.105 187.44 5724.385 188.44 ;
    END
  END Data_PMOS[195]
  PIN Data_PMOS[194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5726.905 187.44 5727.185 188.44 ;
    END
  END Data_PMOS[194]
  PIN Data_PMOS[193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5672.585 187.44 5672.865 188.44 ;
    END
  END Data_PMOS[193]
  PIN Data_PMOS[192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5675.385 187.44 5675.665 188.44 ;
    END
  END Data_PMOS[192]
  PIN Data_PMOS[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5674.825 187.44 5675.105 188.44 ;
    END
  END Data_PMOS[191]
  PIN Data_PMOS[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5670.905 187.44 5671.185 188.44 ;
    END
  END Data_PMOS[190]
  PIN Data_PMOS[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5670.345 187.44 5670.625 188.44 ;
    END
  END Data_PMOS[189]
  PIN Data_PMOS[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5621.065 187.44 5621.345 188.44 ;
    END
  END Data_PMOS[188]
  PIN Data_PMOS[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5648.225 187.44 5648.505 188.44 ;
    END
  END Data_PMOS[187]
  PIN Data_PMOS[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5649.905 187.44 5650.185 188.44 ;
    END
  END Data_PMOS[186]
  PIN Data_PMOS[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5591.385 187.44 5591.665 188.44 ;
    END
  END Data_PMOS[185]
  PIN Data_PMOS[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5593.625 187.44 5593.905 188.44 ;
    END
  END Data_PMOS[184]
  PIN Data_PMOS[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5595.305 187.44 5595.585 188.44 ;
    END
  END Data_PMOS[183]
  PIN Data_PMOS[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5620.505 187.44 5620.785 188.44 ;
    END
  END Data_PMOS[182]
  PIN Data_PMOS[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5621.625 187.44 5621.905 188.44 ;
    END
  END Data_PMOS[181]
  PIN Data_PMOS[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5648.785 187.44 5649.065 188.44 ;
    END
  END Data_PMOS[180]
  PIN Data_PMOS[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5593.065 187.44 5593.345 188.44 ;
    END
  END Data_PMOS[179]
  PIN Data_PMOS[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5594.745 187.44 5595.025 188.44 ;
    END
  END Data_PMOS[178]
  PIN Data_PMOS[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5608.745 187.44 5609.025 188.44 ;
    END
  END Data_PMOS[177]
  PIN Data_PMOS[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5649.345 187.44 5649.625 188.44 ;
    END
  END Data_PMOS[176]
  PIN Data_PMOS[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5619.945 187.44 5620.225 188.44 ;
    END
  END Data_PMOS[175]
  PIN Data_PMOS[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5619.385 187.44 5619.665 188.44 ;
    END
  END Data_PMOS[174]
  PIN Data_PMOS[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5647.665 187.44 5647.945 188.44 ;
    END
  END Data_PMOS[173]
  PIN Data_PMOS[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5594.185 187.44 5594.465 188.44 ;
    END
  END Data_PMOS[172]
  PIN Data_PMOS[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5609.865 187.44 5610.145 188.44 ;
    END
  END Data_PMOS[171]
  PIN Data_PMOS[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5609.305 187.44 5609.585 188.44 ;
    END
  END Data_PMOS[170]
  PIN Data_PMOS[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5592.505 187.44 5592.785 188.44 ;
    END
  END Data_PMOS[169]
  PIN Data_PMOS[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5591.945 187.44 5592.225 188.44 ;
    END
  END Data_PMOS[168]
  PIN Data_PMOS[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5538.745 187.44 5539.025 188.44 ;
    END
  END Data_PMOS[167]
  PIN Data_PMOS[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5540.425 187.44 5540.705 188.44 ;
    END
  END Data_PMOS[166]
  PIN Data_PMOS[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5542.105 187.44 5542.385 188.44 ;
    END
  END Data_PMOS[165]
  PIN Data_PMOS[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5513.545 187.44 5513.825 188.44 ;
    END
  END Data_PMOS[164]
  PIN Data_PMOS[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5515.785 187.44 5516.065 188.44 ;
    END
  END Data_PMOS[163]
  PIN Data_PMOS[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5517.465 187.44 5517.745 188.44 ;
    END
  END Data_PMOS[162]
  PIN Data_PMOS[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5538.185 187.44 5538.465 188.44 ;
    END
  END Data_PMOS[161]
  PIN Data_PMOS[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5539.305 187.44 5539.585 188.44 ;
    END
  END Data_PMOS[160]
  PIN Data_PMOS[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5540.985 187.44 5541.265 188.44 ;
    END
  END Data_PMOS[159]
  PIN Data_PMOS[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5515.225 187.44 5515.505 188.44 ;
    END
  END Data_PMOS[158]
  PIN Data_PMOS[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5516.905 187.44 5517.185 188.44 ;
    END
  END Data_PMOS[157]
  PIN Data_PMOS[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5518.025 187.44 5518.305 188.44 ;
    END
  END Data_PMOS[156]
  PIN Data_PMOS[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5541.545 187.44 5541.825 188.44 ;
    END
  END Data_PMOS[155]
  PIN Data_PMOS[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5537.625 187.44 5537.905 188.44 ;
    END
  END Data_PMOS[154]
  PIN Data_PMOS[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5537.065 187.44 5537.345 188.44 ;
    END
  END Data_PMOS[153]
  PIN Data_PMOS[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5539.865 187.44 5540.145 188.44 ;
    END
  END Data_PMOS[152]
  PIN Data_PMOS[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5516.345 187.44 5516.625 188.44 ;
    END
  END Data_PMOS[151]
  PIN Data_PMOS[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5519.145 187.44 5519.425 188.44 ;
    END
  END Data_PMOS[150]
  PIN Data_PMOS[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5518.585 187.44 5518.865 188.44 ;
    END
  END Data_PMOS[149]
  PIN Data_PMOS[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5514.665 187.44 5514.945 188.44 ;
    END
  END Data_PMOS[148]
  PIN Data_PMOS[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5514.105 187.44 5514.385 188.44 ;
    END
  END Data_PMOS[147]
  PIN Data_PMOS[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5472.665 187.44 5472.945 188.44 ;
    END
  END Data_PMOS[146]
  PIN Data_PMOS[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5474.345 187.44 5474.625 188.44 ;
    END
  END Data_PMOS[145]
  PIN Data_PMOS[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5476.025 187.44 5476.305 188.44 ;
    END
  END Data_PMOS[144]
  PIN Data_PMOS[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5442.425 187.44 5442.705 188.44 ;
    END
  END Data_PMOS[143]
  PIN Data_PMOS[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5444.665 187.44 5444.945 188.44 ;
    END
  END Data_PMOS[142]
  PIN Data_PMOS[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5446.345 187.44 5446.625 188.44 ;
    END
  END Data_PMOS[141]
  PIN Data_PMOS[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5472.105 187.44 5472.385 188.44 ;
    END
  END Data_PMOS[140]
  PIN Data_PMOS[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5473.225 187.44 5473.505 188.44 ;
    END
  END Data_PMOS[139]
  PIN Data_PMOS[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5474.905 187.44 5475.185 188.44 ;
    END
  END Data_PMOS[138]
  PIN Data_PMOS[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5444.105 187.44 5444.385 188.44 ;
    END
  END Data_PMOS[137]
  PIN Data_PMOS[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5445.785 187.44 5446.065 188.44 ;
    END
  END Data_PMOS[136]
  PIN Data_PMOS[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5446.905 187.44 5447.185 188.44 ;
    END
  END Data_PMOS[135]
  PIN Data_PMOS[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5475.465 187.44 5475.745 188.44 ;
    END
  END Data_PMOS[134]
  PIN Data_PMOS[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5471.545 187.44 5471.825 188.44 ;
    END
  END Data_PMOS[133]
  PIN Data_PMOS[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5470.985 187.44 5471.265 188.44 ;
    END
  END Data_PMOS[132]
  PIN Data_PMOS[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5473.785 187.44 5474.065 188.44 ;
    END
  END Data_PMOS[131]
  PIN Data_PMOS[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5445.225 187.44 5445.505 188.44 ;
    END
  END Data_PMOS[130]
  PIN Data_PMOS[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5448.025 187.44 5448.305 188.44 ;
    END
  END Data_PMOS[129]
  PIN Data_PMOS[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5447.465 187.44 5447.745 188.44 ;
    END
  END Data_PMOS[128]
  PIN Data_PMOS[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5443.545 187.44 5443.825 188.44 ;
    END
  END Data_PMOS[127]
  PIN Data_PMOS[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5442.985 187.44 5443.265 188.44 ;
    END
  END Data_PMOS[126]
  PIN Data_PMOS[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5390.905 187.44 5391.185 188.44 ;
    END
  END Data_PMOS[125]
  PIN Data_PMOS[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5392.585 187.44 5392.865 188.44 ;
    END
  END Data_PMOS[124]
  PIN Data_PMOS[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5394.265 187.44 5394.545 188.44 ;
    END
  END Data_PMOS[123]
  PIN Data_PMOS[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5338.265 187.44 5338.545 188.44 ;
    END
  END Data_PMOS[122]
  PIN Data_PMOS[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5340.505 187.44 5340.785 188.44 ;
    END
  END Data_PMOS[121]
  PIN Data_PMOS[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5367.665 187.44 5367.945 188.44 ;
    END
  END Data_PMOS[120]
  PIN Data_PMOS[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5390.345 187.44 5390.625 188.44 ;
    END
  END Data_PMOS[119]
  PIN Data_PMOS[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5391.465 187.44 5391.745 188.44 ;
    END
  END Data_PMOS[118]
  PIN Data_PMOS[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5393.145 187.44 5393.425 188.44 ;
    END
  END Data_PMOS[117]
  PIN Data_PMOS[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5339.945 187.44 5340.225 188.44 ;
    END
  END Data_PMOS[116]
  PIN Data_PMOS[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5367.105 187.44 5367.385 188.44 ;
    END
  END Data_PMOS[115]
  PIN Data_PMOS[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5368.225 187.44 5368.505 188.44 ;
    END
  END Data_PMOS[114]
  PIN Data_PMOS[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5393.705 187.44 5393.985 188.44 ;
    END
  END Data_PMOS[113]
  PIN Data_PMOS[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5389.785 187.44 5390.065 188.44 ;
    END
  END Data_PMOS[112]
  PIN Data_PMOS[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5380.825 187.44 5381.105 188.44 ;
    END
  END Data_PMOS[111]
  PIN Data_PMOS[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5392.025 187.44 5392.305 188.44 ;
    END
  END Data_PMOS[110]
  PIN Data_PMOS[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5341.065 187.44 5341.345 188.44 ;
    END
  END Data_PMOS[109]
  PIN Data_PMOS[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5369.345 187.44 5369.625 188.44 ;
    END
  END Data_PMOS[108]
  PIN Data_PMOS[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5368.785 187.44 5369.065 188.44 ;
    END
  END Data_PMOS[107]
  PIN Data_PMOS[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5339.385 187.44 5339.665 188.44 ;
    END
  END Data_PMOS[106]
  PIN Data_PMOS[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5338.825 187.44 5339.105 188.44 ;
    END
  END Data_PMOS[105]
  PIN Data_PMOS[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5312.505 187.44 5312.785 188.44 ;
    END
  END Data_PMOS[104]
  PIN Data_PMOS[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5314.185 187.44 5314.465 188.44 ;
    END
  END Data_PMOS[103]
  PIN Data_PMOS[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5328.745 187.44 5329.025 188.44 ;
    END
  END Data_PMOS[102]
  PIN Data_PMOS[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5257.065 187.44 5257.345 188.44 ;
    END
  END Data_PMOS[101]
  PIN Data_PMOS[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5259.305 187.44 5259.585 188.44 ;
    END
  END Data_PMOS[100]
  PIN Data_PMOS[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5260.985 187.44 5261.265 188.44 ;
    END
  END Data_PMOS[99]
  PIN Data_PMOS[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5311.945 187.44 5312.225 188.44 ;
    END
  END Data_PMOS[98]
  PIN Data_PMOS[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5313.065 187.44 5313.345 188.44 ;
    END
  END Data_PMOS[97]
  PIN Data_PMOS[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5314.745 187.44 5315.025 188.44 ;
    END
  END Data_PMOS[96]
  PIN Data_PMOS[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5258.745 187.44 5259.025 188.44 ;
    END
  END Data_PMOS[95]
  PIN Data_PMOS[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5260.425 187.44 5260.705 188.44 ;
    END
  END Data_PMOS[94]
  PIN Data_PMOS[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5261.545 187.44 5261.825 188.44 ;
    END
  END Data_PMOS[93]
  PIN Data_PMOS[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5328.185 187.44 5328.465 188.44 ;
    END
  END Data_PMOS[92]
  PIN Data_PMOS[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5311.385 187.44 5311.665 188.44 ;
    END
  END Data_PMOS[91]
  PIN Data_PMOS[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5310.825 187.44 5311.105 188.44 ;
    END
  END Data_PMOS[90]
  PIN Data_PMOS[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5313.625 187.44 5313.905 188.44 ;
    END
  END Data_PMOS[89]
  PIN Data_PMOS[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5259.865 187.44 5260.145 188.44 ;
    END
  END Data_PMOS[88]
  PIN Data_PMOS[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5262.665 187.44 5262.945 188.44 ;
    END
  END Data_PMOS[87]
  PIN Data_PMOS[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5262.105 187.44 5262.385 188.44 ;
    END
  END Data_PMOS[86]
  PIN Data_PMOS[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5258.185 187.44 5258.465 188.44 ;
    END
  END Data_PMOS[85]
  PIN Data_PMOS[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5257.625 187.44 5257.905 188.44 ;
    END
  END Data_PMOS[84]
  PIN Data_PMOS[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5235.785 187.44 5236.065 188.44 ;
    END
  END Data_PMOS[83]
  PIN Data_PMOS[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5237.465 187.44 5237.745 188.44 ;
    END
  END Data_PMOS[82]
  PIN Data_PMOS[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5239.145 187.44 5239.425 188.44 ;
    END
  END Data_PMOS[81]
  PIN Data_PMOS[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5191.545 187.44 5191.825 188.44 ;
    END
  END Data_PMOS[80]
  PIN Data_PMOS[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5193.785 187.44 5194.065 188.44 ;
    END
  END Data_PMOS[79]
  PIN Data_PMOS[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5195.465 187.44 5195.745 188.44 ;
    END
  END Data_PMOS[78]
  PIN Data_PMOS[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5235.225 187.44 5235.505 188.44 ;
    END
  END Data_PMOS[77]
  PIN Data_PMOS[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5236.345 187.44 5236.625 188.44 ;
    END
  END Data_PMOS[76]
  PIN Data_PMOS[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5238.025 187.44 5238.305 188.44 ;
    END
  END Data_PMOS[75]
  PIN Data_PMOS[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5193.225 187.44 5193.505 188.44 ;
    END
  END Data_PMOS[74]
  PIN Data_PMOS[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5194.905 187.44 5195.185 188.44 ;
    END
  END Data_PMOS[73]
  PIN Data_PMOS[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5196.025 187.44 5196.305 188.44 ;
    END
  END Data_PMOS[72]
  PIN Data_PMOS[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5238.585 187.44 5238.865 188.44 ;
    END
  END Data_PMOS[71]
  PIN Data_PMOS[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5234.665 187.44 5234.945 188.44 ;
    END
  END Data_PMOS[70]
  PIN Data_PMOS[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5234.105 187.44 5234.385 188.44 ;
    END
  END Data_PMOS[69]
  PIN Data_PMOS[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5236.905 187.44 5237.185 188.44 ;
    END
  END Data_PMOS[68]
  PIN Data_PMOS[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5194.345 187.44 5194.625 188.44 ;
    END
  END Data_PMOS[67]
  PIN Data_PMOS[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5197.145 187.44 5197.425 188.44 ;
    END
  END Data_PMOS[66]
  PIN Data_PMOS[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5196.585 187.44 5196.865 188.44 ;
    END
  END Data_PMOS[65]
  PIN Data_PMOS[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5192.665 187.44 5192.945 188.44 ;
    END
  END Data_PMOS[64]
  PIN Data_PMOS[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5192.105 187.44 5192.385 188.44 ;
    END
  END Data_PMOS[63]
  PIN Data_PMOS[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5165.785 187.44 5166.065 188.44 ;
    END
  END Data_PMOS[62]
  PIN Data_PMOS[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5167.465 187.44 5167.745 188.44 ;
    END
  END Data_PMOS[61]
  PIN Data_PMOS[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5169.145 187.44 5169.425 188.44 ;
    END
  END Data_PMOS[60]
  PIN Data_PMOS[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5109.785 187.44 5110.065 188.44 ;
    END
  END Data_PMOS[59]
  PIN Data_PMOS[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5112.025 187.44 5112.305 188.44 ;
    END
  END Data_PMOS[58]
  PIN Data_PMOS[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5113.705 187.44 5113.985 188.44 ;
    END
  END Data_PMOS[57]
  PIN Data_PMOS[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5165.225 187.44 5165.505 188.44 ;
    END
  END Data_PMOS[56]
  PIN Data_PMOS[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5166.345 187.44 5166.625 188.44 ;
    END
  END Data_PMOS[55]
  PIN Data_PMOS[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5168.025 187.44 5168.305 188.44 ;
    END
  END Data_PMOS[54]
  PIN Data_PMOS[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5111.465 187.44 5111.745 188.44 ;
    END
  END Data_PMOS[53]
  PIN Data_PMOS[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5113.145 187.44 5113.425 188.44 ;
    END
  END Data_PMOS[52]
  PIN Data_PMOS[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5114.265 187.44 5114.545 188.44 ;
    END
  END Data_PMOS[51]
  PIN Data_PMOS[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5168.585 187.44 5168.865 188.44 ;
    END
  END Data_PMOS[50]
  PIN Data_PMOS[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5164.665 187.44 5164.945 188.44 ;
    END
  END Data_PMOS[49]
  PIN Data_PMOS[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5164.105 187.44 5164.385 188.44 ;
    END
  END Data_PMOS[48]
  PIN Data_PMOS[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5166.905 187.44 5167.185 188.44 ;
    END
  END Data_PMOS[47]
  PIN Data_PMOS[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5112.585 187.44 5112.865 188.44 ;
    END
  END Data_PMOS[46]
  PIN Data_PMOS[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5115.385 187.44 5115.665 188.44 ;
    END
  END Data_PMOS[45]
  PIN Data_PMOS[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5114.825 187.44 5115.105 188.44 ;
    END
  END Data_PMOS[44]
  PIN Data_PMOS[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5110.905 187.44 5111.185 188.44 ;
    END
  END Data_PMOS[43]
  PIN Data_PMOS[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5110.345 187.44 5110.625 188.44 ;
    END
  END Data_PMOS[42]
  PIN Data_PMOS[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5061.065 187.44 5061.345 188.44 ;
    END
  END Data_PMOS[41]
  PIN Data_PMOS[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5088.225 187.44 5088.505 188.44 ;
    END
  END Data_PMOS[40]
  PIN Data_PMOS[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5089.905 187.44 5090.185 188.44 ;
    END
  END Data_PMOS[39]
  PIN Data_PMOS[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5031.385 187.44 5031.665 188.44 ;
    END
  END Data_PMOS[38]
  PIN Data_PMOS[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5033.625 187.44 5033.905 188.44 ;
    END
  END Data_PMOS[37]
  PIN Data_PMOS[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5035.305 187.44 5035.585 188.44 ;
    END
  END Data_PMOS[36]
  PIN Data_PMOS[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5060.505 187.44 5060.785 188.44 ;
    END
  END Data_PMOS[35]
  PIN Data_PMOS[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5061.625 187.44 5061.905 188.44 ;
    END
  END Data_PMOS[34]
  PIN Data_PMOS[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5088.785 187.44 5089.065 188.44 ;
    END
  END Data_PMOS[33]
  PIN Data_PMOS[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5033.065 187.44 5033.345 188.44 ;
    END
  END Data_PMOS[32]
  PIN Data_PMOS[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5034.745 187.44 5035.025 188.44 ;
    END
  END Data_PMOS[31]
  PIN Data_PMOS[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5048.745 187.44 5049.025 188.44 ;
    END
  END Data_PMOS[30]
  PIN Data_PMOS[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5089.345 187.44 5089.625 188.44 ;
    END
  END Data_PMOS[29]
  PIN Data_PMOS[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5059.945 187.44 5060.225 188.44 ;
    END
  END Data_PMOS[28]
  PIN Data_PMOS[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5059.385 187.44 5059.665 188.44 ;
    END
  END Data_PMOS[27]
  PIN Data_PMOS[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5087.665 187.44 5087.945 188.44 ;
    END
  END Data_PMOS[26]
  PIN Data_PMOS[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5034.185 187.44 5034.465 188.44 ;
    END
  END Data_PMOS[25]
  PIN Data_PMOS[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5049.865 187.44 5050.145 188.44 ;
    END
  END Data_PMOS[24]
  PIN Data_PMOS[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5049.305 187.44 5049.585 188.44 ;
    END
  END Data_PMOS[23]
  PIN Data_PMOS[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5032.505 187.44 5032.785 188.44 ;
    END
  END Data_PMOS[22]
  PIN Data_PMOS[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5031.945 187.44 5032.225 188.44 ;
    END
  END Data_PMOS[21]
  PIN Data_PMOS[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4978.745 187.44 4979.025 188.44 ;
    END
  END Data_PMOS[20]
  PIN Data_PMOS[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4980.425 187.44 4980.705 188.44 ;
    END
  END Data_PMOS[19]
  PIN Data_PMOS[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4982.105 187.44 4982.385 188.44 ;
    END
  END Data_PMOS[18]
  PIN Data_PMOS[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4953.545 187.44 4953.825 188.44 ;
    END
  END Data_PMOS[17]
  PIN Data_PMOS[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4955.785 187.44 4956.065 188.44 ;
    END
  END Data_PMOS[16]
  PIN Data_PMOS[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4957.465 187.44 4957.745 188.44 ;
    END
  END Data_PMOS[15]
  PIN Data_PMOS[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4978.185 187.44 4978.465 188.44 ;
    END
  END Data_PMOS[14]
  PIN Data_PMOS[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4979.305 187.44 4979.585 188.44 ;
    END
  END Data_PMOS[13]
  PIN Data_PMOS[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4980.985 187.44 4981.265 188.44 ;
    END
  END Data_PMOS[12]
  PIN Data_PMOS[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4955.225 187.44 4955.505 188.44 ;
    END
  END Data_PMOS[11]
  PIN Data_PMOS[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4956.905 187.44 4957.185 188.44 ;
    END
  END Data_PMOS[10]
  PIN Data_PMOS[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4958.025 187.44 4958.305 188.44 ;
    END
  END Data_PMOS[9]
  PIN Data_PMOS[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4981.545 187.44 4981.825 188.44 ;
    END
  END Data_PMOS[8]
  PIN Data_PMOS[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4977.625 187.44 4977.905 188.44 ;
    END
  END Data_PMOS[7]
  PIN Data_PMOS[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4977.065 187.44 4977.345 188.44 ;
    END
  END Data_PMOS[6]
  PIN Data_PMOS[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4979.865 187.44 4980.145 188.44 ;
    END
  END Data_PMOS[5]
  PIN Data_PMOS[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4956.345 187.44 4956.625 188.44 ;
    END
  END Data_PMOS[4]
  PIN Data_PMOS[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4959.145 187.44 4959.425 188.44 ;
    END
  END Data_PMOS[3]
  PIN Data_PMOS[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4958.585 187.44 4958.865 188.44 ;
    END
  END Data_PMOS[2]
  PIN Data_PMOS[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4954.665 187.44 4954.945 188.44 ;
    END
  END Data_PMOS[1]
  PIN Data_PMOS[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4954.105 187.44 4954.385 188.44 ;
    END
  END Data_PMOS[0]
  PIN Data_COMP[1175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13872.665 187.44 13872.945 188.44 ;
    END
  END Data_COMP[1175]
  PIN Data_COMP[1174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13874.345 187.44 13874.625 188.44 ;
    END
  END Data_COMP[1174]
  PIN Data_COMP[1173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13876.025 187.44 13876.305 188.44 ;
    END
  END Data_COMP[1173]
  PIN Data_COMP[1172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13842.425 187.44 13842.705 188.44 ;
    END
  END Data_COMP[1172]
  PIN Data_COMP[1171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13844.665 187.44 13844.945 188.44 ;
    END
  END Data_COMP[1171]
  PIN Data_COMP[1170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13846.345 187.44 13846.625 188.44 ;
    END
  END Data_COMP[1170]
  PIN Data_COMP[1169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13872.105 187.44 13872.385 188.44 ;
    END
  END Data_COMP[1169]
  PIN Data_COMP[1168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13873.225 187.44 13873.505 188.44 ;
    END
  END Data_COMP[1168]
  PIN Data_COMP[1167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13874.905 187.44 13875.185 188.44 ;
    END
  END Data_COMP[1167]
  PIN Data_COMP[1166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13844.105 187.44 13844.385 188.44 ;
    END
  END Data_COMP[1166]
  PIN Data_COMP[1165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13845.785 187.44 13846.065 188.44 ;
    END
  END Data_COMP[1165]
  PIN Data_COMP[1164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13846.905 187.44 13847.185 188.44 ;
    END
  END Data_COMP[1164]
  PIN Data_COMP[1163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13875.465 187.44 13875.745 188.44 ;
    END
  END Data_COMP[1163]
  PIN Data_COMP[1162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13871.545 187.44 13871.825 188.44 ;
    END
  END Data_COMP[1162]
  PIN Data_COMP[1161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13870.985 187.44 13871.265 188.44 ;
    END
  END Data_COMP[1161]
  PIN Data_COMP[1160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13873.785 187.44 13874.065 188.44 ;
    END
  END Data_COMP[1160]
  PIN Data_COMP[1159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13845.225 187.44 13845.505 188.44 ;
    END
  END Data_COMP[1159]
  PIN Data_COMP[1158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13848.025 187.44 13848.305 188.44 ;
    END
  END Data_COMP[1158]
  PIN Data_COMP[1157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13847.465 187.44 13847.745 188.44 ;
    END
  END Data_COMP[1157]
  PIN Data_COMP[1156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13843.545 187.44 13843.825 188.44 ;
    END
  END Data_COMP[1156]
  PIN Data_COMP[1155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13842.985 187.44 13843.265 188.44 ;
    END
  END Data_COMP[1155]
  PIN Data_COMP[1154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13790.905 187.44 13791.185 188.44 ;
    END
  END Data_COMP[1154]
  PIN Data_COMP[1153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13792.585 187.44 13792.865 188.44 ;
    END
  END Data_COMP[1153]
  PIN Data_COMP[1152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13794.265 187.44 13794.545 188.44 ;
    END
  END Data_COMP[1152]
  PIN Data_COMP[1151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13738.265 187.44 13738.545 188.44 ;
    END
  END Data_COMP[1151]
  PIN Data_COMP[1150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13740.505 187.44 13740.785 188.44 ;
    END
  END Data_COMP[1150]
  PIN Data_COMP[1149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13767.665 187.44 13767.945 188.44 ;
    END
  END Data_COMP[1149]
  PIN Data_COMP[1148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13790.345 187.44 13790.625 188.44 ;
    END
  END Data_COMP[1148]
  PIN Data_COMP[1147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13791.465 187.44 13791.745 188.44 ;
    END
  END Data_COMP[1147]
  PIN Data_COMP[1146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13793.145 187.44 13793.425 188.44 ;
    END
  END Data_COMP[1146]
  PIN Data_COMP[1145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13739.945 187.44 13740.225 188.44 ;
    END
  END Data_COMP[1145]
  PIN Data_COMP[1144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13767.105 187.44 13767.385 188.44 ;
    END
  END Data_COMP[1144]
  PIN Data_COMP[1143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13768.225 187.44 13768.505 188.44 ;
    END
  END Data_COMP[1143]
  PIN Data_COMP[1142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13793.705 187.44 13793.985 188.44 ;
    END
  END Data_COMP[1142]
  PIN Data_COMP[1141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13789.785 187.44 13790.065 188.44 ;
    END
  END Data_COMP[1141]
  PIN Data_COMP[1140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13780.825 187.44 13781.105 188.44 ;
    END
  END Data_COMP[1140]
  PIN Data_COMP[1139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13792.025 187.44 13792.305 188.44 ;
    END
  END Data_COMP[1139]
  PIN Data_COMP[1138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13741.065 187.44 13741.345 188.44 ;
    END
  END Data_COMP[1138]
  PIN Data_COMP[1137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13769.345 187.44 13769.625 188.44 ;
    END
  END Data_COMP[1137]
  PIN Data_COMP[1136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13768.785 187.44 13769.065 188.44 ;
    END
  END Data_COMP[1136]
  PIN Data_COMP[1135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13739.385 187.44 13739.665 188.44 ;
    END
  END Data_COMP[1135]
  PIN Data_COMP[1134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13738.825 187.44 13739.105 188.44 ;
    END
  END Data_COMP[1134]
  PIN Data_COMP[1133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13712.505 187.44 13712.785 188.44 ;
    END
  END Data_COMP[1133]
  PIN Data_COMP[1132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13714.185 187.44 13714.465 188.44 ;
    END
  END Data_COMP[1132]
  PIN Data_COMP[1131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13728.745 187.44 13729.025 188.44 ;
    END
  END Data_COMP[1131]
  PIN Data_COMP[1130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13657.065 187.44 13657.345 188.44 ;
    END
  END Data_COMP[1130]
  PIN Data_COMP[1129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13659.305 187.44 13659.585 188.44 ;
    END
  END Data_COMP[1129]
  PIN Data_COMP[1128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13660.985 187.44 13661.265 188.44 ;
    END
  END Data_COMP[1128]
  PIN Data_COMP[1127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13711.945 187.44 13712.225 188.44 ;
    END
  END Data_COMP[1127]
  PIN Data_COMP[1126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13713.065 187.44 13713.345 188.44 ;
    END
  END Data_COMP[1126]
  PIN Data_COMP[1125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13714.745 187.44 13715.025 188.44 ;
    END
  END Data_COMP[1125]
  PIN Data_COMP[1124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13658.745 187.44 13659.025 188.44 ;
    END
  END Data_COMP[1124]
  PIN Data_COMP[1123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13660.425 187.44 13660.705 188.44 ;
    END
  END Data_COMP[1123]
  PIN Data_COMP[1122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13661.545 187.44 13661.825 188.44 ;
    END
  END Data_COMP[1122]
  PIN Data_COMP[1121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13728.185 187.44 13728.465 188.44 ;
    END
  END Data_COMP[1121]
  PIN Data_COMP[1120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13711.385 187.44 13711.665 188.44 ;
    END
  END Data_COMP[1120]
  PIN Data_COMP[1119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13710.825 187.44 13711.105 188.44 ;
    END
  END Data_COMP[1119]
  PIN Data_COMP[1118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13713.625 187.44 13713.905 188.44 ;
    END
  END Data_COMP[1118]
  PIN Data_COMP[1117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13659.865 187.44 13660.145 188.44 ;
    END
  END Data_COMP[1117]
  PIN Data_COMP[1116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13662.665 187.44 13662.945 188.44 ;
    END
  END Data_COMP[1116]
  PIN Data_COMP[1115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13662.105 187.44 13662.385 188.44 ;
    END
  END Data_COMP[1115]
  PIN Data_COMP[1114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13658.185 187.44 13658.465 188.44 ;
    END
  END Data_COMP[1114]
  PIN Data_COMP[1113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13657.625 187.44 13657.905 188.44 ;
    END
  END Data_COMP[1113]
  PIN Data_COMP[1112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13635.785 187.44 13636.065 188.44 ;
    END
  END Data_COMP[1112]
  PIN Data_COMP[1111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13637.465 187.44 13637.745 188.44 ;
    END
  END Data_COMP[1111]
  PIN Data_COMP[1110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13639.145 187.44 13639.425 188.44 ;
    END
  END Data_COMP[1110]
  PIN Data_COMP[1109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13591.545 187.44 13591.825 188.44 ;
    END
  END Data_COMP[1109]
  PIN Data_COMP[1108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13593.785 187.44 13594.065 188.44 ;
    END
  END Data_COMP[1108]
  PIN Data_COMP[1107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13595.465 187.44 13595.745 188.44 ;
    END
  END Data_COMP[1107]
  PIN Data_COMP[1106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13635.225 187.44 13635.505 188.44 ;
    END
  END Data_COMP[1106]
  PIN Data_COMP[1105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13636.345 187.44 13636.625 188.44 ;
    END
  END Data_COMP[1105]
  PIN Data_COMP[1104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13638.025 187.44 13638.305 188.44 ;
    END
  END Data_COMP[1104]
  PIN Data_COMP[1103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13593.225 187.44 13593.505 188.44 ;
    END
  END Data_COMP[1103]
  PIN Data_COMP[1102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13594.905 187.44 13595.185 188.44 ;
    END
  END Data_COMP[1102]
  PIN Data_COMP[1101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13596.025 187.44 13596.305 188.44 ;
    END
  END Data_COMP[1101]
  PIN Data_COMP[1100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13638.585 187.44 13638.865 188.44 ;
    END
  END Data_COMP[1100]
  PIN Data_COMP[1099]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13634.665 187.44 13634.945 188.44 ;
    END
  END Data_COMP[1099]
  PIN Data_COMP[1098]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13634.105 187.44 13634.385 188.44 ;
    END
  END Data_COMP[1098]
  PIN Data_COMP[1097]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13636.905 187.44 13637.185 188.44 ;
    END
  END Data_COMP[1097]
  PIN Data_COMP[1096]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13594.345 187.44 13594.625 188.44 ;
    END
  END Data_COMP[1096]
  PIN Data_COMP[1095]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13597.145 187.44 13597.425 188.44 ;
    END
  END Data_COMP[1095]
  PIN Data_COMP[1094]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13596.585 187.44 13596.865 188.44 ;
    END
  END Data_COMP[1094]
  PIN Data_COMP[1093]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13592.665 187.44 13592.945 188.44 ;
    END
  END Data_COMP[1093]
  PIN Data_COMP[1092]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13592.105 187.44 13592.385 188.44 ;
    END
  END Data_COMP[1092]
  PIN Data_COMP[1091]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13565.785 187.44 13566.065 188.44 ;
    END
  END Data_COMP[1091]
  PIN Data_COMP[1090]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13567.465 187.44 13567.745 188.44 ;
    END
  END Data_COMP[1090]
  PIN Data_COMP[1089]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13569.145 187.44 13569.425 188.44 ;
    END
  END Data_COMP[1089]
  PIN Data_COMP[1088]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13509.785 187.44 13510.065 188.44 ;
    END
  END Data_COMP[1088]
  PIN Data_COMP[1087]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13512.025 187.44 13512.305 188.44 ;
    END
  END Data_COMP[1087]
  PIN Data_COMP[1086]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13513.705 187.44 13513.985 188.44 ;
    END
  END Data_COMP[1086]
  PIN Data_COMP[1085]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13565.225 187.44 13565.505 188.44 ;
    END
  END Data_COMP[1085]
  PIN Data_COMP[1084]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13566.345 187.44 13566.625 188.44 ;
    END
  END Data_COMP[1084]
  PIN Data_COMP[1083]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13568.025 187.44 13568.305 188.44 ;
    END
  END Data_COMP[1083]
  PIN Data_COMP[1082]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13511.465 187.44 13511.745 188.44 ;
    END
  END Data_COMP[1082]
  PIN Data_COMP[1081]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13513.145 187.44 13513.425 188.44 ;
    END
  END Data_COMP[1081]
  PIN Data_COMP[1080]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13514.265 187.44 13514.545 188.44 ;
    END
  END Data_COMP[1080]
  PIN Data_COMP[1079]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13568.585 187.44 13568.865 188.44 ;
    END
  END Data_COMP[1079]
  PIN Data_COMP[1078]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13564.665 187.44 13564.945 188.44 ;
    END
  END Data_COMP[1078]
  PIN Data_COMP[1077]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13564.105 187.44 13564.385 188.44 ;
    END
  END Data_COMP[1077]
  PIN Data_COMP[1076]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13566.905 187.44 13567.185 188.44 ;
    END
  END Data_COMP[1076]
  PIN Data_COMP[1075]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13512.585 187.44 13512.865 188.44 ;
    END
  END Data_COMP[1075]
  PIN Data_COMP[1074]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13515.385 187.44 13515.665 188.44 ;
    END
  END Data_COMP[1074]
  PIN Data_COMP[1073]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13514.825 187.44 13515.105 188.44 ;
    END
  END Data_COMP[1073]
  PIN Data_COMP[1072]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13510.905 187.44 13511.185 188.44 ;
    END
  END Data_COMP[1072]
  PIN Data_COMP[1071]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13510.345 187.44 13510.625 188.44 ;
    END
  END Data_COMP[1071]
  PIN Data_COMP[1070]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13461.065 187.44 13461.345 188.44 ;
    END
  END Data_COMP[1070]
  PIN Data_COMP[1069]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13488.225 187.44 13488.505 188.44 ;
    END
  END Data_COMP[1069]
  PIN Data_COMP[1068]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13489.905 187.44 13490.185 188.44 ;
    END
  END Data_COMP[1068]
  PIN Data_COMP[1067]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13431.385 187.44 13431.665 188.44 ;
    END
  END Data_COMP[1067]
  PIN Data_COMP[1066]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13433.625 187.44 13433.905 188.44 ;
    END
  END Data_COMP[1066]
  PIN Data_COMP[1065]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13435.305 187.44 13435.585 188.44 ;
    END
  END Data_COMP[1065]
  PIN Data_COMP[1064]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13460.505 187.44 13460.785 188.44 ;
    END
  END Data_COMP[1064]
  PIN Data_COMP[1063]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13461.625 187.44 13461.905 188.44 ;
    END
  END Data_COMP[1063]
  PIN Data_COMP[1062]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13488.785 187.44 13489.065 188.44 ;
    END
  END Data_COMP[1062]
  PIN Data_COMP[1061]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13433.065 187.44 13433.345 188.44 ;
    END
  END Data_COMP[1061]
  PIN Data_COMP[1060]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13434.745 187.44 13435.025 188.44 ;
    END
  END Data_COMP[1060]
  PIN Data_COMP[1059]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13448.745 187.44 13449.025 188.44 ;
    END
  END Data_COMP[1059]
  PIN Data_COMP[1058]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13489.345 187.44 13489.625 188.44 ;
    END
  END Data_COMP[1058]
  PIN Data_COMP[1057]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13459.945 187.44 13460.225 188.44 ;
    END
  END Data_COMP[1057]
  PIN Data_COMP[1056]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13459.385 187.44 13459.665 188.44 ;
    END
  END Data_COMP[1056]
  PIN Data_COMP[1055]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13487.665 187.44 13487.945 188.44 ;
    END
  END Data_COMP[1055]
  PIN Data_COMP[1054]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13434.185 187.44 13434.465 188.44 ;
    END
  END Data_COMP[1054]
  PIN Data_COMP[1053]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13449.865 187.44 13450.145 188.44 ;
    END
  END Data_COMP[1053]
  PIN Data_COMP[1052]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13449.305 187.44 13449.585 188.44 ;
    END
  END Data_COMP[1052]
  PIN Data_COMP[1051]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13432.505 187.44 13432.785 188.44 ;
    END
  END Data_COMP[1051]
  PIN Data_COMP[1050]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13431.945 187.44 13432.225 188.44 ;
    END
  END Data_COMP[1050]
  PIN Data_COMP[1049]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13378.745 187.44 13379.025 188.44 ;
    END
  END Data_COMP[1049]
  PIN Data_COMP[1048]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13380.425 187.44 13380.705 188.44 ;
    END
  END Data_COMP[1048]
  PIN Data_COMP[1047]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13382.105 187.44 13382.385 188.44 ;
    END
  END Data_COMP[1047]
  PIN Data_COMP[1046]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13353.545 187.44 13353.825 188.44 ;
    END
  END Data_COMP[1046]
  PIN Data_COMP[1045]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13355.785 187.44 13356.065 188.44 ;
    END
  END Data_COMP[1045]
  PIN Data_COMP[1044]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13357.465 187.44 13357.745 188.44 ;
    END
  END Data_COMP[1044]
  PIN Data_COMP[1043]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13378.185 187.44 13378.465 188.44 ;
    END
  END Data_COMP[1043]
  PIN Data_COMP[1042]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13379.305 187.44 13379.585 188.44 ;
    END
  END Data_COMP[1042]
  PIN Data_COMP[1041]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13380.985 187.44 13381.265 188.44 ;
    END
  END Data_COMP[1041]
  PIN Data_COMP[1040]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13355.225 187.44 13355.505 188.44 ;
    END
  END Data_COMP[1040]
  PIN Data_COMP[1039]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13356.905 187.44 13357.185 188.44 ;
    END
  END Data_COMP[1039]
  PIN Data_COMP[1038]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13358.025 187.44 13358.305 188.44 ;
    END
  END Data_COMP[1038]
  PIN Data_COMP[1037]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13381.545 187.44 13381.825 188.44 ;
    END
  END Data_COMP[1037]
  PIN Data_COMP[1036]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13377.625 187.44 13377.905 188.44 ;
    END
  END Data_COMP[1036]
  PIN Data_COMP[1035]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13377.065 187.44 13377.345 188.44 ;
    END
  END Data_COMP[1035]
  PIN Data_COMP[1034]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13379.865 187.44 13380.145 188.44 ;
    END
  END Data_COMP[1034]
  PIN Data_COMP[1033]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13356.345 187.44 13356.625 188.44 ;
    END
  END Data_COMP[1033]
  PIN Data_COMP[1032]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13359.145 187.44 13359.425 188.44 ;
    END
  END Data_COMP[1032]
  PIN Data_COMP[1031]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13358.585 187.44 13358.865 188.44 ;
    END
  END Data_COMP[1031]
  PIN Data_COMP[1030]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13354.665 187.44 13354.945 188.44 ;
    END
  END Data_COMP[1030]
  PIN Data_COMP[1029]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13354.105 187.44 13354.385 188.44 ;
    END
  END Data_COMP[1029]
  PIN Data_COMP[1028]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13312.665 187.44 13312.945 188.44 ;
    END
  END Data_COMP[1028]
  PIN Data_COMP[1027]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13314.345 187.44 13314.625 188.44 ;
    END
  END Data_COMP[1027]
  PIN Data_COMP[1026]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13316.025 187.44 13316.305 188.44 ;
    END
  END Data_COMP[1026]
  PIN Data_COMP[1025]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13282.425 187.44 13282.705 188.44 ;
    END
  END Data_COMP[1025]
  PIN Data_COMP[1024]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13284.665 187.44 13284.945 188.44 ;
    END
  END Data_COMP[1024]
  PIN Data_COMP[1023]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13286.345 187.44 13286.625 188.44 ;
    END
  END Data_COMP[1023]
  PIN Data_COMP[1022]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13312.105 187.44 13312.385 188.44 ;
    END
  END Data_COMP[1022]
  PIN Data_COMP[1021]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13313.225 187.44 13313.505 188.44 ;
    END
  END Data_COMP[1021]
  PIN Data_COMP[1020]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13314.905 187.44 13315.185 188.44 ;
    END
  END Data_COMP[1020]
  PIN Data_COMP[1019]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13284.105 187.44 13284.385 188.44 ;
    END
  END Data_COMP[1019]
  PIN Data_COMP[1018]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13285.785 187.44 13286.065 188.44 ;
    END
  END Data_COMP[1018]
  PIN Data_COMP[1017]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13286.905 187.44 13287.185 188.44 ;
    END
  END Data_COMP[1017]
  PIN Data_COMP[1016]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13315.465 187.44 13315.745 188.44 ;
    END
  END Data_COMP[1016]
  PIN Data_COMP[1015]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13311.545 187.44 13311.825 188.44 ;
    END
  END Data_COMP[1015]
  PIN Data_COMP[1014]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13310.985 187.44 13311.265 188.44 ;
    END
  END Data_COMP[1014]
  PIN Data_COMP[1013]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13313.785 187.44 13314.065 188.44 ;
    END
  END Data_COMP[1013]
  PIN Data_COMP[1012]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13285.225 187.44 13285.505 188.44 ;
    END
  END Data_COMP[1012]
  PIN Data_COMP[1011]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13288.025 187.44 13288.305 188.44 ;
    END
  END Data_COMP[1011]
  PIN Data_COMP[1010]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13287.465 187.44 13287.745 188.44 ;
    END
  END Data_COMP[1010]
  PIN Data_COMP[1009]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13283.545 187.44 13283.825 188.44 ;
    END
  END Data_COMP[1009]
  PIN Data_COMP[1008]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13282.985 187.44 13283.265 188.44 ;
    END
  END Data_COMP[1008]
  PIN Data_COMP[1007]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13230.905 187.44 13231.185 188.44 ;
    END
  END Data_COMP[1007]
  PIN Data_COMP[1006]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13232.585 187.44 13232.865 188.44 ;
    END
  END Data_COMP[1006]
  PIN Data_COMP[1005]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13234.265 187.44 13234.545 188.44 ;
    END
  END Data_COMP[1005]
  PIN Data_COMP[1004]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13178.265 187.44 13178.545 188.44 ;
    END
  END Data_COMP[1004]
  PIN Data_COMP[1003]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13180.505 187.44 13180.785 188.44 ;
    END
  END Data_COMP[1003]
  PIN Data_COMP[1002]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13207.665 187.44 13207.945 188.44 ;
    END
  END Data_COMP[1002]
  PIN Data_COMP[1001]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13230.345 187.44 13230.625 188.44 ;
    END
  END Data_COMP[1001]
  PIN Data_COMP[1000]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13231.465 187.44 13231.745 188.44 ;
    END
  END Data_COMP[1000]
  PIN Data_COMP[999]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13233.145 187.44 13233.425 188.44 ;
    END
  END Data_COMP[999]
  PIN Data_COMP[998]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13179.945 187.44 13180.225 188.44 ;
    END
  END Data_COMP[998]
  PIN Data_COMP[997]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13207.105 187.44 13207.385 188.44 ;
    END
  END Data_COMP[997]
  PIN Data_COMP[996]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13208.225 187.44 13208.505 188.44 ;
    END
  END Data_COMP[996]
  PIN Data_COMP[995]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13233.705 187.44 13233.985 188.44 ;
    END
  END Data_COMP[995]
  PIN Data_COMP[994]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13229.785 187.44 13230.065 188.44 ;
    END
  END Data_COMP[994]
  PIN Data_COMP[993]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13220.825 187.44 13221.105 188.44 ;
    END
  END Data_COMP[993]
  PIN Data_COMP[992]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13232.025 187.44 13232.305 188.44 ;
    END
  END Data_COMP[992]
  PIN Data_COMP[991]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13181.065 187.44 13181.345 188.44 ;
    END
  END Data_COMP[991]
  PIN Data_COMP[990]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13209.345 187.44 13209.625 188.44 ;
    END
  END Data_COMP[990]
  PIN Data_COMP[989]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13208.785 187.44 13209.065 188.44 ;
    END
  END Data_COMP[989]
  PIN Data_COMP[988]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13179.385 187.44 13179.665 188.44 ;
    END
  END Data_COMP[988]
  PIN Data_COMP[987]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13178.825 187.44 13179.105 188.44 ;
    END
  END Data_COMP[987]
  PIN Data_COMP[986]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13152.505 187.44 13152.785 188.44 ;
    END
  END Data_COMP[986]
  PIN Data_COMP[985]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13154.185 187.44 13154.465 188.44 ;
    END
  END Data_COMP[985]
  PIN Data_COMP[984]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13168.745 187.44 13169.025 188.44 ;
    END
  END Data_COMP[984]
  PIN Data_COMP[983]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13097.065 187.44 13097.345 188.44 ;
    END
  END Data_COMP[983]
  PIN Data_COMP[982]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13099.305 187.44 13099.585 188.44 ;
    END
  END Data_COMP[982]
  PIN Data_COMP[981]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13100.985 187.44 13101.265 188.44 ;
    END
  END Data_COMP[981]
  PIN Data_COMP[980]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13151.945 187.44 13152.225 188.44 ;
    END
  END Data_COMP[980]
  PIN Data_COMP[979]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13153.065 187.44 13153.345 188.44 ;
    END
  END Data_COMP[979]
  PIN Data_COMP[978]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13154.745 187.44 13155.025 188.44 ;
    END
  END Data_COMP[978]
  PIN Data_COMP[977]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13098.745 187.44 13099.025 188.44 ;
    END
  END Data_COMP[977]
  PIN Data_COMP[976]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13100.425 187.44 13100.705 188.44 ;
    END
  END Data_COMP[976]
  PIN Data_COMP[975]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13101.545 187.44 13101.825 188.44 ;
    END
  END Data_COMP[975]
  PIN Data_COMP[974]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13168.185 187.44 13168.465 188.44 ;
    END
  END Data_COMP[974]
  PIN Data_COMP[973]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13151.385 187.44 13151.665 188.44 ;
    END
  END Data_COMP[973]
  PIN Data_COMP[972]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13150.825 187.44 13151.105 188.44 ;
    END
  END Data_COMP[972]
  PIN Data_COMP[971]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13153.625 187.44 13153.905 188.44 ;
    END
  END Data_COMP[971]
  PIN Data_COMP[970]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13099.865 187.44 13100.145 188.44 ;
    END
  END Data_COMP[970]
  PIN Data_COMP[969]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13102.665 187.44 13102.945 188.44 ;
    END
  END Data_COMP[969]
  PIN Data_COMP[968]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13102.105 187.44 13102.385 188.44 ;
    END
  END Data_COMP[968]
  PIN Data_COMP[967]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13098.185 187.44 13098.465 188.44 ;
    END
  END Data_COMP[967]
  PIN Data_COMP[966]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13097.625 187.44 13097.905 188.44 ;
    END
  END Data_COMP[966]
  PIN Data_COMP[965]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13075.785 187.44 13076.065 188.44 ;
    END
  END Data_COMP[965]
  PIN Data_COMP[964]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13077.465 187.44 13077.745 188.44 ;
    END
  END Data_COMP[964]
  PIN Data_COMP[963]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13079.145 187.44 13079.425 188.44 ;
    END
  END Data_COMP[963]
  PIN Data_COMP[962]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13031.545 187.44 13031.825 188.44 ;
    END
  END Data_COMP[962]
  PIN Data_COMP[961]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13033.785 187.44 13034.065 188.44 ;
    END
  END Data_COMP[961]
  PIN Data_COMP[960]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13035.465 187.44 13035.745 188.44 ;
    END
  END Data_COMP[960]
  PIN Data_COMP[959]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13075.225 187.44 13075.505 188.44 ;
    END
  END Data_COMP[959]
  PIN Data_COMP[958]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13076.345 187.44 13076.625 188.44 ;
    END
  END Data_COMP[958]
  PIN Data_COMP[957]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13078.025 187.44 13078.305 188.44 ;
    END
  END Data_COMP[957]
  PIN Data_COMP[956]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13033.225 187.44 13033.505 188.44 ;
    END
  END Data_COMP[956]
  PIN Data_COMP[955]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13034.905 187.44 13035.185 188.44 ;
    END
  END Data_COMP[955]
  PIN Data_COMP[954]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13036.025 187.44 13036.305 188.44 ;
    END
  END Data_COMP[954]
  PIN Data_COMP[953]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13078.585 187.44 13078.865 188.44 ;
    END
  END Data_COMP[953]
  PIN Data_COMP[952]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13074.665 187.44 13074.945 188.44 ;
    END
  END Data_COMP[952]
  PIN Data_COMP[951]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13074.105 187.44 13074.385 188.44 ;
    END
  END Data_COMP[951]
  PIN Data_COMP[950]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13076.905 187.44 13077.185 188.44 ;
    END
  END Data_COMP[950]
  PIN Data_COMP[949]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13034.345 187.44 13034.625 188.44 ;
    END
  END Data_COMP[949]
  PIN Data_COMP[948]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13037.145 187.44 13037.425 188.44 ;
    END
  END Data_COMP[948]
  PIN Data_COMP[947]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13036.585 187.44 13036.865 188.44 ;
    END
  END Data_COMP[947]
  PIN Data_COMP[946]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13032.665 187.44 13032.945 188.44 ;
    END
  END Data_COMP[946]
  PIN Data_COMP[945]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13032.105 187.44 13032.385 188.44 ;
    END
  END Data_COMP[945]
  PIN Data_COMP[944]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13005.785 187.44 13006.065 188.44 ;
    END
  END Data_COMP[944]
  PIN Data_COMP[943]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13007.465 187.44 13007.745 188.44 ;
    END
  END Data_COMP[943]
  PIN Data_COMP[942]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13009.145 187.44 13009.425 188.44 ;
    END
  END Data_COMP[942]
  PIN Data_COMP[941]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12949.785 187.44 12950.065 188.44 ;
    END
  END Data_COMP[941]
  PIN Data_COMP[940]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12952.025 187.44 12952.305 188.44 ;
    END
  END Data_COMP[940]
  PIN Data_COMP[939]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12953.705 187.44 12953.985 188.44 ;
    END
  END Data_COMP[939]
  PIN Data_COMP[938]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13005.225 187.44 13005.505 188.44 ;
    END
  END Data_COMP[938]
  PIN Data_COMP[937]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13006.345 187.44 13006.625 188.44 ;
    END
  END Data_COMP[937]
  PIN Data_COMP[936]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13008.025 187.44 13008.305 188.44 ;
    END
  END Data_COMP[936]
  PIN Data_COMP[935]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12951.465 187.44 12951.745 188.44 ;
    END
  END Data_COMP[935]
  PIN Data_COMP[934]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12953.145 187.44 12953.425 188.44 ;
    END
  END Data_COMP[934]
  PIN Data_COMP[933]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12954.265 187.44 12954.545 188.44 ;
    END
  END Data_COMP[933]
  PIN Data_COMP[932]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13008.585 187.44 13008.865 188.44 ;
    END
  END Data_COMP[932]
  PIN Data_COMP[931]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13004.665 187.44 13004.945 188.44 ;
    END
  END Data_COMP[931]
  PIN Data_COMP[930]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13004.105 187.44 13004.385 188.44 ;
    END
  END Data_COMP[930]
  PIN Data_COMP[929]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13006.905 187.44 13007.185 188.44 ;
    END
  END Data_COMP[929]
  PIN Data_COMP[928]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12952.585 187.44 12952.865 188.44 ;
    END
  END Data_COMP[928]
  PIN Data_COMP[927]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12955.385 187.44 12955.665 188.44 ;
    END
  END Data_COMP[927]
  PIN Data_COMP[926]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12954.825 187.44 12955.105 188.44 ;
    END
  END Data_COMP[926]
  PIN Data_COMP[925]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12950.905 187.44 12951.185 188.44 ;
    END
  END Data_COMP[925]
  PIN Data_COMP[924]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12950.345 187.44 12950.625 188.44 ;
    END
  END Data_COMP[924]
  PIN Data_COMP[923]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12901.065 187.44 12901.345 188.44 ;
    END
  END Data_COMP[923]
  PIN Data_COMP[922]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12928.225 187.44 12928.505 188.44 ;
    END
  END Data_COMP[922]
  PIN Data_COMP[921]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12929.905 187.44 12930.185 188.44 ;
    END
  END Data_COMP[921]
  PIN Data_COMP[920]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12871.385 187.44 12871.665 188.44 ;
    END
  END Data_COMP[920]
  PIN Data_COMP[919]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12873.625 187.44 12873.905 188.44 ;
    END
  END Data_COMP[919]
  PIN Data_COMP[918]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12875.305 187.44 12875.585 188.44 ;
    END
  END Data_COMP[918]
  PIN Data_COMP[917]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12900.505 187.44 12900.785 188.44 ;
    END
  END Data_COMP[917]
  PIN Data_COMP[916]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12901.625 187.44 12901.905 188.44 ;
    END
  END Data_COMP[916]
  PIN Data_COMP[915]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12928.785 187.44 12929.065 188.44 ;
    END
  END Data_COMP[915]
  PIN Data_COMP[914]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12873.065 187.44 12873.345 188.44 ;
    END
  END Data_COMP[914]
  PIN Data_COMP[913]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12874.745 187.44 12875.025 188.44 ;
    END
  END Data_COMP[913]
  PIN Data_COMP[912]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12888.745 187.44 12889.025 188.44 ;
    END
  END Data_COMP[912]
  PIN Data_COMP[911]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12929.345 187.44 12929.625 188.44 ;
    END
  END Data_COMP[911]
  PIN Data_COMP[910]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12899.945 187.44 12900.225 188.44 ;
    END
  END Data_COMP[910]
  PIN Data_COMP[909]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12899.385 187.44 12899.665 188.44 ;
    END
  END Data_COMP[909]
  PIN Data_COMP[908]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12927.665 187.44 12927.945 188.44 ;
    END
  END Data_COMP[908]
  PIN Data_COMP[907]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12874.185 187.44 12874.465 188.44 ;
    END
  END Data_COMP[907]
  PIN Data_COMP[906]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12889.865 187.44 12890.145 188.44 ;
    END
  END Data_COMP[906]
  PIN Data_COMP[905]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12889.305 187.44 12889.585 188.44 ;
    END
  END Data_COMP[905]
  PIN Data_COMP[904]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12872.505 187.44 12872.785 188.44 ;
    END
  END Data_COMP[904]
  PIN Data_COMP[903]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12871.945 187.44 12872.225 188.44 ;
    END
  END Data_COMP[903]
  PIN Data_COMP[902]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12818.745 187.44 12819.025 188.44 ;
    END
  END Data_COMP[902]
  PIN Data_COMP[901]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12820.425 187.44 12820.705 188.44 ;
    END
  END Data_COMP[901]
  PIN Data_COMP[900]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12822.105 187.44 12822.385 188.44 ;
    END
  END Data_COMP[900]
  PIN Data_COMP[899]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12793.545 187.44 12793.825 188.44 ;
    END
  END Data_COMP[899]
  PIN Data_COMP[898]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12795.785 187.44 12796.065 188.44 ;
    END
  END Data_COMP[898]
  PIN Data_COMP[897]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12797.465 187.44 12797.745 188.44 ;
    END
  END Data_COMP[897]
  PIN Data_COMP[896]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12818.185 187.44 12818.465 188.44 ;
    END
  END Data_COMP[896]
  PIN Data_COMP[895]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12819.305 187.44 12819.585 188.44 ;
    END
  END Data_COMP[895]
  PIN Data_COMP[894]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12820.985 187.44 12821.265 188.44 ;
    END
  END Data_COMP[894]
  PIN Data_COMP[893]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12795.225 187.44 12795.505 188.44 ;
    END
  END Data_COMP[893]
  PIN Data_COMP[892]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12796.905 187.44 12797.185 188.44 ;
    END
  END Data_COMP[892]
  PIN Data_COMP[891]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12798.025 187.44 12798.305 188.44 ;
    END
  END Data_COMP[891]
  PIN Data_COMP[890]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12821.545 187.44 12821.825 188.44 ;
    END
  END Data_COMP[890]
  PIN Data_COMP[889]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12817.625 187.44 12817.905 188.44 ;
    END
  END Data_COMP[889]
  PIN Data_COMP[888]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12817.065 187.44 12817.345 188.44 ;
    END
  END Data_COMP[888]
  PIN Data_COMP[887]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12819.865 187.44 12820.145 188.44 ;
    END
  END Data_COMP[887]
  PIN Data_COMP[886]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12796.345 187.44 12796.625 188.44 ;
    END
  END Data_COMP[886]
  PIN Data_COMP[885]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12799.145 187.44 12799.425 188.44 ;
    END
  END Data_COMP[885]
  PIN Data_COMP[884]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12798.585 187.44 12798.865 188.44 ;
    END
  END Data_COMP[884]
  PIN Data_COMP[883]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12794.665 187.44 12794.945 188.44 ;
    END
  END Data_COMP[883]
  PIN Data_COMP[882]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12794.105 187.44 12794.385 188.44 ;
    END
  END Data_COMP[882]
  PIN Data_COMP[881]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12752.665 187.44 12752.945 188.44 ;
    END
  END Data_COMP[881]
  PIN Data_COMP[880]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12754.345 187.44 12754.625 188.44 ;
    END
  END Data_COMP[880]
  PIN Data_COMP[879]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12756.025 187.44 12756.305 188.44 ;
    END
  END Data_COMP[879]
  PIN Data_COMP[878]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12722.425 187.44 12722.705 188.44 ;
    END
  END Data_COMP[878]
  PIN Data_COMP[877]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12724.665 187.44 12724.945 188.44 ;
    END
  END Data_COMP[877]
  PIN Data_COMP[876]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12726.345 187.44 12726.625 188.44 ;
    END
  END Data_COMP[876]
  PIN Data_COMP[875]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12752.105 187.44 12752.385 188.44 ;
    END
  END Data_COMP[875]
  PIN Data_COMP[874]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12753.225 187.44 12753.505 188.44 ;
    END
  END Data_COMP[874]
  PIN Data_COMP[873]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12754.905 187.44 12755.185 188.44 ;
    END
  END Data_COMP[873]
  PIN Data_COMP[872]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12724.105 187.44 12724.385 188.44 ;
    END
  END Data_COMP[872]
  PIN Data_COMP[871]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12725.785 187.44 12726.065 188.44 ;
    END
  END Data_COMP[871]
  PIN Data_COMP[870]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12726.905 187.44 12727.185 188.44 ;
    END
  END Data_COMP[870]
  PIN Data_COMP[869]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12755.465 187.44 12755.745 188.44 ;
    END
  END Data_COMP[869]
  PIN Data_COMP[868]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12751.545 187.44 12751.825 188.44 ;
    END
  END Data_COMP[868]
  PIN Data_COMP[867]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12750.985 187.44 12751.265 188.44 ;
    END
  END Data_COMP[867]
  PIN Data_COMP[866]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12753.785 187.44 12754.065 188.44 ;
    END
  END Data_COMP[866]
  PIN Data_COMP[865]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12725.225 187.44 12725.505 188.44 ;
    END
  END Data_COMP[865]
  PIN Data_COMP[864]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12728.025 187.44 12728.305 188.44 ;
    END
  END Data_COMP[864]
  PIN Data_COMP[863]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12727.465 187.44 12727.745 188.44 ;
    END
  END Data_COMP[863]
  PIN Data_COMP[862]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12723.545 187.44 12723.825 188.44 ;
    END
  END Data_COMP[862]
  PIN Data_COMP[861]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12722.985 187.44 12723.265 188.44 ;
    END
  END Data_COMP[861]
  PIN Data_COMP[860]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12670.905 187.44 12671.185 188.44 ;
    END
  END Data_COMP[860]
  PIN Data_COMP[859]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12672.585 187.44 12672.865 188.44 ;
    END
  END Data_COMP[859]
  PIN Data_COMP[858]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12674.265 187.44 12674.545 188.44 ;
    END
  END Data_COMP[858]
  PIN Data_COMP[857]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12618.265 187.44 12618.545 188.44 ;
    END
  END Data_COMP[857]
  PIN Data_COMP[856]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12620.505 187.44 12620.785 188.44 ;
    END
  END Data_COMP[856]
  PIN Data_COMP[855]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12647.665 187.44 12647.945 188.44 ;
    END
  END Data_COMP[855]
  PIN Data_COMP[854]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12670.345 187.44 12670.625 188.44 ;
    END
  END Data_COMP[854]
  PIN Data_COMP[853]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12671.465 187.44 12671.745 188.44 ;
    END
  END Data_COMP[853]
  PIN Data_COMP[852]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12673.145 187.44 12673.425 188.44 ;
    END
  END Data_COMP[852]
  PIN Data_COMP[851]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12619.945 187.44 12620.225 188.44 ;
    END
  END Data_COMP[851]
  PIN Data_COMP[850]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12647.105 187.44 12647.385 188.44 ;
    END
  END Data_COMP[850]
  PIN Data_COMP[849]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12648.225 187.44 12648.505 188.44 ;
    END
  END Data_COMP[849]
  PIN Data_COMP[848]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12673.705 187.44 12673.985 188.44 ;
    END
  END Data_COMP[848]
  PIN Data_COMP[847]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12669.785 187.44 12670.065 188.44 ;
    END
  END Data_COMP[847]
  PIN Data_COMP[846]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12660.825 187.44 12661.105 188.44 ;
    END
  END Data_COMP[846]
  PIN Data_COMP[845]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12672.025 187.44 12672.305 188.44 ;
    END
  END Data_COMP[845]
  PIN Data_COMP[844]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12621.065 187.44 12621.345 188.44 ;
    END
  END Data_COMP[844]
  PIN Data_COMP[843]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12649.345 187.44 12649.625 188.44 ;
    END
  END Data_COMP[843]
  PIN Data_COMP[842]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12648.785 187.44 12649.065 188.44 ;
    END
  END Data_COMP[842]
  PIN Data_COMP[841]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12619.385 187.44 12619.665 188.44 ;
    END
  END Data_COMP[841]
  PIN Data_COMP[840]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12618.825 187.44 12619.105 188.44 ;
    END
  END Data_COMP[840]
  PIN Data_COMP[839]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12592.505 187.44 12592.785 188.44 ;
    END
  END Data_COMP[839]
  PIN Data_COMP[838]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12594.185 187.44 12594.465 188.44 ;
    END
  END Data_COMP[838]
  PIN Data_COMP[837]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12608.745 187.44 12609.025 188.44 ;
    END
  END Data_COMP[837]
  PIN Data_COMP[836]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12537.065 187.44 12537.345 188.44 ;
    END
  END Data_COMP[836]
  PIN Data_COMP[835]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12539.305 187.44 12539.585 188.44 ;
    END
  END Data_COMP[835]
  PIN Data_COMP[834]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12540.985 187.44 12541.265 188.44 ;
    END
  END Data_COMP[834]
  PIN Data_COMP[833]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12591.945 187.44 12592.225 188.44 ;
    END
  END Data_COMP[833]
  PIN Data_COMP[832]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12593.065 187.44 12593.345 188.44 ;
    END
  END Data_COMP[832]
  PIN Data_COMP[831]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12594.745 187.44 12595.025 188.44 ;
    END
  END Data_COMP[831]
  PIN Data_COMP[830]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12538.745 187.44 12539.025 188.44 ;
    END
  END Data_COMP[830]
  PIN Data_COMP[829]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12540.425 187.44 12540.705 188.44 ;
    END
  END Data_COMP[829]
  PIN Data_COMP[828]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12541.545 187.44 12541.825 188.44 ;
    END
  END Data_COMP[828]
  PIN Data_COMP[827]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12608.185 187.44 12608.465 188.44 ;
    END
  END Data_COMP[827]
  PIN Data_COMP[826]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12591.385 187.44 12591.665 188.44 ;
    END
  END Data_COMP[826]
  PIN Data_COMP[825]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12590.825 187.44 12591.105 188.44 ;
    END
  END Data_COMP[825]
  PIN Data_COMP[824]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12593.625 187.44 12593.905 188.44 ;
    END
  END Data_COMP[824]
  PIN Data_COMP[823]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12539.865 187.44 12540.145 188.44 ;
    END
  END Data_COMP[823]
  PIN Data_COMP[822]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12542.665 187.44 12542.945 188.44 ;
    END
  END Data_COMP[822]
  PIN Data_COMP[821]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12542.105 187.44 12542.385 188.44 ;
    END
  END Data_COMP[821]
  PIN Data_COMP[820]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12538.185 187.44 12538.465 188.44 ;
    END
  END Data_COMP[820]
  PIN Data_COMP[819]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12537.625 187.44 12537.905 188.44 ;
    END
  END Data_COMP[819]
  PIN Data_COMP[818]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12515.785 187.44 12516.065 188.44 ;
    END
  END Data_COMP[818]
  PIN Data_COMP[817]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12517.465 187.44 12517.745 188.44 ;
    END
  END Data_COMP[817]
  PIN Data_COMP[816]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12519.145 187.44 12519.425 188.44 ;
    END
  END Data_COMP[816]
  PIN Data_COMP[815]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12471.545 187.44 12471.825 188.44 ;
    END
  END Data_COMP[815]
  PIN Data_COMP[814]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12473.785 187.44 12474.065 188.44 ;
    END
  END Data_COMP[814]
  PIN Data_COMP[813]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12475.465 187.44 12475.745 188.44 ;
    END
  END Data_COMP[813]
  PIN Data_COMP[812]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12515.225 187.44 12515.505 188.44 ;
    END
  END Data_COMP[812]
  PIN Data_COMP[811]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12516.345 187.44 12516.625 188.44 ;
    END
  END Data_COMP[811]
  PIN Data_COMP[810]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12518.025 187.44 12518.305 188.44 ;
    END
  END Data_COMP[810]
  PIN Data_COMP[809]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12473.225 187.44 12473.505 188.44 ;
    END
  END Data_COMP[809]
  PIN Data_COMP[808]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12474.905 187.44 12475.185 188.44 ;
    END
  END Data_COMP[808]
  PIN Data_COMP[807]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12476.025 187.44 12476.305 188.44 ;
    END
  END Data_COMP[807]
  PIN Data_COMP[806]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12518.585 187.44 12518.865 188.44 ;
    END
  END Data_COMP[806]
  PIN Data_COMP[805]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12514.665 187.44 12514.945 188.44 ;
    END
  END Data_COMP[805]
  PIN Data_COMP[804]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12514.105 187.44 12514.385 188.44 ;
    END
  END Data_COMP[804]
  PIN Data_COMP[803]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12516.905 187.44 12517.185 188.44 ;
    END
  END Data_COMP[803]
  PIN Data_COMP[802]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12474.345 187.44 12474.625 188.44 ;
    END
  END Data_COMP[802]
  PIN Data_COMP[801]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12477.145 187.44 12477.425 188.44 ;
    END
  END Data_COMP[801]
  PIN Data_COMP[800]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12476.585 187.44 12476.865 188.44 ;
    END
  END Data_COMP[800]
  PIN Data_COMP[799]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12472.665 187.44 12472.945 188.44 ;
    END
  END Data_COMP[799]
  PIN Data_COMP[798]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12472.105 187.44 12472.385 188.44 ;
    END
  END Data_COMP[798]
  PIN Data_COMP[797]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12445.785 187.44 12446.065 188.44 ;
    END
  END Data_COMP[797]
  PIN Data_COMP[796]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12447.465 187.44 12447.745 188.44 ;
    END
  END Data_COMP[796]
  PIN Data_COMP[795]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12449.145 187.44 12449.425 188.44 ;
    END
  END Data_COMP[795]
  PIN Data_COMP[794]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12389.785 187.44 12390.065 188.44 ;
    END
  END Data_COMP[794]
  PIN Data_COMP[793]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12392.025 187.44 12392.305 188.44 ;
    END
  END Data_COMP[793]
  PIN Data_COMP[792]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12393.705 187.44 12393.985 188.44 ;
    END
  END Data_COMP[792]
  PIN Data_COMP[791]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12445.225 187.44 12445.505 188.44 ;
    END
  END Data_COMP[791]
  PIN Data_COMP[790]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12446.345 187.44 12446.625 188.44 ;
    END
  END Data_COMP[790]
  PIN Data_COMP[789]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12448.025 187.44 12448.305 188.44 ;
    END
  END Data_COMP[789]
  PIN Data_COMP[788]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12391.465 187.44 12391.745 188.44 ;
    END
  END Data_COMP[788]
  PIN Data_COMP[787]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12393.145 187.44 12393.425 188.44 ;
    END
  END Data_COMP[787]
  PIN Data_COMP[786]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12394.265 187.44 12394.545 188.44 ;
    END
  END Data_COMP[786]
  PIN Data_COMP[785]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12448.585 187.44 12448.865 188.44 ;
    END
  END Data_COMP[785]
  PIN Data_COMP[784]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12444.665 187.44 12444.945 188.44 ;
    END
  END Data_COMP[784]
  PIN Data_COMP[783]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12444.105 187.44 12444.385 188.44 ;
    END
  END Data_COMP[783]
  PIN Data_COMP[782]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12446.905 187.44 12447.185 188.44 ;
    END
  END Data_COMP[782]
  PIN Data_COMP[781]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12392.585 187.44 12392.865 188.44 ;
    END
  END Data_COMP[781]
  PIN Data_COMP[780]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12395.385 187.44 12395.665 188.44 ;
    END
  END Data_COMP[780]
  PIN Data_COMP[779]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12394.825 187.44 12395.105 188.44 ;
    END
  END Data_COMP[779]
  PIN Data_COMP[778]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12390.905 187.44 12391.185 188.44 ;
    END
  END Data_COMP[778]
  PIN Data_COMP[777]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12390.345 187.44 12390.625 188.44 ;
    END
  END Data_COMP[777]
  PIN Data_COMP[776]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12341.065 187.44 12341.345 188.44 ;
    END
  END Data_COMP[776]
  PIN Data_COMP[775]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12368.225 187.44 12368.505 188.44 ;
    END
  END Data_COMP[775]
  PIN Data_COMP[774]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12369.905 187.44 12370.185 188.44 ;
    END
  END Data_COMP[774]
  PIN Data_COMP[773]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12311.385 187.44 12311.665 188.44 ;
    END
  END Data_COMP[773]
  PIN Data_COMP[772]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12313.625 187.44 12313.905 188.44 ;
    END
  END Data_COMP[772]
  PIN Data_COMP[771]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12315.305 187.44 12315.585 188.44 ;
    END
  END Data_COMP[771]
  PIN Data_COMP[770]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12340.505 187.44 12340.785 188.44 ;
    END
  END Data_COMP[770]
  PIN Data_COMP[769]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12341.625 187.44 12341.905 188.44 ;
    END
  END Data_COMP[769]
  PIN Data_COMP[768]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12368.785 187.44 12369.065 188.44 ;
    END
  END Data_COMP[768]
  PIN Data_COMP[767]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12313.065 187.44 12313.345 188.44 ;
    END
  END Data_COMP[767]
  PIN Data_COMP[766]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12314.745 187.44 12315.025 188.44 ;
    END
  END Data_COMP[766]
  PIN Data_COMP[765]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12328.745 187.44 12329.025 188.44 ;
    END
  END Data_COMP[765]
  PIN Data_COMP[764]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12369.345 187.44 12369.625 188.44 ;
    END
  END Data_COMP[764]
  PIN Data_COMP[763]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12339.945 187.44 12340.225 188.44 ;
    END
  END Data_COMP[763]
  PIN Data_COMP[762]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12339.385 187.44 12339.665 188.44 ;
    END
  END Data_COMP[762]
  PIN Data_COMP[761]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12367.665 187.44 12367.945 188.44 ;
    END
  END Data_COMP[761]
  PIN Data_COMP[760]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12314.185 187.44 12314.465 188.44 ;
    END
  END Data_COMP[760]
  PIN Data_COMP[759]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12329.865 187.44 12330.145 188.44 ;
    END
  END Data_COMP[759]
  PIN Data_COMP[758]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12329.305 187.44 12329.585 188.44 ;
    END
  END Data_COMP[758]
  PIN Data_COMP[757]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12312.505 187.44 12312.785 188.44 ;
    END
  END Data_COMP[757]
  PIN Data_COMP[756]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12311.945 187.44 12312.225 188.44 ;
    END
  END Data_COMP[756]
  PIN Data_COMP[755]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12258.745 187.44 12259.025 188.44 ;
    END
  END Data_COMP[755]
  PIN Data_COMP[754]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12260.425 187.44 12260.705 188.44 ;
    END
  END Data_COMP[754]
  PIN Data_COMP[753]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12262.105 187.44 12262.385 188.44 ;
    END
  END Data_COMP[753]
  PIN Data_COMP[752]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12233.545 187.44 12233.825 188.44 ;
    END
  END Data_COMP[752]
  PIN Data_COMP[751]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12235.785 187.44 12236.065 188.44 ;
    END
  END Data_COMP[751]
  PIN Data_COMP[750]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12237.465 187.44 12237.745 188.44 ;
    END
  END Data_COMP[750]
  PIN Data_COMP[749]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12258.185 187.44 12258.465 188.44 ;
    END
  END Data_COMP[749]
  PIN Data_COMP[748]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12259.305 187.44 12259.585 188.44 ;
    END
  END Data_COMP[748]
  PIN Data_COMP[747]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12260.985 187.44 12261.265 188.44 ;
    END
  END Data_COMP[747]
  PIN Data_COMP[746]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12235.225 187.44 12235.505 188.44 ;
    END
  END Data_COMP[746]
  PIN Data_COMP[745]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12236.905 187.44 12237.185 188.44 ;
    END
  END Data_COMP[745]
  PIN Data_COMP[744]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12238.025 187.44 12238.305 188.44 ;
    END
  END Data_COMP[744]
  PIN Data_COMP[743]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12261.545 187.44 12261.825 188.44 ;
    END
  END Data_COMP[743]
  PIN Data_COMP[742]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12257.625 187.44 12257.905 188.44 ;
    END
  END Data_COMP[742]
  PIN Data_COMP[741]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12257.065 187.44 12257.345 188.44 ;
    END
  END Data_COMP[741]
  PIN Data_COMP[740]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12259.865 187.44 12260.145 188.44 ;
    END
  END Data_COMP[740]
  PIN Data_COMP[739]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12236.345 187.44 12236.625 188.44 ;
    END
  END Data_COMP[739]
  PIN Data_COMP[738]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12239.145 187.44 12239.425 188.44 ;
    END
  END Data_COMP[738]
  PIN Data_COMP[737]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12238.585 187.44 12238.865 188.44 ;
    END
  END Data_COMP[737]
  PIN Data_COMP[736]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12234.665 187.44 12234.945 188.44 ;
    END
  END Data_COMP[736]
  PIN Data_COMP[735]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12234.105 187.44 12234.385 188.44 ;
    END
  END Data_COMP[735]
  PIN Data_COMP[734]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12192.665 187.44 12192.945 188.44 ;
    END
  END Data_COMP[734]
  PIN Data_COMP[733]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12194.345 187.44 12194.625 188.44 ;
    END
  END Data_COMP[733]
  PIN Data_COMP[732]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12196.025 187.44 12196.305 188.44 ;
    END
  END Data_COMP[732]
  PIN Data_COMP[731]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12162.425 187.44 12162.705 188.44 ;
    END
  END Data_COMP[731]
  PIN Data_COMP[730]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12164.665 187.44 12164.945 188.44 ;
    END
  END Data_COMP[730]
  PIN Data_COMP[729]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12166.345 187.44 12166.625 188.44 ;
    END
  END Data_COMP[729]
  PIN Data_COMP[728]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12192.105 187.44 12192.385 188.44 ;
    END
  END Data_COMP[728]
  PIN Data_COMP[727]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12193.225 187.44 12193.505 188.44 ;
    END
  END Data_COMP[727]
  PIN Data_COMP[726]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12194.905 187.44 12195.185 188.44 ;
    END
  END Data_COMP[726]
  PIN Data_COMP[725]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12164.105 187.44 12164.385 188.44 ;
    END
  END Data_COMP[725]
  PIN Data_COMP[724]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12165.785 187.44 12166.065 188.44 ;
    END
  END Data_COMP[724]
  PIN Data_COMP[723]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12166.905 187.44 12167.185 188.44 ;
    END
  END Data_COMP[723]
  PIN Data_COMP[722]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12195.465 187.44 12195.745 188.44 ;
    END
  END Data_COMP[722]
  PIN Data_COMP[721]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12191.545 187.44 12191.825 188.44 ;
    END
  END Data_COMP[721]
  PIN Data_COMP[720]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12190.985 187.44 12191.265 188.44 ;
    END
  END Data_COMP[720]
  PIN Data_COMP[719]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12193.785 187.44 12194.065 188.44 ;
    END
  END Data_COMP[719]
  PIN Data_COMP[718]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12165.225 187.44 12165.505 188.44 ;
    END
  END Data_COMP[718]
  PIN Data_COMP[717]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12168.025 187.44 12168.305 188.44 ;
    END
  END Data_COMP[717]
  PIN Data_COMP[716]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12167.465 187.44 12167.745 188.44 ;
    END
  END Data_COMP[716]
  PIN Data_COMP[715]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12163.545 187.44 12163.825 188.44 ;
    END
  END Data_COMP[715]
  PIN Data_COMP[714]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12162.985 187.44 12163.265 188.44 ;
    END
  END Data_COMP[714]
  PIN Data_COMP[713]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12110.905 187.44 12111.185 188.44 ;
    END
  END Data_COMP[713]
  PIN Data_COMP[712]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12112.585 187.44 12112.865 188.44 ;
    END
  END Data_COMP[712]
  PIN Data_COMP[711]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12114.265 187.44 12114.545 188.44 ;
    END
  END Data_COMP[711]
  PIN Data_COMP[710]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12058.265 187.44 12058.545 188.44 ;
    END
  END Data_COMP[710]
  PIN Data_COMP[709]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12060.505 187.44 12060.785 188.44 ;
    END
  END Data_COMP[709]
  PIN Data_COMP[708]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12087.665 187.44 12087.945 188.44 ;
    END
  END Data_COMP[708]
  PIN Data_COMP[707]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12110.345 187.44 12110.625 188.44 ;
    END
  END Data_COMP[707]
  PIN Data_COMP[706]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12111.465 187.44 12111.745 188.44 ;
    END
  END Data_COMP[706]
  PIN Data_COMP[705]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12113.145 187.44 12113.425 188.44 ;
    END
  END Data_COMP[705]
  PIN Data_COMP[704]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12059.945 187.44 12060.225 188.44 ;
    END
  END Data_COMP[704]
  PIN Data_COMP[703]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12087.105 187.44 12087.385 188.44 ;
    END
  END Data_COMP[703]
  PIN Data_COMP[702]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12088.225 187.44 12088.505 188.44 ;
    END
  END Data_COMP[702]
  PIN Data_COMP[701]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12113.705 187.44 12113.985 188.44 ;
    END
  END Data_COMP[701]
  PIN Data_COMP[700]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12109.785 187.44 12110.065 188.44 ;
    END
  END Data_COMP[700]
  PIN Data_COMP[699]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12100.825 187.44 12101.105 188.44 ;
    END
  END Data_COMP[699]
  PIN Data_COMP[698]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12112.025 187.44 12112.305 188.44 ;
    END
  END Data_COMP[698]
  PIN Data_COMP[697]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12061.065 187.44 12061.345 188.44 ;
    END
  END Data_COMP[697]
  PIN Data_COMP[696]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12089.345 187.44 12089.625 188.44 ;
    END
  END Data_COMP[696]
  PIN Data_COMP[695]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12088.785 187.44 12089.065 188.44 ;
    END
  END Data_COMP[695]
  PIN Data_COMP[694]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12059.385 187.44 12059.665 188.44 ;
    END
  END Data_COMP[694]
  PIN Data_COMP[693]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12058.825 187.44 12059.105 188.44 ;
    END
  END Data_COMP[693]
  PIN Data_COMP[692]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12032.505 187.44 12032.785 188.44 ;
    END
  END Data_COMP[692]
  PIN Data_COMP[691]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12034.185 187.44 12034.465 188.44 ;
    END
  END Data_COMP[691]
  PIN Data_COMP[690]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12048.745 187.44 12049.025 188.44 ;
    END
  END Data_COMP[690]
  PIN Data_COMP[689]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11977.065 187.44 11977.345 188.44 ;
    END
  END Data_COMP[689]
  PIN Data_COMP[688]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11979.305 187.44 11979.585 188.44 ;
    END
  END Data_COMP[688]
  PIN Data_COMP[687]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11980.985 187.44 11981.265 188.44 ;
    END
  END Data_COMP[687]
  PIN Data_COMP[686]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12031.945 187.44 12032.225 188.44 ;
    END
  END Data_COMP[686]
  PIN Data_COMP[685]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12033.065 187.44 12033.345 188.44 ;
    END
  END Data_COMP[685]
  PIN Data_COMP[684]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12034.745 187.44 12035.025 188.44 ;
    END
  END Data_COMP[684]
  PIN Data_COMP[683]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11978.745 187.44 11979.025 188.44 ;
    END
  END Data_COMP[683]
  PIN Data_COMP[682]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11980.425 187.44 11980.705 188.44 ;
    END
  END Data_COMP[682]
  PIN Data_COMP[681]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11981.545 187.44 11981.825 188.44 ;
    END
  END Data_COMP[681]
  PIN Data_COMP[680]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12048.185 187.44 12048.465 188.44 ;
    END
  END Data_COMP[680]
  PIN Data_COMP[679]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12031.385 187.44 12031.665 188.44 ;
    END
  END Data_COMP[679]
  PIN Data_COMP[678]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12030.825 187.44 12031.105 188.44 ;
    END
  END Data_COMP[678]
  PIN Data_COMP[677]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12033.625 187.44 12033.905 188.44 ;
    END
  END Data_COMP[677]
  PIN Data_COMP[676]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11979.865 187.44 11980.145 188.44 ;
    END
  END Data_COMP[676]
  PIN Data_COMP[675]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11982.665 187.44 11982.945 188.44 ;
    END
  END Data_COMP[675]
  PIN Data_COMP[674]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11982.105 187.44 11982.385 188.44 ;
    END
  END Data_COMP[674]
  PIN Data_COMP[673]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11978.185 187.44 11978.465 188.44 ;
    END
  END Data_COMP[673]
  PIN Data_COMP[672]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11977.625 187.44 11977.905 188.44 ;
    END
  END Data_COMP[672]
  PIN Data_COMP[671]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11955.785 187.44 11956.065 188.44 ;
    END
  END Data_COMP[671]
  PIN Data_COMP[670]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11957.465 187.44 11957.745 188.44 ;
    END
  END Data_COMP[670]
  PIN Data_COMP[669]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11959.145 187.44 11959.425 188.44 ;
    END
  END Data_COMP[669]
  PIN Data_COMP[668]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11911.545 187.44 11911.825 188.44 ;
    END
  END Data_COMP[668]
  PIN Data_COMP[667]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11913.785 187.44 11914.065 188.44 ;
    END
  END Data_COMP[667]
  PIN Data_COMP[666]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11915.465 187.44 11915.745 188.44 ;
    END
  END Data_COMP[666]
  PIN Data_COMP[665]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11955.225 187.44 11955.505 188.44 ;
    END
  END Data_COMP[665]
  PIN Data_COMP[664]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11956.345 187.44 11956.625 188.44 ;
    END
  END Data_COMP[664]
  PIN Data_COMP[663]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11958.025 187.44 11958.305 188.44 ;
    END
  END Data_COMP[663]
  PIN Data_COMP[662]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11913.225 187.44 11913.505 188.44 ;
    END
  END Data_COMP[662]
  PIN Data_COMP[661]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11914.905 187.44 11915.185 188.44 ;
    END
  END Data_COMP[661]
  PIN Data_COMP[660]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11916.025 187.44 11916.305 188.44 ;
    END
  END Data_COMP[660]
  PIN Data_COMP[659]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11958.585 187.44 11958.865 188.44 ;
    END
  END Data_COMP[659]
  PIN Data_COMP[658]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11954.665 187.44 11954.945 188.44 ;
    END
  END Data_COMP[658]
  PIN Data_COMP[657]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11954.105 187.44 11954.385 188.44 ;
    END
  END Data_COMP[657]
  PIN Data_COMP[656]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11956.905 187.44 11957.185 188.44 ;
    END
  END Data_COMP[656]
  PIN Data_COMP[655]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11914.345 187.44 11914.625 188.44 ;
    END
  END Data_COMP[655]
  PIN Data_COMP[654]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11917.145 187.44 11917.425 188.44 ;
    END
  END Data_COMP[654]
  PIN Data_COMP[653]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11916.585 187.44 11916.865 188.44 ;
    END
  END Data_COMP[653]
  PIN Data_COMP[652]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11912.665 187.44 11912.945 188.44 ;
    END
  END Data_COMP[652]
  PIN Data_COMP[651]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11912.105 187.44 11912.385 188.44 ;
    END
  END Data_COMP[651]
  PIN Data_COMP[650]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11885.785 187.44 11886.065 188.44 ;
    END
  END Data_COMP[650]
  PIN Data_COMP[649]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11887.465 187.44 11887.745 188.44 ;
    END
  END Data_COMP[649]
  PIN Data_COMP[648]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11889.145 187.44 11889.425 188.44 ;
    END
  END Data_COMP[648]
  PIN Data_COMP[647]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11829.785 187.44 11830.065 188.44 ;
    END
  END Data_COMP[647]
  PIN Data_COMP[646]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11832.025 187.44 11832.305 188.44 ;
    END
  END Data_COMP[646]
  PIN Data_COMP[645]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11833.705 187.44 11833.985 188.44 ;
    END
  END Data_COMP[645]
  PIN Data_COMP[644]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11885.225 187.44 11885.505 188.44 ;
    END
  END Data_COMP[644]
  PIN Data_COMP[643]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11886.345 187.44 11886.625 188.44 ;
    END
  END Data_COMP[643]
  PIN Data_COMP[642]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11888.025 187.44 11888.305 188.44 ;
    END
  END Data_COMP[642]
  PIN Data_COMP[641]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11831.465 187.44 11831.745 188.44 ;
    END
  END Data_COMP[641]
  PIN Data_COMP[640]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11833.145 187.44 11833.425 188.44 ;
    END
  END Data_COMP[640]
  PIN Data_COMP[639]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11834.265 187.44 11834.545 188.44 ;
    END
  END Data_COMP[639]
  PIN Data_COMP[638]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11888.585 187.44 11888.865 188.44 ;
    END
  END Data_COMP[638]
  PIN Data_COMP[637]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11884.665 187.44 11884.945 188.44 ;
    END
  END Data_COMP[637]
  PIN Data_COMP[636]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11884.105 187.44 11884.385 188.44 ;
    END
  END Data_COMP[636]
  PIN Data_COMP[635]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11886.905 187.44 11887.185 188.44 ;
    END
  END Data_COMP[635]
  PIN Data_COMP[634]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11832.585 187.44 11832.865 188.44 ;
    END
  END Data_COMP[634]
  PIN Data_COMP[633]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11835.385 187.44 11835.665 188.44 ;
    END
  END Data_COMP[633]
  PIN Data_COMP[632]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11834.825 187.44 11835.105 188.44 ;
    END
  END Data_COMP[632]
  PIN Data_COMP[631]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11830.905 187.44 11831.185 188.44 ;
    END
  END Data_COMP[631]
  PIN Data_COMP[630]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11830.345 187.44 11830.625 188.44 ;
    END
  END Data_COMP[630]
  PIN Data_COMP[629]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11781.065 187.44 11781.345 188.44 ;
    END
  END Data_COMP[629]
  PIN Data_COMP[628]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11808.225 187.44 11808.505 188.44 ;
    END
  END Data_COMP[628]
  PIN Data_COMP[627]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11809.905 187.44 11810.185 188.44 ;
    END
  END Data_COMP[627]
  PIN Data_COMP[626]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11751.385 187.44 11751.665 188.44 ;
    END
  END Data_COMP[626]
  PIN Data_COMP[625]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11753.625 187.44 11753.905 188.44 ;
    END
  END Data_COMP[625]
  PIN Data_COMP[624]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11755.305 187.44 11755.585 188.44 ;
    END
  END Data_COMP[624]
  PIN Data_COMP[623]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11780.505 187.44 11780.785 188.44 ;
    END
  END Data_COMP[623]
  PIN Data_COMP[622]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11781.625 187.44 11781.905 188.44 ;
    END
  END Data_COMP[622]
  PIN Data_COMP[621]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11808.785 187.44 11809.065 188.44 ;
    END
  END Data_COMP[621]
  PIN Data_COMP[620]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11753.065 187.44 11753.345 188.44 ;
    END
  END Data_COMP[620]
  PIN Data_COMP[619]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11754.745 187.44 11755.025 188.44 ;
    END
  END Data_COMP[619]
  PIN Data_COMP[618]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11768.745 187.44 11769.025 188.44 ;
    END
  END Data_COMP[618]
  PIN Data_COMP[617]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11809.345 187.44 11809.625 188.44 ;
    END
  END Data_COMP[617]
  PIN Data_COMP[616]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11779.945 187.44 11780.225 188.44 ;
    END
  END Data_COMP[616]
  PIN Data_COMP[615]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11779.385 187.44 11779.665 188.44 ;
    END
  END Data_COMP[615]
  PIN Data_COMP[614]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11807.665 187.44 11807.945 188.44 ;
    END
  END Data_COMP[614]
  PIN Data_COMP[613]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11754.185 187.44 11754.465 188.44 ;
    END
  END Data_COMP[613]
  PIN Data_COMP[612]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11769.865 187.44 11770.145 188.44 ;
    END
  END Data_COMP[612]
  PIN Data_COMP[611]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11769.305 187.44 11769.585 188.44 ;
    END
  END Data_COMP[611]
  PIN Data_COMP[610]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11752.505 187.44 11752.785 188.44 ;
    END
  END Data_COMP[610]
  PIN Data_COMP[609]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11751.945 187.44 11752.225 188.44 ;
    END
  END Data_COMP[609]
  PIN Data_COMP[608]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11698.745 187.44 11699.025 188.44 ;
    END
  END Data_COMP[608]
  PIN Data_COMP[607]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11700.425 187.44 11700.705 188.44 ;
    END
  END Data_COMP[607]
  PIN Data_COMP[606]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11702.105 187.44 11702.385 188.44 ;
    END
  END Data_COMP[606]
  PIN Data_COMP[605]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11673.545 187.44 11673.825 188.44 ;
    END
  END Data_COMP[605]
  PIN Data_COMP[604]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11675.785 187.44 11676.065 188.44 ;
    END
  END Data_COMP[604]
  PIN Data_COMP[603]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11677.465 187.44 11677.745 188.44 ;
    END
  END Data_COMP[603]
  PIN Data_COMP[602]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11698.185 187.44 11698.465 188.44 ;
    END
  END Data_COMP[602]
  PIN Data_COMP[601]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11699.305 187.44 11699.585 188.44 ;
    END
  END Data_COMP[601]
  PIN Data_COMP[600]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11700.985 187.44 11701.265 188.44 ;
    END
  END Data_COMP[600]
  PIN Data_COMP[599]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11675.225 187.44 11675.505 188.44 ;
    END
  END Data_COMP[599]
  PIN Data_COMP[598]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11676.905 187.44 11677.185 188.44 ;
    END
  END Data_COMP[598]
  PIN Data_COMP[597]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11678.025 187.44 11678.305 188.44 ;
    END
  END Data_COMP[597]
  PIN Data_COMP[596]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11701.545 187.44 11701.825 188.44 ;
    END
  END Data_COMP[596]
  PIN Data_COMP[595]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11697.625 187.44 11697.905 188.44 ;
    END
  END Data_COMP[595]
  PIN Data_COMP[594]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11697.065 187.44 11697.345 188.44 ;
    END
  END Data_COMP[594]
  PIN Data_COMP[593]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11699.865 187.44 11700.145 188.44 ;
    END
  END Data_COMP[593]
  PIN Data_COMP[592]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11676.345 187.44 11676.625 188.44 ;
    END
  END Data_COMP[592]
  PIN Data_COMP[591]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11679.145 187.44 11679.425 188.44 ;
    END
  END Data_COMP[591]
  PIN Data_COMP[590]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11678.585 187.44 11678.865 188.44 ;
    END
  END Data_COMP[590]
  PIN Data_COMP[589]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11674.665 187.44 11674.945 188.44 ;
    END
  END Data_COMP[589]
  PIN Data_COMP[588]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11674.105 187.44 11674.385 188.44 ;
    END
  END Data_COMP[588]
  PIN Data_COMP[587]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11632.665 187.44 11632.945 188.44 ;
    END
  END Data_COMP[587]
  PIN Data_COMP[586]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11634.345 187.44 11634.625 188.44 ;
    END
  END Data_COMP[586]
  PIN Data_COMP[585]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11636.025 187.44 11636.305 188.44 ;
    END
  END Data_COMP[585]
  PIN Data_COMP[584]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11602.425 187.44 11602.705 188.44 ;
    END
  END Data_COMP[584]
  PIN Data_COMP[583]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11604.665 187.44 11604.945 188.44 ;
    END
  END Data_COMP[583]
  PIN Data_COMP[582]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11606.345 187.44 11606.625 188.44 ;
    END
  END Data_COMP[582]
  PIN Data_COMP[581]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11632.105 187.44 11632.385 188.44 ;
    END
  END Data_COMP[581]
  PIN Data_COMP[580]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11633.225 187.44 11633.505 188.44 ;
    END
  END Data_COMP[580]
  PIN Data_COMP[579]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11634.905 187.44 11635.185 188.44 ;
    END
  END Data_COMP[579]
  PIN Data_COMP[578]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11604.105 187.44 11604.385 188.44 ;
    END
  END Data_COMP[578]
  PIN Data_COMP[577]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11605.785 187.44 11606.065 188.44 ;
    END
  END Data_COMP[577]
  PIN Data_COMP[576]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11606.905 187.44 11607.185 188.44 ;
    END
  END Data_COMP[576]
  PIN Data_COMP[575]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11635.465 187.44 11635.745 188.44 ;
    END
  END Data_COMP[575]
  PIN Data_COMP[574]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11631.545 187.44 11631.825 188.44 ;
    END
  END Data_COMP[574]
  PIN Data_COMP[573]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11630.985 187.44 11631.265 188.44 ;
    END
  END Data_COMP[573]
  PIN Data_COMP[572]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11633.785 187.44 11634.065 188.44 ;
    END
  END Data_COMP[572]
  PIN Data_COMP[571]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11605.225 187.44 11605.505 188.44 ;
    END
  END Data_COMP[571]
  PIN Data_COMP[570]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11608.025 187.44 11608.305 188.44 ;
    END
  END Data_COMP[570]
  PIN Data_COMP[569]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11607.465 187.44 11607.745 188.44 ;
    END
  END Data_COMP[569]
  PIN Data_COMP[568]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11603.545 187.44 11603.825 188.44 ;
    END
  END Data_COMP[568]
  PIN Data_COMP[567]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11602.985 187.44 11603.265 188.44 ;
    END
  END Data_COMP[567]
  PIN Data_COMP[566]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11550.905 187.44 11551.185 188.44 ;
    END
  END Data_COMP[566]
  PIN Data_COMP[565]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11552.585 187.44 11552.865 188.44 ;
    END
  END Data_COMP[565]
  PIN Data_COMP[564]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11554.265 187.44 11554.545 188.44 ;
    END
  END Data_COMP[564]
  PIN Data_COMP[563]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11498.265 187.44 11498.545 188.44 ;
    END
  END Data_COMP[563]
  PIN Data_COMP[562]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11500.505 187.44 11500.785 188.44 ;
    END
  END Data_COMP[562]
  PIN Data_COMP[561]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11527.665 187.44 11527.945 188.44 ;
    END
  END Data_COMP[561]
  PIN Data_COMP[560]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11550.345 187.44 11550.625 188.44 ;
    END
  END Data_COMP[560]
  PIN Data_COMP[559]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11551.465 187.44 11551.745 188.44 ;
    END
  END Data_COMP[559]
  PIN Data_COMP[558]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11553.145 187.44 11553.425 188.44 ;
    END
  END Data_COMP[558]
  PIN Data_COMP[557]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11499.945 187.44 11500.225 188.44 ;
    END
  END Data_COMP[557]
  PIN Data_COMP[556]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11527.105 187.44 11527.385 188.44 ;
    END
  END Data_COMP[556]
  PIN Data_COMP[555]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11528.225 187.44 11528.505 188.44 ;
    END
  END Data_COMP[555]
  PIN Data_COMP[554]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11553.705 187.44 11553.985 188.44 ;
    END
  END Data_COMP[554]
  PIN Data_COMP[553]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11549.785 187.44 11550.065 188.44 ;
    END
  END Data_COMP[553]
  PIN Data_COMP[552]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11540.825 187.44 11541.105 188.44 ;
    END
  END Data_COMP[552]
  PIN Data_COMP[551]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11552.025 187.44 11552.305 188.44 ;
    END
  END Data_COMP[551]
  PIN Data_COMP[550]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11501.065 187.44 11501.345 188.44 ;
    END
  END Data_COMP[550]
  PIN Data_COMP[549]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11529.345 187.44 11529.625 188.44 ;
    END
  END Data_COMP[549]
  PIN Data_COMP[548]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11528.785 187.44 11529.065 188.44 ;
    END
  END Data_COMP[548]
  PIN Data_COMP[547]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11499.385 187.44 11499.665 188.44 ;
    END
  END Data_COMP[547]
  PIN Data_COMP[546]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11498.825 187.44 11499.105 188.44 ;
    END
  END Data_COMP[546]
  PIN Data_COMP[545]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11472.505 187.44 11472.785 188.44 ;
    END
  END Data_COMP[545]
  PIN Data_COMP[544]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11474.185 187.44 11474.465 188.44 ;
    END
  END Data_COMP[544]
  PIN Data_COMP[543]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11488.745 187.44 11489.025 188.44 ;
    END
  END Data_COMP[543]
  PIN Data_COMP[542]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11417.065 187.44 11417.345 188.44 ;
    END
  END Data_COMP[542]
  PIN Data_COMP[541]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11419.305 187.44 11419.585 188.44 ;
    END
  END Data_COMP[541]
  PIN Data_COMP[540]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11420.985 187.44 11421.265 188.44 ;
    END
  END Data_COMP[540]
  PIN Data_COMP[539]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11471.945 187.44 11472.225 188.44 ;
    END
  END Data_COMP[539]
  PIN Data_COMP[538]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11473.065 187.44 11473.345 188.44 ;
    END
  END Data_COMP[538]
  PIN Data_COMP[537]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11474.745 187.44 11475.025 188.44 ;
    END
  END Data_COMP[537]
  PIN Data_COMP[536]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11418.745 187.44 11419.025 188.44 ;
    END
  END Data_COMP[536]
  PIN Data_COMP[535]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11420.425 187.44 11420.705 188.44 ;
    END
  END Data_COMP[535]
  PIN Data_COMP[534]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11421.545 187.44 11421.825 188.44 ;
    END
  END Data_COMP[534]
  PIN Data_COMP[533]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11488.185 187.44 11488.465 188.44 ;
    END
  END Data_COMP[533]
  PIN Data_COMP[532]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11471.385 187.44 11471.665 188.44 ;
    END
  END Data_COMP[532]
  PIN Data_COMP[531]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11470.825 187.44 11471.105 188.44 ;
    END
  END Data_COMP[531]
  PIN Data_COMP[530]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11473.625 187.44 11473.905 188.44 ;
    END
  END Data_COMP[530]
  PIN Data_COMP[529]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11419.865 187.44 11420.145 188.44 ;
    END
  END Data_COMP[529]
  PIN Data_COMP[528]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11422.665 187.44 11422.945 188.44 ;
    END
  END Data_COMP[528]
  PIN Data_COMP[527]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11422.105 187.44 11422.385 188.44 ;
    END
  END Data_COMP[527]
  PIN Data_COMP[526]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11418.185 187.44 11418.465 188.44 ;
    END
  END Data_COMP[526]
  PIN Data_COMP[525]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11417.625 187.44 11417.905 188.44 ;
    END
  END Data_COMP[525]
  PIN Data_COMP[524]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11395.785 187.44 11396.065 188.44 ;
    END
  END Data_COMP[524]
  PIN Data_COMP[523]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11397.465 187.44 11397.745 188.44 ;
    END
  END Data_COMP[523]
  PIN Data_COMP[522]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11399.145 187.44 11399.425 188.44 ;
    END
  END Data_COMP[522]
  PIN Data_COMP[521]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11351.545 187.44 11351.825 188.44 ;
    END
  END Data_COMP[521]
  PIN Data_COMP[520]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11353.785 187.44 11354.065 188.44 ;
    END
  END Data_COMP[520]
  PIN Data_COMP[519]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11355.465 187.44 11355.745 188.44 ;
    END
  END Data_COMP[519]
  PIN Data_COMP[518]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11395.225 187.44 11395.505 188.44 ;
    END
  END Data_COMP[518]
  PIN Data_COMP[517]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11396.345 187.44 11396.625 188.44 ;
    END
  END Data_COMP[517]
  PIN Data_COMP[516]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11398.025 187.44 11398.305 188.44 ;
    END
  END Data_COMP[516]
  PIN Data_COMP[515]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11353.225 187.44 11353.505 188.44 ;
    END
  END Data_COMP[515]
  PIN Data_COMP[514]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11354.905 187.44 11355.185 188.44 ;
    END
  END Data_COMP[514]
  PIN Data_COMP[513]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11356.025 187.44 11356.305 188.44 ;
    END
  END Data_COMP[513]
  PIN Data_COMP[512]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11398.585 187.44 11398.865 188.44 ;
    END
  END Data_COMP[512]
  PIN Data_COMP[511]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11394.665 187.44 11394.945 188.44 ;
    END
  END Data_COMP[511]
  PIN Data_COMP[510]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11394.105 187.44 11394.385 188.44 ;
    END
  END Data_COMP[510]
  PIN Data_COMP[509]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11396.905 187.44 11397.185 188.44 ;
    END
  END Data_COMP[509]
  PIN Data_COMP[508]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11354.345 187.44 11354.625 188.44 ;
    END
  END Data_COMP[508]
  PIN Data_COMP[507]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11357.145 187.44 11357.425 188.44 ;
    END
  END Data_COMP[507]
  PIN Data_COMP[506]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11356.585 187.44 11356.865 188.44 ;
    END
  END Data_COMP[506]
  PIN Data_COMP[505]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11352.665 187.44 11352.945 188.44 ;
    END
  END Data_COMP[505]
  PIN Data_COMP[504]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11352.105 187.44 11352.385 188.44 ;
    END
  END Data_COMP[504]
  PIN Data_COMP[503]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11325.785 187.44 11326.065 188.44 ;
    END
  END Data_COMP[503]
  PIN Data_COMP[502]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11327.465 187.44 11327.745 188.44 ;
    END
  END Data_COMP[502]
  PIN Data_COMP[501]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11329.145 187.44 11329.425 188.44 ;
    END
  END Data_COMP[501]
  PIN Data_COMP[500]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11269.785 187.44 11270.065 188.44 ;
    END
  END Data_COMP[500]
  PIN Data_COMP[499]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11272.025 187.44 11272.305 188.44 ;
    END
  END Data_COMP[499]
  PIN Data_COMP[498]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11273.705 187.44 11273.985 188.44 ;
    END
  END Data_COMP[498]
  PIN Data_COMP[497]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11325.225 187.44 11325.505 188.44 ;
    END
  END Data_COMP[497]
  PIN Data_COMP[496]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11326.345 187.44 11326.625 188.44 ;
    END
  END Data_COMP[496]
  PIN Data_COMP[495]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11328.025 187.44 11328.305 188.44 ;
    END
  END Data_COMP[495]
  PIN Data_COMP[494]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11271.465 187.44 11271.745 188.44 ;
    END
  END Data_COMP[494]
  PIN Data_COMP[493]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11273.145 187.44 11273.425 188.44 ;
    END
  END Data_COMP[493]
  PIN Data_COMP[492]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11274.265 187.44 11274.545 188.44 ;
    END
  END Data_COMP[492]
  PIN Data_COMP[491]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11328.585 187.44 11328.865 188.44 ;
    END
  END Data_COMP[491]
  PIN Data_COMP[490]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11324.665 187.44 11324.945 188.44 ;
    END
  END Data_COMP[490]
  PIN Data_COMP[489]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11324.105 187.44 11324.385 188.44 ;
    END
  END Data_COMP[489]
  PIN Data_COMP[488]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11326.905 187.44 11327.185 188.44 ;
    END
  END Data_COMP[488]
  PIN Data_COMP[487]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11272.585 187.44 11272.865 188.44 ;
    END
  END Data_COMP[487]
  PIN Data_COMP[486]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11275.385 187.44 11275.665 188.44 ;
    END
  END Data_COMP[486]
  PIN Data_COMP[485]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11274.825 187.44 11275.105 188.44 ;
    END
  END Data_COMP[485]
  PIN Data_COMP[484]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11270.905 187.44 11271.185 188.44 ;
    END
  END Data_COMP[484]
  PIN Data_COMP[483]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11270.345 187.44 11270.625 188.44 ;
    END
  END Data_COMP[483]
  PIN Data_COMP[482]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11221.065 187.44 11221.345 188.44 ;
    END
  END Data_COMP[482]
  PIN Data_COMP[481]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11248.225 187.44 11248.505 188.44 ;
    END
  END Data_COMP[481]
  PIN Data_COMP[480]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11249.905 187.44 11250.185 188.44 ;
    END
  END Data_COMP[480]
  PIN Data_COMP[479]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11191.385 187.44 11191.665 188.44 ;
    END
  END Data_COMP[479]
  PIN Data_COMP[478]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11193.625 187.44 11193.905 188.44 ;
    END
  END Data_COMP[478]
  PIN Data_COMP[477]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11195.305 187.44 11195.585 188.44 ;
    END
  END Data_COMP[477]
  PIN Data_COMP[476]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11220.505 187.44 11220.785 188.44 ;
    END
  END Data_COMP[476]
  PIN Data_COMP[475]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11221.625 187.44 11221.905 188.44 ;
    END
  END Data_COMP[475]
  PIN Data_COMP[474]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11248.785 187.44 11249.065 188.44 ;
    END
  END Data_COMP[474]
  PIN Data_COMP[473]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11193.065 187.44 11193.345 188.44 ;
    END
  END Data_COMP[473]
  PIN Data_COMP[472]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11194.745 187.44 11195.025 188.44 ;
    END
  END Data_COMP[472]
  PIN Data_COMP[471]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11208.745 187.44 11209.025 188.44 ;
    END
  END Data_COMP[471]
  PIN Data_COMP[470]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11249.345 187.44 11249.625 188.44 ;
    END
  END Data_COMP[470]
  PIN Data_COMP[469]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11219.945 187.44 11220.225 188.44 ;
    END
  END Data_COMP[469]
  PIN Data_COMP[468]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11219.385 187.44 11219.665 188.44 ;
    END
  END Data_COMP[468]
  PIN Data_COMP[467]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11247.665 187.44 11247.945 188.44 ;
    END
  END Data_COMP[467]
  PIN Data_COMP[466]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11194.185 187.44 11194.465 188.44 ;
    END
  END Data_COMP[466]
  PIN Data_COMP[465]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11209.865 187.44 11210.145 188.44 ;
    END
  END Data_COMP[465]
  PIN Data_COMP[464]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11209.305 187.44 11209.585 188.44 ;
    END
  END Data_COMP[464]
  PIN Data_COMP[463]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11192.505 187.44 11192.785 188.44 ;
    END
  END Data_COMP[463]
  PIN Data_COMP[462]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11191.945 187.44 11192.225 188.44 ;
    END
  END Data_COMP[462]
  PIN Data_COMP[461]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11138.745 187.44 11139.025 188.44 ;
    END
  END Data_COMP[461]
  PIN Data_COMP[460]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11140.425 187.44 11140.705 188.44 ;
    END
  END Data_COMP[460]
  PIN Data_COMP[459]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11142.105 187.44 11142.385 188.44 ;
    END
  END Data_COMP[459]
  PIN Data_COMP[458]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11113.545 187.44 11113.825 188.44 ;
    END
  END Data_COMP[458]
  PIN Data_COMP[457]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11115.785 187.44 11116.065 188.44 ;
    END
  END Data_COMP[457]
  PIN Data_COMP[456]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11117.465 187.44 11117.745 188.44 ;
    END
  END Data_COMP[456]
  PIN Data_COMP[455]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11138.185 187.44 11138.465 188.44 ;
    END
  END Data_COMP[455]
  PIN Data_COMP[454]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11139.305 187.44 11139.585 188.44 ;
    END
  END Data_COMP[454]
  PIN Data_COMP[453]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11140.985 187.44 11141.265 188.44 ;
    END
  END Data_COMP[453]
  PIN Data_COMP[452]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11115.225 187.44 11115.505 188.44 ;
    END
  END Data_COMP[452]
  PIN Data_COMP[451]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11116.905 187.44 11117.185 188.44 ;
    END
  END Data_COMP[451]
  PIN Data_COMP[450]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11118.025 187.44 11118.305 188.44 ;
    END
  END Data_COMP[450]
  PIN Data_COMP[449]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11141.545 187.44 11141.825 188.44 ;
    END
  END Data_COMP[449]
  PIN Data_COMP[448]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11137.625 187.44 11137.905 188.44 ;
    END
  END Data_COMP[448]
  PIN Data_COMP[447]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11137.065 187.44 11137.345 188.44 ;
    END
  END Data_COMP[447]
  PIN Data_COMP[446]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11139.865 187.44 11140.145 188.44 ;
    END
  END Data_COMP[446]
  PIN Data_COMP[445]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11116.345 187.44 11116.625 188.44 ;
    END
  END Data_COMP[445]
  PIN Data_COMP[444]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11119.145 187.44 11119.425 188.44 ;
    END
  END Data_COMP[444]
  PIN Data_COMP[443]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11118.585 187.44 11118.865 188.44 ;
    END
  END Data_COMP[443]
  PIN Data_COMP[442]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11114.665 187.44 11114.945 188.44 ;
    END
  END Data_COMP[442]
  PIN Data_COMP[441]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11114.105 187.44 11114.385 188.44 ;
    END
  END Data_COMP[441]
  PIN Data_COMP[440]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11072.665 187.44 11072.945 188.44 ;
    END
  END Data_COMP[440]
  PIN Data_COMP[439]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11074.345 187.44 11074.625 188.44 ;
    END
  END Data_COMP[439]
  PIN Data_COMP[438]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11076.025 187.44 11076.305 188.44 ;
    END
  END Data_COMP[438]
  PIN Data_COMP[437]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11042.425 187.44 11042.705 188.44 ;
    END
  END Data_COMP[437]
  PIN Data_COMP[436]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11044.665 187.44 11044.945 188.44 ;
    END
  END Data_COMP[436]
  PIN Data_COMP[435]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11046.345 187.44 11046.625 188.44 ;
    END
  END Data_COMP[435]
  PIN Data_COMP[434]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11072.105 187.44 11072.385 188.44 ;
    END
  END Data_COMP[434]
  PIN Data_COMP[433]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11073.225 187.44 11073.505 188.44 ;
    END
  END Data_COMP[433]
  PIN Data_COMP[432]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11074.905 187.44 11075.185 188.44 ;
    END
  END Data_COMP[432]
  PIN Data_COMP[431]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11044.105 187.44 11044.385 188.44 ;
    END
  END Data_COMP[431]
  PIN Data_COMP[430]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11045.785 187.44 11046.065 188.44 ;
    END
  END Data_COMP[430]
  PIN Data_COMP[429]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11046.905 187.44 11047.185 188.44 ;
    END
  END Data_COMP[429]
  PIN Data_COMP[428]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11075.465 187.44 11075.745 188.44 ;
    END
  END Data_COMP[428]
  PIN Data_COMP[427]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11071.545 187.44 11071.825 188.44 ;
    END
  END Data_COMP[427]
  PIN Data_COMP[426]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11070.985 187.44 11071.265 188.44 ;
    END
  END Data_COMP[426]
  PIN Data_COMP[425]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11073.785 187.44 11074.065 188.44 ;
    END
  END Data_COMP[425]
  PIN Data_COMP[424]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11045.225 187.44 11045.505 188.44 ;
    END
  END Data_COMP[424]
  PIN Data_COMP[423]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11048.025 187.44 11048.305 188.44 ;
    END
  END Data_COMP[423]
  PIN Data_COMP[422]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11047.465 187.44 11047.745 188.44 ;
    END
  END Data_COMP[422]
  PIN Data_COMP[421]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11043.545 187.44 11043.825 188.44 ;
    END
  END Data_COMP[421]
  PIN Data_COMP[420]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11042.985 187.44 11043.265 188.44 ;
    END
  END Data_COMP[420]
  PIN Data_COMP[419]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10990.905 187.44 10991.185 188.44 ;
    END
  END Data_COMP[419]
  PIN Data_COMP[418]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10992.585 187.44 10992.865 188.44 ;
    END
  END Data_COMP[418]
  PIN Data_COMP[417]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10994.265 187.44 10994.545 188.44 ;
    END
  END Data_COMP[417]
  PIN Data_COMP[416]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10938.265 187.44 10938.545 188.44 ;
    END
  END Data_COMP[416]
  PIN Data_COMP[415]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10940.505 187.44 10940.785 188.44 ;
    END
  END Data_COMP[415]
  PIN Data_COMP[414]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10967.665 187.44 10967.945 188.44 ;
    END
  END Data_COMP[414]
  PIN Data_COMP[413]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10990.345 187.44 10990.625 188.44 ;
    END
  END Data_COMP[413]
  PIN Data_COMP[412]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10991.465 187.44 10991.745 188.44 ;
    END
  END Data_COMP[412]
  PIN Data_COMP[411]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10993.145 187.44 10993.425 188.44 ;
    END
  END Data_COMP[411]
  PIN Data_COMP[410]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10939.945 187.44 10940.225 188.44 ;
    END
  END Data_COMP[410]
  PIN Data_COMP[409]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10967.105 187.44 10967.385 188.44 ;
    END
  END Data_COMP[409]
  PIN Data_COMP[408]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10968.225 187.44 10968.505 188.44 ;
    END
  END Data_COMP[408]
  PIN Data_COMP[407]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10993.705 187.44 10993.985 188.44 ;
    END
  END Data_COMP[407]
  PIN Data_COMP[406]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10989.785 187.44 10990.065 188.44 ;
    END
  END Data_COMP[406]
  PIN Data_COMP[405]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10980.825 187.44 10981.105 188.44 ;
    END
  END Data_COMP[405]
  PIN Data_COMP[404]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10992.025 187.44 10992.305 188.44 ;
    END
  END Data_COMP[404]
  PIN Data_COMP[403]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10941.065 187.44 10941.345 188.44 ;
    END
  END Data_COMP[403]
  PIN Data_COMP[402]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10969.345 187.44 10969.625 188.44 ;
    END
  END Data_COMP[402]
  PIN Data_COMP[401]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10968.785 187.44 10969.065 188.44 ;
    END
  END Data_COMP[401]
  PIN Data_COMP[400]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10939.385 187.44 10939.665 188.44 ;
    END
  END Data_COMP[400]
  PIN Data_COMP[399]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10938.825 187.44 10939.105 188.44 ;
    END
  END Data_COMP[399]
  PIN Data_COMP[398]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10912.505 187.44 10912.785 188.44 ;
    END
  END Data_COMP[398]
  PIN Data_COMP[397]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10914.185 187.44 10914.465 188.44 ;
    END
  END Data_COMP[397]
  PIN Data_COMP[396]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10928.745 187.44 10929.025 188.44 ;
    END
  END Data_COMP[396]
  PIN Data_COMP[395]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10857.065 187.44 10857.345 188.44 ;
    END
  END Data_COMP[395]
  PIN Data_COMP[394]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10859.305 187.44 10859.585 188.44 ;
    END
  END Data_COMP[394]
  PIN Data_COMP[393]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10860.985 187.44 10861.265 188.44 ;
    END
  END Data_COMP[393]
  PIN Data_COMP[392]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10911.945 187.44 10912.225 188.44 ;
    END
  END Data_COMP[392]
  PIN Data_COMP[391]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10913.065 187.44 10913.345 188.44 ;
    END
  END Data_COMP[391]
  PIN Data_COMP[390]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10914.745 187.44 10915.025 188.44 ;
    END
  END Data_COMP[390]
  PIN Data_COMP[389]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10858.745 187.44 10859.025 188.44 ;
    END
  END Data_COMP[389]
  PIN Data_COMP[388]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10860.425 187.44 10860.705 188.44 ;
    END
  END Data_COMP[388]
  PIN Data_COMP[387]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10861.545 187.44 10861.825 188.44 ;
    END
  END Data_COMP[387]
  PIN Data_COMP[386]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10928.185 187.44 10928.465 188.44 ;
    END
  END Data_COMP[386]
  PIN Data_COMP[385]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10911.385 187.44 10911.665 188.44 ;
    END
  END Data_COMP[385]
  PIN Data_COMP[384]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10910.825 187.44 10911.105 188.44 ;
    END
  END Data_COMP[384]
  PIN Data_COMP[383]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10913.625 187.44 10913.905 188.44 ;
    END
  END Data_COMP[383]
  PIN Data_COMP[382]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10859.865 187.44 10860.145 188.44 ;
    END
  END Data_COMP[382]
  PIN Data_COMP[381]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10862.665 187.44 10862.945 188.44 ;
    END
  END Data_COMP[381]
  PIN Data_COMP[380]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10862.105 187.44 10862.385 188.44 ;
    END
  END Data_COMP[380]
  PIN Data_COMP[379]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10858.185 187.44 10858.465 188.44 ;
    END
  END Data_COMP[379]
  PIN Data_COMP[378]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10857.625 187.44 10857.905 188.44 ;
    END
  END Data_COMP[378]
  PIN Data_COMP[377]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10835.785 187.44 10836.065 188.44 ;
    END
  END Data_COMP[377]
  PIN Data_COMP[376]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10837.465 187.44 10837.745 188.44 ;
    END
  END Data_COMP[376]
  PIN Data_COMP[375]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10839.145 187.44 10839.425 188.44 ;
    END
  END Data_COMP[375]
  PIN Data_COMP[374]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10791.545 187.44 10791.825 188.44 ;
    END
  END Data_COMP[374]
  PIN Data_COMP[373]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10793.785 187.44 10794.065 188.44 ;
    END
  END Data_COMP[373]
  PIN Data_COMP[372]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10795.465 187.44 10795.745 188.44 ;
    END
  END Data_COMP[372]
  PIN Data_COMP[371]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10835.225 187.44 10835.505 188.44 ;
    END
  END Data_COMP[371]
  PIN Data_COMP[370]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10836.345 187.44 10836.625 188.44 ;
    END
  END Data_COMP[370]
  PIN Data_COMP[369]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10838.025 187.44 10838.305 188.44 ;
    END
  END Data_COMP[369]
  PIN Data_COMP[368]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10793.225 187.44 10793.505 188.44 ;
    END
  END Data_COMP[368]
  PIN Data_COMP[367]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10794.905 187.44 10795.185 188.44 ;
    END
  END Data_COMP[367]
  PIN Data_COMP[366]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10796.025 187.44 10796.305 188.44 ;
    END
  END Data_COMP[366]
  PIN Data_COMP[365]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10838.585 187.44 10838.865 188.44 ;
    END
  END Data_COMP[365]
  PIN Data_COMP[364]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10834.665 187.44 10834.945 188.44 ;
    END
  END Data_COMP[364]
  PIN Data_COMP[363]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10834.105 187.44 10834.385 188.44 ;
    END
  END Data_COMP[363]
  PIN Data_COMP[362]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10836.905 187.44 10837.185 188.44 ;
    END
  END Data_COMP[362]
  PIN Data_COMP[361]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10794.345 187.44 10794.625 188.44 ;
    END
  END Data_COMP[361]
  PIN Data_COMP[360]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10797.145 187.44 10797.425 188.44 ;
    END
  END Data_COMP[360]
  PIN Data_COMP[359]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10796.585 187.44 10796.865 188.44 ;
    END
  END Data_COMP[359]
  PIN Data_COMP[358]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10792.665 187.44 10792.945 188.44 ;
    END
  END Data_COMP[358]
  PIN Data_COMP[357]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10792.105 187.44 10792.385 188.44 ;
    END
  END Data_COMP[357]
  PIN Data_COMP[356]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10765.785 187.44 10766.065 188.44 ;
    END
  END Data_COMP[356]
  PIN Data_COMP[355]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10767.465 187.44 10767.745 188.44 ;
    END
  END Data_COMP[355]
  PIN Data_COMP[354]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10769.145 187.44 10769.425 188.44 ;
    END
  END Data_COMP[354]
  PIN Data_COMP[353]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10709.785 187.44 10710.065 188.44 ;
    END
  END Data_COMP[353]
  PIN Data_COMP[352]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10712.025 187.44 10712.305 188.44 ;
    END
  END Data_COMP[352]
  PIN Data_COMP[351]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10713.705 187.44 10713.985 188.44 ;
    END
  END Data_COMP[351]
  PIN Data_COMP[350]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10765.225 187.44 10765.505 188.44 ;
    END
  END Data_COMP[350]
  PIN Data_COMP[349]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10766.345 187.44 10766.625 188.44 ;
    END
  END Data_COMP[349]
  PIN Data_COMP[348]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10768.025 187.44 10768.305 188.44 ;
    END
  END Data_COMP[348]
  PIN Data_COMP[347]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10711.465 187.44 10711.745 188.44 ;
    END
  END Data_COMP[347]
  PIN Data_COMP[346]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10713.145 187.44 10713.425 188.44 ;
    END
  END Data_COMP[346]
  PIN Data_COMP[345]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10714.265 187.44 10714.545 188.44 ;
    END
  END Data_COMP[345]
  PIN Data_COMP[344]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10768.585 187.44 10768.865 188.44 ;
    END
  END Data_COMP[344]
  PIN Data_COMP[343]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10764.665 187.44 10764.945 188.44 ;
    END
  END Data_COMP[343]
  PIN Data_COMP[342]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10764.105 187.44 10764.385 188.44 ;
    END
  END Data_COMP[342]
  PIN Data_COMP[341]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10766.905 187.44 10767.185 188.44 ;
    END
  END Data_COMP[341]
  PIN Data_COMP[340]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10712.585 187.44 10712.865 188.44 ;
    END
  END Data_COMP[340]
  PIN Data_COMP[339]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10715.385 187.44 10715.665 188.44 ;
    END
  END Data_COMP[339]
  PIN Data_COMP[338]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10714.825 187.44 10715.105 188.44 ;
    END
  END Data_COMP[338]
  PIN Data_COMP[337]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10710.905 187.44 10711.185 188.44 ;
    END
  END Data_COMP[337]
  PIN Data_COMP[336]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10710.345 187.44 10710.625 188.44 ;
    END
  END Data_COMP[336]
  PIN Data_COMP[335]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10661.065 187.44 10661.345 188.44 ;
    END
  END Data_COMP[335]
  PIN Data_COMP[334]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10688.225 187.44 10688.505 188.44 ;
    END
  END Data_COMP[334]
  PIN Data_COMP[333]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10689.905 187.44 10690.185 188.44 ;
    END
  END Data_COMP[333]
  PIN Data_COMP[332]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10631.385 187.44 10631.665 188.44 ;
    END
  END Data_COMP[332]
  PIN Data_COMP[331]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10633.625 187.44 10633.905 188.44 ;
    END
  END Data_COMP[331]
  PIN Data_COMP[330]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10635.305 187.44 10635.585 188.44 ;
    END
  END Data_COMP[330]
  PIN Data_COMP[329]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10660.505 187.44 10660.785 188.44 ;
    END
  END Data_COMP[329]
  PIN Data_COMP[328]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10661.625 187.44 10661.905 188.44 ;
    END
  END Data_COMP[328]
  PIN Data_COMP[327]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10688.785 187.44 10689.065 188.44 ;
    END
  END Data_COMP[327]
  PIN Data_COMP[326]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10633.065 187.44 10633.345 188.44 ;
    END
  END Data_COMP[326]
  PIN Data_COMP[325]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10634.745 187.44 10635.025 188.44 ;
    END
  END Data_COMP[325]
  PIN Data_COMP[324]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10648.745 187.44 10649.025 188.44 ;
    END
  END Data_COMP[324]
  PIN Data_COMP[323]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10689.345 187.44 10689.625 188.44 ;
    END
  END Data_COMP[323]
  PIN Data_COMP[322]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10659.945 187.44 10660.225 188.44 ;
    END
  END Data_COMP[322]
  PIN Data_COMP[321]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10659.385 187.44 10659.665 188.44 ;
    END
  END Data_COMP[321]
  PIN Data_COMP[320]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10687.665 187.44 10687.945 188.44 ;
    END
  END Data_COMP[320]
  PIN Data_COMP[319]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10634.185 187.44 10634.465 188.44 ;
    END
  END Data_COMP[319]
  PIN Data_COMP[318]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10649.865 187.44 10650.145 188.44 ;
    END
  END Data_COMP[318]
  PIN Data_COMP[317]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10649.305 187.44 10649.585 188.44 ;
    END
  END Data_COMP[317]
  PIN Data_COMP[316]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10632.505 187.44 10632.785 188.44 ;
    END
  END Data_COMP[316]
  PIN Data_COMP[315]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10631.945 187.44 10632.225 188.44 ;
    END
  END Data_COMP[315]
  PIN Data_COMP[314]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10578.745 187.44 10579.025 188.44 ;
    END
  END Data_COMP[314]
  PIN Data_COMP[313]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10580.425 187.44 10580.705 188.44 ;
    END
  END Data_COMP[313]
  PIN Data_COMP[312]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10582.105 187.44 10582.385 188.44 ;
    END
  END Data_COMP[312]
  PIN Data_COMP[311]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10553.545 187.44 10553.825 188.44 ;
    END
  END Data_COMP[311]
  PIN Data_COMP[310]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10555.785 187.44 10556.065 188.44 ;
    END
  END Data_COMP[310]
  PIN Data_COMP[309]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10557.465 187.44 10557.745 188.44 ;
    END
  END Data_COMP[309]
  PIN Data_COMP[308]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10578.185 187.44 10578.465 188.44 ;
    END
  END Data_COMP[308]
  PIN Data_COMP[307]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10579.305 187.44 10579.585 188.44 ;
    END
  END Data_COMP[307]
  PIN Data_COMP[306]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10580.985 187.44 10581.265 188.44 ;
    END
  END Data_COMP[306]
  PIN Data_COMP[305]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10555.225 187.44 10555.505 188.44 ;
    END
  END Data_COMP[305]
  PIN Data_COMP[304]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10556.905 187.44 10557.185 188.44 ;
    END
  END Data_COMP[304]
  PIN Data_COMP[303]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10558.025 187.44 10558.305 188.44 ;
    END
  END Data_COMP[303]
  PIN Data_COMP[302]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10581.545 187.44 10581.825 188.44 ;
    END
  END Data_COMP[302]
  PIN Data_COMP[301]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10577.625 187.44 10577.905 188.44 ;
    END
  END Data_COMP[301]
  PIN Data_COMP[300]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10577.065 187.44 10577.345 188.44 ;
    END
  END Data_COMP[300]
  PIN Data_COMP[299]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10579.865 187.44 10580.145 188.44 ;
    END
  END Data_COMP[299]
  PIN Data_COMP[298]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10556.345 187.44 10556.625 188.44 ;
    END
  END Data_COMP[298]
  PIN Data_COMP[297]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10559.145 187.44 10559.425 188.44 ;
    END
  END Data_COMP[297]
  PIN Data_COMP[296]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10558.585 187.44 10558.865 188.44 ;
    END
  END Data_COMP[296]
  PIN Data_COMP[295]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10554.665 187.44 10554.945 188.44 ;
    END
  END Data_COMP[295]
  PIN Data_COMP[294]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10554.105 187.44 10554.385 188.44 ;
    END
  END Data_COMP[294]
  PIN Data_COMP[293]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10512.665 187.44 10512.945 188.44 ;
    END
  END Data_COMP[293]
  PIN Data_COMP[292]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10514.345 187.44 10514.625 188.44 ;
    END
  END Data_COMP[292]
  PIN Data_COMP[291]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10516.025 187.44 10516.305 188.44 ;
    END
  END Data_COMP[291]
  PIN Data_COMP[290]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10482.425 187.44 10482.705 188.44 ;
    END
  END Data_COMP[290]
  PIN Data_COMP[289]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10484.665 187.44 10484.945 188.44 ;
    END
  END Data_COMP[289]
  PIN Data_COMP[288]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10486.345 187.44 10486.625 188.44 ;
    END
  END Data_COMP[288]
  PIN Data_COMP[287]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10512.105 187.44 10512.385 188.44 ;
    END
  END Data_COMP[287]
  PIN Data_COMP[286]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10513.225 187.44 10513.505 188.44 ;
    END
  END Data_COMP[286]
  PIN Data_COMP[285]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10514.905 187.44 10515.185 188.44 ;
    END
  END Data_COMP[285]
  PIN Data_COMP[284]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10484.105 187.44 10484.385 188.44 ;
    END
  END Data_COMP[284]
  PIN Data_COMP[283]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10485.785 187.44 10486.065 188.44 ;
    END
  END Data_COMP[283]
  PIN Data_COMP[282]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10486.905 187.44 10487.185 188.44 ;
    END
  END Data_COMP[282]
  PIN Data_COMP[281]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10515.465 187.44 10515.745 188.44 ;
    END
  END Data_COMP[281]
  PIN Data_COMP[280]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10511.545 187.44 10511.825 188.44 ;
    END
  END Data_COMP[280]
  PIN Data_COMP[279]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10510.985 187.44 10511.265 188.44 ;
    END
  END Data_COMP[279]
  PIN Data_COMP[278]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10513.785 187.44 10514.065 188.44 ;
    END
  END Data_COMP[278]
  PIN Data_COMP[277]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10485.225 187.44 10485.505 188.44 ;
    END
  END Data_COMP[277]
  PIN Data_COMP[276]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10488.025 187.44 10488.305 188.44 ;
    END
  END Data_COMP[276]
  PIN Data_COMP[275]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10487.465 187.44 10487.745 188.44 ;
    END
  END Data_COMP[275]
  PIN Data_COMP[274]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10483.545 187.44 10483.825 188.44 ;
    END
  END Data_COMP[274]
  PIN Data_COMP[273]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10482.985 187.44 10483.265 188.44 ;
    END
  END Data_COMP[273]
  PIN Data_COMP[272]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10430.905 187.44 10431.185 188.44 ;
    END
  END Data_COMP[272]
  PIN Data_COMP[271]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10432.585 187.44 10432.865 188.44 ;
    END
  END Data_COMP[271]
  PIN Data_COMP[270]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10434.265 187.44 10434.545 188.44 ;
    END
  END Data_COMP[270]
  PIN Data_COMP[269]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10378.265 187.44 10378.545 188.44 ;
    END
  END Data_COMP[269]
  PIN Data_COMP[268]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10380.505 187.44 10380.785 188.44 ;
    END
  END Data_COMP[268]
  PIN Data_COMP[267]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10407.665 187.44 10407.945 188.44 ;
    END
  END Data_COMP[267]
  PIN Data_COMP[266]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10430.345 187.44 10430.625 188.44 ;
    END
  END Data_COMP[266]
  PIN Data_COMP[265]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10431.465 187.44 10431.745 188.44 ;
    END
  END Data_COMP[265]
  PIN Data_COMP[264]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10433.145 187.44 10433.425 188.44 ;
    END
  END Data_COMP[264]
  PIN Data_COMP[263]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10379.945 187.44 10380.225 188.44 ;
    END
  END Data_COMP[263]
  PIN Data_COMP[262]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10407.105 187.44 10407.385 188.44 ;
    END
  END Data_COMP[262]
  PIN Data_COMP[261]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10408.225 187.44 10408.505 188.44 ;
    END
  END Data_COMP[261]
  PIN Data_COMP[260]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10433.705 187.44 10433.985 188.44 ;
    END
  END Data_COMP[260]
  PIN Data_COMP[259]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10429.785 187.44 10430.065 188.44 ;
    END
  END Data_COMP[259]
  PIN Data_COMP[258]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10420.825 187.44 10421.105 188.44 ;
    END
  END Data_COMP[258]
  PIN Data_COMP[257]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10432.025 187.44 10432.305 188.44 ;
    END
  END Data_COMP[257]
  PIN Data_COMP[256]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10381.065 187.44 10381.345 188.44 ;
    END
  END Data_COMP[256]
  PIN Data_COMP[255]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10409.345 187.44 10409.625 188.44 ;
    END
  END Data_COMP[255]
  PIN Data_COMP[254]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10408.785 187.44 10409.065 188.44 ;
    END
  END Data_COMP[254]
  PIN Data_COMP[253]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10379.385 187.44 10379.665 188.44 ;
    END
  END Data_COMP[253]
  PIN Data_COMP[252]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10378.825 187.44 10379.105 188.44 ;
    END
  END Data_COMP[252]
  PIN Data_COMP[251]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10352.505 187.44 10352.785 188.44 ;
    END
  END Data_COMP[251]
  PIN Data_COMP[250]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10354.185 187.44 10354.465 188.44 ;
    END
  END Data_COMP[250]
  PIN Data_COMP[249]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10368.745 187.44 10369.025 188.44 ;
    END
  END Data_COMP[249]
  PIN Data_COMP[248]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10297.065 187.44 10297.345 188.44 ;
    END
  END Data_COMP[248]
  PIN Data_COMP[247]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10299.305 187.44 10299.585 188.44 ;
    END
  END Data_COMP[247]
  PIN Data_COMP[246]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10300.985 187.44 10301.265 188.44 ;
    END
  END Data_COMP[246]
  PIN Data_COMP[245]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10351.945 187.44 10352.225 188.44 ;
    END
  END Data_COMP[245]
  PIN Data_COMP[244]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10353.065 187.44 10353.345 188.44 ;
    END
  END Data_COMP[244]
  PIN Data_COMP[243]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10354.745 187.44 10355.025 188.44 ;
    END
  END Data_COMP[243]
  PIN Data_COMP[242]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10298.745 187.44 10299.025 188.44 ;
    END
  END Data_COMP[242]
  PIN Data_COMP[241]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10300.425 187.44 10300.705 188.44 ;
    END
  END Data_COMP[241]
  PIN Data_COMP[240]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10301.545 187.44 10301.825 188.44 ;
    END
  END Data_COMP[240]
  PIN Data_COMP[239]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10368.185 187.44 10368.465 188.44 ;
    END
  END Data_COMP[239]
  PIN Data_COMP[238]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10351.385 187.44 10351.665 188.44 ;
    END
  END Data_COMP[238]
  PIN Data_COMP[237]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10350.825 187.44 10351.105 188.44 ;
    END
  END Data_COMP[237]
  PIN Data_COMP[236]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10353.625 187.44 10353.905 188.44 ;
    END
  END Data_COMP[236]
  PIN Data_COMP[235]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10299.865 187.44 10300.145 188.44 ;
    END
  END Data_COMP[235]
  PIN Data_COMP[234]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10302.665 187.44 10302.945 188.44 ;
    END
  END Data_COMP[234]
  PIN Data_COMP[233]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10302.105 187.44 10302.385 188.44 ;
    END
  END Data_COMP[233]
  PIN Data_COMP[232]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10298.185 187.44 10298.465 188.44 ;
    END
  END Data_COMP[232]
  PIN Data_COMP[231]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10297.625 187.44 10297.905 188.44 ;
    END
  END Data_COMP[231]
  PIN Data_COMP[230]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10275.785 187.44 10276.065 188.44 ;
    END
  END Data_COMP[230]
  PIN Data_COMP[229]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10277.465 187.44 10277.745 188.44 ;
    END
  END Data_COMP[229]
  PIN Data_COMP[228]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10279.145 187.44 10279.425 188.44 ;
    END
  END Data_COMP[228]
  PIN Data_COMP[227]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10231.545 187.44 10231.825 188.44 ;
    END
  END Data_COMP[227]
  PIN Data_COMP[226]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10233.785 187.44 10234.065 188.44 ;
    END
  END Data_COMP[226]
  PIN Data_COMP[225]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10235.465 187.44 10235.745 188.44 ;
    END
  END Data_COMP[225]
  PIN Data_COMP[224]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10275.225 187.44 10275.505 188.44 ;
    END
  END Data_COMP[224]
  PIN Data_COMP[223]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10276.345 187.44 10276.625 188.44 ;
    END
  END Data_COMP[223]
  PIN Data_COMP[222]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10278.025 187.44 10278.305 188.44 ;
    END
  END Data_COMP[222]
  PIN Data_COMP[221]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10233.225 187.44 10233.505 188.44 ;
    END
  END Data_COMP[221]
  PIN Data_COMP[220]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10234.905 187.44 10235.185 188.44 ;
    END
  END Data_COMP[220]
  PIN Data_COMP[219]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10236.025 187.44 10236.305 188.44 ;
    END
  END Data_COMP[219]
  PIN Data_COMP[218]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10278.585 187.44 10278.865 188.44 ;
    END
  END Data_COMP[218]
  PIN Data_COMP[217]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10274.665 187.44 10274.945 188.44 ;
    END
  END Data_COMP[217]
  PIN Data_COMP[216]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10274.105 187.44 10274.385 188.44 ;
    END
  END Data_COMP[216]
  PIN Data_COMP[215]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10276.905 187.44 10277.185 188.44 ;
    END
  END Data_COMP[215]
  PIN Data_COMP[214]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10234.345 187.44 10234.625 188.44 ;
    END
  END Data_COMP[214]
  PIN Data_COMP[213]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10237.145 187.44 10237.425 188.44 ;
    END
  END Data_COMP[213]
  PIN Data_COMP[212]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10236.585 187.44 10236.865 188.44 ;
    END
  END Data_COMP[212]
  PIN Data_COMP[211]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10232.665 187.44 10232.945 188.44 ;
    END
  END Data_COMP[211]
  PIN Data_COMP[210]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10232.105 187.44 10232.385 188.44 ;
    END
  END Data_COMP[210]
  PIN Data_COMP[209]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10205.785 187.44 10206.065 188.44 ;
    END
  END Data_COMP[209]
  PIN Data_COMP[208]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10207.465 187.44 10207.745 188.44 ;
    END
  END Data_COMP[208]
  PIN Data_COMP[207]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10209.145 187.44 10209.425 188.44 ;
    END
  END Data_COMP[207]
  PIN Data_COMP[206]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10149.785 187.44 10150.065 188.44 ;
    END
  END Data_COMP[206]
  PIN Data_COMP[205]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10152.025 187.44 10152.305 188.44 ;
    END
  END Data_COMP[205]
  PIN Data_COMP[204]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10153.705 187.44 10153.985 188.44 ;
    END
  END Data_COMP[204]
  PIN Data_COMP[203]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10205.225 187.44 10205.505 188.44 ;
    END
  END Data_COMP[203]
  PIN Data_COMP[202]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10206.345 187.44 10206.625 188.44 ;
    END
  END Data_COMP[202]
  PIN Data_COMP[201]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10208.025 187.44 10208.305 188.44 ;
    END
  END Data_COMP[201]
  PIN Data_COMP[200]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10151.465 187.44 10151.745 188.44 ;
    END
  END Data_COMP[200]
  PIN Data_COMP[199]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10153.145 187.44 10153.425 188.44 ;
    END
  END Data_COMP[199]
  PIN Data_COMP[198]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10154.265 187.44 10154.545 188.44 ;
    END
  END Data_COMP[198]
  PIN Data_COMP[197]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10208.585 187.44 10208.865 188.44 ;
    END
  END Data_COMP[197]
  PIN Data_COMP[196]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10204.665 187.44 10204.945 188.44 ;
    END
  END Data_COMP[196]
  PIN Data_COMP[195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10204.105 187.44 10204.385 188.44 ;
    END
  END Data_COMP[195]
  PIN Data_COMP[194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10206.905 187.44 10207.185 188.44 ;
    END
  END Data_COMP[194]
  PIN Data_COMP[193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10152.585 187.44 10152.865 188.44 ;
    END
  END Data_COMP[193]
  PIN Data_COMP[192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10155.385 187.44 10155.665 188.44 ;
    END
  END Data_COMP[192]
  PIN Data_COMP[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10154.825 187.44 10155.105 188.44 ;
    END
  END Data_COMP[191]
  PIN Data_COMP[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10150.905 187.44 10151.185 188.44 ;
    END
  END Data_COMP[190]
  PIN Data_COMP[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10150.345 187.44 10150.625 188.44 ;
    END
  END Data_COMP[189]
  PIN Data_COMP[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10101.065 187.44 10101.345 188.44 ;
    END
  END Data_COMP[188]
  PIN Data_COMP[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10128.225 187.44 10128.505 188.44 ;
    END
  END Data_COMP[187]
  PIN Data_COMP[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10129.905 187.44 10130.185 188.44 ;
    END
  END Data_COMP[186]
  PIN Data_COMP[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10071.385 187.44 10071.665 188.44 ;
    END
  END Data_COMP[185]
  PIN Data_COMP[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10073.625 187.44 10073.905 188.44 ;
    END
  END Data_COMP[184]
  PIN Data_COMP[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10075.305 187.44 10075.585 188.44 ;
    END
  END Data_COMP[183]
  PIN Data_COMP[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10100.505 187.44 10100.785 188.44 ;
    END
  END Data_COMP[182]
  PIN Data_COMP[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10101.625 187.44 10101.905 188.44 ;
    END
  END Data_COMP[181]
  PIN Data_COMP[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10128.785 187.44 10129.065 188.44 ;
    END
  END Data_COMP[180]
  PIN Data_COMP[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10073.065 187.44 10073.345 188.44 ;
    END
  END Data_COMP[179]
  PIN Data_COMP[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10074.745 187.44 10075.025 188.44 ;
    END
  END Data_COMP[178]
  PIN Data_COMP[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10088.745 187.44 10089.025 188.44 ;
    END
  END Data_COMP[177]
  PIN Data_COMP[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10129.345 187.44 10129.625 188.44 ;
    END
  END Data_COMP[176]
  PIN Data_COMP[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10099.945 187.44 10100.225 188.44 ;
    END
  END Data_COMP[175]
  PIN Data_COMP[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10099.385 187.44 10099.665 188.44 ;
    END
  END Data_COMP[174]
  PIN Data_COMP[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10127.665 187.44 10127.945 188.44 ;
    END
  END Data_COMP[173]
  PIN Data_COMP[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10074.185 187.44 10074.465 188.44 ;
    END
  END Data_COMP[172]
  PIN Data_COMP[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10089.865 187.44 10090.145 188.44 ;
    END
  END Data_COMP[171]
  PIN Data_COMP[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10089.305 187.44 10089.585 188.44 ;
    END
  END Data_COMP[170]
  PIN Data_COMP[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10072.505 187.44 10072.785 188.44 ;
    END
  END Data_COMP[169]
  PIN Data_COMP[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10071.945 187.44 10072.225 188.44 ;
    END
  END Data_COMP[168]
  PIN Data_COMP[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10018.745 187.44 10019.025 188.44 ;
    END
  END Data_COMP[167]
  PIN Data_COMP[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10020.425 187.44 10020.705 188.44 ;
    END
  END Data_COMP[166]
  PIN Data_COMP[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10022.105 187.44 10022.385 188.44 ;
    END
  END Data_COMP[165]
  PIN Data_COMP[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9993.545 187.44 9993.825 188.44 ;
    END
  END Data_COMP[164]
  PIN Data_COMP[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9995.785 187.44 9996.065 188.44 ;
    END
  END Data_COMP[163]
  PIN Data_COMP[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9997.465 187.44 9997.745 188.44 ;
    END
  END Data_COMP[162]
  PIN Data_COMP[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10018.185 187.44 10018.465 188.44 ;
    END
  END Data_COMP[161]
  PIN Data_COMP[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10019.305 187.44 10019.585 188.44 ;
    END
  END Data_COMP[160]
  PIN Data_COMP[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10020.985 187.44 10021.265 188.44 ;
    END
  END Data_COMP[159]
  PIN Data_COMP[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9995.225 187.44 9995.505 188.44 ;
    END
  END Data_COMP[158]
  PIN Data_COMP[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9996.905 187.44 9997.185 188.44 ;
    END
  END Data_COMP[157]
  PIN Data_COMP[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9998.025 187.44 9998.305 188.44 ;
    END
  END Data_COMP[156]
  PIN Data_COMP[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10021.545 187.44 10021.825 188.44 ;
    END
  END Data_COMP[155]
  PIN Data_COMP[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10017.625 187.44 10017.905 188.44 ;
    END
  END Data_COMP[154]
  PIN Data_COMP[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10017.065 187.44 10017.345 188.44 ;
    END
  END Data_COMP[153]
  PIN Data_COMP[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10019.865 187.44 10020.145 188.44 ;
    END
  END Data_COMP[152]
  PIN Data_COMP[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9996.345 187.44 9996.625 188.44 ;
    END
  END Data_COMP[151]
  PIN Data_COMP[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9999.145 187.44 9999.425 188.44 ;
    END
  END Data_COMP[150]
  PIN Data_COMP[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9998.585 187.44 9998.865 188.44 ;
    END
  END Data_COMP[149]
  PIN Data_COMP[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9994.665 187.44 9994.945 188.44 ;
    END
  END Data_COMP[148]
  PIN Data_COMP[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9994.105 187.44 9994.385 188.44 ;
    END
  END Data_COMP[147]
  PIN Data_COMP[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9952.665 187.44 9952.945 188.44 ;
    END
  END Data_COMP[146]
  PIN Data_COMP[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9954.345 187.44 9954.625 188.44 ;
    END
  END Data_COMP[145]
  PIN Data_COMP[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9956.025 187.44 9956.305 188.44 ;
    END
  END Data_COMP[144]
  PIN Data_COMP[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9922.425 187.44 9922.705 188.44 ;
    END
  END Data_COMP[143]
  PIN Data_COMP[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9924.665 187.44 9924.945 188.44 ;
    END
  END Data_COMP[142]
  PIN Data_COMP[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9926.345 187.44 9926.625 188.44 ;
    END
  END Data_COMP[141]
  PIN Data_COMP[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9952.105 187.44 9952.385 188.44 ;
    END
  END Data_COMP[140]
  PIN Data_COMP[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9953.225 187.44 9953.505 188.44 ;
    END
  END Data_COMP[139]
  PIN Data_COMP[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9954.905 187.44 9955.185 188.44 ;
    END
  END Data_COMP[138]
  PIN Data_COMP[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9924.105 187.44 9924.385 188.44 ;
    END
  END Data_COMP[137]
  PIN Data_COMP[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9925.785 187.44 9926.065 188.44 ;
    END
  END Data_COMP[136]
  PIN Data_COMP[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9926.905 187.44 9927.185 188.44 ;
    END
  END Data_COMP[135]
  PIN Data_COMP[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9955.465 187.44 9955.745 188.44 ;
    END
  END Data_COMP[134]
  PIN Data_COMP[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9951.545 187.44 9951.825 188.44 ;
    END
  END Data_COMP[133]
  PIN Data_COMP[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9950.985 187.44 9951.265 188.44 ;
    END
  END Data_COMP[132]
  PIN Data_COMP[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9953.785 187.44 9954.065 188.44 ;
    END
  END Data_COMP[131]
  PIN Data_COMP[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9925.225 187.44 9925.505 188.44 ;
    END
  END Data_COMP[130]
  PIN Data_COMP[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9928.025 187.44 9928.305 188.44 ;
    END
  END Data_COMP[129]
  PIN Data_COMP[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9927.465 187.44 9927.745 188.44 ;
    END
  END Data_COMP[128]
  PIN Data_COMP[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9923.545 187.44 9923.825 188.44 ;
    END
  END Data_COMP[127]
  PIN Data_COMP[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9922.985 187.44 9923.265 188.44 ;
    END
  END Data_COMP[126]
  PIN Data_COMP[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9870.905 187.44 9871.185 188.44 ;
    END
  END Data_COMP[125]
  PIN Data_COMP[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9872.585 187.44 9872.865 188.44 ;
    END
  END Data_COMP[124]
  PIN Data_COMP[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9874.265 187.44 9874.545 188.44 ;
    END
  END Data_COMP[123]
  PIN Data_COMP[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9818.265 187.44 9818.545 188.44 ;
    END
  END Data_COMP[122]
  PIN Data_COMP[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9820.505 187.44 9820.785 188.44 ;
    END
  END Data_COMP[121]
  PIN Data_COMP[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9847.665 187.44 9847.945 188.44 ;
    END
  END Data_COMP[120]
  PIN Data_COMP[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9870.345 187.44 9870.625 188.44 ;
    END
  END Data_COMP[119]
  PIN Data_COMP[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9871.465 187.44 9871.745 188.44 ;
    END
  END Data_COMP[118]
  PIN Data_COMP[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9873.145 187.44 9873.425 188.44 ;
    END
  END Data_COMP[117]
  PIN Data_COMP[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9819.945 187.44 9820.225 188.44 ;
    END
  END Data_COMP[116]
  PIN Data_COMP[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9847.105 187.44 9847.385 188.44 ;
    END
  END Data_COMP[115]
  PIN Data_COMP[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9848.225 187.44 9848.505 188.44 ;
    END
  END Data_COMP[114]
  PIN Data_COMP[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9873.705 187.44 9873.985 188.44 ;
    END
  END Data_COMP[113]
  PIN Data_COMP[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9869.785 187.44 9870.065 188.44 ;
    END
  END Data_COMP[112]
  PIN Data_COMP[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9860.825 187.44 9861.105 188.44 ;
    END
  END Data_COMP[111]
  PIN Data_COMP[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9872.025 187.44 9872.305 188.44 ;
    END
  END Data_COMP[110]
  PIN Data_COMP[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9821.065 187.44 9821.345 188.44 ;
    END
  END Data_COMP[109]
  PIN Data_COMP[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9849.345 187.44 9849.625 188.44 ;
    END
  END Data_COMP[108]
  PIN Data_COMP[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9848.785 187.44 9849.065 188.44 ;
    END
  END Data_COMP[107]
  PIN Data_COMP[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9819.385 187.44 9819.665 188.44 ;
    END
  END Data_COMP[106]
  PIN Data_COMP[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9818.825 187.44 9819.105 188.44 ;
    END
  END Data_COMP[105]
  PIN Data_COMP[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9792.505 187.44 9792.785 188.44 ;
    END
  END Data_COMP[104]
  PIN Data_COMP[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9794.185 187.44 9794.465 188.44 ;
    END
  END Data_COMP[103]
  PIN Data_COMP[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9808.745 187.44 9809.025 188.44 ;
    END
  END Data_COMP[102]
  PIN Data_COMP[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9737.065 187.44 9737.345 188.44 ;
    END
  END Data_COMP[101]
  PIN Data_COMP[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9739.305 187.44 9739.585 188.44 ;
    END
  END Data_COMP[100]
  PIN Data_COMP[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9740.985 187.44 9741.265 188.44 ;
    END
  END Data_COMP[99]
  PIN Data_COMP[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9791.945 187.44 9792.225 188.44 ;
    END
  END Data_COMP[98]
  PIN Data_COMP[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9793.065 187.44 9793.345 188.44 ;
    END
  END Data_COMP[97]
  PIN Data_COMP[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9794.745 187.44 9795.025 188.44 ;
    END
  END Data_COMP[96]
  PIN Data_COMP[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9738.745 187.44 9739.025 188.44 ;
    END
  END Data_COMP[95]
  PIN Data_COMP[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9740.425 187.44 9740.705 188.44 ;
    END
  END Data_COMP[94]
  PIN Data_COMP[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9741.545 187.44 9741.825 188.44 ;
    END
  END Data_COMP[93]
  PIN Data_COMP[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9808.185 187.44 9808.465 188.44 ;
    END
  END Data_COMP[92]
  PIN Data_COMP[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9791.385 187.44 9791.665 188.44 ;
    END
  END Data_COMP[91]
  PIN Data_COMP[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9790.825 187.44 9791.105 188.44 ;
    END
  END Data_COMP[90]
  PIN Data_COMP[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9793.625 187.44 9793.905 188.44 ;
    END
  END Data_COMP[89]
  PIN Data_COMP[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9739.865 187.44 9740.145 188.44 ;
    END
  END Data_COMP[88]
  PIN Data_COMP[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9742.665 187.44 9742.945 188.44 ;
    END
  END Data_COMP[87]
  PIN Data_COMP[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9742.105 187.44 9742.385 188.44 ;
    END
  END Data_COMP[86]
  PIN Data_COMP[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9738.185 187.44 9738.465 188.44 ;
    END
  END Data_COMP[85]
  PIN Data_COMP[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9737.625 187.44 9737.905 188.44 ;
    END
  END Data_COMP[84]
  PIN Data_COMP[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9715.785 187.44 9716.065 188.44 ;
    END
  END Data_COMP[83]
  PIN Data_COMP[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9717.465 187.44 9717.745 188.44 ;
    END
  END Data_COMP[82]
  PIN Data_COMP[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9719.145 187.44 9719.425 188.44 ;
    END
  END Data_COMP[81]
  PIN Data_COMP[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9671.545 187.44 9671.825 188.44 ;
    END
  END Data_COMP[80]
  PIN Data_COMP[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9673.785 187.44 9674.065 188.44 ;
    END
  END Data_COMP[79]
  PIN Data_COMP[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9675.465 187.44 9675.745 188.44 ;
    END
  END Data_COMP[78]
  PIN Data_COMP[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9715.225 187.44 9715.505 188.44 ;
    END
  END Data_COMP[77]
  PIN Data_COMP[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9716.345 187.44 9716.625 188.44 ;
    END
  END Data_COMP[76]
  PIN Data_COMP[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9718.025 187.44 9718.305 188.44 ;
    END
  END Data_COMP[75]
  PIN Data_COMP[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9673.225 187.44 9673.505 188.44 ;
    END
  END Data_COMP[74]
  PIN Data_COMP[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9674.905 187.44 9675.185 188.44 ;
    END
  END Data_COMP[73]
  PIN Data_COMP[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9676.025 187.44 9676.305 188.44 ;
    END
  END Data_COMP[72]
  PIN Data_COMP[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9718.585 187.44 9718.865 188.44 ;
    END
  END Data_COMP[71]
  PIN Data_COMP[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9714.665 187.44 9714.945 188.44 ;
    END
  END Data_COMP[70]
  PIN Data_COMP[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9714.105 187.44 9714.385 188.44 ;
    END
  END Data_COMP[69]
  PIN Data_COMP[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9716.905 187.44 9717.185 188.44 ;
    END
  END Data_COMP[68]
  PIN Data_COMP[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9674.345 187.44 9674.625 188.44 ;
    END
  END Data_COMP[67]
  PIN Data_COMP[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9677.145 187.44 9677.425 188.44 ;
    END
  END Data_COMP[66]
  PIN Data_COMP[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9676.585 187.44 9676.865 188.44 ;
    END
  END Data_COMP[65]
  PIN Data_COMP[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9672.665 187.44 9672.945 188.44 ;
    END
  END Data_COMP[64]
  PIN Data_COMP[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9672.105 187.44 9672.385 188.44 ;
    END
  END Data_COMP[63]
  PIN Data_COMP[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9645.785 187.44 9646.065 188.44 ;
    END
  END Data_COMP[62]
  PIN Data_COMP[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9647.465 187.44 9647.745 188.44 ;
    END
  END Data_COMP[61]
  PIN Data_COMP[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9649.145 187.44 9649.425 188.44 ;
    END
  END Data_COMP[60]
  PIN Data_COMP[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9589.785 187.44 9590.065 188.44 ;
    END
  END Data_COMP[59]
  PIN Data_COMP[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9592.025 187.44 9592.305 188.44 ;
    END
  END Data_COMP[58]
  PIN Data_COMP[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9593.705 187.44 9593.985 188.44 ;
    END
  END Data_COMP[57]
  PIN Data_COMP[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9645.225 187.44 9645.505 188.44 ;
    END
  END Data_COMP[56]
  PIN Data_COMP[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9646.345 187.44 9646.625 188.44 ;
    END
  END Data_COMP[55]
  PIN Data_COMP[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9648.025 187.44 9648.305 188.44 ;
    END
  END Data_COMP[54]
  PIN Data_COMP[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9591.465 187.44 9591.745 188.44 ;
    END
  END Data_COMP[53]
  PIN Data_COMP[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9593.145 187.44 9593.425 188.44 ;
    END
  END Data_COMP[52]
  PIN Data_COMP[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9594.265 187.44 9594.545 188.44 ;
    END
  END Data_COMP[51]
  PIN Data_COMP[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9648.585 187.44 9648.865 188.44 ;
    END
  END Data_COMP[50]
  PIN Data_COMP[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9644.665 187.44 9644.945 188.44 ;
    END
  END Data_COMP[49]
  PIN Data_COMP[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9644.105 187.44 9644.385 188.44 ;
    END
  END Data_COMP[48]
  PIN Data_COMP[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9646.905 187.44 9647.185 188.44 ;
    END
  END Data_COMP[47]
  PIN Data_COMP[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9592.585 187.44 9592.865 188.44 ;
    END
  END Data_COMP[46]
  PIN Data_COMP[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9595.385 187.44 9595.665 188.44 ;
    END
  END Data_COMP[45]
  PIN Data_COMP[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9594.825 187.44 9595.105 188.44 ;
    END
  END Data_COMP[44]
  PIN Data_COMP[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9590.905 187.44 9591.185 188.44 ;
    END
  END Data_COMP[43]
  PIN Data_COMP[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9590.345 187.44 9590.625 188.44 ;
    END
  END Data_COMP[42]
  PIN Data_COMP[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9541.065 187.44 9541.345 188.44 ;
    END
  END Data_COMP[41]
  PIN Data_COMP[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9568.225 187.44 9568.505 188.44 ;
    END
  END Data_COMP[40]
  PIN Data_COMP[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9569.905 187.44 9570.185 188.44 ;
    END
  END Data_COMP[39]
  PIN Data_COMP[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9511.385 187.44 9511.665 188.44 ;
    END
  END Data_COMP[38]
  PIN Data_COMP[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9513.625 187.44 9513.905 188.44 ;
    END
  END Data_COMP[37]
  PIN Data_COMP[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9515.305 187.44 9515.585 188.44 ;
    END
  END Data_COMP[36]
  PIN Data_COMP[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9540.505 187.44 9540.785 188.44 ;
    END
  END Data_COMP[35]
  PIN Data_COMP[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9541.625 187.44 9541.905 188.44 ;
    END
  END Data_COMP[34]
  PIN Data_COMP[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9568.785 187.44 9569.065 188.44 ;
    END
  END Data_COMP[33]
  PIN Data_COMP[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9513.065 187.44 9513.345 188.44 ;
    END
  END Data_COMP[32]
  PIN Data_COMP[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9514.745 187.44 9515.025 188.44 ;
    END
  END Data_COMP[31]
  PIN Data_COMP[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9528.745 187.44 9529.025 188.44 ;
    END
  END Data_COMP[30]
  PIN Data_COMP[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9569.345 187.44 9569.625 188.44 ;
    END
  END Data_COMP[29]
  PIN Data_COMP[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9539.945 187.44 9540.225 188.44 ;
    END
  END Data_COMP[28]
  PIN Data_COMP[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9539.385 187.44 9539.665 188.44 ;
    END
  END Data_COMP[27]
  PIN Data_COMP[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9567.665 187.44 9567.945 188.44 ;
    END
  END Data_COMP[26]
  PIN Data_COMP[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9514.185 187.44 9514.465 188.44 ;
    END
  END Data_COMP[25]
  PIN Data_COMP[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9529.865 187.44 9530.145 188.44 ;
    END
  END Data_COMP[24]
  PIN Data_COMP[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9529.305 187.44 9529.585 188.44 ;
    END
  END Data_COMP[23]
  PIN Data_COMP[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9512.505 187.44 9512.785 188.44 ;
    END
  END Data_COMP[22]
  PIN Data_COMP[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9511.945 187.44 9512.225 188.44 ;
    END
  END Data_COMP[21]
  PIN Data_COMP[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9458.745 187.44 9459.025 188.44 ;
    END
  END Data_COMP[20]
  PIN Data_COMP[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9460.425 187.44 9460.705 188.44 ;
    END
  END Data_COMP[19]
  PIN Data_COMP[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9462.105 187.44 9462.385 188.44 ;
    END
  END Data_COMP[18]
  PIN Data_COMP[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9433.545 187.44 9433.825 188.44 ;
    END
  END Data_COMP[17]
  PIN Data_COMP[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9435.785 187.44 9436.065 188.44 ;
    END
  END Data_COMP[16]
  PIN Data_COMP[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9437.465 187.44 9437.745 188.44 ;
    END
  END Data_COMP[15]
  PIN Data_COMP[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9458.185 187.44 9458.465 188.44 ;
    END
  END Data_COMP[14]
  PIN Data_COMP[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9459.305 187.44 9459.585 188.44 ;
    END
  END Data_COMP[13]
  PIN Data_COMP[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9460.985 187.44 9461.265 188.44 ;
    END
  END Data_COMP[12]
  PIN Data_COMP[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9435.225 187.44 9435.505 188.44 ;
    END
  END Data_COMP[11]
  PIN Data_COMP[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9436.905 187.44 9437.185 188.44 ;
    END
  END Data_COMP[10]
  PIN Data_COMP[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9438.025 187.44 9438.305 188.44 ;
    END
  END Data_COMP[9]
  PIN Data_COMP[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9461.545 187.44 9461.825 188.44 ;
    END
  END Data_COMP[8]
  PIN Data_COMP[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9457.625 187.44 9457.905 188.44 ;
    END
  END Data_COMP[7]
  PIN Data_COMP[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9457.065 187.44 9457.345 188.44 ;
    END
  END Data_COMP[6]
  PIN Data_COMP[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9459.865 187.44 9460.145 188.44 ;
    END
  END Data_COMP[5]
  PIN Data_COMP[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9436.345 187.44 9436.625 188.44 ;
    END
  END Data_COMP[4]
  PIN Data_COMP[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9439.145 187.44 9439.425 188.44 ;
    END
  END Data_COMP[3]
  PIN Data_COMP[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9438.585 187.44 9438.865 188.44 ;
    END
  END Data_COMP[2]
  PIN Data_COMP[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9434.665 187.44 9434.945 188.44 ;
    END
  END Data_COMP[1]
  PIN Data_COMP[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9434.105 187.44 9434.385 188.44 ;
    END
  END Data_COMP[0]
  PIN nTOK_PMOS[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9388.745 187.44 9389.025 188.44 ;
    END
  END nTOK_PMOS[55]
  PIN nTOK_PMOS[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9298.585 187.44 9298.865 188.44 ;
    END
  END nTOK_PMOS[54]
  PIN nTOK_PMOS[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9228.585 187.44 9228.865 188.44 ;
    END
  END nTOK_PMOS[53]
  PIN nTOK_PMOS[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9149.905 187.44 9150.185 188.44 ;
    END
  END nTOK_PMOS[52]
  PIN nTOK_PMOS[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9042.665 187.44 9042.945 188.44 ;
    END
  END nTOK_PMOS[51]
  PIN nTOK_PMOS[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8977.145 187.44 8977.425 188.44 ;
    END
  END nTOK_PMOS[50]
  PIN nTOK_PMOS[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8894.825 187.44 8895.105 188.44 ;
    END
  END nTOK_PMOS[49]
  PIN nTOK_PMOS[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8828.745 187.44 8829.025 188.44 ;
    END
  END nTOK_PMOS[48]
  PIN nTOK_PMOS[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8738.585 187.44 8738.865 188.44 ;
    END
  END nTOK_PMOS[47]
  PIN nTOK_PMOS[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8668.585 187.44 8668.865 188.44 ;
    END
  END nTOK_PMOS[46]
  PIN nTOK_PMOS[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8589.905 187.44 8590.185 188.44 ;
    END
  END nTOK_PMOS[45]
  PIN nTOK_PMOS[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8482.665 187.44 8482.945 188.44 ;
    END
  END nTOK_PMOS[44]
  PIN nTOK_PMOS[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8417.145 187.44 8417.425 188.44 ;
    END
  END nTOK_PMOS[43]
  PIN nTOK_PMOS[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8334.825 187.44 8335.105 188.44 ;
    END
  END nTOK_PMOS[42]
  PIN nTOK_PMOS[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8268.745 187.44 8269.025 188.44 ;
    END
  END nTOK_PMOS[41]
  PIN nTOK_PMOS[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8178.585 187.44 8178.865 188.44 ;
    END
  END nTOK_PMOS[40]
  PIN nTOK_PMOS[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8108.585 187.44 8108.865 188.44 ;
    END
  END nTOK_PMOS[39]
  PIN nTOK_PMOS[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8029.905 187.44 8030.185 188.44 ;
    END
  END nTOK_PMOS[38]
  PIN nTOK_PMOS[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7922.665 187.44 7922.945 188.44 ;
    END
  END nTOK_PMOS[37]
  PIN nTOK_PMOS[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7857.145 187.44 7857.425 188.44 ;
    END
  END nTOK_PMOS[36]
  PIN nTOK_PMOS[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7774.825 187.44 7775.105 188.44 ;
    END
  END nTOK_PMOS[35]
  PIN nTOK_PMOS[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7708.745 187.44 7709.025 188.44 ;
    END
  END nTOK_PMOS[34]
  PIN nTOK_PMOS[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7618.585 187.44 7618.865 188.44 ;
    END
  END nTOK_PMOS[33]
  PIN nTOK_PMOS[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7548.585 187.44 7548.865 188.44 ;
    END
  END nTOK_PMOS[32]
  PIN nTOK_PMOS[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7469.905 187.44 7470.185 188.44 ;
    END
  END nTOK_PMOS[31]
  PIN nTOK_PMOS[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7362.665 187.44 7362.945 188.44 ;
    END
  END nTOK_PMOS[30]
  PIN nTOK_PMOS[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7297.145 187.44 7297.425 188.44 ;
    END
  END nTOK_PMOS[29]
  PIN nTOK_PMOS[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7214.825 187.44 7215.105 188.44 ;
    END
  END nTOK_PMOS[28]
  PIN nTOK_PMOS[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7148.745 187.44 7149.025 188.44 ;
    END
  END nTOK_PMOS[27]
  PIN nTOK_PMOS[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7058.585 187.44 7058.865 188.44 ;
    END
  END nTOK_PMOS[26]
  PIN nTOK_PMOS[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6988.585 187.44 6988.865 188.44 ;
    END
  END nTOK_PMOS[25]
  PIN nTOK_PMOS[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6909.905 187.44 6910.185 188.44 ;
    END
  END nTOK_PMOS[24]
  PIN nTOK_PMOS[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6802.665 187.44 6802.945 188.44 ;
    END
  END nTOK_PMOS[23]
  PIN nTOK_PMOS[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6737.145 187.44 6737.425 188.44 ;
    END
  END nTOK_PMOS[22]
  PIN nTOK_PMOS[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6654.825 187.44 6655.105 188.44 ;
    END
  END nTOK_PMOS[21]
  PIN nTOK_PMOS[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6588.745 187.44 6589.025 188.44 ;
    END
  END nTOK_PMOS[20]
  PIN nTOK_PMOS[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6498.585 187.44 6498.865 188.44 ;
    END
  END nTOK_PMOS[19]
  PIN nTOK_PMOS[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6428.585 187.44 6428.865 188.44 ;
    END
  END nTOK_PMOS[18]
  PIN nTOK_PMOS[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6349.905 187.44 6350.185 188.44 ;
    END
  END nTOK_PMOS[17]
  PIN nTOK_PMOS[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6242.665 187.44 6242.945 188.44 ;
    END
  END nTOK_PMOS[16]
  PIN nTOK_PMOS[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6177.145 187.44 6177.425 188.44 ;
    END
  END nTOK_PMOS[15]
  PIN nTOK_PMOS[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6094.825 187.44 6095.105 188.44 ;
    END
  END nTOK_PMOS[14]
  PIN nTOK_PMOS[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6028.745 187.44 6029.025 188.44 ;
    END
  END nTOK_PMOS[13]
  PIN nTOK_PMOS[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5938.585 187.44 5938.865 188.44 ;
    END
  END nTOK_PMOS[12]
  PIN nTOK_PMOS[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5868.585 187.44 5868.865 188.44 ;
    END
  END nTOK_PMOS[11]
  PIN nTOK_PMOS[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5789.905 187.44 5790.185 188.44 ;
    END
  END nTOK_PMOS[10]
  PIN nTOK_PMOS[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5682.665 187.44 5682.945 188.44 ;
    END
  END nTOK_PMOS[9]
  PIN nTOK_PMOS[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5617.145 187.44 5617.425 188.44 ;
    END
  END nTOK_PMOS[8]
  PIN nTOK_PMOS[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5534.825 187.44 5535.105 188.44 ;
    END
  END nTOK_PMOS[7]
  PIN nTOK_PMOS[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5468.745 187.44 5469.025 188.44 ;
    END
  END nTOK_PMOS[6]
  PIN nTOK_PMOS[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5378.585 187.44 5378.865 188.44 ;
    END
  END nTOK_PMOS[5]
  PIN nTOK_PMOS[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5308.585 187.44 5308.865 188.44 ;
    END
  END nTOK_PMOS[4]
  PIN nTOK_PMOS[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5229.905 187.44 5230.185 188.44 ;
    END
  END nTOK_PMOS[3]
  PIN nTOK_PMOS[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5122.665 187.44 5122.945 188.44 ;
    END
  END nTOK_PMOS[2]
  PIN nTOK_PMOS[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5057.145 187.44 5057.425 188.44 ;
    END
  END nTOK_PMOS[1]
  PIN nTOK_PMOS[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4974.825 187.44 4975.105 188.44 ;
    END
  END nTOK_PMOS[0]
  PIN Data_HV[1175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18352.665 187.44 18352.945 188.44 ;
    END
  END Data_HV[1175]
  PIN Data_HV[1174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18354.345 187.44 18354.625 188.44 ;
    END
  END Data_HV[1174]
  PIN Data_HV[1173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18356.025 187.44 18356.305 188.44 ;
    END
  END Data_HV[1173]
  PIN Data_HV[1172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18322.425 187.44 18322.705 188.44 ;
    END
  END Data_HV[1172]
  PIN Data_HV[1171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18324.665 187.44 18324.945 188.44 ;
    END
  END Data_HV[1171]
  PIN Data_HV[1170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18326.345 187.44 18326.625 188.44 ;
    END
  END Data_HV[1170]
  PIN Data_HV[1169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18352.105 187.44 18352.385 188.44 ;
    END
  END Data_HV[1169]
  PIN Data_HV[1168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18353.225 187.44 18353.505 188.44 ;
    END
  END Data_HV[1168]
  PIN Data_HV[1167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18354.905 187.44 18355.185 188.44 ;
    END
  END Data_HV[1167]
  PIN Data_HV[1166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18324.105 187.44 18324.385 188.44 ;
    END
  END Data_HV[1166]
  PIN Data_HV[1165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18325.785 187.44 18326.065 188.44 ;
    END
  END Data_HV[1165]
  PIN Data_HV[1164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18326.905 187.44 18327.185 188.44 ;
    END
  END Data_HV[1164]
  PIN Data_HV[1163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18355.465 187.44 18355.745 188.44 ;
    END
  END Data_HV[1163]
  PIN Data_HV[1162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18351.545 187.44 18351.825 188.44 ;
    END
  END Data_HV[1162]
  PIN Data_HV[1161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18350.985 187.44 18351.265 188.44 ;
    END
  END Data_HV[1161]
  PIN Data_HV[1160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18353.785 187.44 18354.065 188.44 ;
    END
  END Data_HV[1160]
  PIN Data_HV[1159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18325.225 187.44 18325.505 188.44 ;
    END
  END Data_HV[1159]
  PIN Data_HV[1158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18328.025 187.44 18328.305 188.44 ;
    END
  END Data_HV[1158]
  PIN Data_HV[1157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18327.465 187.44 18327.745 188.44 ;
    END
  END Data_HV[1157]
  PIN Data_HV[1156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18323.545 187.44 18323.825 188.44 ;
    END
  END Data_HV[1156]
  PIN Data_HV[1155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18322.985 187.44 18323.265 188.44 ;
    END
  END Data_HV[1155]
  PIN Data_HV[1154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18270.905 187.44 18271.185 188.44 ;
    END
  END Data_HV[1154]
  PIN Data_HV[1153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18272.585 187.44 18272.865 188.44 ;
    END
  END Data_HV[1153]
  PIN Data_HV[1152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18274.265 187.44 18274.545 188.44 ;
    END
  END Data_HV[1152]
  PIN Data_HV[1151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18218.265 187.44 18218.545 188.44 ;
    END
  END Data_HV[1151]
  PIN Data_HV[1150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18220.505 187.44 18220.785 188.44 ;
    END
  END Data_HV[1150]
  PIN Data_HV[1149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18247.665 187.44 18247.945 188.44 ;
    END
  END Data_HV[1149]
  PIN Data_HV[1148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18270.345 187.44 18270.625 188.44 ;
    END
  END Data_HV[1148]
  PIN Data_HV[1147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18271.465 187.44 18271.745 188.44 ;
    END
  END Data_HV[1147]
  PIN Data_HV[1146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18273.145 187.44 18273.425 188.44 ;
    END
  END Data_HV[1146]
  PIN Data_HV[1145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18219.945 187.44 18220.225 188.44 ;
    END
  END Data_HV[1145]
  PIN Data_HV[1144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18247.105 187.44 18247.385 188.44 ;
    END
  END Data_HV[1144]
  PIN Data_HV[1143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18248.225 187.44 18248.505 188.44 ;
    END
  END Data_HV[1143]
  PIN Data_HV[1142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18273.705 187.44 18273.985 188.44 ;
    END
  END Data_HV[1142]
  PIN Data_HV[1141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18269.785 187.44 18270.065 188.44 ;
    END
  END Data_HV[1141]
  PIN Data_HV[1140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18260.825 187.44 18261.105 188.44 ;
    END
  END Data_HV[1140]
  PIN Data_HV[1139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18272.025 187.44 18272.305 188.44 ;
    END
  END Data_HV[1139]
  PIN Data_HV[1138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18221.065 187.44 18221.345 188.44 ;
    END
  END Data_HV[1138]
  PIN Data_HV[1137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18249.345 187.44 18249.625 188.44 ;
    END
  END Data_HV[1137]
  PIN Data_HV[1136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18248.785 187.44 18249.065 188.44 ;
    END
  END Data_HV[1136]
  PIN Data_HV[1135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18219.385 187.44 18219.665 188.44 ;
    END
  END Data_HV[1135]
  PIN Data_HV[1134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18218.825 187.44 18219.105 188.44 ;
    END
  END Data_HV[1134]
  PIN Data_HV[1133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18192.505 187.44 18192.785 188.44 ;
    END
  END Data_HV[1133]
  PIN Data_HV[1132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18194.185 187.44 18194.465 188.44 ;
    END
  END Data_HV[1132]
  PIN Data_HV[1131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18208.745 187.44 18209.025 188.44 ;
    END
  END Data_HV[1131]
  PIN Data_HV[1130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18137.065 187.44 18137.345 188.44 ;
    END
  END Data_HV[1130]
  PIN Data_HV[1129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18139.305 187.44 18139.585 188.44 ;
    END
  END Data_HV[1129]
  PIN Data_HV[1128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18140.985 187.44 18141.265 188.44 ;
    END
  END Data_HV[1128]
  PIN Data_HV[1127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18191.945 187.44 18192.225 188.44 ;
    END
  END Data_HV[1127]
  PIN Data_HV[1126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18193.065 187.44 18193.345 188.44 ;
    END
  END Data_HV[1126]
  PIN Data_HV[1125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18194.745 187.44 18195.025 188.44 ;
    END
  END Data_HV[1125]
  PIN Data_HV[1124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18138.745 187.44 18139.025 188.44 ;
    END
  END Data_HV[1124]
  PIN Data_HV[1123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18140.425 187.44 18140.705 188.44 ;
    END
  END Data_HV[1123]
  PIN Data_HV[1122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18141.545 187.44 18141.825 188.44 ;
    END
  END Data_HV[1122]
  PIN Data_HV[1121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18208.185 187.44 18208.465 188.44 ;
    END
  END Data_HV[1121]
  PIN Data_HV[1120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18191.385 187.44 18191.665 188.44 ;
    END
  END Data_HV[1120]
  PIN Data_HV[1119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18190.825 187.44 18191.105 188.44 ;
    END
  END Data_HV[1119]
  PIN Data_HV[1118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18193.625 187.44 18193.905 188.44 ;
    END
  END Data_HV[1118]
  PIN Data_HV[1117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18139.865 187.44 18140.145 188.44 ;
    END
  END Data_HV[1117]
  PIN Data_HV[1116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18142.665 187.44 18142.945 188.44 ;
    END
  END Data_HV[1116]
  PIN Data_HV[1115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18142.105 187.44 18142.385 188.44 ;
    END
  END Data_HV[1115]
  PIN Data_HV[1114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18138.185 187.44 18138.465 188.44 ;
    END
  END Data_HV[1114]
  PIN Data_HV[1113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18137.625 187.44 18137.905 188.44 ;
    END
  END Data_HV[1113]
  PIN Data_HV[1112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18115.785 187.44 18116.065 188.44 ;
    END
  END Data_HV[1112]
  PIN Data_HV[1111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18117.465 187.44 18117.745 188.44 ;
    END
  END Data_HV[1111]
  PIN Data_HV[1110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18119.145 187.44 18119.425 188.44 ;
    END
  END Data_HV[1110]
  PIN Data_HV[1109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18071.545 187.44 18071.825 188.44 ;
    END
  END Data_HV[1109]
  PIN Data_HV[1108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18073.785 187.44 18074.065 188.44 ;
    END
  END Data_HV[1108]
  PIN Data_HV[1107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18075.465 187.44 18075.745 188.44 ;
    END
  END Data_HV[1107]
  PIN Data_HV[1106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18115.225 187.44 18115.505 188.44 ;
    END
  END Data_HV[1106]
  PIN Data_HV[1105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18116.345 187.44 18116.625 188.44 ;
    END
  END Data_HV[1105]
  PIN Data_HV[1104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18118.025 187.44 18118.305 188.44 ;
    END
  END Data_HV[1104]
  PIN Data_HV[1103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18073.225 187.44 18073.505 188.44 ;
    END
  END Data_HV[1103]
  PIN Data_HV[1102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18074.905 187.44 18075.185 188.44 ;
    END
  END Data_HV[1102]
  PIN Data_HV[1101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18076.025 187.44 18076.305 188.44 ;
    END
  END Data_HV[1101]
  PIN Data_HV[1100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18118.585 187.44 18118.865 188.44 ;
    END
  END Data_HV[1100]
  PIN Data_HV[1099]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18114.665 187.44 18114.945 188.44 ;
    END
  END Data_HV[1099]
  PIN Data_HV[1098]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18114.105 187.44 18114.385 188.44 ;
    END
  END Data_HV[1098]
  PIN Data_HV[1097]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18116.905 187.44 18117.185 188.44 ;
    END
  END Data_HV[1097]
  PIN Data_HV[1096]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18074.345 187.44 18074.625 188.44 ;
    END
  END Data_HV[1096]
  PIN Data_HV[1095]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18077.145 187.44 18077.425 188.44 ;
    END
  END Data_HV[1095]
  PIN Data_HV[1094]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18076.585 187.44 18076.865 188.44 ;
    END
  END Data_HV[1094]
  PIN Data_HV[1093]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18072.665 187.44 18072.945 188.44 ;
    END
  END Data_HV[1093]
  PIN Data_HV[1092]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18072.105 187.44 18072.385 188.44 ;
    END
  END Data_HV[1092]
  PIN Data_HV[1091]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18045.785 187.44 18046.065 188.44 ;
    END
  END Data_HV[1091]
  PIN Data_HV[1090]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18047.465 187.44 18047.745 188.44 ;
    END
  END Data_HV[1090]
  PIN Data_HV[1089]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18049.145 187.44 18049.425 188.44 ;
    END
  END Data_HV[1089]
  PIN Data_HV[1088]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17989.785 187.44 17990.065 188.44 ;
    END
  END Data_HV[1088]
  PIN Data_HV[1087]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17992.025 187.44 17992.305 188.44 ;
    END
  END Data_HV[1087]
  PIN Data_HV[1086]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17993.705 187.44 17993.985 188.44 ;
    END
  END Data_HV[1086]
  PIN Data_HV[1085]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18045.225 187.44 18045.505 188.44 ;
    END
  END Data_HV[1085]
  PIN Data_HV[1084]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18046.345 187.44 18046.625 188.44 ;
    END
  END Data_HV[1084]
  PIN Data_HV[1083]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18048.025 187.44 18048.305 188.44 ;
    END
  END Data_HV[1083]
  PIN Data_HV[1082]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17991.465 187.44 17991.745 188.44 ;
    END
  END Data_HV[1082]
  PIN Data_HV[1081]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17993.145 187.44 17993.425 188.44 ;
    END
  END Data_HV[1081]
  PIN Data_HV[1080]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17994.265 187.44 17994.545 188.44 ;
    END
  END Data_HV[1080]
  PIN Data_HV[1079]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18048.585 187.44 18048.865 188.44 ;
    END
  END Data_HV[1079]
  PIN Data_HV[1078]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18044.665 187.44 18044.945 188.44 ;
    END
  END Data_HV[1078]
  PIN Data_HV[1077]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18044.105 187.44 18044.385 188.44 ;
    END
  END Data_HV[1077]
  PIN Data_HV[1076]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18046.905 187.44 18047.185 188.44 ;
    END
  END Data_HV[1076]
  PIN Data_HV[1075]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17992.585 187.44 17992.865 188.44 ;
    END
  END Data_HV[1075]
  PIN Data_HV[1074]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17995.385 187.44 17995.665 188.44 ;
    END
  END Data_HV[1074]
  PIN Data_HV[1073]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17994.825 187.44 17995.105 188.44 ;
    END
  END Data_HV[1073]
  PIN Data_HV[1072]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17990.905 187.44 17991.185 188.44 ;
    END
  END Data_HV[1072]
  PIN Data_HV[1071]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17990.345 187.44 17990.625 188.44 ;
    END
  END Data_HV[1071]
  PIN Data_HV[1070]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17941.065 187.44 17941.345 188.44 ;
    END
  END Data_HV[1070]
  PIN Data_HV[1069]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17968.225 187.44 17968.505 188.44 ;
    END
  END Data_HV[1069]
  PIN Data_HV[1068]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17969.905 187.44 17970.185 188.44 ;
    END
  END Data_HV[1068]
  PIN Data_HV[1067]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17911.385 187.44 17911.665 188.44 ;
    END
  END Data_HV[1067]
  PIN Data_HV[1066]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17913.625 187.44 17913.905 188.44 ;
    END
  END Data_HV[1066]
  PIN Data_HV[1065]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17915.305 187.44 17915.585 188.44 ;
    END
  END Data_HV[1065]
  PIN Data_HV[1064]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17940.505 187.44 17940.785 188.44 ;
    END
  END Data_HV[1064]
  PIN Data_HV[1063]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17941.625 187.44 17941.905 188.44 ;
    END
  END Data_HV[1063]
  PIN Data_HV[1062]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17968.785 187.44 17969.065 188.44 ;
    END
  END Data_HV[1062]
  PIN Data_HV[1061]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17913.065 187.44 17913.345 188.44 ;
    END
  END Data_HV[1061]
  PIN Data_HV[1060]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17914.745 187.44 17915.025 188.44 ;
    END
  END Data_HV[1060]
  PIN Data_HV[1059]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17928.745 187.44 17929.025 188.44 ;
    END
  END Data_HV[1059]
  PIN Data_HV[1058]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17969.345 187.44 17969.625 188.44 ;
    END
  END Data_HV[1058]
  PIN Data_HV[1057]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17939.945 187.44 17940.225 188.44 ;
    END
  END Data_HV[1057]
  PIN Data_HV[1056]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17939.385 187.44 17939.665 188.44 ;
    END
  END Data_HV[1056]
  PIN Data_HV[1055]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17967.665 187.44 17967.945 188.44 ;
    END
  END Data_HV[1055]
  PIN Data_HV[1054]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17914.185 187.44 17914.465 188.44 ;
    END
  END Data_HV[1054]
  PIN Data_HV[1053]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17929.865 187.44 17930.145 188.44 ;
    END
  END Data_HV[1053]
  PIN Data_HV[1052]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17929.305 187.44 17929.585 188.44 ;
    END
  END Data_HV[1052]
  PIN Data_HV[1051]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17912.505 187.44 17912.785 188.44 ;
    END
  END Data_HV[1051]
  PIN Data_HV[1050]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17911.945 187.44 17912.225 188.44 ;
    END
  END Data_HV[1050]
  PIN Data_HV[1049]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17858.745 187.44 17859.025 188.44 ;
    END
  END Data_HV[1049]
  PIN Data_HV[1048]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17860.425 187.44 17860.705 188.44 ;
    END
  END Data_HV[1048]
  PIN Data_HV[1047]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17862.105 187.44 17862.385 188.44 ;
    END
  END Data_HV[1047]
  PIN Data_HV[1046]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17833.545 187.44 17833.825 188.44 ;
    END
  END Data_HV[1046]
  PIN Data_HV[1045]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17835.785 187.44 17836.065 188.44 ;
    END
  END Data_HV[1045]
  PIN Data_HV[1044]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17837.465 187.44 17837.745 188.44 ;
    END
  END Data_HV[1044]
  PIN Data_HV[1043]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17858.185 187.44 17858.465 188.44 ;
    END
  END Data_HV[1043]
  PIN Data_HV[1042]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17859.305 187.44 17859.585 188.44 ;
    END
  END Data_HV[1042]
  PIN Data_HV[1041]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17860.985 187.44 17861.265 188.44 ;
    END
  END Data_HV[1041]
  PIN Data_HV[1040]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17835.225 187.44 17835.505 188.44 ;
    END
  END Data_HV[1040]
  PIN Data_HV[1039]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17836.905 187.44 17837.185 188.44 ;
    END
  END Data_HV[1039]
  PIN Data_HV[1038]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17838.025 187.44 17838.305 188.44 ;
    END
  END Data_HV[1038]
  PIN Data_HV[1037]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17861.545 187.44 17861.825 188.44 ;
    END
  END Data_HV[1037]
  PIN Data_HV[1036]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17857.625 187.44 17857.905 188.44 ;
    END
  END Data_HV[1036]
  PIN Data_HV[1035]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17857.065 187.44 17857.345 188.44 ;
    END
  END Data_HV[1035]
  PIN Data_HV[1034]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17859.865 187.44 17860.145 188.44 ;
    END
  END Data_HV[1034]
  PIN Data_HV[1033]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17836.345 187.44 17836.625 188.44 ;
    END
  END Data_HV[1033]
  PIN Data_HV[1032]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17839.145 187.44 17839.425 188.44 ;
    END
  END Data_HV[1032]
  PIN Data_HV[1031]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17838.585 187.44 17838.865 188.44 ;
    END
  END Data_HV[1031]
  PIN Data_HV[1030]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17834.665 187.44 17834.945 188.44 ;
    END
  END Data_HV[1030]
  PIN Data_HV[1029]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17834.105 187.44 17834.385 188.44 ;
    END
  END Data_HV[1029]
  PIN Data_HV[1028]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17792.665 187.44 17792.945 188.44 ;
    END
  END Data_HV[1028]
  PIN Data_HV[1027]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17794.345 187.44 17794.625 188.44 ;
    END
  END Data_HV[1027]
  PIN Data_HV[1026]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17796.025 187.44 17796.305 188.44 ;
    END
  END Data_HV[1026]
  PIN Data_HV[1025]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17762.425 187.44 17762.705 188.44 ;
    END
  END Data_HV[1025]
  PIN Data_HV[1024]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17764.665 187.44 17764.945 188.44 ;
    END
  END Data_HV[1024]
  PIN Data_HV[1023]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17766.345 187.44 17766.625 188.44 ;
    END
  END Data_HV[1023]
  PIN Data_HV[1022]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17792.105 187.44 17792.385 188.44 ;
    END
  END Data_HV[1022]
  PIN Data_HV[1021]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17793.225 187.44 17793.505 188.44 ;
    END
  END Data_HV[1021]
  PIN Data_HV[1020]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17794.905 187.44 17795.185 188.44 ;
    END
  END Data_HV[1020]
  PIN Data_HV[1019]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17764.105 187.44 17764.385 188.44 ;
    END
  END Data_HV[1019]
  PIN Data_HV[1018]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17765.785 187.44 17766.065 188.44 ;
    END
  END Data_HV[1018]
  PIN Data_HV[1017]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17766.905 187.44 17767.185 188.44 ;
    END
  END Data_HV[1017]
  PIN Data_HV[1016]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17795.465 187.44 17795.745 188.44 ;
    END
  END Data_HV[1016]
  PIN Data_HV[1015]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17791.545 187.44 17791.825 188.44 ;
    END
  END Data_HV[1015]
  PIN Data_HV[1014]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17790.985 187.44 17791.265 188.44 ;
    END
  END Data_HV[1014]
  PIN Data_HV[1013]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17793.785 187.44 17794.065 188.44 ;
    END
  END Data_HV[1013]
  PIN Data_HV[1012]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17765.225 187.44 17765.505 188.44 ;
    END
  END Data_HV[1012]
  PIN Data_HV[1011]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17768.025 187.44 17768.305 188.44 ;
    END
  END Data_HV[1011]
  PIN Data_HV[1010]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17767.465 187.44 17767.745 188.44 ;
    END
  END Data_HV[1010]
  PIN Data_HV[1009]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17763.545 187.44 17763.825 188.44 ;
    END
  END Data_HV[1009]
  PIN Data_HV[1008]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17762.985 187.44 17763.265 188.44 ;
    END
  END Data_HV[1008]
  PIN Data_HV[1007]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17710.905 187.44 17711.185 188.44 ;
    END
  END Data_HV[1007]
  PIN Data_HV[1006]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17712.585 187.44 17712.865 188.44 ;
    END
  END Data_HV[1006]
  PIN Data_HV[1005]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17714.265 187.44 17714.545 188.44 ;
    END
  END Data_HV[1005]
  PIN Data_HV[1004]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17658.265 187.44 17658.545 188.44 ;
    END
  END Data_HV[1004]
  PIN Data_HV[1003]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17660.505 187.44 17660.785 188.44 ;
    END
  END Data_HV[1003]
  PIN Data_HV[1002]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17687.665 187.44 17687.945 188.44 ;
    END
  END Data_HV[1002]
  PIN Data_HV[1001]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17710.345 187.44 17710.625 188.44 ;
    END
  END Data_HV[1001]
  PIN Data_HV[1000]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17711.465 187.44 17711.745 188.44 ;
    END
  END Data_HV[1000]
  PIN Data_HV[999]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17713.145 187.44 17713.425 188.44 ;
    END
  END Data_HV[999]
  PIN Data_HV[998]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17659.945 187.44 17660.225 188.44 ;
    END
  END Data_HV[998]
  PIN Data_HV[997]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17687.105 187.44 17687.385 188.44 ;
    END
  END Data_HV[997]
  PIN Data_HV[996]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17688.225 187.44 17688.505 188.44 ;
    END
  END Data_HV[996]
  PIN Data_HV[995]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17713.705 187.44 17713.985 188.44 ;
    END
  END Data_HV[995]
  PIN Data_HV[994]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17709.785 187.44 17710.065 188.44 ;
    END
  END Data_HV[994]
  PIN Data_HV[993]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17700.825 187.44 17701.105 188.44 ;
    END
  END Data_HV[993]
  PIN Data_HV[992]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17712.025 187.44 17712.305 188.44 ;
    END
  END Data_HV[992]
  PIN Data_HV[991]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17661.065 187.44 17661.345 188.44 ;
    END
  END Data_HV[991]
  PIN Data_HV[990]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17689.345 187.44 17689.625 188.44 ;
    END
  END Data_HV[990]
  PIN Data_HV[989]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17688.785 187.44 17689.065 188.44 ;
    END
  END Data_HV[989]
  PIN Data_HV[988]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17659.385 187.44 17659.665 188.44 ;
    END
  END Data_HV[988]
  PIN Data_HV[987]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17658.825 187.44 17659.105 188.44 ;
    END
  END Data_HV[987]
  PIN Data_HV[986]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17632.505 187.44 17632.785 188.44 ;
    END
  END Data_HV[986]
  PIN Data_HV[985]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17634.185 187.44 17634.465 188.44 ;
    END
  END Data_HV[985]
  PIN Data_HV[984]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17648.745 187.44 17649.025 188.44 ;
    END
  END Data_HV[984]
  PIN Data_HV[983]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17577.065 187.44 17577.345 188.44 ;
    END
  END Data_HV[983]
  PIN Data_HV[982]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17579.305 187.44 17579.585 188.44 ;
    END
  END Data_HV[982]
  PIN Data_HV[981]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17580.985 187.44 17581.265 188.44 ;
    END
  END Data_HV[981]
  PIN Data_HV[980]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17631.945 187.44 17632.225 188.44 ;
    END
  END Data_HV[980]
  PIN Data_HV[979]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17633.065 187.44 17633.345 188.44 ;
    END
  END Data_HV[979]
  PIN Data_HV[978]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17634.745 187.44 17635.025 188.44 ;
    END
  END Data_HV[978]
  PIN Data_HV[977]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17578.745 187.44 17579.025 188.44 ;
    END
  END Data_HV[977]
  PIN Data_HV[976]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17580.425 187.44 17580.705 188.44 ;
    END
  END Data_HV[976]
  PIN Data_HV[975]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17581.545 187.44 17581.825 188.44 ;
    END
  END Data_HV[975]
  PIN Data_HV[974]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17648.185 187.44 17648.465 188.44 ;
    END
  END Data_HV[974]
  PIN Data_HV[973]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17631.385 187.44 17631.665 188.44 ;
    END
  END Data_HV[973]
  PIN Data_HV[972]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17630.825 187.44 17631.105 188.44 ;
    END
  END Data_HV[972]
  PIN Data_HV[971]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17633.625 187.44 17633.905 188.44 ;
    END
  END Data_HV[971]
  PIN Data_HV[970]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17579.865 187.44 17580.145 188.44 ;
    END
  END Data_HV[970]
  PIN Data_HV[969]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17582.665 187.44 17582.945 188.44 ;
    END
  END Data_HV[969]
  PIN Data_HV[968]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17582.105 187.44 17582.385 188.44 ;
    END
  END Data_HV[968]
  PIN Data_HV[967]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17578.185 187.44 17578.465 188.44 ;
    END
  END Data_HV[967]
  PIN Data_HV[966]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17577.625 187.44 17577.905 188.44 ;
    END
  END Data_HV[966]
  PIN Data_HV[965]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17555.785 187.44 17556.065 188.44 ;
    END
  END Data_HV[965]
  PIN Data_HV[964]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17557.465 187.44 17557.745 188.44 ;
    END
  END Data_HV[964]
  PIN Data_HV[963]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17559.145 187.44 17559.425 188.44 ;
    END
  END Data_HV[963]
  PIN Data_HV[962]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17511.545 187.44 17511.825 188.44 ;
    END
  END Data_HV[962]
  PIN Data_HV[961]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17513.785 187.44 17514.065 188.44 ;
    END
  END Data_HV[961]
  PIN Data_HV[960]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17515.465 187.44 17515.745 188.44 ;
    END
  END Data_HV[960]
  PIN Data_HV[959]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17555.225 187.44 17555.505 188.44 ;
    END
  END Data_HV[959]
  PIN Data_HV[958]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17556.345 187.44 17556.625 188.44 ;
    END
  END Data_HV[958]
  PIN Data_HV[957]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17558.025 187.44 17558.305 188.44 ;
    END
  END Data_HV[957]
  PIN Data_HV[956]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17513.225 187.44 17513.505 188.44 ;
    END
  END Data_HV[956]
  PIN Data_HV[955]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17514.905 187.44 17515.185 188.44 ;
    END
  END Data_HV[955]
  PIN Data_HV[954]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17516.025 187.44 17516.305 188.44 ;
    END
  END Data_HV[954]
  PIN Data_HV[953]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17558.585 187.44 17558.865 188.44 ;
    END
  END Data_HV[953]
  PIN Data_HV[952]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17554.665 187.44 17554.945 188.44 ;
    END
  END Data_HV[952]
  PIN Data_HV[951]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17554.105 187.44 17554.385 188.44 ;
    END
  END Data_HV[951]
  PIN Data_HV[950]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17556.905 187.44 17557.185 188.44 ;
    END
  END Data_HV[950]
  PIN Data_HV[949]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17514.345 187.44 17514.625 188.44 ;
    END
  END Data_HV[949]
  PIN Data_HV[948]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17517.145 187.44 17517.425 188.44 ;
    END
  END Data_HV[948]
  PIN Data_HV[947]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17516.585 187.44 17516.865 188.44 ;
    END
  END Data_HV[947]
  PIN Data_HV[946]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17512.665 187.44 17512.945 188.44 ;
    END
  END Data_HV[946]
  PIN Data_HV[945]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17512.105 187.44 17512.385 188.44 ;
    END
  END Data_HV[945]
  PIN Data_HV[944]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17485.785 187.44 17486.065 188.44 ;
    END
  END Data_HV[944]
  PIN Data_HV[943]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17487.465 187.44 17487.745 188.44 ;
    END
  END Data_HV[943]
  PIN Data_HV[942]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17489.145 187.44 17489.425 188.44 ;
    END
  END Data_HV[942]
  PIN Data_HV[941]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17429.785 187.44 17430.065 188.44 ;
    END
  END Data_HV[941]
  PIN Data_HV[940]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17432.025 187.44 17432.305 188.44 ;
    END
  END Data_HV[940]
  PIN Data_HV[939]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17433.705 187.44 17433.985 188.44 ;
    END
  END Data_HV[939]
  PIN Data_HV[938]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17485.225 187.44 17485.505 188.44 ;
    END
  END Data_HV[938]
  PIN Data_HV[937]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17486.345 187.44 17486.625 188.44 ;
    END
  END Data_HV[937]
  PIN Data_HV[936]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17488.025 187.44 17488.305 188.44 ;
    END
  END Data_HV[936]
  PIN Data_HV[935]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17431.465 187.44 17431.745 188.44 ;
    END
  END Data_HV[935]
  PIN Data_HV[934]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17433.145 187.44 17433.425 188.44 ;
    END
  END Data_HV[934]
  PIN Data_HV[933]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17434.265 187.44 17434.545 188.44 ;
    END
  END Data_HV[933]
  PIN Data_HV[932]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17488.585 187.44 17488.865 188.44 ;
    END
  END Data_HV[932]
  PIN Data_HV[931]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17484.665 187.44 17484.945 188.44 ;
    END
  END Data_HV[931]
  PIN Data_HV[930]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17484.105 187.44 17484.385 188.44 ;
    END
  END Data_HV[930]
  PIN Data_HV[929]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17486.905 187.44 17487.185 188.44 ;
    END
  END Data_HV[929]
  PIN Data_HV[928]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17432.585 187.44 17432.865 188.44 ;
    END
  END Data_HV[928]
  PIN Data_HV[927]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17435.385 187.44 17435.665 188.44 ;
    END
  END Data_HV[927]
  PIN Data_HV[926]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17434.825 187.44 17435.105 188.44 ;
    END
  END Data_HV[926]
  PIN Data_HV[925]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17430.905 187.44 17431.185 188.44 ;
    END
  END Data_HV[925]
  PIN Data_HV[924]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17430.345 187.44 17430.625 188.44 ;
    END
  END Data_HV[924]
  PIN Data_HV[923]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17381.065 187.44 17381.345 188.44 ;
    END
  END Data_HV[923]
  PIN Data_HV[922]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17408.225 187.44 17408.505 188.44 ;
    END
  END Data_HV[922]
  PIN Data_HV[921]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17409.905 187.44 17410.185 188.44 ;
    END
  END Data_HV[921]
  PIN Data_HV[920]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17351.385 187.44 17351.665 188.44 ;
    END
  END Data_HV[920]
  PIN Data_HV[919]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17353.625 187.44 17353.905 188.44 ;
    END
  END Data_HV[919]
  PIN Data_HV[918]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17355.305 187.44 17355.585 188.44 ;
    END
  END Data_HV[918]
  PIN Data_HV[917]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17380.505 187.44 17380.785 188.44 ;
    END
  END Data_HV[917]
  PIN Data_HV[916]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17381.625 187.44 17381.905 188.44 ;
    END
  END Data_HV[916]
  PIN Data_HV[915]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17408.785 187.44 17409.065 188.44 ;
    END
  END Data_HV[915]
  PIN Data_HV[914]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17353.065 187.44 17353.345 188.44 ;
    END
  END Data_HV[914]
  PIN Data_HV[913]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17354.745 187.44 17355.025 188.44 ;
    END
  END Data_HV[913]
  PIN Data_HV[912]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17368.745 187.44 17369.025 188.44 ;
    END
  END Data_HV[912]
  PIN Data_HV[911]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17409.345 187.44 17409.625 188.44 ;
    END
  END Data_HV[911]
  PIN Data_HV[910]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17379.945 187.44 17380.225 188.44 ;
    END
  END Data_HV[910]
  PIN Data_HV[909]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17379.385 187.44 17379.665 188.44 ;
    END
  END Data_HV[909]
  PIN Data_HV[908]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17407.665 187.44 17407.945 188.44 ;
    END
  END Data_HV[908]
  PIN Data_HV[907]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17354.185 187.44 17354.465 188.44 ;
    END
  END Data_HV[907]
  PIN Data_HV[906]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17369.865 187.44 17370.145 188.44 ;
    END
  END Data_HV[906]
  PIN Data_HV[905]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17369.305 187.44 17369.585 188.44 ;
    END
  END Data_HV[905]
  PIN Data_HV[904]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17352.505 187.44 17352.785 188.44 ;
    END
  END Data_HV[904]
  PIN Data_HV[903]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17351.945 187.44 17352.225 188.44 ;
    END
  END Data_HV[903]
  PIN Data_HV[902]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17298.745 187.44 17299.025 188.44 ;
    END
  END Data_HV[902]
  PIN Data_HV[901]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17300.425 187.44 17300.705 188.44 ;
    END
  END Data_HV[901]
  PIN Data_HV[900]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17302.105 187.44 17302.385 188.44 ;
    END
  END Data_HV[900]
  PIN Data_HV[899]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17273.545 187.44 17273.825 188.44 ;
    END
  END Data_HV[899]
  PIN Data_HV[898]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17275.785 187.44 17276.065 188.44 ;
    END
  END Data_HV[898]
  PIN Data_HV[897]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17277.465 187.44 17277.745 188.44 ;
    END
  END Data_HV[897]
  PIN Data_HV[896]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17298.185 187.44 17298.465 188.44 ;
    END
  END Data_HV[896]
  PIN Data_HV[895]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17299.305 187.44 17299.585 188.44 ;
    END
  END Data_HV[895]
  PIN Data_HV[894]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17300.985 187.44 17301.265 188.44 ;
    END
  END Data_HV[894]
  PIN Data_HV[893]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17275.225 187.44 17275.505 188.44 ;
    END
  END Data_HV[893]
  PIN Data_HV[892]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17276.905 187.44 17277.185 188.44 ;
    END
  END Data_HV[892]
  PIN Data_HV[891]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17278.025 187.44 17278.305 188.44 ;
    END
  END Data_HV[891]
  PIN Data_HV[890]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17301.545 187.44 17301.825 188.44 ;
    END
  END Data_HV[890]
  PIN Data_HV[889]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17297.625 187.44 17297.905 188.44 ;
    END
  END Data_HV[889]
  PIN Data_HV[888]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17297.065 187.44 17297.345 188.44 ;
    END
  END Data_HV[888]
  PIN Data_HV[887]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17299.865 187.44 17300.145 188.44 ;
    END
  END Data_HV[887]
  PIN Data_HV[886]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17276.345 187.44 17276.625 188.44 ;
    END
  END Data_HV[886]
  PIN Data_HV[885]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17279.145 187.44 17279.425 188.44 ;
    END
  END Data_HV[885]
  PIN Data_HV[884]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17278.585 187.44 17278.865 188.44 ;
    END
  END Data_HV[884]
  PIN Data_HV[883]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17274.665 187.44 17274.945 188.44 ;
    END
  END Data_HV[883]
  PIN Data_HV[882]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17274.105 187.44 17274.385 188.44 ;
    END
  END Data_HV[882]
  PIN Data_HV[881]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17232.665 187.44 17232.945 188.44 ;
    END
  END Data_HV[881]
  PIN Data_HV[880]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17234.345 187.44 17234.625 188.44 ;
    END
  END Data_HV[880]
  PIN Data_HV[879]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17236.025 187.44 17236.305 188.44 ;
    END
  END Data_HV[879]
  PIN Data_HV[878]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17202.425 187.44 17202.705 188.44 ;
    END
  END Data_HV[878]
  PIN Data_HV[877]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17204.665 187.44 17204.945 188.44 ;
    END
  END Data_HV[877]
  PIN Data_HV[876]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17206.345 187.44 17206.625 188.44 ;
    END
  END Data_HV[876]
  PIN Data_HV[875]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17232.105 187.44 17232.385 188.44 ;
    END
  END Data_HV[875]
  PIN Data_HV[874]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17233.225 187.44 17233.505 188.44 ;
    END
  END Data_HV[874]
  PIN Data_HV[873]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17234.905 187.44 17235.185 188.44 ;
    END
  END Data_HV[873]
  PIN Data_HV[872]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17204.105 187.44 17204.385 188.44 ;
    END
  END Data_HV[872]
  PIN Data_HV[871]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17205.785 187.44 17206.065 188.44 ;
    END
  END Data_HV[871]
  PIN Data_HV[870]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17206.905 187.44 17207.185 188.44 ;
    END
  END Data_HV[870]
  PIN Data_HV[869]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17235.465 187.44 17235.745 188.44 ;
    END
  END Data_HV[869]
  PIN Data_HV[868]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17231.545 187.44 17231.825 188.44 ;
    END
  END Data_HV[868]
  PIN Data_HV[867]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17230.985 187.44 17231.265 188.44 ;
    END
  END Data_HV[867]
  PIN Data_HV[866]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17233.785 187.44 17234.065 188.44 ;
    END
  END Data_HV[866]
  PIN Data_HV[865]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17205.225 187.44 17205.505 188.44 ;
    END
  END Data_HV[865]
  PIN Data_HV[864]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17208.025 187.44 17208.305 188.44 ;
    END
  END Data_HV[864]
  PIN Data_HV[863]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17207.465 187.44 17207.745 188.44 ;
    END
  END Data_HV[863]
  PIN Data_HV[862]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17203.545 187.44 17203.825 188.44 ;
    END
  END Data_HV[862]
  PIN Data_HV[861]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17202.985 187.44 17203.265 188.44 ;
    END
  END Data_HV[861]
  PIN Data_HV[860]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17150.905 187.44 17151.185 188.44 ;
    END
  END Data_HV[860]
  PIN Data_HV[859]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17152.585 187.44 17152.865 188.44 ;
    END
  END Data_HV[859]
  PIN Data_HV[858]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17154.265 187.44 17154.545 188.44 ;
    END
  END Data_HV[858]
  PIN Data_HV[857]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17098.265 187.44 17098.545 188.44 ;
    END
  END Data_HV[857]
  PIN Data_HV[856]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17100.505 187.44 17100.785 188.44 ;
    END
  END Data_HV[856]
  PIN Data_HV[855]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17127.665 187.44 17127.945 188.44 ;
    END
  END Data_HV[855]
  PIN Data_HV[854]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17150.345 187.44 17150.625 188.44 ;
    END
  END Data_HV[854]
  PIN Data_HV[853]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17151.465 187.44 17151.745 188.44 ;
    END
  END Data_HV[853]
  PIN Data_HV[852]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17153.145 187.44 17153.425 188.44 ;
    END
  END Data_HV[852]
  PIN Data_HV[851]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17099.945 187.44 17100.225 188.44 ;
    END
  END Data_HV[851]
  PIN Data_HV[850]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17127.105 187.44 17127.385 188.44 ;
    END
  END Data_HV[850]
  PIN Data_HV[849]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17128.225 187.44 17128.505 188.44 ;
    END
  END Data_HV[849]
  PIN Data_HV[848]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17153.705 187.44 17153.985 188.44 ;
    END
  END Data_HV[848]
  PIN Data_HV[847]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17149.785 187.44 17150.065 188.44 ;
    END
  END Data_HV[847]
  PIN Data_HV[846]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17140.825 187.44 17141.105 188.44 ;
    END
  END Data_HV[846]
  PIN Data_HV[845]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17152.025 187.44 17152.305 188.44 ;
    END
  END Data_HV[845]
  PIN Data_HV[844]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17101.065 187.44 17101.345 188.44 ;
    END
  END Data_HV[844]
  PIN Data_HV[843]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17129.345 187.44 17129.625 188.44 ;
    END
  END Data_HV[843]
  PIN Data_HV[842]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17128.785 187.44 17129.065 188.44 ;
    END
  END Data_HV[842]
  PIN Data_HV[841]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17099.385 187.44 17099.665 188.44 ;
    END
  END Data_HV[841]
  PIN Data_HV[840]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17098.825 187.44 17099.105 188.44 ;
    END
  END Data_HV[840]
  PIN Data_HV[839]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17072.505 187.44 17072.785 188.44 ;
    END
  END Data_HV[839]
  PIN Data_HV[838]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17074.185 187.44 17074.465 188.44 ;
    END
  END Data_HV[838]
  PIN Data_HV[837]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17088.745 187.44 17089.025 188.44 ;
    END
  END Data_HV[837]
  PIN Data_HV[836]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17017.065 187.44 17017.345 188.44 ;
    END
  END Data_HV[836]
  PIN Data_HV[835]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17019.305 187.44 17019.585 188.44 ;
    END
  END Data_HV[835]
  PIN Data_HV[834]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17020.985 187.44 17021.265 188.44 ;
    END
  END Data_HV[834]
  PIN Data_HV[833]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17071.945 187.44 17072.225 188.44 ;
    END
  END Data_HV[833]
  PIN Data_HV[832]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17073.065 187.44 17073.345 188.44 ;
    END
  END Data_HV[832]
  PIN Data_HV[831]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17074.745 187.44 17075.025 188.44 ;
    END
  END Data_HV[831]
  PIN Data_HV[830]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17018.745 187.44 17019.025 188.44 ;
    END
  END Data_HV[830]
  PIN Data_HV[829]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17020.425 187.44 17020.705 188.44 ;
    END
  END Data_HV[829]
  PIN Data_HV[828]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17021.545 187.44 17021.825 188.44 ;
    END
  END Data_HV[828]
  PIN Data_HV[827]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17088.185 187.44 17088.465 188.44 ;
    END
  END Data_HV[827]
  PIN Data_HV[826]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17071.385 187.44 17071.665 188.44 ;
    END
  END Data_HV[826]
  PIN Data_HV[825]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17070.825 187.44 17071.105 188.44 ;
    END
  END Data_HV[825]
  PIN Data_HV[824]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17073.625 187.44 17073.905 188.44 ;
    END
  END Data_HV[824]
  PIN Data_HV[823]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17019.865 187.44 17020.145 188.44 ;
    END
  END Data_HV[823]
  PIN Data_HV[822]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17022.665 187.44 17022.945 188.44 ;
    END
  END Data_HV[822]
  PIN Data_HV[821]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17022.105 187.44 17022.385 188.44 ;
    END
  END Data_HV[821]
  PIN Data_HV[820]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17018.185 187.44 17018.465 188.44 ;
    END
  END Data_HV[820]
  PIN Data_HV[819]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17017.625 187.44 17017.905 188.44 ;
    END
  END Data_HV[819]
  PIN Data_HV[818]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16995.785 187.44 16996.065 188.44 ;
    END
  END Data_HV[818]
  PIN Data_HV[817]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16997.465 187.44 16997.745 188.44 ;
    END
  END Data_HV[817]
  PIN Data_HV[816]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16999.145 187.44 16999.425 188.44 ;
    END
  END Data_HV[816]
  PIN Data_HV[815]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16951.545 187.44 16951.825 188.44 ;
    END
  END Data_HV[815]
  PIN Data_HV[814]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16953.785 187.44 16954.065 188.44 ;
    END
  END Data_HV[814]
  PIN Data_HV[813]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16955.465 187.44 16955.745 188.44 ;
    END
  END Data_HV[813]
  PIN Data_HV[812]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16995.225 187.44 16995.505 188.44 ;
    END
  END Data_HV[812]
  PIN Data_HV[811]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16996.345 187.44 16996.625 188.44 ;
    END
  END Data_HV[811]
  PIN Data_HV[810]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16998.025 187.44 16998.305 188.44 ;
    END
  END Data_HV[810]
  PIN Data_HV[809]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16953.225 187.44 16953.505 188.44 ;
    END
  END Data_HV[809]
  PIN Data_HV[808]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16954.905 187.44 16955.185 188.44 ;
    END
  END Data_HV[808]
  PIN Data_HV[807]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16956.025 187.44 16956.305 188.44 ;
    END
  END Data_HV[807]
  PIN Data_HV[806]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16998.585 187.44 16998.865 188.44 ;
    END
  END Data_HV[806]
  PIN Data_HV[805]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16994.665 187.44 16994.945 188.44 ;
    END
  END Data_HV[805]
  PIN Data_HV[804]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16994.105 187.44 16994.385 188.44 ;
    END
  END Data_HV[804]
  PIN Data_HV[803]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16996.905 187.44 16997.185 188.44 ;
    END
  END Data_HV[803]
  PIN Data_HV[802]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16954.345 187.44 16954.625 188.44 ;
    END
  END Data_HV[802]
  PIN Data_HV[801]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16957.145 187.44 16957.425 188.44 ;
    END
  END Data_HV[801]
  PIN Data_HV[800]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16956.585 187.44 16956.865 188.44 ;
    END
  END Data_HV[800]
  PIN Data_HV[799]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16952.665 187.44 16952.945 188.44 ;
    END
  END Data_HV[799]
  PIN Data_HV[798]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16952.105 187.44 16952.385 188.44 ;
    END
  END Data_HV[798]
  PIN Data_HV[797]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16925.785 187.44 16926.065 188.44 ;
    END
  END Data_HV[797]
  PIN Data_HV[796]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16927.465 187.44 16927.745 188.44 ;
    END
  END Data_HV[796]
  PIN Data_HV[795]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16929.145 187.44 16929.425 188.44 ;
    END
  END Data_HV[795]
  PIN Data_HV[794]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16869.785 187.44 16870.065 188.44 ;
    END
  END Data_HV[794]
  PIN Data_HV[793]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16872.025 187.44 16872.305 188.44 ;
    END
  END Data_HV[793]
  PIN Data_HV[792]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16873.705 187.44 16873.985 188.44 ;
    END
  END Data_HV[792]
  PIN Data_HV[791]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16925.225 187.44 16925.505 188.44 ;
    END
  END Data_HV[791]
  PIN Data_HV[790]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16926.345 187.44 16926.625 188.44 ;
    END
  END Data_HV[790]
  PIN Data_HV[789]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16928.025 187.44 16928.305 188.44 ;
    END
  END Data_HV[789]
  PIN Data_HV[788]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16871.465 187.44 16871.745 188.44 ;
    END
  END Data_HV[788]
  PIN Data_HV[787]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16873.145 187.44 16873.425 188.44 ;
    END
  END Data_HV[787]
  PIN Data_HV[786]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16874.265 187.44 16874.545 188.44 ;
    END
  END Data_HV[786]
  PIN Data_HV[785]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16928.585 187.44 16928.865 188.44 ;
    END
  END Data_HV[785]
  PIN Data_HV[784]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16924.665 187.44 16924.945 188.44 ;
    END
  END Data_HV[784]
  PIN Data_HV[783]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16924.105 187.44 16924.385 188.44 ;
    END
  END Data_HV[783]
  PIN Data_HV[782]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16926.905 187.44 16927.185 188.44 ;
    END
  END Data_HV[782]
  PIN Data_HV[781]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16872.585 187.44 16872.865 188.44 ;
    END
  END Data_HV[781]
  PIN Data_HV[780]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16875.385 187.44 16875.665 188.44 ;
    END
  END Data_HV[780]
  PIN Data_HV[779]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16874.825 187.44 16875.105 188.44 ;
    END
  END Data_HV[779]
  PIN Data_HV[778]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16870.905 187.44 16871.185 188.44 ;
    END
  END Data_HV[778]
  PIN Data_HV[777]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16870.345 187.44 16870.625 188.44 ;
    END
  END Data_HV[777]
  PIN Data_HV[776]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16821.065 187.44 16821.345 188.44 ;
    END
  END Data_HV[776]
  PIN Data_HV[775]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16848.225 187.44 16848.505 188.44 ;
    END
  END Data_HV[775]
  PIN Data_HV[774]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16849.905 187.44 16850.185 188.44 ;
    END
  END Data_HV[774]
  PIN Data_HV[773]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16791.385 187.44 16791.665 188.44 ;
    END
  END Data_HV[773]
  PIN Data_HV[772]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16793.625 187.44 16793.905 188.44 ;
    END
  END Data_HV[772]
  PIN Data_HV[771]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16795.305 187.44 16795.585 188.44 ;
    END
  END Data_HV[771]
  PIN Data_HV[770]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16820.505 187.44 16820.785 188.44 ;
    END
  END Data_HV[770]
  PIN Data_HV[769]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16821.625 187.44 16821.905 188.44 ;
    END
  END Data_HV[769]
  PIN Data_HV[768]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16848.785 187.44 16849.065 188.44 ;
    END
  END Data_HV[768]
  PIN Data_HV[767]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16793.065 187.44 16793.345 188.44 ;
    END
  END Data_HV[767]
  PIN Data_HV[766]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16794.745 187.44 16795.025 188.44 ;
    END
  END Data_HV[766]
  PIN Data_HV[765]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16808.745 187.44 16809.025 188.44 ;
    END
  END Data_HV[765]
  PIN Data_HV[764]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16849.345 187.44 16849.625 188.44 ;
    END
  END Data_HV[764]
  PIN Data_HV[763]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16819.945 187.44 16820.225 188.44 ;
    END
  END Data_HV[763]
  PIN Data_HV[762]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16819.385 187.44 16819.665 188.44 ;
    END
  END Data_HV[762]
  PIN Data_HV[761]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16847.665 187.44 16847.945 188.44 ;
    END
  END Data_HV[761]
  PIN Data_HV[760]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16794.185 187.44 16794.465 188.44 ;
    END
  END Data_HV[760]
  PIN Data_HV[759]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16809.865 187.44 16810.145 188.44 ;
    END
  END Data_HV[759]
  PIN Data_HV[758]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16809.305 187.44 16809.585 188.44 ;
    END
  END Data_HV[758]
  PIN Data_HV[757]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16792.505 187.44 16792.785 188.44 ;
    END
  END Data_HV[757]
  PIN Data_HV[756]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16791.945 187.44 16792.225 188.44 ;
    END
  END Data_HV[756]
  PIN Data_HV[755]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16738.745 187.44 16739.025 188.44 ;
    END
  END Data_HV[755]
  PIN Data_HV[754]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16740.425 187.44 16740.705 188.44 ;
    END
  END Data_HV[754]
  PIN Data_HV[753]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16742.105 187.44 16742.385 188.44 ;
    END
  END Data_HV[753]
  PIN Data_HV[752]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16713.545 187.44 16713.825 188.44 ;
    END
  END Data_HV[752]
  PIN Data_HV[751]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16715.785 187.44 16716.065 188.44 ;
    END
  END Data_HV[751]
  PIN Data_HV[750]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16717.465 187.44 16717.745 188.44 ;
    END
  END Data_HV[750]
  PIN Data_HV[749]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16738.185 187.44 16738.465 188.44 ;
    END
  END Data_HV[749]
  PIN Data_HV[748]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16739.305 187.44 16739.585 188.44 ;
    END
  END Data_HV[748]
  PIN Data_HV[747]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16740.985 187.44 16741.265 188.44 ;
    END
  END Data_HV[747]
  PIN Data_HV[746]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16715.225 187.44 16715.505 188.44 ;
    END
  END Data_HV[746]
  PIN Data_HV[745]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16716.905 187.44 16717.185 188.44 ;
    END
  END Data_HV[745]
  PIN Data_HV[744]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16718.025 187.44 16718.305 188.44 ;
    END
  END Data_HV[744]
  PIN Data_HV[743]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16741.545 187.44 16741.825 188.44 ;
    END
  END Data_HV[743]
  PIN Data_HV[742]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16737.625 187.44 16737.905 188.44 ;
    END
  END Data_HV[742]
  PIN Data_HV[741]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16737.065 187.44 16737.345 188.44 ;
    END
  END Data_HV[741]
  PIN Data_HV[740]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16739.865 187.44 16740.145 188.44 ;
    END
  END Data_HV[740]
  PIN Data_HV[739]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16716.345 187.44 16716.625 188.44 ;
    END
  END Data_HV[739]
  PIN Data_HV[738]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16719.145 187.44 16719.425 188.44 ;
    END
  END Data_HV[738]
  PIN Data_HV[737]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16718.585 187.44 16718.865 188.44 ;
    END
  END Data_HV[737]
  PIN Data_HV[736]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16714.665 187.44 16714.945 188.44 ;
    END
  END Data_HV[736]
  PIN Data_HV[735]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16714.105 187.44 16714.385 188.44 ;
    END
  END Data_HV[735]
  PIN Data_HV[734]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16672.665 187.44 16672.945 188.44 ;
    END
  END Data_HV[734]
  PIN Data_HV[733]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16674.345 187.44 16674.625 188.44 ;
    END
  END Data_HV[733]
  PIN Data_HV[732]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16676.025 187.44 16676.305 188.44 ;
    END
  END Data_HV[732]
  PIN Data_HV[731]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16642.425 187.44 16642.705 188.44 ;
    END
  END Data_HV[731]
  PIN Data_HV[730]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16644.665 187.44 16644.945 188.44 ;
    END
  END Data_HV[730]
  PIN Data_HV[729]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16646.345 187.44 16646.625 188.44 ;
    END
  END Data_HV[729]
  PIN Data_HV[728]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16672.105 187.44 16672.385 188.44 ;
    END
  END Data_HV[728]
  PIN Data_HV[727]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16673.225 187.44 16673.505 188.44 ;
    END
  END Data_HV[727]
  PIN Data_HV[726]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16674.905 187.44 16675.185 188.44 ;
    END
  END Data_HV[726]
  PIN Data_HV[725]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16644.105 187.44 16644.385 188.44 ;
    END
  END Data_HV[725]
  PIN Data_HV[724]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16645.785 187.44 16646.065 188.44 ;
    END
  END Data_HV[724]
  PIN Data_HV[723]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16646.905 187.44 16647.185 188.44 ;
    END
  END Data_HV[723]
  PIN Data_HV[722]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16675.465 187.44 16675.745 188.44 ;
    END
  END Data_HV[722]
  PIN Data_HV[721]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16671.545 187.44 16671.825 188.44 ;
    END
  END Data_HV[721]
  PIN Data_HV[720]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16670.985 187.44 16671.265 188.44 ;
    END
  END Data_HV[720]
  PIN Data_HV[719]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16673.785 187.44 16674.065 188.44 ;
    END
  END Data_HV[719]
  PIN Data_HV[718]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16645.225 187.44 16645.505 188.44 ;
    END
  END Data_HV[718]
  PIN Data_HV[717]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16648.025 187.44 16648.305 188.44 ;
    END
  END Data_HV[717]
  PIN Data_HV[716]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16647.465 187.44 16647.745 188.44 ;
    END
  END Data_HV[716]
  PIN Data_HV[715]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16643.545 187.44 16643.825 188.44 ;
    END
  END Data_HV[715]
  PIN Data_HV[714]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16642.985 187.44 16643.265 188.44 ;
    END
  END Data_HV[714]
  PIN Data_HV[713]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16590.905 187.44 16591.185 188.44 ;
    END
  END Data_HV[713]
  PIN Data_HV[712]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16592.585 187.44 16592.865 188.44 ;
    END
  END Data_HV[712]
  PIN Data_HV[711]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16594.265 187.44 16594.545 188.44 ;
    END
  END Data_HV[711]
  PIN Data_HV[710]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16538.265 187.44 16538.545 188.44 ;
    END
  END Data_HV[710]
  PIN Data_HV[709]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16540.505 187.44 16540.785 188.44 ;
    END
  END Data_HV[709]
  PIN Data_HV[708]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16567.665 187.44 16567.945 188.44 ;
    END
  END Data_HV[708]
  PIN Data_HV[707]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16590.345 187.44 16590.625 188.44 ;
    END
  END Data_HV[707]
  PIN Data_HV[706]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16591.465 187.44 16591.745 188.44 ;
    END
  END Data_HV[706]
  PIN Data_HV[705]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16593.145 187.44 16593.425 188.44 ;
    END
  END Data_HV[705]
  PIN Data_HV[704]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16539.945 187.44 16540.225 188.44 ;
    END
  END Data_HV[704]
  PIN Data_HV[703]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16567.105 187.44 16567.385 188.44 ;
    END
  END Data_HV[703]
  PIN Data_HV[702]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16568.225 187.44 16568.505 188.44 ;
    END
  END Data_HV[702]
  PIN Data_HV[701]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16593.705 187.44 16593.985 188.44 ;
    END
  END Data_HV[701]
  PIN Data_HV[700]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16589.785 187.44 16590.065 188.44 ;
    END
  END Data_HV[700]
  PIN Data_HV[699]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16580.825 187.44 16581.105 188.44 ;
    END
  END Data_HV[699]
  PIN Data_HV[698]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16592.025 187.44 16592.305 188.44 ;
    END
  END Data_HV[698]
  PIN Data_HV[697]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16541.065 187.44 16541.345 188.44 ;
    END
  END Data_HV[697]
  PIN Data_HV[696]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16569.345 187.44 16569.625 188.44 ;
    END
  END Data_HV[696]
  PIN Data_HV[695]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16568.785 187.44 16569.065 188.44 ;
    END
  END Data_HV[695]
  PIN Data_HV[694]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16539.385 187.44 16539.665 188.44 ;
    END
  END Data_HV[694]
  PIN Data_HV[693]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16538.825 187.44 16539.105 188.44 ;
    END
  END Data_HV[693]
  PIN Data_HV[692]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16512.505 187.44 16512.785 188.44 ;
    END
  END Data_HV[692]
  PIN Data_HV[691]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16514.185 187.44 16514.465 188.44 ;
    END
  END Data_HV[691]
  PIN Data_HV[690]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16528.745 187.44 16529.025 188.44 ;
    END
  END Data_HV[690]
  PIN Data_HV[689]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16457.065 187.44 16457.345 188.44 ;
    END
  END Data_HV[689]
  PIN Data_HV[688]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16459.305 187.44 16459.585 188.44 ;
    END
  END Data_HV[688]
  PIN Data_HV[687]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16460.985 187.44 16461.265 188.44 ;
    END
  END Data_HV[687]
  PIN Data_HV[686]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16511.945 187.44 16512.225 188.44 ;
    END
  END Data_HV[686]
  PIN Data_HV[685]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16513.065 187.44 16513.345 188.44 ;
    END
  END Data_HV[685]
  PIN Data_HV[684]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16514.745 187.44 16515.025 188.44 ;
    END
  END Data_HV[684]
  PIN Data_HV[683]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16458.745 187.44 16459.025 188.44 ;
    END
  END Data_HV[683]
  PIN Data_HV[682]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16460.425 187.44 16460.705 188.44 ;
    END
  END Data_HV[682]
  PIN Data_HV[681]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16461.545 187.44 16461.825 188.44 ;
    END
  END Data_HV[681]
  PIN Data_HV[680]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16528.185 187.44 16528.465 188.44 ;
    END
  END Data_HV[680]
  PIN Data_HV[679]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16511.385 187.44 16511.665 188.44 ;
    END
  END Data_HV[679]
  PIN Data_HV[678]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16510.825 187.44 16511.105 188.44 ;
    END
  END Data_HV[678]
  PIN Data_HV[677]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16513.625 187.44 16513.905 188.44 ;
    END
  END Data_HV[677]
  PIN Data_HV[676]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16459.865 187.44 16460.145 188.44 ;
    END
  END Data_HV[676]
  PIN Data_HV[675]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16462.665 187.44 16462.945 188.44 ;
    END
  END Data_HV[675]
  PIN Data_HV[674]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16462.105 187.44 16462.385 188.44 ;
    END
  END Data_HV[674]
  PIN Data_HV[673]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16458.185 187.44 16458.465 188.44 ;
    END
  END Data_HV[673]
  PIN Data_HV[672]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16457.625 187.44 16457.905 188.44 ;
    END
  END Data_HV[672]
  PIN Data_HV[671]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16435.785 187.44 16436.065 188.44 ;
    END
  END Data_HV[671]
  PIN Data_HV[670]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16437.465 187.44 16437.745 188.44 ;
    END
  END Data_HV[670]
  PIN Data_HV[669]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16439.145 187.44 16439.425 188.44 ;
    END
  END Data_HV[669]
  PIN Data_HV[668]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16391.545 187.44 16391.825 188.44 ;
    END
  END Data_HV[668]
  PIN Data_HV[667]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16393.785 187.44 16394.065 188.44 ;
    END
  END Data_HV[667]
  PIN Data_HV[666]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16395.465 187.44 16395.745 188.44 ;
    END
  END Data_HV[666]
  PIN Data_HV[665]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16435.225 187.44 16435.505 188.44 ;
    END
  END Data_HV[665]
  PIN Data_HV[664]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16436.345 187.44 16436.625 188.44 ;
    END
  END Data_HV[664]
  PIN Data_HV[663]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16438.025 187.44 16438.305 188.44 ;
    END
  END Data_HV[663]
  PIN Data_HV[662]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16393.225 187.44 16393.505 188.44 ;
    END
  END Data_HV[662]
  PIN Data_HV[661]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16394.905 187.44 16395.185 188.44 ;
    END
  END Data_HV[661]
  PIN Data_HV[660]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16396.025 187.44 16396.305 188.44 ;
    END
  END Data_HV[660]
  PIN Data_HV[659]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16438.585 187.44 16438.865 188.44 ;
    END
  END Data_HV[659]
  PIN Data_HV[658]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16434.665 187.44 16434.945 188.44 ;
    END
  END Data_HV[658]
  PIN Data_HV[657]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16434.105 187.44 16434.385 188.44 ;
    END
  END Data_HV[657]
  PIN Data_HV[656]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16436.905 187.44 16437.185 188.44 ;
    END
  END Data_HV[656]
  PIN Data_HV[655]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16394.345 187.44 16394.625 188.44 ;
    END
  END Data_HV[655]
  PIN Data_HV[654]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16397.145 187.44 16397.425 188.44 ;
    END
  END Data_HV[654]
  PIN Data_HV[653]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16396.585 187.44 16396.865 188.44 ;
    END
  END Data_HV[653]
  PIN Data_HV[652]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16392.665 187.44 16392.945 188.44 ;
    END
  END Data_HV[652]
  PIN Data_HV[651]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16392.105 187.44 16392.385 188.44 ;
    END
  END Data_HV[651]
  PIN Data_HV[650]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16365.785 187.44 16366.065 188.44 ;
    END
  END Data_HV[650]
  PIN Data_HV[649]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16367.465 187.44 16367.745 188.44 ;
    END
  END Data_HV[649]
  PIN Data_HV[648]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16369.145 187.44 16369.425 188.44 ;
    END
  END Data_HV[648]
  PIN Data_HV[647]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16309.785 187.44 16310.065 188.44 ;
    END
  END Data_HV[647]
  PIN Data_HV[646]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16312.025 187.44 16312.305 188.44 ;
    END
  END Data_HV[646]
  PIN Data_HV[645]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16313.705 187.44 16313.985 188.44 ;
    END
  END Data_HV[645]
  PIN Data_HV[644]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16365.225 187.44 16365.505 188.44 ;
    END
  END Data_HV[644]
  PIN Data_HV[643]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16366.345 187.44 16366.625 188.44 ;
    END
  END Data_HV[643]
  PIN Data_HV[642]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16368.025 187.44 16368.305 188.44 ;
    END
  END Data_HV[642]
  PIN Data_HV[641]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16311.465 187.44 16311.745 188.44 ;
    END
  END Data_HV[641]
  PIN Data_HV[640]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16313.145 187.44 16313.425 188.44 ;
    END
  END Data_HV[640]
  PIN Data_HV[639]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16314.265 187.44 16314.545 188.44 ;
    END
  END Data_HV[639]
  PIN Data_HV[638]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16368.585 187.44 16368.865 188.44 ;
    END
  END Data_HV[638]
  PIN Data_HV[637]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16364.665 187.44 16364.945 188.44 ;
    END
  END Data_HV[637]
  PIN Data_HV[636]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16364.105 187.44 16364.385 188.44 ;
    END
  END Data_HV[636]
  PIN Data_HV[635]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16366.905 187.44 16367.185 188.44 ;
    END
  END Data_HV[635]
  PIN Data_HV[634]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16312.585 187.44 16312.865 188.44 ;
    END
  END Data_HV[634]
  PIN Data_HV[633]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16315.385 187.44 16315.665 188.44 ;
    END
  END Data_HV[633]
  PIN Data_HV[632]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16314.825 187.44 16315.105 188.44 ;
    END
  END Data_HV[632]
  PIN Data_HV[631]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16310.905 187.44 16311.185 188.44 ;
    END
  END Data_HV[631]
  PIN Data_HV[630]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16310.345 187.44 16310.625 188.44 ;
    END
  END Data_HV[630]
  PIN Data_HV[629]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16261.065 187.44 16261.345 188.44 ;
    END
  END Data_HV[629]
  PIN Data_HV[628]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16288.225 187.44 16288.505 188.44 ;
    END
  END Data_HV[628]
  PIN Data_HV[627]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16289.905 187.44 16290.185 188.44 ;
    END
  END Data_HV[627]
  PIN Data_HV[626]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16231.385 187.44 16231.665 188.44 ;
    END
  END Data_HV[626]
  PIN Data_HV[625]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16233.625 187.44 16233.905 188.44 ;
    END
  END Data_HV[625]
  PIN Data_HV[624]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16235.305 187.44 16235.585 188.44 ;
    END
  END Data_HV[624]
  PIN Data_HV[623]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16260.505 187.44 16260.785 188.44 ;
    END
  END Data_HV[623]
  PIN Data_HV[622]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16261.625 187.44 16261.905 188.44 ;
    END
  END Data_HV[622]
  PIN Data_HV[621]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16288.785 187.44 16289.065 188.44 ;
    END
  END Data_HV[621]
  PIN Data_HV[620]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16233.065 187.44 16233.345 188.44 ;
    END
  END Data_HV[620]
  PIN Data_HV[619]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16234.745 187.44 16235.025 188.44 ;
    END
  END Data_HV[619]
  PIN Data_HV[618]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16248.745 187.44 16249.025 188.44 ;
    END
  END Data_HV[618]
  PIN Data_HV[617]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16289.345 187.44 16289.625 188.44 ;
    END
  END Data_HV[617]
  PIN Data_HV[616]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16259.945 187.44 16260.225 188.44 ;
    END
  END Data_HV[616]
  PIN Data_HV[615]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16259.385 187.44 16259.665 188.44 ;
    END
  END Data_HV[615]
  PIN Data_HV[614]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16287.665 187.44 16287.945 188.44 ;
    END
  END Data_HV[614]
  PIN Data_HV[613]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16234.185 187.44 16234.465 188.44 ;
    END
  END Data_HV[613]
  PIN Data_HV[612]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16249.865 187.44 16250.145 188.44 ;
    END
  END Data_HV[612]
  PIN Data_HV[611]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16249.305 187.44 16249.585 188.44 ;
    END
  END Data_HV[611]
  PIN Data_HV[610]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16232.505 187.44 16232.785 188.44 ;
    END
  END Data_HV[610]
  PIN Data_HV[609]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16231.945 187.44 16232.225 188.44 ;
    END
  END Data_HV[609]
  PIN Data_HV[608]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16178.745 187.44 16179.025 188.44 ;
    END
  END Data_HV[608]
  PIN Data_HV[607]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16180.425 187.44 16180.705 188.44 ;
    END
  END Data_HV[607]
  PIN Data_HV[606]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16182.105 187.44 16182.385 188.44 ;
    END
  END Data_HV[606]
  PIN Data_HV[605]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16153.545 187.44 16153.825 188.44 ;
    END
  END Data_HV[605]
  PIN Data_HV[604]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16155.785 187.44 16156.065 188.44 ;
    END
  END Data_HV[604]
  PIN Data_HV[603]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16157.465 187.44 16157.745 188.44 ;
    END
  END Data_HV[603]
  PIN Data_HV[602]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16178.185 187.44 16178.465 188.44 ;
    END
  END Data_HV[602]
  PIN Data_HV[601]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16179.305 187.44 16179.585 188.44 ;
    END
  END Data_HV[601]
  PIN Data_HV[600]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16180.985 187.44 16181.265 188.44 ;
    END
  END Data_HV[600]
  PIN Data_HV[599]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16155.225 187.44 16155.505 188.44 ;
    END
  END Data_HV[599]
  PIN Data_HV[598]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16156.905 187.44 16157.185 188.44 ;
    END
  END Data_HV[598]
  PIN Data_HV[597]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16158.025 187.44 16158.305 188.44 ;
    END
  END Data_HV[597]
  PIN Data_HV[596]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16181.545 187.44 16181.825 188.44 ;
    END
  END Data_HV[596]
  PIN Data_HV[595]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16177.625 187.44 16177.905 188.44 ;
    END
  END Data_HV[595]
  PIN Data_HV[594]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16177.065 187.44 16177.345 188.44 ;
    END
  END Data_HV[594]
  PIN Data_HV[593]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16179.865 187.44 16180.145 188.44 ;
    END
  END Data_HV[593]
  PIN Data_HV[592]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16156.345 187.44 16156.625 188.44 ;
    END
  END Data_HV[592]
  PIN Data_HV[591]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16159.145 187.44 16159.425 188.44 ;
    END
  END Data_HV[591]
  PIN Data_HV[590]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16158.585 187.44 16158.865 188.44 ;
    END
  END Data_HV[590]
  PIN Data_HV[589]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16154.665 187.44 16154.945 188.44 ;
    END
  END Data_HV[589]
  PIN Data_HV[588]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16154.105 187.44 16154.385 188.44 ;
    END
  END Data_HV[588]
  PIN Data_HV[587]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16112.665 187.44 16112.945 188.44 ;
    END
  END Data_HV[587]
  PIN Data_HV[586]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16114.345 187.44 16114.625 188.44 ;
    END
  END Data_HV[586]
  PIN Data_HV[585]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16116.025 187.44 16116.305 188.44 ;
    END
  END Data_HV[585]
  PIN Data_HV[584]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16082.425 187.44 16082.705 188.44 ;
    END
  END Data_HV[584]
  PIN Data_HV[583]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16084.665 187.44 16084.945 188.44 ;
    END
  END Data_HV[583]
  PIN Data_HV[582]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16086.345 187.44 16086.625 188.44 ;
    END
  END Data_HV[582]
  PIN Data_HV[581]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16112.105 187.44 16112.385 188.44 ;
    END
  END Data_HV[581]
  PIN Data_HV[580]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16113.225 187.44 16113.505 188.44 ;
    END
  END Data_HV[580]
  PIN Data_HV[579]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16114.905 187.44 16115.185 188.44 ;
    END
  END Data_HV[579]
  PIN Data_HV[578]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16084.105 187.44 16084.385 188.44 ;
    END
  END Data_HV[578]
  PIN Data_HV[577]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16085.785 187.44 16086.065 188.44 ;
    END
  END Data_HV[577]
  PIN Data_HV[576]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16086.905 187.44 16087.185 188.44 ;
    END
  END Data_HV[576]
  PIN Data_HV[575]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16115.465 187.44 16115.745 188.44 ;
    END
  END Data_HV[575]
  PIN Data_HV[574]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16111.545 187.44 16111.825 188.44 ;
    END
  END Data_HV[574]
  PIN Data_HV[573]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16110.985 187.44 16111.265 188.44 ;
    END
  END Data_HV[573]
  PIN Data_HV[572]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16113.785 187.44 16114.065 188.44 ;
    END
  END Data_HV[572]
  PIN Data_HV[571]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16085.225 187.44 16085.505 188.44 ;
    END
  END Data_HV[571]
  PIN Data_HV[570]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16088.025 187.44 16088.305 188.44 ;
    END
  END Data_HV[570]
  PIN Data_HV[569]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16087.465 187.44 16087.745 188.44 ;
    END
  END Data_HV[569]
  PIN Data_HV[568]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16083.545 187.44 16083.825 188.44 ;
    END
  END Data_HV[568]
  PIN Data_HV[567]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16082.985 187.44 16083.265 188.44 ;
    END
  END Data_HV[567]
  PIN Data_HV[566]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16030.905 187.44 16031.185 188.44 ;
    END
  END Data_HV[566]
  PIN Data_HV[565]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16032.585 187.44 16032.865 188.44 ;
    END
  END Data_HV[565]
  PIN Data_HV[564]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16034.265 187.44 16034.545 188.44 ;
    END
  END Data_HV[564]
  PIN Data_HV[563]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15978.265 187.44 15978.545 188.44 ;
    END
  END Data_HV[563]
  PIN Data_HV[562]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15980.505 187.44 15980.785 188.44 ;
    END
  END Data_HV[562]
  PIN Data_HV[561]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16007.665 187.44 16007.945 188.44 ;
    END
  END Data_HV[561]
  PIN Data_HV[560]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16030.345 187.44 16030.625 188.44 ;
    END
  END Data_HV[560]
  PIN Data_HV[559]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16031.465 187.44 16031.745 188.44 ;
    END
  END Data_HV[559]
  PIN Data_HV[558]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16033.145 187.44 16033.425 188.44 ;
    END
  END Data_HV[558]
  PIN Data_HV[557]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15979.945 187.44 15980.225 188.44 ;
    END
  END Data_HV[557]
  PIN Data_HV[556]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16007.105 187.44 16007.385 188.44 ;
    END
  END Data_HV[556]
  PIN Data_HV[555]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16008.225 187.44 16008.505 188.44 ;
    END
  END Data_HV[555]
  PIN Data_HV[554]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16033.705 187.44 16033.985 188.44 ;
    END
  END Data_HV[554]
  PIN Data_HV[553]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16029.785 187.44 16030.065 188.44 ;
    END
  END Data_HV[553]
  PIN Data_HV[552]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16020.825 187.44 16021.105 188.44 ;
    END
  END Data_HV[552]
  PIN Data_HV[551]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16032.025 187.44 16032.305 188.44 ;
    END
  END Data_HV[551]
  PIN Data_HV[550]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15981.065 187.44 15981.345 188.44 ;
    END
  END Data_HV[550]
  PIN Data_HV[549]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16009.345 187.44 16009.625 188.44 ;
    END
  END Data_HV[549]
  PIN Data_HV[548]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16008.785 187.44 16009.065 188.44 ;
    END
  END Data_HV[548]
  PIN Data_HV[547]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15979.385 187.44 15979.665 188.44 ;
    END
  END Data_HV[547]
  PIN Data_HV[546]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15978.825 187.44 15979.105 188.44 ;
    END
  END Data_HV[546]
  PIN Data_HV[545]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15952.505 187.44 15952.785 188.44 ;
    END
  END Data_HV[545]
  PIN Data_HV[544]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15954.185 187.44 15954.465 188.44 ;
    END
  END Data_HV[544]
  PIN Data_HV[543]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15968.745 187.44 15969.025 188.44 ;
    END
  END Data_HV[543]
  PIN Data_HV[542]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15897.065 187.44 15897.345 188.44 ;
    END
  END Data_HV[542]
  PIN Data_HV[541]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15899.305 187.44 15899.585 188.44 ;
    END
  END Data_HV[541]
  PIN Data_HV[540]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15900.985 187.44 15901.265 188.44 ;
    END
  END Data_HV[540]
  PIN Data_HV[539]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15951.945 187.44 15952.225 188.44 ;
    END
  END Data_HV[539]
  PIN Data_HV[538]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15953.065 187.44 15953.345 188.44 ;
    END
  END Data_HV[538]
  PIN Data_HV[537]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15954.745 187.44 15955.025 188.44 ;
    END
  END Data_HV[537]
  PIN Data_HV[536]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15898.745 187.44 15899.025 188.44 ;
    END
  END Data_HV[536]
  PIN Data_HV[535]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15900.425 187.44 15900.705 188.44 ;
    END
  END Data_HV[535]
  PIN Data_HV[534]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15901.545 187.44 15901.825 188.44 ;
    END
  END Data_HV[534]
  PIN Data_HV[533]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15968.185 187.44 15968.465 188.44 ;
    END
  END Data_HV[533]
  PIN Data_HV[532]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15951.385 187.44 15951.665 188.44 ;
    END
  END Data_HV[532]
  PIN Data_HV[531]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15950.825 187.44 15951.105 188.44 ;
    END
  END Data_HV[531]
  PIN Data_HV[530]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15953.625 187.44 15953.905 188.44 ;
    END
  END Data_HV[530]
  PIN Data_HV[529]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15899.865 187.44 15900.145 188.44 ;
    END
  END Data_HV[529]
  PIN Data_HV[528]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15902.665 187.44 15902.945 188.44 ;
    END
  END Data_HV[528]
  PIN Data_HV[527]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15902.105 187.44 15902.385 188.44 ;
    END
  END Data_HV[527]
  PIN Data_HV[526]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15898.185 187.44 15898.465 188.44 ;
    END
  END Data_HV[526]
  PIN Data_HV[525]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15897.625 187.44 15897.905 188.44 ;
    END
  END Data_HV[525]
  PIN Data_HV[524]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15875.785 187.44 15876.065 188.44 ;
    END
  END Data_HV[524]
  PIN Data_HV[523]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15877.465 187.44 15877.745 188.44 ;
    END
  END Data_HV[523]
  PIN Data_HV[522]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15879.145 187.44 15879.425 188.44 ;
    END
  END Data_HV[522]
  PIN Data_HV[521]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15831.545 187.44 15831.825 188.44 ;
    END
  END Data_HV[521]
  PIN Data_HV[520]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15833.785 187.44 15834.065 188.44 ;
    END
  END Data_HV[520]
  PIN Data_HV[519]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15835.465 187.44 15835.745 188.44 ;
    END
  END Data_HV[519]
  PIN Data_HV[518]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15875.225 187.44 15875.505 188.44 ;
    END
  END Data_HV[518]
  PIN Data_HV[517]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15876.345 187.44 15876.625 188.44 ;
    END
  END Data_HV[517]
  PIN Data_HV[516]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15878.025 187.44 15878.305 188.44 ;
    END
  END Data_HV[516]
  PIN Data_HV[515]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15833.225 187.44 15833.505 188.44 ;
    END
  END Data_HV[515]
  PIN Data_HV[514]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15834.905 187.44 15835.185 188.44 ;
    END
  END Data_HV[514]
  PIN Data_HV[513]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15836.025 187.44 15836.305 188.44 ;
    END
  END Data_HV[513]
  PIN Data_HV[512]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15878.585 187.44 15878.865 188.44 ;
    END
  END Data_HV[512]
  PIN Data_HV[511]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15874.665 187.44 15874.945 188.44 ;
    END
  END Data_HV[511]
  PIN Data_HV[510]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15874.105 187.44 15874.385 188.44 ;
    END
  END Data_HV[510]
  PIN Data_HV[509]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15876.905 187.44 15877.185 188.44 ;
    END
  END Data_HV[509]
  PIN Data_HV[508]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15834.345 187.44 15834.625 188.44 ;
    END
  END Data_HV[508]
  PIN Data_HV[507]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15837.145 187.44 15837.425 188.44 ;
    END
  END Data_HV[507]
  PIN Data_HV[506]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15836.585 187.44 15836.865 188.44 ;
    END
  END Data_HV[506]
  PIN Data_HV[505]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15832.665 187.44 15832.945 188.44 ;
    END
  END Data_HV[505]
  PIN Data_HV[504]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15832.105 187.44 15832.385 188.44 ;
    END
  END Data_HV[504]
  PIN Data_HV[503]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15805.785 187.44 15806.065 188.44 ;
    END
  END Data_HV[503]
  PIN Data_HV[502]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15807.465 187.44 15807.745 188.44 ;
    END
  END Data_HV[502]
  PIN Data_HV[501]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15809.145 187.44 15809.425 188.44 ;
    END
  END Data_HV[501]
  PIN Data_HV[500]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15749.785 187.44 15750.065 188.44 ;
    END
  END Data_HV[500]
  PIN Data_HV[499]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15752.025 187.44 15752.305 188.44 ;
    END
  END Data_HV[499]
  PIN Data_HV[498]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15753.705 187.44 15753.985 188.44 ;
    END
  END Data_HV[498]
  PIN Data_HV[497]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15805.225 187.44 15805.505 188.44 ;
    END
  END Data_HV[497]
  PIN Data_HV[496]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15806.345 187.44 15806.625 188.44 ;
    END
  END Data_HV[496]
  PIN Data_HV[495]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15808.025 187.44 15808.305 188.44 ;
    END
  END Data_HV[495]
  PIN Data_HV[494]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15751.465 187.44 15751.745 188.44 ;
    END
  END Data_HV[494]
  PIN Data_HV[493]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15753.145 187.44 15753.425 188.44 ;
    END
  END Data_HV[493]
  PIN Data_HV[492]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15754.265 187.44 15754.545 188.44 ;
    END
  END Data_HV[492]
  PIN Data_HV[491]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15808.585 187.44 15808.865 188.44 ;
    END
  END Data_HV[491]
  PIN Data_HV[490]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15804.665 187.44 15804.945 188.44 ;
    END
  END Data_HV[490]
  PIN Data_HV[489]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15804.105 187.44 15804.385 188.44 ;
    END
  END Data_HV[489]
  PIN Data_HV[488]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15806.905 187.44 15807.185 188.44 ;
    END
  END Data_HV[488]
  PIN Data_HV[487]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15752.585 187.44 15752.865 188.44 ;
    END
  END Data_HV[487]
  PIN Data_HV[486]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15755.385 187.44 15755.665 188.44 ;
    END
  END Data_HV[486]
  PIN Data_HV[485]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15754.825 187.44 15755.105 188.44 ;
    END
  END Data_HV[485]
  PIN Data_HV[484]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15750.905 187.44 15751.185 188.44 ;
    END
  END Data_HV[484]
  PIN Data_HV[483]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15750.345 187.44 15750.625 188.44 ;
    END
  END Data_HV[483]
  PIN Data_HV[482]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15701.065 187.44 15701.345 188.44 ;
    END
  END Data_HV[482]
  PIN Data_HV[481]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15728.225 187.44 15728.505 188.44 ;
    END
  END Data_HV[481]
  PIN Data_HV[480]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15729.905 187.44 15730.185 188.44 ;
    END
  END Data_HV[480]
  PIN Data_HV[479]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15671.385 187.44 15671.665 188.44 ;
    END
  END Data_HV[479]
  PIN Data_HV[478]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15673.625 187.44 15673.905 188.44 ;
    END
  END Data_HV[478]
  PIN Data_HV[477]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15675.305 187.44 15675.585 188.44 ;
    END
  END Data_HV[477]
  PIN Data_HV[476]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15700.505 187.44 15700.785 188.44 ;
    END
  END Data_HV[476]
  PIN Data_HV[475]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15701.625 187.44 15701.905 188.44 ;
    END
  END Data_HV[475]
  PIN Data_HV[474]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15728.785 187.44 15729.065 188.44 ;
    END
  END Data_HV[474]
  PIN Data_HV[473]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15673.065 187.44 15673.345 188.44 ;
    END
  END Data_HV[473]
  PIN Data_HV[472]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15674.745 187.44 15675.025 188.44 ;
    END
  END Data_HV[472]
  PIN Data_HV[471]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15688.745 187.44 15689.025 188.44 ;
    END
  END Data_HV[471]
  PIN Data_HV[470]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15729.345 187.44 15729.625 188.44 ;
    END
  END Data_HV[470]
  PIN Data_HV[469]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15699.945 187.44 15700.225 188.44 ;
    END
  END Data_HV[469]
  PIN Data_HV[468]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15699.385 187.44 15699.665 188.44 ;
    END
  END Data_HV[468]
  PIN Data_HV[467]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15727.665 187.44 15727.945 188.44 ;
    END
  END Data_HV[467]
  PIN Data_HV[466]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15674.185 187.44 15674.465 188.44 ;
    END
  END Data_HV[466]
  PIN Data_HV[465]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15689.865 187.44 15690.145 188.44 ;
    END
  END Data_HV[465]
  PIN Data_HV[464]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15689.305 187.44 15689.585 188.44 ;
    END
  END Data_HV[464]
  PIN Data_HV[463]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15672.505 187.44 15672.785 188.44 ;
    END
  END Data_HV[463]
  PIN Data_HV[462]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15671.945 187.44 15672.225 188.44 ;
    END
  END Data_HV[462]
  PIN Data_HV[461]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15618.745 187.44 15619.025 188.44 ;
    END
  END Data_HV[461]
  PIN Data_HV[460]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15620.425 187.44 15620.705 188.44 ;
    END
  END Data_HV[460]
  PIN Data_HV[459]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15622.105 187.44 15622.385 188.44 ;
    END
  END Data_HV[459]
  PIN Data_HV[458]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15593.545 187.44 15593.825 188.44 ;
    END
  END Data_HV[458]
  PIN Data_HV[457]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15595.785 187.44 15596.065 188.44 ;
    END
  END Data_HV[457]
  PIN Data_HV[456]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15597.465 187.44 15597.745 188.44 ;
    END
  END Data_HV[456]
  PIN Data_HV[455]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15618.185 187.44 15618.465 188.44 ;
    END
  END Data_HV[455]
  PIN Data_HV[454]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15619.305 187.44 15619.585 188.44 ;
    END
  END Data_HV[454]
  PIN Data_HV[453]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15620.985 187.44 15621.265 188.44 ;
    END
  END Data_HV[453]
  PIN Data_HV[452]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15595.225 187.44 15595.505 188.44 ;
    END
  END Data_HV[452]
  PIN Data_HV[451]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15596.905 187.44 15597.185 188.44 ;
    END
  END Data_HV[451]
  PIN Data_HV[450]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15598.025 187.44 15598.305 188.44 ;
    END
  END Data_HV[450]
  PIN Data_HV[449]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15621.545 187.44 15621.825 188.44 ;
    END
  END Data_HV[449]
  PIN Data_HV[448]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15617.625 187.44 15617.905 188.44 ;
    END
  END Data_HV[448]
  PIN Data_HV[447]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15617.065 187.44 15617.345 188.44 ;
    END
  END Data_HV[447]
  PIN Data_HV[446]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15619.865 187.44 15620.145 188.44 ;
    END
  END Data_HV[446]
  PIN Data_HV[445]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15596.345 187.44 15596.625 188.44 ;
    END
  END Data_HV[445]
  PIN Data_HV[444]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15599.145 187.44 15599.425 188.44 ;
    END
  END Data_HV[444]
  PIN Data_HV[443]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15598.585 187.44 15598.865 188.44 ;
    END
  END Data_HV[443]
  PIN Data_HV[442]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15594.665 187.44 15594.945 188.44 ;
    END
  END Data_HV[442]
  PIN Data_HV[441]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15594.105 187.44 15594.385 188.44 ;
    END
  END Data_HV[441]
  PIN Data_HV[440]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15552.665 187.44 15552.945 188.44 ;
    END
  END Data_HV[440]
  PIN Data_HV[439]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15554.345 187.44 15554.625 188.44 ;
    END
  END Data_HV[439]
  PIN Data_HV[438]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15556.025 187.44 15556.305 188.44 ;
    END
  END Data_HV[438]
  PIN Data_HV[437]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15522.425 187.44 15522.705 188.44 ;
    END
  END Data_HV[437]
  PIN Data_HV[436]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15524.665 187.44 15524.945 188.44 ;
    END
  END Data_HV[436]
  PIN Data_HV[435]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15526.345 187.44 15526.625 188.44 ;
    END
  END Data_HV[435]
  PIN Data_HV[434]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15552.105 187.44 15552.385 188.44 ;
    END
  END Data_HV[434]
  PIN Data_HV[433]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15553.225 187.44 15553.505 188.44 ;
    END
  END Data_HV[433]
  PIN Data_HV[432]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15554.905 187.44 15555.185 188.44 ;
    END
  END Data_HV[432]
  PIN Data_HV[431]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15524.105 187.44 15524.385 188.44 ;
    END
  END Data_HV[431]
  PIN Data_HV[430]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15525.785 187.44 15526.065 188.44 ;
    END
  END Data_HV[430]
  PIN Data_HV[429]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15526.905 187.44 15527.185 188.44 ;
    END
  END Data_HV[429]
  PIN Data_HV[428]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15555.465 187.44 15555.745 188.44 ;
    END
  END Data_HV[428]
  PIN Data_HV[427]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15551.545 187.44 15551.825 188.44 ;
    END
  END Data_HV[427]
  PIN Data_HV[426]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15550.985 187.44 15551.265 188.44 ;
    END
  END Data_HV[426]
  PIN Data_HV[425]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15553.785 187.44 15554.065 188.44 ;
    END
  END Data_HV[425]
  PIN Data_HV[424]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15525.225 187.44 15525.505 188.44 ;
    END
  END Data_HV[424]
  PIN Data_HV[423]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15528.025 187.44 15528.305 188.44 ;
    END
  END Data_HV[423]
  PIN Data_HV[422]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15527.465 187.44 15527.745 188.44 ;
    END
  END Data_HV[422]
  PIN Data_HV[421]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15523.545 187.44 15523.825 188.44 ;
    END
  END Data_HV[421]
  PIN Data_HV[420]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15522.985 187.44 15523.265 188.44 ;
    END
  END Data_HV[420]
  PIN Data_HV[419]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15470.905 187.44 15471.185 188.44 ;
    END
  END Data_HV[419]
  PIN Data_HV[418]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15472.585 187.44 15472.865 188.44 ;
    END
  END Data_HV[418]
  PIN Data_HV[417]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15474.265 187.44 15474.545 188.44 ;
    END
  END Data_HV[417]
  PIN Data_HV[416]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15418.265 187.44 15418.545 188.44 ;
    END
  END Data_HV[416]
  PIN Data_HV[415]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15420.505 187.44 15420.785 188.44 ;
    END
  END Data_HV[415]
  PIN Data_HV[414]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15447.665 187.44 15447.945 188.44 ;
    END
  END Data_HV[414]
  PIN Data_HV[413]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15470.345 187.44 15470.625 188.44 ;
    END
  END Data_HV[413]
  PIN Data_HV[412]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15471.465 187.44 15471.745 188.44 ;
    END
  END Data_HV[412]
  PIN Data_HV[411]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15473.145 187.44 15473.425 188.44 ;
    END
  END Data_HV[411]
  PIN Data_HV[410]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15419.945 187.44 15420.225 188.44 ;
    END
  END Data_HV[410]
  PIN Data_HV[409]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15447.105 187.44 15447.385 188.44 ;
    END
  END Data_HV[409]
  PIN Data_HV[408]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15448.225 187.44 15448.505 188.44 ;
    END
  END Data_HV[408]
  PIN Data_HV[407]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15473.705 187.44 15473.985 188.44 ;
    END
  END Data_HV[407]
  PIN Data_HV[406]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15469.785 187.44 15470.065 188.44 ;
    END
  END Data_HV[406]
  PIN Data_HV[405]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15460.825 187.44 15461.105 188.44 ;
    END
  END Data_HV[405]
  PIN Data_HV[404]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15472.025 187.44 15472.305 188.44 ;
    END
  END Data_HV[404]
  PIN Data_HV[403]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15421.065 187.44 15421.345 188.44 ;
    END
  END Data_HV[403]
  PIN Data_HV[402]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15449.345 187.44 15449.625 188.44 ;
    END
  END Data_HV[402]
  PIN Data_HV[401]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15448.785 187.44 15449.065 188.44 ;
    END
  END Data_HV[401]
  PIN Data_HV[400]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15419.385 187.44 15419.665 188.44 ;
    END
  END Data_HV[400]
  PIN Data_HV[399]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15418.825 187.44 15419.105 188.44 ;
    END
  END Data_HV[399]
  PIN Data_HV[398]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15392.505 187.44 15392.785 188.44 ;
    END
  END Data_HV[398]
  PIN Data_HV[397]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15394.185 187.44 15394.465 188.44 ;
    END
  END Data_HV[397]
  PIN Data_HV[396]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15408.745 187.44 15409.025 188.44 ;
    END
  END Data_HV[396]
  PIN Data_HV[395]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15337.065 187.44 15337.345 188.44 ;
    END
  END Data_HV[395]
  PIN Data_HV[394]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15339.305 187.44 15339.585 188.44 ;
    END
  END Data_HV[394]
  PIN Data_HV[393]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15340.985 187.44 15341.265 188.44 ;
    END
  END Data_HV[393]
  PIN Data_HV[392]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15391.945 187.44 15392.225 188.44 ;
    END
  END Data_HV[392]
  PIN Data_HV[391]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15393.065 187.44 15393.345 188.44 ;
    END
  END Data_HV[391]
  PIN Data_HV[390]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15394.745 187.44 15395.025 188.44 ;
    END
  END Data_HV[390]
  PIN Data_HV[389]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15338.745 187.44 15339.025 188.44 ;
    END
  END Data_HV[389]
  PIN Data_HV[388]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15340.425 187.44 15340.705 188.44 ;
    END
  END Data_HV[388]
  PIN Data_HV[387]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15341.545 187.44 15341.825 188.44 ;
    END
  END Data_HV[387]
  PIN Data_HV[386]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15408.185 187.44 15408.465 188.44 ;
    END
  END Data_HV[386]
  PIN Data_HV[385]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15391.385 187.44 15391.665 188.44 ;
    END
  END Data_HV[385]
  PIN Data_HV[384]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15390.825 187.44 15391.105 188.44 ;
    END
  END Data_HV[384]
  PIN Data_HV[383]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15393.625 187.44 15393.905 188.44 ;
    END
  END Data_HV[383]
  PIN Data_HV[382]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15339.865 187.44 15340.145 188.44 ;
    END
  END Data_HV[382]
  PIN Data_HV[381]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15342.665 187.44 15342.945 188.44 ;
    END
  END Data_HV[381]
  PIN Data_HV[380]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15342.105 187.44 15342.385 188.44 ;
    END
  END Data_HV[380]
  PIN Data_HV[379]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15338.185 187.44 15338.465 188.44 ;
    END
  END Data_HV[379]
  PIN Data_HV[378]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15337.625 187.44 15337.905 188.44 ;
    END
  END Data_HV[378]
  PIN Data_HV[377]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15315.785 187.44 15316.065 188.44 ;
    END
  END Data_HV[377]
  PIN Data_HV[376]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15317.465 187.44 15317.745 188.44 ;
    END
  END Data_HV[376]
  PIN Data_HV[375]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15319.145 187.44 15319.425 188.44 ;
    END
  END Data_HV[375]
  PIN Data_HV[374]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15271.545 187.44 15271.825 188.44 ;
    END
  END Data_HV[374]
  PIN Data_HV[373]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15273.785 187.44 15274.065 188.44 ;
    END
  END Data_HV[373]
  PIN Data_HV[372]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15275.465 187.44 15275.745 188.44 ;
    END
  END Data_HV[372]
  PIN Data_HV[371]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15315.225 187.44 15315.505 188.44 ;
    END
  END Data_HV[371]
  PIN Data_HV[370]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15316.345 187.44 15316.625 188.44 ;
    END
  END Data_HV[370]
  PIN Data_HV[369]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15318.025 187.44 15318.305 188.44 ;
    END
  END Data_HV[369]
  PIN Data_HV[368]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15273.225 187.44 15273.505 188.44 ;
    END
  END Data_HV[368]
  PIN Data_HV[367]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15274.905 187.44 15275.185 188.44 ;
    END
  END Data_HV[367]
  PIN Data_HV[366]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15276.025 187.44 15276.305 188.44 ;
    END
  END Data_HV[366]
  PIN Data_HV[365]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15318.585 187.44 15318.865 188.44 ;
    END
  END Data_HV[365]
  PIN Data_HV[364]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15314.665 187.44 15314.945 188.44 ;
    END
  END Data_HV[364]
  PIN Data_HV[363]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15314.105 187.44 15314.385 188.44 ;
    END
  END Data_HV[363]
  PIN Data_HV[362]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15316.905 187.44 15317.185 188.44 ;
    END
  END Data_HV[362]
  PIN Data_HV[361]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15274.345 187.44 15274.625 188.44 ;
    END
  END Data_HV[361]
  PIN Data_HV[360]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15277.145 187.44 15277.425 188.44 ;
    END
  END Data_HV[360]
  PIN Data_HV[359]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15276.585 187.44 15276.865 188.44 ;
    END
  END Data_HV[359]
  PIN Data_HV[358]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15272.665 187.44 15272.945 188.44 ;
    END
  END Data_HV[358]
  PIN Data_HV[357]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15272.105 187.44 15272.385 188.44 ;
    END
  END Data_HV[357]
  PIN Data_HV[356]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15245.785 187.44 15246.065 188.44 ;
    END
  END Data_HV[356]
  PIN Data_HV[355]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15247.465 187.44 15247.745 188.44 ;
    END
  END Data_HV[355]
  PIN Data_HV[354]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15249.145 187.44 15249.425 188.44 ;
    END
  END Data_HV[354]
  PIN Data_HV[353]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15189.785 187.44 15190.065 188.44 ;
    END
  END Data_HV[353]
  PIN Data_HV[352]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15192.025 187.44 15192.305 188.44 ;
    END
  END Data_HV[352]
  PIN Data_HV[351]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15193.705 187.44 15193.985 188.44 ;
    END
  END Data_HV[351]
  PIN Data_HV[350]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15245.225 187.44 15245.505 188.44 ;
    END
  END Data_HV[350]
  PIN Data_HV[349]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15246.345 187.44 15246.625 188.44 ;
    END
  END Data_HV[349]
  PIN Data_HV[348]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15248.025 187.44 15248.305 188.44 ;
    END
  END Data_HV[348]
  PIN Data_HV[347]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15191.465 187.44 15191.745 188.44 ;
    END
  END Data_HV[347]
  PIN Data_HV[346]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15193.145 187.44 15193.425 188.44 ;
    END
  END Data_HV[346]
  PIN Data_HV[345]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15194.265 187.44 15194.545 188.44 ;
    END
  END Data_HV[345]
  PIN Data_HV[344]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15248.585 187.44 15248.865 188.44 ;
    END
  END Data_HV[344]
  PIN Data_HV[343]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15244.665 187.44 15244.945 188.44 ;
    END
  END Data_HV[343]
  PIN Data_HV[342]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15244.105 187.44 15244.385 188.44 ;
    END
  END Data_HV[342]
  PIN Data_HV[341]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15246.905 187.44 15247.185 188.44 ;
    END
  END Data_HV[341]
  PIN Data_HV[340]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15192.585 187.44 15192.865 188.44 ;
    END
  END Data_HV[340]
  PIN Data_HV[339]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15195.385 187.44 15195.665 188.44 ;
    END
  END Data_HV[339]
  PIN Data_HV[338]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15194.825 187.44 15195.105 188.44 ;
    END
  END Data_HV[338]
  PIN Data_HV[337]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15190.905 187.44 15191.185 188.44 ;
    END
  END Data_HV[337]
  PIN Data_HV[336]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15190.345 187.44 15190.625 188.44 ;
    END
  END Data_HV[336]
  PIN Data_HV[335]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15141.065 187.44 15141.345 188.44 ;
    END
  END Data_HV[335]
  PIN Data_HV[334]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15168.225 187.44 15168.505 188.44 ;
    END
  END Data_HV[334]
  PIN Data_HV[333]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15169.905 187.44 15170.185 188.44 ;
    END
  END Data_HV[333]
  PIN Data_HV[332]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15111.385 187.44 15111.665 188.44 ;
    END
  END Data_HV[332]
  PIN Data_HV[331]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15113.625 187.44 15113.905 188.44 ;
    END
  END Data_HV[331]
  PIN Data_HV[330]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15115.305 187.44 15115.585 188.44 ;
    END
  END Data_HV[330]
  PIN Data_HV[329]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15140.505 187.44 15140.785 188.44 ;
    END
  END Data_HV[329]
  PIN Data_HV[328]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15141.625 187.44 15141.905 188.44 ;
    END
  END Data_HV[328]
  PIN Data_HV[327]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15168.785 187.44 15169.065 188.44 ;
    END
  END Data_HV[327]
  PIN Data_HV[326]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15113.065 187.44 15113.345 188.44 ;
    END
  END Data_HV[326]
  PIN Data_HV[325]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15114.745 187.44 15115.025 188.44 ;
    END
  END Data_HV[325]
  PIN Data_HV[324]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15128.745 187.44 15129.025 188.44 ;
    END
  END Data_HV[324]
  PIN Data_HV[323]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15169.345 187.44 15169.625 188.44 ;
    END
  END Data_HV[323]
  PIN Data_HV[322]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15139.945 187.44 15140.225 188.44 ;
    END
  END Data_HV[322]
  PIN Data_HV[321]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15139.385 187.44 15139.665 188.44 ;
    END
  END Data_HV[321]
  PIN Data_HV[320]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15167.665 187.44 15167.945 188.44 ;
    END
  END Data_HV[320]
  PIN Data_HV[319]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15114.185 187.44 15114.465 188.44 ;
    END
  END Data_HV[319]
  PIN Data_HV[318]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15129.865 187.44 15130.145 188.44 ;
    END
  END Data_HV[318]
  PIN Data_HV[317]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15129.305 187.44 15129.585 188.44 ;
    END
  END Data_HV[317]
  PIN Data_HV[316]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15112.505 187.44 15112.785 188.44 ;
    END
  END Data_HV[316]
  PIN Data_HV[315]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15111.945 187.44 15112.225 188.44 ;
    END
  END Data_HV[315]
  PIN Data_HV[314]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15058.745 187.44 15059.025 188.44 ;
    END
  END Data_HV[314]
  PIN Data_HV[313]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15060.425 187.44 15060.705 188.44 ;
    END
  END Data_HV[313]
  PIN Data_HV[312]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15062.105 187.44 15062.385 188.44 ;
    END
  END Data_HV[312]
  PIN Data_HV[311]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15033.545 187.44 15033.825 188.44 ;
    END
  END Data_HV[311]
  PIN Data_HV[310]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15035.785 187.44 15036.065 188.44 ;
    END
  END Data_HV[310]
  PIN Data_HV[309]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15037.465 187.44 15037.745 188.44 ;
    END
  END Data_HV[309]
  PIN Data_HV[308]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15058.185 187.44 15058.465 188.44 ;
    END
  END Data_HV[308]
  PIN Data_HV[307]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15059.305 187.44 15059.585 188.44 ;
    END
  END Data_HV[307]
  PIN Data_HV[306]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15060.985 187.44 15061.265 188.44 ;
    END
  END Data_HV[306]
  PIN Data_HV[305]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15035.225 187.44 15035.505 188.44 ;
    END
  END Data_HV[305]
  PIN Data_HV[304]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15036.905 187.44 15037.185 188.44 ;
    END
  END Data_HV[304]
  PIN Data_HV[303]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15038.025 187.44 15038.305 188.44 ;
    END
  END Data_HV[303]
  PIN Data_HV[302]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15061.545 187.44 15061.825 188.44 ;
    END
  END Data_HV[302]
  PIN Data_HV[301]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15057.625 187.44 15057.905 188.44 ;
    END
  END Data_HV[301]
  PIN Data_HV[300]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15057.065 187.44 15057.345 188.44 ;
    END
  END Data_HV[300]
  PIN Data_HV[299]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15059.865 187.44 15060.145 188.44 ;
    END
  END Data_HV[299]
  PIN Data_HV[298]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15036.345 187.44 15036.625 188.44 ;
    END
  END Data_HV[298]
  PIN Data_HV[297]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15039.145 187.44 15039.425 188.44 ;
    END
  END Data_HV[297]
  PIN Data_HV[296]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15038.585 187.44 15038.865 188.44 ;
    END
  END Data_HV[296]
  PIN Data_HV[295]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15034.665 187.44 15034.945 188.44 ;
    END
  END Data_HV[295]
  PIN Data_HV[294]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15034.105 187.44 15034.385 188.44 ;
    END
  END Data_HV[294]
  PIN Data_HV[293]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14992.665 187.44 14992.945 188.44 ;
    END
  END Data_HV[293]
  PIN Data_HV[292]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14994.345 187.44 14994.625 188.44 ;
    END
  END Data_HV[292]
  PIN Data_HV[291]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14996.025 187.44 14996.305 188.44 ;
    END
  END Data_HV[291]
  PIN Data_HV[290]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14962.425 187.44 14962.705 188.44 ;
    END
  END Data_HV[290]
  PIN Data_HV[289]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14964.665 187.44 14964.945 188.44 ;
    END
  END Data_HV[289]
  PIN Data_HV[288]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14966.345 187.44 14966.625 188.44 ;
    END
  END Data_HV[288]
  PIN Data_HV[287]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14992.105 187.44 14992.385 188.44 ;
    END
  END Data_HV[287]
  PIN Data_HV[286]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14993.225 187.44 14993.505 188.44 ;
    END
  END Data_HV[286]
  PIN Data_HV[285]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14994.905 187.44 14995.185 188.44 ;
    END
  END Data_HV[285]
  PIN Data_HV[284]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14964.105 187.44 14964.385 188.44 ;
    END
  END Data_HV[284]
  PIN Data_HV[283]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14965.785 187.44 14966.065 188.44 ;
    END
  END Data_HV[283]
  PIN Data_HV[282]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14966.905 187.44 14967.185 188.44 ;
    END
  END Data_HV[282]
  PIN Data_HV[281]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14995.465 187.44 14995.745 188.44 ;
    END
  END Data_HV[281]
  PIN Data_HV[280]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14991.545 187.44 14991.825 188.44 ;
    END
  END Data_HV[280]
  PIN Data_HV[279]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14990.985 187.44 14991.265 188.44 ;
    END
  END Data_HV[279]
  PIN Data_HV[278]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14993.785 187.44 14994.065 188.44 ;
    END
  END Data_HV[278]
  PIN Data_HV[277]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14965.225 187.44 14965.505 188.44 ;
    END
  END Data_HV[277]
  PIN Data_HV[276]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14968.025 187.44 14968.305 188.44 ;
    END
  END Data_HV[276]
  PIN Data_HV[275]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14967.465 187.44 14967.745 188.44 ;
    END
  END Data_HV[275]
  PIN Data_HV[274]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14963.545 187.44 14963.825 188.44 ;
    END
  END Data_HV[274]
  PIN Data_HV[273]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14962.985 187.44 14963.265 188.44 ;
    END
  END Data_HV[273]
  PIN Data_HV[272]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14910.905 187.44 14911.185 188.44 ;
    END
  END Data_HV[272]
  PIN Data_HV[271]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14912.585 187.44 14912.865 188.44 ;
    END
  END Data_HV[271]
  PIN Data_HV[270]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14914.265 187.44 14914.545 188.44 ;
    END
  END Data_HV[270]
  PIN Data_HV[269]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14858.265 187.44 14858.545 188.44 ;
    END
  END Data_HV[269]
  PIN Data_HV[268]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14860.505 187.44 14860.785 188.44 ;
    END
  END Data_HV[268]
  PIN Data_HV[267]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14887.665 187.44 14887.945 188.44 ;
    END
  END Data_HV[267]
  PIN Data_HV[266]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14910.345 187.44 14910.625 188.44 ;
    END
  END Data_HV[266]
  PIN Data_HV[265]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14911.465 187.44 14911.745 188.44 ;
    END
  END Data_HV[265]
  PIN Data_HV[264]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14913.145 187.44 14913.425 188.44 ;
    END
  END Data_HV[264]
  PIN Data_HV[263]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14859.945 187.44 14860.225 188.44 ;
    END
  END Data_HV[263]
  PIN Data_HV[262]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14887.105 187.44 14887.385 188.44 ;
    END
  END Data_HV[262]
  PIN Data_HV[261]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14888.225 187.44 14888.505 188.44 ;
    END
  END Data_HV[261]
  PIN Data_HV[260]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14913.705 187.44 14913.985 188.44 ;
    END
  END Data_HV[260]
  PIN Data_HV[259]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14909.785 187.44 14910.065 188.44 ;
    END
  END Data_HV[259]
  PIN Data_HV[258]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14900.825 187.44 14901.105 188.44 ;
    END
  END Data_HV[258]
  PIN Data_HV[257]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14912.025 187.44 14912.305 188.44 ;
    END
  END Data_HV[257]
  PIN Data_HV[256]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14861.065 187.44 14861.345 188.44 ;
    END
  END Data_HV[256]
  PIN Data_HV[255]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14889.345 187.44 14889.625 188.44 ;
    END
  END Data_HV[255]
  PIN Data_HV[254]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14888.785 187.44 14889.065 188.44 ;
    END
  END Data_HV[254]
  PIN Data_HV[253]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14859.385 187.44 14859.665 188.44 ;
    END
  END Data_HV[253]
  PIN Data_HV[252]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14858.825 187.44 14859.105 188.44 ;
    END
  END Data_HV[252]
  PIN Data_HV[251]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14832.505 187.44 14832.785 188.44 ;
    END
  END Data_HV[251]
  PIN Data_HV[250]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14834.185 187.44 14834.465 188.44 ;
    END
  END Data_HV[250]
  PIN Data_HV[249]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14848.745 187.44 14849.025 188.44 ;
    END
  END Data_HV[249]
  PIN Data_HV[248]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14777.065 187.44 14777.345 188.44 ;
    END
  END Data_HV[248]
  PIN Data_HV[247]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14779.305 187.44 14779.585 188.44 ;
    END
  END Data_HV[247]
  PIN Data_HV[246]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14780.985 187.44 14781.265 188.44 ;
    END
  END Data_HV[246]
  PIN Data_HV[245]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14831.945 187.44 14832.225 188.44 ;
    END
  END Data_HV[245]
  PIN Data_HV[244]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14833.065 187.44 14833.345 188.44 ;
    END
  END Data_HV[244]
  PIN Data_HV[243]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14834.745 187.44 14835.025 188.44 ;
    END
  END Data_HV[243]
  PIN Data_HV[242]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14778.745 187.44 14779.025 188.44 ;
    END
  END Data_HV[242]
  PIN Data_HV[241]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14780.425 187.44 14780.705 188.44 ;
    END
  END Data_HV[241]
  PIN Data_HV[240]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14781.545 187.44 14781.825 188.44 ;
    END
  END Data_HV[240]
  PIN Data_HV[239]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14848.185 187.44 14848.465 188.44 ;
    END
  END Data_HV[239]
  PIN Data_HV[238]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14831.385 187.44 14831.665 188.44 ;
    END
  END Data_HV[238]
  PIN Data_HV[237]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14830.825 187.44 14831.105 188.44 ;
    END
  END Data_HV[237]
  PIN Data_HV[236]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14833.625 187.44 14833.905 188.44 ;
    END
  END Data_HV[236]
  PIN Data_HV[235]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14779.865 187.44 14780.145 188.44 ;
    END
  END Data_HV[235]
  PIN Data_HV[234]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14782.665 187.44 14782.945 188.44 ;
    END
  END Data_HV[234]
  PIN Data_HV[233]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14782.105 187.44 14782.385 188.44 ;
    END
  END Data_HV[233]
  PIN Data_HV[232]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14778.185 187.44 14778.465 188.44 ;
    END
  END Data_HV[232]
  PIN Data_HV[231]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14777.625 187.44 14777.905 188.44 ;
    END
  END Data_HV[231]
  PIN Data_HV[230]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14755.785 187.44 14756.065 188.44 ;
    END
  END Data_HV[230]
  PIN Data_HV[229]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14757.465 187.44 14757.745 188.44 ;
    END
  END Data_HV[229]
  PIN Data_HV[228]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14759.145 187.44 14759.425 188.44 ;
    END
  END Data_HV[228]
  PIN Data_HV[227]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14711.545 187.44 14711.825 188.44 ;
    END
  END Data_HV[227]
  PIN Data_HV[226]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14713.785 187.44 14714.065 188.44 ;
    END
  END Data_HV[226]
  PIN Data_HV[225]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14715.465 187.44 14715.745 188.44 ;
    END
  END Data_HV[225]
  PIN Data_HV[224]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14755.225 187.44 14755.505 188.44 ;
    END
  END Data_HV[224]
  PIN Data_HV[223]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14756.345 187.44 14756.625 188.44 ;
    END
  END Data_HV[223]
  PIN Data_HV[222]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14758.025 187.44 14758.305 188.44 ;
    END
  END Data_HV[222]
  PIN Data_HV[221]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14713.225 187.44 14713.505 188.44 ;
    END
  END Data_HV[221]
  PIN Data_HV[220]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14714.905 187.44 14715.185 188.44 ;
    END
  END Data_HV[220]
  PIN Data_HV[219]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14716.025 187.44 14716.305 188.44 ;
    END
  END Data_HV[219]
  PIN Data_HV[218]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14758.585 187.44 14758.865 188.44 ;
    END
  END Data_HV[218]
  PIN Data_HV[217]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14754.665 187.44 14754.945 188.44 ;
    END
  END Data_HV[217]
  PIN Data_HV[216]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14754.105 187.44 14754.385 188.44 ;
    END
  END Data_HV[216]
  PIN Data_HV[215]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14756.905 187.44 14757.185 188.44 ;
    END
  END Data_HV[215]
  PIN Data_HV[214]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14714.345 187.44 14714.625 188.44 ;
    END
  END Data_HV[214]
  PIN Data_HV[213]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14717.145 187.44 14717.425 188.44 ;
    END
  END Data_HV[213]
  PIN Data_HV[212]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14716.585 187.44 14716.865 188.44 ;
    END
  END Data_HV[212]
  PIN Data_HV[211]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14712.665 187.44 14712.945 188.44 ;
    END
  END Data_HV[211]
  PIN Data_HV[210]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14712.105 187.44 14712.385 188.44 ;
    END
  END Data_HV[210]
  PIN Data_HV[209]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14685.785 187.44 14686.065 188.44 ;
    END
  END Data_HV[209]
  PIN Data_HV[208]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14687.465 187.44 14687.745 188.44 ;
    END
  END Data_HV[208]
  PIN Data_HV[207]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14689.145 187.44 14689.425 188.44 ;
    END
  END Data_HV[207]
  PIN Data_HV[206]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14629.785 187.44 14630.065 188.44 ;
    END
  END Data_HV[206]
  PIN Data_HV[205]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14632.025 187.44 14632.305 188.44 ;
    END
  END Data_HV[205]
  PIN Data_HV[204]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14633.705 187.44 14633.985 188.44 ;
    END
  END Data_HV[204]
  PIN Data_HV[203]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14685.225 187.44 14685.505 188.44 ;
    END
  END Data_HV[203]
  PIN Data_HV[202]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14686.345 187.44 14686.625 188.44 ;
    END
  END Data_HV[202]
  PIN Data_HV[201]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14688.025 187.44 14688.305 188.44 ;
    END
  END Data_HV[201]
  PIN Data_HV[200]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14631.465 187.44 14631.745 188.44 ;
    END
  END Data_HV[200]
  PIN Data_HV[199]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14633.145 187.44 14633.425 188.44 ;
    END
  END Data_HV[199]
  PIN Data_HV[198]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14634.265 187.44 14634.545 188.44 ;
    END
  END Data_HV[198]
  PIN Data_HV[197]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14688.585 187.44 14688.865 188.44 ;
    END
  END Data_HV[197]
  PIN Data_HV[196]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14684.665 187.44 14684.945 188.44 ;
    END
  END Data_HV[196]
  PIN Data_HV[195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14684.105 187.44 14684.385 188.44 ;
    END
  END Data_HV[195]
  PIN Data_HV[194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14686.905 187.44 14687.185 188.44 ;
    END
  END Data_HV[194]
  PIN Data_HV[193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14632.585 187.44 14632.865 188.44 ;
    END
  END Data_HV[193]
  PIN Data_HV[192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14635.385 187.44 14635.665 188.44 ;
    END
  END Data_HV[192]
  PIN Data_HV[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14634.825 187.44 14635.105 188.44 ;
    END
  END Data_HV[191]
  PIN Data_HV[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14630.905 187.44 14631.185 188.44 ;
    END
  END Data_HV[190]
  PIN Data_HV[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14630.345 187.44 14630.625 188.44 ;
    END
  END Data_HV[189]
  PIN Data_HV[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14581.065 187.44 14581.345 188.44 ;
    END
  END Data_HV[188]
  PIN Data_HV[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14608.225 187.44 14608.505 188.44 ;
    END
  END Data_HV[187]
  PIN Data_HV[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14609.905 187.44 14610.185 188.44 ;
    END
  END Data_HV[186]
  PIN Data_HV[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14551.385 187.44 14551.665 188.44 ;
    END
  END Data_HV[185]
  PIN Data_HV[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14553.625 187.44 14553.905 188.44 ;
    END
  END Data_HV[184]
  PIN Data_HV[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14555.305 187.44 14555.585 188.44 ;
    END
  END Data_HV[183]
  PIN Data_HV[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14580.505 187.44 14580.785 188.44 ;
    END
  END Data_HV[182]
  PIN Data_HV[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14581.625 187.44 14581.905 188.44 ;
    END
  END Data_HV[181]
  PIN Data_HV[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14608.785 187.44 14609.065 188.44 ;
    END
  END Data_HV[180]
  PIN Data_HV[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14553.065 187.44 14553.345 188.44 ;
    END
  END Data_HV[179]
  PIN Data_HV[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14554.745 187.44 14555.025 188.44 ;
    END
  END Data_HV[178]
  PIN Data_HV[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14568.745 187.44 14569.025 188.44 ;
    END
  END Data_HV[177]
  PIN Data_HV[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14609.345 187.44 14609.625 188.44 ;
    END
  END Data_HV[176]
  PIN Data_HV[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14579.945 187.44 14580.225 188.44 ;
    END
  END Data_HV[175]
  PIN Data_HV[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14579.385 187.44 14579.665 188.44 ;
    END
  END Data_HV[174]
  PIN Data_HV[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14607.665 187.44 14607.945 188.44 ;
    END
  END Data_HV[173]
  PIN Data_HV[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14554.185 187.44 14554.465 188.44 ;
    END
  END Data_HV[172]
  PIN Data_HV[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14569.865 187.44 14570.145 188.44 ;
    END
  END Data_HV[171]
  PIN Data_HV[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14569.305 187.44 14569.585 188.44 ;
    END
  END Data_HV[170]
  PIN Data_HV[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14552.505 187.44 14552.785 188.44 ;
    END
  END Data_HV[169]
  PIN Data_HV[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14551.945 187.44 14552.225 188.44 ;
    END
  END Data_HV[168]
  PIN Data_HV[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14498.745 187.44 14499.025 188.44 ;
    END
  END Data_HV[167]
  PIN Data_HV[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14500.425 187.44 14500.705 188.44 ;
    END
  END Data_HV[166]
  PIN Data_HV[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14502.105 187.44 14502.385 188.44 ;
    END
  END Data_HV[165]
  PIN Data_HV[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14473.545 187.44 14473.825 188.44 ;
    END
  END Data_HV[164]
  PIN Data_HV[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14475.785 187.44 14476.065 188.44 ;
    END
  END Data_HV[163]
  PIN Data_HV[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14477.465 187.44 14477.745 188.44 ;
    END
  END Data_HV[162]
  PIN Data_HV[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14498.185 187.44 14498.465 188.44 ;
    END
  END Data_HV[161]
  PIN Data_HV[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14499.305 187.44 14499.585 188.44 ;
    END
  END Data_HV[160]
  PIN Data_HV[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14500.985 187.44 14501.265 188.44 ;
    END
  END Data_HV[159]
  PIN Data_HV[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14475.225 187.44 14475.505 188.44 ;
    END
  END Data_HV[158]
  PIN Data_HV[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14476.905 187.44 14477.185 188.44 ;
    END
  END Data_HV[157]
  PIN Data_HV[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14478.025 187.44 14478.305 188.44 ;
    END
  END Data_HV[156]
  PIN Data_HV[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14501.545 187.44 14501.825 188.44 ;
    END
  END Data_HV[155]
  PIN Data_HV[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14497.625 187.44 14497.905 188.44 ;
    END
  END Data_HV[154]
  PIN Data_HV[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14497.065 187.44 14497.345 188.44 ;
    END
  END Data_HV[153]
  PIN Data_HV[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14499.865 187.44 14500.145 188.44 ;
    END
  END Data_HV[152]
  PIN Data_HV[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14476.345 187.44 14476.625 188.44 ;
    END
  END Data_HV[151]
  PIN Data_HV[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14479.145 187.44 14479.425 188.44 ;
    END
  END Data_HV[150]
  PIN Data_HV[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14478.585 187.44 14478.865 188.44 ;
    END
  END Data_HV[149]
  PIN Data_HV[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14474.665 187.44 14474.945 188.44 ;
    END
  END Data_HV[148]
  PIN Data_HV[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14474.105 187.44 14474.385 188.44 ;
    END
  END Data_HV[147]
  PIN Data_HV[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14432.665 187.44 14432.945 188.44 ;
    END
  END Data_HV[146]
  PIN Data_HV[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14434.345 187.44 14434.625 188.44 ;
    END
  END Data_HV[145]
  PIN Data_HV[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14436.025 187.44 14436.305 188.44 ;
    END
  END Data_HV[144]
  PIN Data_HV[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14402.425 187.44 14402.705 188.44 ;
    END
  END Data_HV[143]
  PIN Data_HV[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14404.665 187.44 14404.945 188.44 ;
    END
  END Data_HV[142]
  PIN Data_HV[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14406.345 187.44 14406.625 188.44 ;
    END
  END Data_HV[141]
  PIN Data_HV[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14432.105 187.44 14432.385 188.44 ;
    END
  END Data_HV[140]
  PIN Data_HV[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14433.225 187.44 14433.505 188.44 ;
    END
  END Data_HV[139]
  PIN Data_HV[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14434.905 187.44 14435.185 188.44 ;
    END
  END Data_HV[138]
  PIN Data_HV[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14404.105 187.44 14404.385 188.44 ;
    END
  END Data_HV[137]
  PIN Data_HV[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14405.785 187.44 14406.065 188.44 ;
    END
  END Data_HV[136]
  PIN Data_HV[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14406.905 187.44 14407.185 188.44 ;
    END
  END Data_HV[135]
  PIN Data_HV[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14435.465 187.44 14435.745 188.44 ;
    END
  END Data_HV[134]
  PIN Data_HV[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14431.545 187.44 14431.825 188.44 ;
    END
  END Data_HV[133]
  PIN Data_HV[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14430.985 187.44 14431.265 188.44 ;
    END
  END Data_HV[132]
  PIN Data_HV[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14433.785 187.44 14434.065 188.44 ;
    END
  END Data_HV[131]
  PIN Data_HV[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14405.225 187.44 14405.505 188.44 ;
    END
  END Data_HV[130]
  PIN Data_HV[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14408.025 187.44 14408.305 188.44 ;
    END
  END Data_HV[129]
  PIN Data_HV[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14407.465 187.44 14407.745 188.44 ;
    END
  END Data_HV[128]
  PIN Data_HV[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14403.545 187.44 14403.825 188.44 ;
    END
  END Data_HV[127]
  PIN Data_HV[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14402.985 187.44 14403.265 188.44 ;
    END
  END Data_HV[126]
  PIN Data_HV[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14350.905 187.44 14351.185 188.44 ;
    END
  END Data_HV[125]
  PIN Data_HV[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14352.585 187.44 14352.865 188.44 ;
    END
  END Data_HV[124]
  PIN Data_HV[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14354.265 187.44 14354.545 188.44 ;
    END
  END Data_HV[123]
  PIN Data_HV[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14298.265 187.44 14298.545 188.44 ;
    END
  END Data_HV[122]
  PIN Data_HV[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14300.505 187.44 14300.785 188.44 ;
    END
  END Data_HV[121]
  PIN Data_HV[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14327.665 187.44 14327.945 188.44 ;
    END
  END Data_HV[120]
  PIN Data_HV[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14350.345 187.44 14350.625 188.44 ;
    END
  END Data_HV[119]
  PIN Data_HV[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14351.465 187.44 14351.745 188.44 ;
    END
  END Data_HV[118]
  PIN Data_HV[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14353.145 187.44 14353.425 188.44 ;
    END
  END Data_HV[117]
  PIN Data_HV[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14299.945 187.44 14300.225 188.44 ;
    END
  END Data_HV[116]
  PIN Data_HV[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14327.105 187.44 14327.385 188.44 ;
    END
  END Data_HV[115]
  PIN Data_HV[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14328.225 187.44 14328.505 188.44 ;
    END
  END Data_HV[114]
  PIN Data_HV[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14353.705 187.44 14353.985 188.44 ;
    END
  END Data_HV[113]
  PIN Data_HV[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14349.785 187.44 14350.065 188.44 ;
    END
  END Data_HV[112]
  PIN Data_HV[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14340.825 187.44 14341.105 188.44 ;
    END
  END Data_HV[111]
  PIN Data_HV[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14352.025 187.44 14352.305 188.44 ;
    END
  END Data_HV[110]
  PIN Data_HV[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14301.065 187.44 14301.345 188.44 ;
    END
  END Data_HV[109]
  PIN Data_HV[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14329.345 187.44 14329.625 188.44 ;
    END
  END Data_HV[108]
  PIN Data_HV[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14328.785 187.44 14329.065 188.44 ;
    END
  END Data_HV[107]
  PIN Data_HV[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14299.385 187.44 14299.665 188.44 ;
    END
  END Data_HV[106]
  PIN Data_HV[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14298.825 187.44 14299.105 188.44 ;
    END
  END Data_HV[105]
  PIN Data_HV[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14272.505 187.44 14272.785 188.44 ;
    END
  END Data_HV[104]
  PIN Data_HV[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14274.185 187.44 14274.465 188.44 ;
    END
  END Data_HV[103]
  PIN Data_HV[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14288.745 187.44 14289.025 188.44 ;
    END
  END Data_HV[102]
  PIN Data_HV[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14217.065 187.44 14217.345 188.44 ;
    END
  END Data_HV[101]
  PIN Data_HV[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14219.305 187.44 14219.585 188.44 ;
    END
  END Data_HV[100]
  PIN Data_HV[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14220.985 187.44 14221.265 188.44 ;
    END
  END Data_HV[99]
  PIN Data_HV[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14271.945 187.44 14272.225 188.44 ;
    END
  END Data_HV[98]
  PIN Data_HV[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14273.065 187.44 14273.345 188.44 ;
    END
  END Data_HV[97]
  PIN Data_HV[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14274.745 187.44 14275.025 188.44 ;
    END
  END Data_HV[96]
  PIN Data_HV[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14218.745 187.44 14219.025 188.44 ;
    END
  END Data_HV[95]
  PIN Data_HV[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14220.425 187.44 14220.705 188.44 ;
    END
  END Data_HV[94]
  PIN Data_HV[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14221.545 187.44 14221.825 188.44 ;
    END
  END Data_HV[93]
  PIN Data_HV[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14288.185 187.44 14288.465 188.44 ;
    END
  END Data_HV[92]
  PIN Data_HV[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14271.385 187.44 14271.665 188.44 ;
    END
  END Data_HV[91]
  PIN Data_HV[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14270.825 187.44 14271.105 188.44 ;
    END
  END Data_HV[90]
  PIN Data_HV[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14273.625 187.44 14273.905 188.44 ;
    END
  END Data_HV[89]
  PIN Data_HV[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14219.865 187.44 14220.145 188.44 ;
    END
  END Data_HV[88]
  PIN Data_HV[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14222.665 187.44 14222.945 188.44 ;
    END
  END Data_HV[87]
  PIN Data_HV[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14222.105 187.44 14222.385 188.44 ;
    END
  END Data_HV[86]
  PIN Data_HV[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14218.185 187.44 14218.465 188.44 ;
    END
  END Data_HV[85]
  PIN Data_HV[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14217.625 187.44 14217.905 188.44 ;
    END
  END Data_HV[84]
  PIN Data_HV[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14195.785 187.44 14196.065 188.44 ;
    END
  END Data_HV[83]
  PIN Data_HV[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14197.465 187.44 14197.745 188.44 ;
    END
  END Data_HV[82]
  PIN Data_HV[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14199.145 187.44 14199.425 188.44 ;
    END
  END Data_HV[81]
  PIN Data_HV[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14151.545 187.44 14151.825 188.44 ;
    END
  END Data_HV[80]
  PIN Data_HV[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14153.785 187.44 14154.065 188.44 ;
    END
  END Data_HV[79]
  PIN Data_HV[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14155.465 187.44 14155.745 188.44 ;
    END
  END Data_HV[78]
  PIN Data_HV[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14195.225 187.44 14195.505 188.44 ;
    END
  END Data_HV[77]
  PIN Data_HV[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14196.345 187.44 14196.625 188.44 ;
    END
  END Data_HV[76]
  PIN Data_HV[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14198.025 187.44 14198.305 188.44 ;
    END
  END Data_HV[75]
  PIN Data_HV[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14153.225 187.44 14153.505 188.44 ;
    END
  END Data_HV[74]
  PIN Data_HV[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14154.905 187.44 14155.185 188.44 ;
    END
  END Data_HV[73]
  PIN Data_HV[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14156.025 187.44 14156.305 188.44 ;
    END
  END Data_HV[72]
  PIN Data_HV[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14198.585 187.44 14198.865 188.44 ;
    END
  END Data_HV[71]
  PIN Data_HV[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14194.665 187.44 14194.945 188.44 ;
    END
  END Data_HV[70]
  PIN Data_HV[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14194.105 187.44 14194.385 188.44 ;
    END
  END Data_HV[69]
  PIN Data_HV[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14196.905 187.44 14197.185 188.44 ;
    END
  END Data_HV[68]
  PIN Data_HV[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14154.345 187.44 14154.625 188.44 ;
    END
  END Data_HV[67]
  PIN Data_HV[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14157.145 187.44 14157.425 188.44 ;
    END
  END Data_HV[66]
  PIN Data_HV[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14156.585 187.44 14156.865 188.44 ;
    END
  END Data_HV[65]
  PIN Data_HV[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14152.665 187.44 14152.945 188.44 ;
    END
  END Data_HV[64]
  PIN Data_HV[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14152.105 187.44 14152.385 188.44 ;
    END
  END Data_HV[63]
  PIN Data_HV[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14125.785 187.44 14126.065 188.44 ;
    END
  END Data_HV[62]
  PIN Data_HV[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14127.465 187.44 14127.745 188.44 ;
    END
  END Data_HV[61]
  PIN Data_HV[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14129.145 187.44 14129.425 188.44 ;
    END
  END Data_HV[60]
  PIN Data_HV[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14069.785 187.44 14070.065 188.44 ;
    END
  END Data_HV[59]
  PIN Data_HV[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14072.025 187.44 14072.305 188.44 ;
    END
  END Data_HV[58]
  PIN Data_HV[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14073.705 187.44 14073.985 188.44 ;
    END
  END Data_HV[57]
  PIN Data_HV[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14125.225 187.44 14125.505 188.44 ;
    END
  END Data_HV[56]
  PIN Data_HV[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14126.345 187.44 14126.625 188.44 ;
    END
  END Data_HV[55]
  PIN Data_HV[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14128.025 187.44 14128.305 188.44 ;
    END
  END Data_HV[54]
  PIN Data_HV[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14071.465 187.44 14071.745 188.44 ;
    END
  END Data_HV[53]
  PIN Data_HV[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14073.145 187.44 14073.425 188.44 ;
    END
  END Data_HV[52]
  PIN Data_HV[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14074.265 187.44 14074.545 188.44 ;
    END
  END Data_HV[51]
  PIN Data_HV[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14128.585 187.44 14128.865 188.44 ;
    END
  END Data_HV[50]
  PIN Data_HV[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14124.665 187.44 14124.945 188.44 ;
    END
  END Data_HV[49]
  PIN Data_HV[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14124.105 187.44 14124.385 188.44 ;
    END
  END Data_HV[48]
  PIN Data_HV[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14126.905 187.44 14127.185 188.44 ;
    END
  END Data_HV[47]
  PIN Data_HV[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14072.585 187.44 14072.865 188.44 ;
    END
  END Data_HV[46]
  PIN Data_HV[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14075.385 187.44 14075.665 188.44 ;
    END
  END Data_HV[45]
  PIN Data_HV[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14074.825 187.44 14075.105 188.44 ;
    END
  END Data_HV[44]
  PIN Data_HV[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14070.905 187.44 14071.185 188.44 ;
    END
  END Data_HV[43]
  PIN Data_HV[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14070.345 187.44 14070.625 188.44 ;
    END
  END Data_HV[42]
  PIN Data_HV[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14021.065 187.44 14021.345 188.44 ;
    END
  END Data_HV[41]
  PIN Data_HV[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14048.225 187.44 14048.505 188.44 ;
    END
  END Data_HV[40]
  PIN Data_HV[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14049.905 187.44 14050.185 188.44 ;
    END
  END Data_HV[39]
  PIN Data_HV[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13991.385 187.44 13991.665 188.44 ;
    END
  END Data_HV[38]
  PIN Data_HV[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13993.625 187.44 13993.905 188.44 ;
    END
  END Data_HV[37]
  PIN Data_HV[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13995.305 187.44 13995.585 188.44 ;
    END
  END Data_HV[36]
  PIN Data_HV[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14020.505 187.44 14020.785 188.44 ;
    END
  END Data_HV[35]
  PIN Data_HV[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14021.625 187.44 14021.905 188.44 ;
    END
  END Data_HV[34]
  PIN Data_HV[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14048.785 187.44 14049.065 188.44 ;
    END
  END Data_HV[33]
  PIN Data_HV[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13993.065 187.44 13993.345 188.44 ;
    END
  END Data_HV[32]
  PIN Data_HV[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13994.745 187.44 13995.025 188.44 ;
    END
  END Data_HV[31]
  PIN Data_HV[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14008.745 187.44 14009.025 188.44 ;
    END
  END Data_HV[30]
  PIN Data_HV[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14049.345 187.44 14049.625 188.44 ;
    END
  END Data_HV[29]
  PIN Data_HV[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14019.945 187.44 14020.225 188.44 ;
    END
  END Data_HV[28]
  PIN Data_HV[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14019.385 187.44 14019.665 188.44 ;
    END
  END Data_HV[27]
  PIN Data_HV[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14047.665 187.44 14047.945 188.44 ;
    END
  END Data_HV[26]
  PIN Data_HV[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13994.185 187.44 13994.465 188.44 ;
    END
  END Data_HV[25]
  PIN Data_HV[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14009.865 187.44 14010.145 188.44 ;
    END
  END Data_HV[24]
  PIN Data_HV[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14009.305 187.44 14009.585 188.44 ;
    END
  END Data_HV[23]
  PIN Data_HV[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13992.505 187.44 13992.785 188.44 ;
    END
  END Data_HV[22]
  PIN Data_HV[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13991.945 187.44 13992.225 188.44 ;
    END
  END Data_HV[21]
  PIN Data_HV[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13938.745 187.44 13939.025 188.44 ;
    END
  END Data_HV[20]
  PIN Data_HV[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13940.425 187.44 13940.705 188.44 ;
    END
  END Data_HV[19]
  PIN Data_HV[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13942.105 187.44 13942.385 188.44 ;
    END
  END Data_HV[18]
  PIN Data_HV[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13913.545 187.44 13913.825 188.44 ;
    END
  END Data_HV[17]
  PIN Data_HV[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13915.785 187.44 13916.065 188.44 ;
    END
  END Data_HV[16]
  PIN Data_HV[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13917.465 187.44 13917.745 188.44 ;
    END
  END Data_HV[15]
  PIN Data_HV[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13938.185 187.44 13938.465 188.44 ;
    END
  END Data_HV[14]
  PIN Data_HV[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13939.305 187.44 13939.585 188.44 ;
    END
  END Data_HV[13]
  PIN Data_HV[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13940.985 187.44 13941.265 188.44 ;
    END
  END Data_HV[12]
  PIN Data_HV[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13915.225 187.44 13915.505 188.44 ;
    END
  END Data_HV[11]
  PIN Data_HV[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13916.905 187.44 13917.185 188.44 ;
    END
  END Data_HV[10]
  PIN Data_HV[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13918.025 187.44 13918.305 188.44 ;
    END
  END Data_HV[9]
  PIN Data_HV[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13941.545 187.44 13941.825 188.44 ;
    END
  END Data_HV[8]
  PIN Data_HV[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13937.625 187.44 13937.905 188.44 ;
    END
  END Data_HV[7]
  PIN Data_HV[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13937.065 187.44 13937.345 188.44 ;
    END
  END Data_HV[6]
  PIN Data_HV[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13939.865 187.44 13940.145 188.44 ;
    END
  END Data_HV[5]
  PIN Data_HV[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13916.345 187.44 13916.625 188.44 ;
    END
  END Data_HV[4]
  PIN Data_HV[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13919.145 187.44 13919.425 188.44 ;
    END
  END Data_HV[3]
  PIN Data_HV[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13918.585 187.44 13918.865 188.44 ;
    END
  END Data_HV[2]
  PIN Data_HV[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13914.665 187.44 13914.945 188.44 ;
    END
  END Data_HV[1]
  PIN Data_HV[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13914.105 187.44 13914.385 188.44 ;
    END
  END Data_HV[0]
  PIN nTOK_COMP[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13868.745 187.44 13869.025 188.44 ;
    END
  END nTOK_COMP[55]
  PIN nTOK_COMP[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13778.585 187.44 13778.865 188.44 ;
    END
  END nTOK_COMP[54]
  PIN nTOK_COMP[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13708.585 187.44 13708.865 188.44 ;
    END
  END nTOK_COMP[53]
  PIN nTOK_COMP[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13629.905 187.44 13630.185 188.44 ;
    END
  END nTOK_COMP[52]
  PIN nTOK_COMP[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13522.665 187.44 13522.945 188.44 ;
    END
  END nTOK_COMP[51]
  PIN nTOK_COMP[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13457.145 187.44 13457.425 188.44 ;
    END
  END nTOK_COMP[50]
  PIN nTOK_COMP[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13374.825 187.44 13375.105 188.44 ;
    END
  END nTOK_COMP[49]
  PIN nTOK_COMP[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13308.745 187.44 13309.025 188.44 ;
    END
  END nTOK_COMP[48]
  PIN nTOK_COMP[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13218.585 187.44 13218.865 188.44 ;
    END
  END nTOK_COMP[47]
  PIN nTOK_COMP[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13148.585 187.44 13148.865 188.44 ;
    END
  END nTOK_COMP[46]
  PIN nTOK_COMP[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13069.905 187.44 13070.185 188.44 ;
    END
  END nTOK_COMP[45]
  PIN nTOK_COMP[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12962.665 187.44 12962.945 188.44 ;
    END
  END nTOK_COMP[44]
  PIN nTOK_COMP[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12897.145 187.44 12897.425 188.44 ;
    END
  END nTOK_COMP[43]
  PIN nTOK_COMP[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12814.825 187.44 12815.105 188.44 ;
    END
  END nTOK_COMP[42]
  PIN nTOK_COMP[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12748.745 187.44 12749.025 188.44 ;
    END
  END nTOK_COMP[41]
  PIN nTOK_COMP[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12658.585 187.44 12658.865 188.44 ;
    END
  END nTOK_COMP[40]
  PIN nTOK_COMP[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12588.585 187.44 12588.865 188.44 ;
    END
  END nTOK_COMP[39]
  PIN nTOK_COMP[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12509.905 187.44 12510.185 188.44 ;
    END
  END nTOK_COMP[38]
  PIN nTOK_COMP[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12402.665 187.44 12402.945 188.44 ;
    END
  END nTOK_COMP[37]
  PIN nTOK_COMP[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12337.145 187.44 12337.425 188.44 ;
    END
  END nTOK_COMP[36]
  PIN nTOK_COMP[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12254.825 187.44 12255.105 188.44 ;
    END
  END nTOK_COMP[35]
  PIN nTOK_COMP[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12188.745 187.44 12189.025 188.44 ;
    END
  END nTOK_COMP[34]
  PIN nTOK_COMP[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12098.585 187.44 12098.865 188.44 ;
    END
  END nTOK_COMP[33]
  PIN nTOK_COMP[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12028.585 187.44 12028.865 188.44 ;
    END
  END nTOK_COMP[32]
  PIN nTOK_COMP[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11949.905 187.44 11950.185 188.44 ;
    END
  END nTOK_COMP[31]
  PIN nTOK_COMP[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11842.665 187.44 11842.945 188.44 ;
    END
  END nTOK_COMP[30]
  PIN nTOK_COMP[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11777.145 187.44 11777.425 188.44 ;
    END
  END nTOK_COMP[29]
  PIN nTOK_COMP[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11694.825 187.44 11695.105 188.44 ;
    END
  END nTOK_COMP[28]
  PIN nTOK_COMP[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11628.745 187.44 11629.025 188.44 ;
    END
  END nTOK_COMP[27]
  PIN nTOK_COMP[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11538.585 187.44 11538.865 188.44 ;
    END
  END nTOK_COMP[26]
  PIN nTOK_COMP[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11468.585 187.44 11468.865 188.44 ;
    END
  END nTOK_COMP[25]
  PIN nTOK_COMP[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11389.905 187.44 11390.185 188.44 ;
    END
  END nTOK_COMP[24]
  PIN nTOK_COMP[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11282.665 187.44 11282.945 188.44 ;
    END
  END nTOK_COMP[23]
  PIN nTOK_COMP[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11217.145 187.44 11217.425 188.44 ;
    END
  END nTOK_COMP[22]
  PIN nTOK_COMP[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11134.825 187.44 11135.105 188.44 ;
    END
  END nTOK_COMP[21]
  PIN nTOK_COMP[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11068.745 187.44 11069.025 188.44 ;
    END
  END nTOK_COMP[20]
  PIN nTOK_COMP[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10978.585 187.44 10978.865 188.44 ;
    END
  END nTOK_COMP[19]
  PIN nTOK_COMP[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10908.585 187.44 10908.865 188.44 ;
    END
  END nTOK_COMP[18]
  PIN nTOK_COMP[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10829.905 187.44 10830.185 188.44 ;
    END
  END nTOK_COMP[17]
  PIN nTOK_COMP[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10722.665 187.44 10722.945 188.44 ;
    END
  END nTOK_COMP[16]
  PIN nTOK_COMP[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10657.145 187.44 10657.425 188.44 ;
    END
  END nTOK_COMP[15]
  PIN nTOK_COMP[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10574.825 187.44 10575.105 188.44 ;
    END
  END nTOK_COMP[14]
  PIN nTOK_COMP[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10508.745 187.44 10509.025 188.44 ;
    END
  END nTOK_COMP[13]
  PIN nTOK_COMP[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10418.585 187.44 10418.865 188.44 ;
    END
  END nTOK_COMP[12]
  PIN nTOK_COMP[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10348.585 187.44 10348.865 188.44 ;
    END
  END nTOK_COMP[11]
  PIN nTOK_COMP[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10269.905 187.44 10270.185 188.44 ;
    END
  END nTOK_COMP[10]
  PIN nTOK_COMP[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10162.665 187.44 10162.945 188.44 ;
    END
  END nTOK_COMP[9]
  PIN nTOK_COMP[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10097.145 187.44 10097.425 188.44 ;
    END
  END nTOK_COMP[8]
  PIN nTOK_COMP[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10014.825 187.44 10015.105 188.44 ;
    END
  END nTOK_COMP[7]
  PIN nTOK_COMP[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9948.745 187.44 9949.025 188.44 ;
    END
  END nTOK_COMP[6]
  PIN nTOK_COMP[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9858.585 187.44 9858.865 188.44 ;
    END
  END nTOK_COMP[5]
  PIN nTOK_COMP[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9788.585 187.44 9788.865 188.44 ;
    END
  END nTOK_COMP[4]
  PIN nTOK_COMP[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9709.905 187.44 9710.185 188.44 ;
    END
  END nTOK_COMP[3]
  PIN nTOK_COMP[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9602.665 187.44 9602.945 188.44 ;
    END
  END nTOK_COMP[2]
  PIN nTOK_COMP[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9537.145 187.44 9537.425 188.44 ;
    END
  END nTOK_COMP[1]
  PIN nTOK_COMP[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9454.825 187.44 9455.105 188.44 ;
    END
  END nTOK_COMP[0]
  PIN nTOK_HV[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18348.745 187.44 18349.025 188.44 ;
    END
  END nTOK_HV[55]
  PIN nTOK_HV[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18258.585 187.44 18258.865 188.44 ;
    END
  END nTOK_HV[54]
  PIN nTOK_HV[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18188.585 187.44 18188.865 188.44 ;
    END
  END nTOK_HV[53]
  PIN nTOK_HV[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18109.905 187.44 18110.185 188.44 ;
    END
  END nTOK_HV[52]
  PIN nTOK_HV[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18002.665 187.44 18002.945 188.44 ;
    END
  END nTOK_HV[51]
  PIN nTOK_HV[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17937.145 187.44 17937.425 188.44 ;
    END
  END nTOK_HV[50]
  PIN nTOK_HV[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17854.825 187.44 17855.105 188.44 ;
    END
  END nTOK_HV[49]
  PIN nTOK_HV[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17788.745 187.44 17789.025 188.44 ;
    END
  END nTOK_HV[48]
  PIN nTOK_HV[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17698.585 187.44 17698.865 188.44 ;
    END
  END nTOK_HV[47]
  PIN nTOK_HV[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17628.585 187.44 17628.865 188.44 ;
    END
  END nTOK_HV[46]
  PIN nTOK_HV[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17549.905 187.44 17550.185 188.44 ;
    END
  END nTOK_HV[45]
  PIN nTOK_HV[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17442.665 187.44 17442.945 188.44 ;
    END
  END nTOK_HV[44]
  PIN nTOK_HV[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17377.145 187.44 17377.425 188.44 ;
    END
  END nTOK_HV[43]
  PIN nTOK_HV[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17294.825 187.44 17295.105 188.44 ;
    END
  END nTOK_HV[42]
  PIN nTOK_HV[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17228.745 187.44 17229.025 188.44 ;
    END
  END nTOK_HV[41]
  PIN nTOK_HV[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17138.585 187.44 17138.865 188.44 ;
    END
  END nTOK_HV[40]
  PIN nTOK_HV[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17068.585 187.44 17068.865 188.44 ;
    END
  END nTOK_HV[39]
  PIN nTOK_HV[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16989.905 187.44 16990.185 188.44 ;
    END
  END nTOK_HV[38]
  PIN nTOK_HV[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16882.665 187.44 16882.945 188.44 ;
    END
  END nTOK_HV[37]
  PIN nTOK_HV[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16817.145 187.44 16817.425 188.44 ;
    END
  END nTOK_HV[36]
  PIN nTOK_HV[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16734.825 187.44 16735.105 188.44 ;
    END
  END nTOK_HV[35]
  PIN nTOK_HV[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16668.745 187.44 16669.025 188.44 ;
    END
  END nTOK_HV[34]
  PIN nTOK_HV[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16578.585 187.44 16578.865 188.44 ;
    END
  END nTOK_HV[33]
  PIN nTOK_HV[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16508.585 187.44 16508.865 188.44 ;
    END
  END nTOK_HV[32]
  PIN nTOK_HV[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16429.905 187.44 16430.185 188.44 ;
    END
  END nTOK_HV[31]
  PIN nTOK_HV[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16322.665 187.44 16322.945 188.44 ;
    END
  END nTOK_HV[30]
  PIN nTOK_HV[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16257.145 187.44 16257.425 188.44 ;
    END
  END nTOK_HV[29]
  PIN nTOK_HV[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16174.825 187.44 16175.105 188.44 ;
    END
  END nTOK_HV[28]
  PIN nTOK_HV[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16108.745 187.44 16109.025 188.44 ;
    END
  END nTOK_HV[27]
  PIN nTOK_HV[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16018.585 187.44 16018.865 188.44 ;
    END
  END nTOK_HV[26]
  PIN nTOK_HV[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15948.585 187.44 15948.865 188.44 ;
    END
  END nTOK_HV[25]
  PIN nTOK_HV[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15869.905 187.44 15870.185 188.44 ;
    END
  END nTOK_HV[24]
  PIN nTOK_HV[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15762.665 187.44 15762.945 188.44 ;
    END
  END nTOK_HV[23]
  PIN nTOK_HV[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15697.145 187.44 15697.425 188.44 ;
    END
  END nTOK_HV[22]
  PIN nTOK_HV[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15614.825 187.44 15615.105 188.44 ;
    END
  END nTOK_HV[21]
  PIN nTOK_HV[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15548.745 187.44 15549.025 188.44 ;
    END
  END nTOK_HV[20]
  PIN nTOK_HV[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15458.585 187.44 15458.865 188.44 ;
    END
  END nTOK_HV[19]
  PIN nTOK_HV[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15388.585 187.44 15388.865 188.44 ;
    END
  END nTOK_HV[18]
  PIN nTOK_HV[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15309.905 187.44 15310.185 188.44 ;
    END
  END nTOK_HV[17]
  PIN nTOK_HV[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15202.665 187.44 15202.945 188.44 ;
    END
  END nTOK_HV[16]
  PIN nTOK_HV[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15137.145 187.44 15137.425 188.44 ;
    END
  END nTOK_HV[15]
  PIN nTOK_HV[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15054.825 187.44 15055.105 188.44 ;
    END
  END nTOK_HV[14]
  PIN nTOK_HV[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14988.745 187.44 14989.025 188.44 ;
    END
  END nTOK_HV[13]
  PIN nTOK_HV[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14898.585 187.44 14898.865 188.44 ;
    END
  END nTOK_HV[12]
  PIN nTOK_HV[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14828.585 187.44 14828.865 188.44 ;
    END
  END nTOK_HV[11]
  PIN nTOK_HV[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14749.905 187.44 14750.185 188.44 ;
    END
  END nTOK_HV[10]
  PIN nTOK_HV[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14642.665 187.44 14642.945 188.44 ;
    END
  END nTOK_HV[9]
  PIN nTOK_HV[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14577.145 187.44 14577.425 188.44 ;
    END
  END nTOK_HV[8]
  PIN nTOK_HV[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14494.825 187.44 14495.105 188.44 ;
    END
  END nTOK_HV[7]
  PIN nTOK_HV[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14428.745 187.44 14429.025 188.44 ;
    END
  END nTOK_HV[6]
  PIN nTOK_HV[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14338.585 187.44 14338.865 188.44 ;
    END
  END nTOK_HV[5]
  PIN nTOK_HV[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14268.585 187.44 14268.865 188.44 ;
    END
  END nTOK_HV[4]
  PIN nTOK_HV[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14189.905 187.44 14190.185 188.44 ;
    END
  END nTOK_HV[3]
  PIN nTOK_HV[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14082.665 187.44 14082.945 188.44 ;
    END
  END nTOK_HV[2]
  PIN nTOK_HV[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14017.145 187.44 14017.425 188.44 ;
    END
  END nTOK_HV[1]
  PIN nTOK_HV[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13934.825 187.44 13935.105 188.44 ;
    END
  END nTOK_HV[0]
  PIN OUTA_MON_L[3]
    DIRECTION OUTPUT ;
    USE ANALOG ;
    PORT
      LAYER M4 ;
        RECT 326.66 8582.095 327.66 8583.515 ;
    END
  END OUTA_MON_L[3]
  PIN OUTA_MON_L[2]
    DIRECTION OUTPUT ;
    USE ANALOG ;
    PORT
      LAYER M4 ;
        RECT 326.66 8543.58 327.66 8545 ;
    END
  END OUTA_MON_L[2]
  PIN OUTA_MON_L[1]
    DIRECTION OUTPUT ;
    USE ANALOG ;
    PORT
      LAYER M4 ;
        RECT 326.66 8510.095 327.66 8511.515 ;
    END
  END OUTA_MON_L[1]
  PIN OUTA_MON_L[0]
    DIRECTION OUTPUT ;
    USE ANALOG ;
    PORT
      LAYER M4 ;
        RECT 326.66 8471.58 327.66 8473 ;
    END
  END OUTA_MON_L[0]
  PIN OUTA_MON_R[3]
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER M4 ;
        RECT 18489.46 8582.095 18490.46 8583.515 ;
    END
  END OUTA_MON_R[3]
  PIN OUTA_MON_R[2]
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER M4 ;
        RECT 18489.46 8543.58 18490.46 8545 ;
    END
  END OUTA_MON_R[2]
  PIN OUTA_MON_R[1]
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER M4 ;
        RECT 18489.46 8510.095 18490.46 8511.515 ;
    END
  END OUTA_MON_R[1]
  PIN OUTA_MON_R[0]
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER M4 ;
        RECT 18489.46 8471.58 18490.46 8473 ;
    END
  END OUTA_MON_R[0]
  PIN DIG_MON_PMOS[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9398.265 187.44 9398.545 188.44 ;
    END
  END DIG_MON_PMOS[111]
  PIN DIG_MON_PMOS[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9320.985 187.44 9321.265 188.44 ;
    END
  END DIG_MON_PMOS[110]
  PIN DIG_MON_PMOS[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9316.505 187.44 9316.785 188.44 ;
    END
  END DIG_MON_PMOS[109]
  PIN DIG_MON_PMOS[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9255.465 187.44 9255.745 188.44 ;
    END
  END DIG_MON_PMOS[108]
  PIN DIG_MON_PMOS[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9250.985 187.44 9251.265 188.44 ;
    END
  END DIG_MON_PMOS[107]
  PIN DIG_MON_PMOS[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9174.265 187.44 9174.545 188.44 ;
    END
  END DIG_MON_PMOS[106]
  PIN DIG_MON_PMOS[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9169.785 187.44 9170.065 188.44 ;
    END
  END DIG_MON_PMOS[105]
  PIN DIG_MON_PMOS[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9108.745 187.44 9109.025 188.44 ;
    END
  END DIG_MON_PMOS[104]
  PIN DIG_MON_PMOS[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9091.385 187.44 9091.665 188.44 ;
    END
  END DIG_MON_PMOS[103]
  PIN DIG_MON_PMOS[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9018.585 187.44 9018.865 188.44 ;
    END
  END DIG_MON_PMOS[102]
  PIN DIG_MON_PMOS[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9014.105 187.44 9014.385 188.44 ;
    END
  END DIG_MON_PMOS[101]
  PIN DIG_MON_PMOS[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8948.585 187.44 8948.865 188.44 ;
    END
  END DIG_MON_PMOS[100]
  PIN DIG_MON_PMOS[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8944.105 187.44 8944.385 188.44 ;
    END
  END DIG_MON_PMOS[99]
  PIN DIG_MON_PMOS[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8868.785 187.44 8869.065 188.44 ;
    END
  END DIG_MON_PMOS[98]
  PIN DIG_MON_PMOS[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8838.265 187.44 8838.545 188.44 ;
    END
  END DIG_MON_PMOS[97]
  PIN DIG_MON_PMOS[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8760.985 187.44 8761.265 188.44 ;
    END
  END DIG_MON_PMOS[96]
  PIN DIG_MON_PMOS[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8756.505 187.44 8756.785 188.44 ;
    END
  END DIG_MON_PMOS[95]
  PIN DIG_MON_PMOS[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8695.465 187.44 8695.745 188.44 ;
    END
  END DIG_MON_PMOS[94]
  PIN DIG_MON_PMOS[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8690.985 187.44 8691.265 188.44 ;
    END
  END DIG_MON_PMOS[93]
  PIN DIG_MON_PMOS[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8614.265 187.44 8614.545 188.44 ;
    END
  END DIG_MON_PMOS[92]
  PIN DIG_MON_PMOS[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8609.785 187.44 8610.065 188.44 ;
    END
  END DIG_MON_PMOS[91]
  PIN DIG_MON_PMOS[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8548.745 187.44 8549.025 188.44 ;
    END
  END DIG_MON_PMOS[90]
  PIN DIG_MON_PMOS[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8531.385 187.44 8531.665 188.44 ;
    END
  END DIG_MON_PMOS[89]
  PIN DIG_MON_PMOS[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8458.585 187.44 8458.865 188.44 ;
    END
  END DIG_MON_PMOS[88]
  PIN DIG_MON_PMOS[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8454.105 187.44 8454.385 188.44 ;
    END
  END DIG_MON_PMOS[87]
  PIN DIG_MON_PMOS[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8388.585 187.44 8388.865 188.44 ;
    END
  END DIG_MON_PMOS[86]
  PIN DIG_MON_PMOS[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8384.105 187.44 8384.385 188.44 ;
    END
  END DIG_MON_PMOS[85]
  PIN DIG_MON_PMOS[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8308.785 187.44 8309.065 188.44 ;
    END
  END DIG_MON_PMOS[84]
  PIN DIG_MON_PMOS[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8278.265 187.44 8278.545 188.44 ;
    END
  END DIG_MON_PMOS[83]
  PIN DIG_MON_PMOS[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8200.985 187.44 8201.265 188.44 ;
    END
  END DIG_MON_PMOS[82]
  PIN DIG_MON_PMOS[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8196.505 187.44 8196.785 188.44 ;
    END
  END DIG_MON_PMOS[81]
  PIN DIG_MON_PMOS[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8135.465 187.44 8135.745 188.44 ;
    END
  END DIG_MON_PMOS[80]
  PIN DIG_MON_PMOS[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8130.985 187.44 8131.265 188.44 ;
    END
  END DIG_MON_PMOS[79]
  PIN DIG_MON_PMOS[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8054.265 187.44 8054.545 188.44 ;
    END
  END DIG_MON_PMOS[78]
  PIN DIG_MON_PMOS[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8049.785 187.44 8050.065 188.44 ;
    END
  END DIG_MON_PMOS[77]
  PIN DIG_MON_PMOS[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7988.745 187.44 7989.025 188.44 ;
    END
  END DIG_MON_PMOS[76]
  PIN DIG_MON_PMOS[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7971.385 187.44 7971.665 188.44 ;
    END
  END DIG_MON_PMOS[75]
  PIN DIG_MON_PMOS[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7898.585 187.44 7898.865 188.44 ;
    END
  END DIG_MON_PMOS[74]
  PIN DIG_MON_PMOS[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7894.105 187.44 7894.385 188.44 ;
    END
  END DIG_MON_PMOS[73]
  PIN DIG_MON_PMOS[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7828.585 187.44 7828.865 188.44 ;
    END
  END DIG_MON_PMOS[72]
  PIN DIG_MON_PMOS[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7824.105 187.44 7824.385 188.44 ;
    END
  END DIG_MON_PMOS[71]
  PIN DIG_MON_PMOS[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7748.785 187.44 7749.065 188.44 ;
    END
  END DIG_MON_PMOS[70]
  PIN DIG_MON_PMOS[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7718.265 187.44 7718.545 188.44 ;
    END
  END DIG_MON_PMOS[69]
  PIN DIG_MON_PMOS[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7640.985 187.44 7641.265 188.44 ;
    END
  END DIG_MON_PMOS[68]
  PIN DIG_MON_PMOS[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7636.505 187.44 7636.785 188.44 ;
    END
  END DIG_MON_PMOS[67]
  PIN DIG_MON_PMOS[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7575.465 187.44 7575.745 188.44 ;
    END
  END DIG_MON_PMOS[66]
  PIN DIG_MON_PMOS[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7570.985 187.44 7571.265 188.44 ;
    END
  END DIG_MON_PMOS[65]
  PIN DIG_MON_PMOS[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7494.265 187.44 7494.545 188.44 ;
    END
  END DIG_MON_PMOS[64]
  PIN DIG_MON_PMOS[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7489.785 187.44 7490.065 188.44 ;
    END
  END DIG_MON_PMOS[63]
  PIN DIG_MON_PMOS[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7428.745 187.44 7429.025 188.44 ;
    END
  END DIG_MON_PMOS[62]
  PIN DIG_MON_PMOS[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7411.385 187.44 7411.665 188.44 ;
    END
  END DIG_MON_PMOS[61]
  PIN DIG_MON_PMOS[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7338.585 187.44 7338.865 188.44 ;
    END
  END DIG_MON_PMOS[60]
  PIN DIG_MON_PMOS[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7334.105 187.44 7334.385 188.44 ;
    END
  END DIG_MON_PMOS[59]
  PIN DIG_MON_PMOS[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7268.585 187.44 7268.865 188.44 ;
    END
  END DIG_MON_PMOS[58]
  PIN DIG_MON_PMOS[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7264.105 187.44 7264.385 188.44 ;
    END
  END DIG_MON_PMOS[57]
  PIN DIG_MON_PMOS[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7188.785 187.44 7189.065 188.44 ;
    END
  END DIG_MON_PMOS[56]
  PIN DIG_MON_PMOS[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7158.265 187.44 7158.545 188.44 ;
    END
  END DIG_MON_PMOS[55]
  PIN DIG_MON_PMOS[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7080.985 187.44 7081.265 188.44 ;
    END
  END DIG_MON_PMOS[54]
  PIN DIG_MON_PMOS[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7076.505 187.44 7076.785 188.44 ;
    END
  END DIG_MON_PMOS[53]
  PIN DIG_MON_PMOS[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7015.465 187.44 7015.745 188.44 ;
    END
  END DIG_MON_PMOS[52]
  PIN DIG_MON_PMOS[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7010.985 187.44 7011.265 188.44 ;
    END
  END DIG_MON_PMOS[51]
  PIN DIG_MON_PMOS[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6934.265 187.44 6934.545 188.44 ;
    END
  END DIG_MON_PMOS[50]
  PIN DIG_MON_PMOS[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6929.785 187.44 6930.065 188.44 ;
    END
  END DIG_MON_PMOS[49]
  PIN DIG_MON_PMOS[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6868.745 187.44 6869.025 188.44 ;
    END
  END DIG_MON_PMOS[48]
  PIN DIG_MON_PMOS[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6851.385 187.44 6851.665 188.44 ;
    END
  END DIG_MON_PMOS[47]
  PIN DIG_MON_PMOS[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6778.585 187.44 6778.865 188.44 ;
    END
  END DIG_MON_PMOS[46]
  PIN DIG_MON_PMOS[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6774.105 187.44 6774.385 188.44 ;
    END
  END DIG_MON_PMOS[45]
  PIN DIG_MON_PMOS[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6708.585 187.44 6708.865 188.44 ;
    END
  END DIG_MON_PMOS[44]
  PIN DIG_MON_PMOS[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6704.105 187.44 6704.385 188.44 ;
    END
  END DIG_MON_PMOS[43]
  PIN DIG_MON_PMOS[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6628.785 187.44 6629.065 188.44 ;
    END
  END DIG_MON_PMOS[42]
  PIN DIG_MON_PMOS[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6598.265 187.44 6598.545 188.44 ;
    END
  END DIG_MON_PMOS[41]
  PIN DIG_MON_PMOS[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6520.985 187.44 6521.265 188.44 ;
    END
  END DIG_MON_PMOS[40]
  PIN DIG_MON_PMOS[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6516.505 187.44 6516.785 188.44 ;
    END
  END DIG_MON_PMOS[39]
  PIN DIG_MON_PMOS[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6455.465 187.44 6455.745 188.44 ;
    END
  END DIG_MON_PMOS[38]
  PIN DIG_MON_PMOS[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6450.985 187.44 6451.265 188.44 ;
    END
  END DIG_MON_PMOS[37]
  PIN DIG_MON_PMOS[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6374.265 187.44 6374.545 188.44 ;
    END
  END DIG_MON_PMOS[36]
  PIN DIG_MON_PMOS[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6369.785 187.44 6370.065 188.44 ;
    END
  END DIG_MON_PMOS[35]
  PIN DIG_MON_PMOS[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6308.745 187.44 6309.025 188.44 ;
    END
  END DIG_MON_PMOS[34]
  PIN DIG_MON_PMOS[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6291.385 187.44 6291.665 188.44 ;
    END
  END DIG_MON_PMOS[33]
  PIN DIG_MON_PMOS[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6218.585 187.44 6218.865 188.44 ;
    END
  END DIG_MON_PMOS[32]
  PIN DIG_MON_PMOS[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6214.105 187.44 6214.385 188.44 ;
    END
  END DIG_MON_PMOS[31]
  PIN DIG_MON_PMOS[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6148.585 187.44 6148.865 188.44 ;
    END
  END DIG_MON_PMOS[30]
  PIN DIG_MON_PMOS[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6144.105 187.44 6144.385 188.44 ;
    END
  END DIG_MON_PMOS[29]
  PIN DIG_MON_PMOS[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6068.785 187.44 6069.065 188.44 ;
    END
  END DIG_MON_PMOS[28]
  PIN DIG_MON_PMOS[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6038.265 187.44 6038.545 188.44 ;
    END
  END DIG_MON_PMOS[27]
  PIN DIG_MON_PMOS[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5960.985 187.44 5961.265 188.44 ;
    END
  END DIG_MON_PMOS[26]
  PIN DIG_MON_PMOS[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5956.505 187.44 5956.785 188.44 ;
    END
  END DIG_MON_PMOS[25]
  PIN DIG_MON_PMOS[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5895.465 187.44 5895.745 188.44 ;
    END
  END DIG_MON_PMOS[24]
  PIN DIG_MON_PMOS[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5890.985 187.44 5891.265 188.44 ;
    END
  END DIG_MON_PMOS[23]
  PIN DIG_MON_PMOS[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5814.265 187.44 5814.545 188.44 ;
    END
  END DIG_MON_PMOS[22]
  PIN DIG_MON_PMOS[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5809.785 187.44 5810.065 188.44 ;
    END
  END DIG_MON_PMOS[21]
  PIN DIG_MON_PMOS[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5748.745 187.44 5749.025 188.44 ;
    END
  END DIG_MON_PMOS[20]
  PIN DIG_MON_PMOS[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5731.385 187.44 5731.665 188.44 ;
    END
  END DIG_MON_PMOS[19]
  PIN DIG_MON_PMOS[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5658.585 187.44 5658.865 188.44 ;
    END
  END DIG_MON_PMOS[18]
  PIN DIG_MON_PMOS[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5654.105 187.44 5654.385 188.44 ;
    END
  END DIG_MON_PMOS[17]
  PIN DIG_MON_PMOS[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5588.585 187.44 5588.865 188.44 ;
    END
  END DIG_MON_PMOS[16]
  PIN DIG_MON_PMOS[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5584.105 187.44 5584.385 188.44 ;
    END
  END DIG_MON_PMOS[15]
  PIN DIG_MON_PMOS[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5508.785 187.44 5509.065 188.44 ;
    END
  END DIG_MON_PMOS[14]
  PIN DIG_MON_PMOS[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5478.265 187.44 5478.545 188.44 ;
    END
  END DIG_MON_PMOS[13]
  PIN DIG_MON_PMOS[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5400.985 187.44 5401.265 188.44 ;
    END
  END DIG_MON_PMOS[12]
  PIN DIG_MON_PMOS[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5396.505 187.44 5396.785 188.44 ;
    END
  END DIG_MON_PMOS[11]
  PIN DIG_MON_PMOS[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5335.465 187.44 5335.745 188.44 ;
    END
  END DIG_MON_PMOS[10]
  PIN DIG_MON_PMOS[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5330.985 187.44 5331.265 188.44 ;
    END
  END DIG_MON_PMOS[9]
  PIN DIG_MON_PMOS[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5254.265 187.44 5254.545 188.44 ;
    END
  END DIG_MON_PMOS[8]
  PIN DIG_MON_PMOS[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5249.785 187.44 5250.065 188.44 ;
    END
  END DIG_MON_PMOS[7]
  PIN DIG_MON_PMOS[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5188.745 187.44 5189.025 188.44 ;
    END
  END DIG_MON_PMOS[6]
  PIN DIG_MON_PMOS[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5171.385 187.44 5171.665 188.44 ;
    END
  END DIG_MON_PMOS[5]
  PIN DIG_MON_PMOS[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5098.585 187.44 5098.865 188.44 ;
    END
  END DIG_MON_PMOS[4]
  PIN DIG_MON_PMOS[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5094.105 187.44 5094.385 188.44 ;
    END
  END DIG_MON_PMOS[3]
  PIN DIG_MON_PMOS[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5028.585 187.44 5028.865 188.44 ;
    END
  END DIG_MON_PMOS[2]
  PIN DIG_MON_PMOS[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5024.105 187.44 5024.385 188.44 ;
    END
  END DIG_MON_PMOS[1]
  PIN DIG_MON_PMOS[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4948.785 187.44 4949.065 188.44 ;
    END
  END DIG_MON_PMOS[0]
  PIN DIG_MON_COMP[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13878.265 187.44 13878.545 188.44 ;
    END
  END DIG_MON_COMP[111]
  PIN DIG_MON_COMP[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13800.985 187.44 13801.265 188.44 ;
    END
  END DIG_MON_COMP[110]
  PIN DIG_MON_COMP[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13796.505 187.44 13796.785 188.44 ;
    END
  END DIG_MON_COMP[109]
  PIN DIG_MON_COMP[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13735.465 187.44 13735.745 188.44 ;
    END
  END DIG_MON_COMP[108]
  PIN DIG_MON_COMP[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13730.985 187.44 13731.265 188.44 ;
    END
  END DIG_MON_COMP[107]
  PIN DIG_MON_COMP[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13654.265 187.44 13654.545 188.44 ;
    END
  END DIG_MON_COMP[106]
  PIN DIG_MON_COMP[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13649.785 187.44 13650.065 188.44 ;
    END
  END DIG_MON_COMP[105]
  PIN DIG_MON_COMP[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13588.745 187.44 13589.025 188.44 ;
    END
  END DIG_MON_COMP[104]
  PIN DIG_MON_COMP[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13571.385 187.44 13571.665 188.44 ;
    END
  END DIG_MON_COMP[103]
  PIN DIG_MON_COMP[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13498.585 187.44 13498.865 188.44 ;
    END
  END DIG_MON_COMP[102]
  PIN DIG_MON_COMP[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13494.105 187.44 13494.385 188.44 ;
    END
  END DIG_MON_COMP[101]
  PIN DIG_MON_COMP[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13428.585 187.44 13428.865 188.44 ;
    END
  END DIG_MON_COMP[100]
  PIN DIG_MON_COMP[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13424.105 187.44 13424.385 188.44 ;
    END
  END DIG_MON_COMP[99]
  PIN DIG_MON_COMP[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13348.785 187.44 13349.065 188.44 ;
    END
  END DIG_MON_COMP[98]
  PIN DIG_MON_COMP[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13318.265 187.44 13318.545 188.44 ;
    END
  END DIG_MON_COMP[97]
  PIN DIG_MON_COMP[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13240.985 187.44 13241.265 188.44 ;
    END
  END DIG_MON_COMP[96]
  PIN DIG_MON_COMP[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13236.505 187.44 13236.785 188.44 ;
    END
  END DIG_MON_COMP[95]
  PIN DIG_MON_COMP[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13175.465 187.44 13175.745 188.44 ;
    END
  END DIG_MON_COMP[94]
  PIN DIG_MON_COMP[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13170.985 187.44 13171.265 188.44 ;
    END
  END DIG_MON_COMP[93]
  PIN DIG_MON_COMP[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13094.265 187.44 13094.545 188.44 ;
    END
  END DIG_MON_COMP[92]
  PIN DIG_MON_COMP[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13089.785 187.44 13090.065 188.44 ;
    END
  END DIG_MON_COMP[91]
  PIN DIG_MON_COMP[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13028.745 187.44 13029.025 188.44 ;
    END
  END DIG_MON_COMP[90]
  PIN DIG_MON_COMP[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13011.385 187.44 13011.665 188.44 ;
    END
  END DIG_MON_COMP[89]
  PIN DIG_MON_COMP[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12938.585 187.44 12938.865 188.44 ;
    END
  END DIG_MON_COMP[88]
  PIN DIG_MON_COMP[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12934.105 187.44 12934.385 188.44 ;
    END
  END DIG_MON_COMP[87]
  PIN DIG_MON_COMP[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12868.585 187.44 12868.865 188.44 ;
    END
  END DIG_MON_COMP[86]
  PIN DIG_MON_COMP[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12864.105 187.44 12864.385 188.44 ;
    END
  END DIG_MON_COMP[85]
  PIN DIG_MON_COMP[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12788.785 187.44 12789.065 188.44 ;
    END
  END DIG_MON_COMP[84]
  PIN DIG_MON_COMP[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12758.265 187.44 12758.545 188.44 ;
    END
  END DIG_MON_COMP[83]
  PIN DIG_MON_COMP[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12680.985 187.44 12681.265 188.44 ;
    END
  END DIG_MON_COMP[82]
  PIN DIG_MON_COMP[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12676.505 187.44 12676.785 188.44 ;
    END
  END DIG_MON_COMP[81]
  PIN DIG_MON_COMP[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12615.465 187.44 12615.745 188.44 ;
    END
  END DIG_MON_COMP[80]
  PIN DIG_MON_COMP[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12610.985 187.44 12611.265 188.44 ;
    END
  END DIG_MON_COMP[79]
  PIN DIG_MON_COMP[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12534.265 187.44 12534.545 188.44 ;
    END
  END DIG_MON_COMP[78]
  PIN DIG_MON_COMP[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12529.785 187.44 12530.065 188.44 ;
    END
  END DIG_MON_COMP[77]
  PIN DIG_MON_COMP[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12468.745 187.44 12469.025 188.44 ;
    END
  END DIG_MON_COMP[76]
  PIN DIG_MON_COMP[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12451.385 187.44 12451.665 188.44 ;
    END
  END DIG_MON_COMP[75]
  PIN DIG_MON_COMP[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12378.585 187.44 12378.865 188.44 ;
    END
  END DIG_MON_COMP[74]
  PIN DIG_MON_COMP[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12374.105 187.44 12374.385 188.44 ;
    END
  END DIG_MON_COMP[73]
  PIN DIG_MON_COMP[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12308.585 187.44 12308.865 188.44 ;
    END
  END DIG_MON_COMP[72]
  PIN DIG_MON_COMP[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12304.105 187.44 12304.385 188.44 ;
    END
  END DIG_MON_COMP[71]
  PIN DIG_MON_COMP[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12228.785 187.44 12229.065 188.44 ;
    END
  END DIG_MON_COMP[70]
  PIN DIG_MON_COMP[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12198.265 187.44 12198.545 188.44 ;
    END
  END DIG_MON_COMP[69]
  PIN DIG_MON_COMP[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12120.985 187.44 12121.265 188.44 ;
    END
  END DIG_MON_COMP[68]
  PIN DIG_MON_COMP[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12116.505 187.44 12116.785 188.44 ;
    END
  END DIG_MON_COMP[67]
  PIN DIG_MON_COMP[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12055.465 187.44 12055.745 188.44 ;
    END
  END DIG_MON_COMP[66]
  PIN DIG_MON_COMP[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12050.985 187.44 12051.265 188.44 ;
    END
  END DIG_MON_COMP[65]
  PIN DIG_MON_COMP[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11974.265 187.44 11974.545 188.44 ;
    END
  END DIG_MON_COMP[64]
  PIN DIG_MON_COMP[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11969.785 187.44 11970.065 188.44 ;
    END
  END DIG_MON_COMP[63]
  PIN DIG_MON_COMP[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11908.745 187.44 11909.025 188.44 ;
    END
  END DIG_MON_COMP[62]
  PIN DIG_MON_COMP[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11891.385 187.44 11891.665 188.44 ;
    END
  END DIG_MON_COMP[61]
  PIN DIG_MON_COMP[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11818.585 187.44 11818.865 188.44 ;
    END
  END DIG_MON_COMP[60]
  PIN DIG_MON_COMP[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11814.105 187.44 11814.385 188.44 ;
    END
  END DIG_MON_COMP[59]
  PIN DIG_MON_COMP[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11748.585 187.44 11748.865 188.44 ;
    END
  END DIG_MON_COMP[58]
  PIN DIG_MON_COMP[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11744.105 187.44 11744.385 188.44 ;
    END
  END DIG_MON_COMP[57]
  PIN DIG_MON_COMP[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11668.785 187.44 11669.065 188.44 ;
    END
  END DIG_MON_COMP[56]
  PIN DIG_MON_COMP[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11638.265 187.44 11638.545 188.44 ;
    END
  END DIG_MON_COMP[55]
  PIN DIG_MON_COMP[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11560.985 187.44 11561.265 188.44 ;
    END
  END DIG_MON_COMP[54]
  PIN DIG_MON_COMP[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11556.505 187.44 11556.785 188.44 ;
    END
  END DIG_MON_COMP[53]
  PIN DIG_MON_COMP[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11495.465 187.44 11495.745 188.44 ;
    END
  END DIG_MON_COMP[52]
  PIN DIG_MON_COMP[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11490.985 187.44 11491.265 188.44 ;
    END
  END DIG_MON_COMP[51]
  PIN DIG_MON_COMP[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11414.265 187.44 11414.545 188.44 ;
    END
  END DIG_MON_COMP[50]
  PIN DIG_MON_COMP[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11409.785 187.44 11410.065 188.44 ;
    END
  END DIG_MON_COMP[49]
  PIN DIG_MON_COMP[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11348.745 187.44 11349.025 188.44 ;
    END
  END DIG_MON_COMP[48]
  PIN DIG_MON_COMP[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11331.385 187.44 11331.665 188.44 ;
    END
  END DIG_MON_COMP[47]
  PIN DIG_MON_COMP[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11258.585 187.44 11258.865 188.44 ;
    END
  END DIG_MON_COMP[46]
  PIN DIG_MON_COMP[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11254.105 187.44 11254.385 188.44 ;
    END
  END DIG_MON_COMP[45]
  PIN DIG_MON_COMP[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11188.585 187.44 11188.865 188.44 ;
    END
  END DIG_MON_COMP[44]
  PIN DIG_MON_COMP[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11184.105 187.44 11184.385 188.44 ;
    END
  END DIG_MON_COMP[43]
  PIN DIG_MON_COMP[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11108.785 187.44 11109.065 188.44 ;
    END
  END DIG_MON_COMP[42]
  PIN DIG_MON_COMP[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11078.265 187.44 11078.545 188.44 ;
    END
  END DIG_MON_COMP[41]
  PIN DIG_MON_COMP[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11000.985 187.44 11001.265 188.44 ;
    END
  END DIG_MON_COMP[40]
  PIN DIG_MON_COMP[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10996.505 187.44 10996.785 188.44 ;
    END
  END DIG_MON_COMP[39]
  PIN DIG_MON_COMP[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10935.465 187.44 10935.745 188.44 ;
    END
  END DIG_MON_COMP[38]
  PIN DIG_MON_COMP[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10930.985 187.44 10931.265 188.44 ;
    END
  END DIG_MON_COMP[37]
  PIN DIG_MON_COMP[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10854.265 187.44 10854.545 188.44 ;
    END
  END DIG_MON_COMP[36]
  PIN DIG_MON_COMP[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10849.785 187.44 10850.065 188.44 ;
    END
  END DIG_MON_COMP[35]
  PIN DIG_MON_COMP[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10788.745 187.44 10789.025 188.44 ;
    END
  END DIG_MON_COMP[34]
  PIN DIG_MON_COMP[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10771.385 187.44 10771.665 188.44 ;
    END
  END DIG_MON_COMP[33]
  PIN DIG_MON_COMP[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10698.585 187.44 10698.865 188.44 ;
    END
  END DIG_MON_COMP[32]
  PIN DIG_MON_COMP[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10694.105 187.44 10694.385 188.44 ;
    END
  END DIG_MON_COMP[31]
  PIN DIG_MON_COMP[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10628.585 187.44 10628.865 188.44 ;
    END
  END DIG_MON_COMP[30]
  PIN DIG_MON_COMP[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10624.105 187.44 10624.385 188.44 ;
    END
  END DIG_MON_COMP[29]
  PIN DIG_MON_COMP[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10548.785 187.44 10549.065 188.44 ;
    END
  END DIG_MON_COMP[28]
  PIN DIG_MON_COMP[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10518.265 187.44 10518.545 188.44 ;
    END
  END DIG_MON_COMP[27]
  PIN DIG_MON_COMP[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10440.985 187.44 10441.265 188.44 ;
    END
  END DIG_MON_COMP[26]
  PIN DIG_MON_COMP[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10436.505 187.44 10436.785 188.44 ;
    END
  END DIG_MON_COMP[25]
  PIN DIG_MON_COMP[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10375.465 187.44 10375.745 188.44 ;
    END
  END DIG_MON_COMP[24]
  PIN DIG_MON_COMP[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10370.985 187.44 10371.265 188.44 ;
    END
  END DIG_MON_COMP[23]
  PIN DIG_MON_COMP[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10294.265 187.44 10294.545 188.44 ;
    END
  END DIG_MON_COMP[22]
  PIN DIG_MON_COMP[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10289.785 187.44 10290.065 188.44 ;
    END
  END DIG_MON_COMP[21]
  PIN DIG_MON_COMP[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10228.745 187.44 10229.025 188.44 ;
    END
  END DIG_MON_COMP[20]
  PIN DIG_MON_COMP[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10211.385 187.44 10211.665 188.44 ;
    END
  END DIG_MON_COMP[19]
  PIN DIG_MON_COMP[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10138.585 187.44 10138.865 188.44 ;
    END
  END DIG_MON_COMP[18]
  PIN DIG_MON_COMP[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10134.105 187.44 10134.385 188.44 ;
    END
  END DIG_MON_COMP[17]
  PIN DIG_MON_COMP[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10068.585 187.44 10068.865 188.44 ;
    END
  END DIG_MON_COMP[16]
  PIN DIG_MON_COMP[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10064.105 187.44 10064.385 188.44 ;
    END
  END DIG_MON_COMP[15]
  PIN DIG_MON_COMP[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9988.785 187.44 9989.065 188.44 ;
    END
  END DIG_MON_COMP[14]
  PIN DIG_MON_COMP[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9958.265 187.44 9958.545 188.44 ;
    END
  END DIG_MON_COMP[13]
  PIN DIG_MON_COMP[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9880.985 187.44 9881.265 188.44 ;
    END
  END DIG_MON_COMP[12]
  PIN DIG_MON_COMP[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9876.505 187.44 9876.785 188.44 ;
    END
  END DIG_MON_COMP[11]
  PIN DIG_MON_COMP[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9815.465 187.44 9815.745 188.44 ;
    END
  END DIG_MON_COMP[10]
  PIN DIG_MON_COMP[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9810.985 187.44 9811.265 188.44 ;
    END
  END DIG_MON_COMP[9]
  PIN DIG_MON_COMP[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9734.265 187.44 9734.545 188.44 ;
    END
  END DIG_MON_COMP[8]
  PIN DIG_MON_COMP[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9729.785 187.44 9730.065 188.44 ;
    END
  END DIG_MON_COMP[7]
  PIN DIG_MON_COMP[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9668.745 187.44 9669.025 188.44 ;
    END
  END DIG_MON_COMP[6]
  PIN DIG_MON_COMP[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9651.385 187.44 9651.665 188.44 ;
    END
  END DIG_MON_COMP[5]
  PIN DIG_MON_COMP[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9578.585 187.44 9578.865 188.44 ;
    END
  END DIG_MON_COMP[4]
  PIN DIG_MON_COMP[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9574.105 187.44 9574.385 188.44 ;
    END
  END DIG_MON_COMP[3]
  PIN DIG_MON_COMP[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9508.585 187.44 9508.865 188.44 ;
    END
  END DIG_MON_COMP[2]
  PIN DIG_MON_COMP[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9504.105 187.44 9504.385 188.44 ;
    END
  END DIG_MON_COMP[1]
  PIN DIG_MON_COMP[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9428.785 187.44 9429.065 188.44 ;
    END
  END DIG_MON_COMP[0]
  PIN DIG_MON_HV[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18358.265 187.44 18358.545 188.44 ;
    END
  END DIG_MON_HV[111]
  PIN DIG_MON_HV[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18280.985 187.44 18281.265 188.44 ;
    END
  END DIG_MON_HV[110]
  PIN DIG_MON_HV[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18276.505 187.44 18276.785 188.44 ;
    END
  END DIG_MON_HV[109]
  PIN DIG_MON_HV[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18215.465 187.44 18215.745 188.44 ;
    END
  END DIG_MON_HV[108]
  PIN DIG_MON_HV[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18210.985 187.44 18211.265 188.44 ;
    END
  END DIG_MON_HV[107]
  PIN DIG_MON_HV[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18134.265 187.44 18134.545 188.44 ;
    END
  END DIG_MON_HV[106]
  PIN DIG_MON_HV[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18129.785 187.44 18130.065 188.44 ;
    END
  END DIG_MON_HV[105]
  PIN DIG_MON_HV[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18068.745 187.44 18069.025 188.44 ;
    END
  END DIG_MON_HV[104]
  PIN DIG_MON_HV[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18051.385 187.44 18051.665 188.44 ;
    END
  END DIG_MON_HV[103]
  PIN DIG_MON_HV[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17978.585 187.44 17978.865 188.44 ;
    END
  END DIG_MON_HV[102]
  PIN DIG_MON_HV[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17974.105 187.44 17974.385 188.44 ;
    END
  END DIG_MON_HV[101]
  PIN DIG_MON_HV[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17908.585 187.44 17908.865 188.44 ;
    END
  END DIG_MON_HV[100]
  PIN DIG_MON_HV[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17904.105 187.44 17904.385 188.44 ;
    END
  END DIG_MON_HV[99]
  PIN DIG_MON_HV[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17828.785 187.44 17829.065 188.44 ;
    END
  END DIG_MON_HV[98]
  PIN DIG_MON_HV[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17798.265 187.44 17798.545 188.44 ;
    END
  END DIG_MON_HV[97]
  PIN DIG_MON_HV[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17720.985 187.44 17721.265 188.44 ;
    END
  END DIG_MON_HV[96]
  PIN DIG_MON_HV[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17716.505 187.44 17716.785 188.44 ;
    END
  END DIG_MON_HV[95]
  PIN DIG_MON_HV[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17655.465 187.44 17655.745 188.44 ;
    END
  END DIG_MON_HV[94]
  PIN DIG_MON_HV[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17650.985 187.44 17651.265 188.44 ;
    END
  END DIG_MON_HV[93]
  PIN DIG_MON_HV[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17574.265 187.44 17574.545 188.44 ;
    END
  END DIG_MON_HV[92]
  PIN DIG_MON_HV[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17569.785 187.44 17570.065 188.44 ;
    END
  END DIG_MON_HV[91]
  PIN DIG_MON_HV[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17508.745 187.44 17509.025 188.44 ;
    END
  END DIG_MON_HV[90]
  PIN DIG_MON_HV[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17491.385 187.44 17491.665 188.44 ;
    END
  END DIG_MON_HV[89]
  PIN DIG_MON_HV[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17418.585 187.44 17418.865 188.44 ;
    END
  END DIG_MON_HV[88]
  PIN DIG_MON_HV[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17414.105 187.44 17414.385 188.44 ;
    END
  END DIG_MON_HV[87]
  PIN DIG_MON_HV[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17348.585 187.44 17348.865 188.44 ;
    END
  END DIG_MON_HV[86]
  PIN DIG_MON_HV[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17344.105 187.44 17344.385 188.44 ;
    END
  END DIG_MON_HV[85]
  PIN DIG_MON_HV[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17268.785 187.44 17269.065 188.44 ;
    END
  END DIG_MON_HV[84]
  PIN DIG_MON_HV[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17238.265 187.44 17238.545 188.44 ;
    END
  END DIG_MON_HV[83]
  PIN DIG_MON_HV[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17160.985 187.44 17161.265 188.44 ;
    END
  END DIG_MON_HV[82]
  PIN DIG_MON_HV[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17156.505 187.44 17156.785 188.44 ;
    END
  END DIG_MON_HV[81]
  PIN DIG_MON_HV[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17095.465 187.44 17095.745 188.44 ;
    END
  END DIG_MON_HV[80]
  PIN DIG_MON_HV[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17090.985 187.44 17091.265 188.44 ;
    END
  END DIG_MON_HV[79]
  PIN DIG_MON_HV[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17014.265 187.44 17014.545 188.44 ;
    END
  END DIG_MON_HV[78]
  PIN DIG_MON_HV[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17009.785 187.44 17010.065 188.44 ;
    END
  END DIG_MON_HV[77]
  PIN DIG_MON_HV[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16948.745 187.44 16949.025 188.44 ;
    END
  END DIG_MON_HV[76]
  PIN DIG_MON_HV[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16931.385 187.44 16931.665 188.44 ;
    END
  END DIG_MON_HV[75]
  PIN DIG_MON_HV[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16858.585 187.44 16858.865 188.44 ;
    END
  END DIG_MON_HV[74]
  PIN DIG_MON_HV[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16854.105 187.44 16854.385 188.44 ;
    END
  END DIG_MON_HV[73]
  PIN DIG_MON_HV[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16788.585 187.44 16788.865 188.44 ;
    END
  END DIG_MON_HV[72]
  PIN DIG_MON_HV[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16784.105 187.44 16784.385 188.44 ;
    END
  END DIG_MON_HV[71]
  PIN DIG_MON_HV[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16708.785 187.44 16709.065 188.44 ;
    END
  END DIG_MON_HV[70]
  PIN DIG_MON_HV[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16678.265 187.44 16678.545 188.44 ;
    END
  END DIG_MON_HV[69]
  PIN DIG_MON_HV[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16600.985 187.44 16601.265 188.44 ;
    END
  END DIG_MON_HV[68]
  PIN DIG_MON_HV[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16596.505 187.44 16596.785 188.44 ;
    END
  END DIG_MON_HV[67]
  PIN DIG_MON_HV[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16535.465 187.44 16535.745 188.44 ;
    END
  END DIG_MON_HV[66]
  PIN DIG_MON_HV[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16530.985 187.44 16531.265 188.44 ;
    END
  END DIG_MON_HV[65]
  PIN DIG_MON_HV[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16454.265 187.44 16454.545 188.44 ;
    END
  END DIG_MON_HV[64]
  PIN DIG_MON_HV[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16449.785 187.44 16450.065 188.44 ;
    END
  END DIG_MON_HV[63]
  PIN DIG_MON_HV[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16388.745 187.44 16389.025 188.44 ;
    END
  END DIG_MON_HV[62]
  PIN DIG_MON_HV[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16371.385 187.44 16371.665 188.44 ;
    END
  END DIG_MON_HV[61]
  PIN DIG_MON_HV[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16298.585 187.44 16298.865 188.44 ;
    END
  END DIG_MON_HV[60]
  PIN DIG_MON_HV[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16294.105 187.44 16294.385 188.44 ;
    END
  END DIG_MON_HV[59]
  PIN DIG_MON_HV[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16228.585 187.44 16228.865 188.44 ;
    END
  END DIG_MON_HV[58]
  PIN DIG_MON_HV[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16224.105 187.44 16224.385 188.44 ;
    END
  END DIG_MON_HV[57]
  PIN DIG_MON_HV[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16148.785 187.44 16149.065 188.44 ;
    END
  END DIG_MON_HV[56]
  PIN DIG_MON_HV[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16118.265 187.44 16118.545 188.44 ;
    END
  END DIG_MON_HV[55]
  PIN DIG_MON_HV[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16040.985 187.44 16041.265 188.44 ;
    END
  END DIG_MON_HV[54]
  PIN DIG_MON_HV[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16036.505 187.44 16036.785 188.44 ;
    END
  END DIG_MON_HV[53]
  PIN DIG_MON_HV[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15975.465 187.44 15975.745 188.44 ;
    END
  END DIG_MON_HV[52]
  PIN DIG_MON_HV[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15970.985 187.44 15971.265 188.44 ;
    END
  END DIG_MON_HV[51]
  PIN DIG_MON_HV[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15894.265 187.44 15894.545 188.44 ;
    END
  END DIG_MON_HV[50]
  PIN DIG_MON_HV[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15889.785 187.44 15890.065 188.44 ;
    END
  END DIG_MON_HV[49]
  PIN DIG_MON_HV[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15828.745 187.44 15829.025 188.44 ;
    END
  END DIG_MON_HV[48]
  PIN DIG_MON_HV[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15811.385 187.44 15811.665 188.44 ;
    END
  END DIG_MON_HV[47]
  PIN DIG_MON_HV[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15738.585 187.44 15738.865 188.44 ;
    END
  END DIG_MON_HV[46]
  PIN DIG_MON_HV[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15734.105 187.44 15734.385 188.44 ;
    END
  END DIG_MON_HV[45]
  PIN DIG_MON_HV[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15668.585 187.44 15668.865 188.44 ;
    END
  END DIG_MON_HV[44]
  PIN DIG_MON_HV[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15664.105 187.44 15664.385 188.44 ;
    END
  END DIG_MON_HV[43]
  PIN DIG_MON_HV[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15588.785 187.44 15589.065 188.44 ;
    END
  END DIG_MON_HV[42]
  PIN DIG_MON_HV[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15558.265 187.44 15558.545 188.44 ;
    END
  END DIG_MON_HV[41]
  PIN DIG_MON_HV[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15480.985 187.44 15481.265 188.44 ;
    END
  END DIG_MON_HV[40]
  PIN DIG_MON_HV[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15476.505 187.44 15476.785 188.44 ;
    END
  END DIG_MON_HV[39]
  PIN DIG_MON_HV[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15415.465 187.44 15415.745 188.44 ;
    END
  END DIG_MON_HV[38]
  PIN DIG_MON_HV[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15410.985 187.44 15411.265 188.44 ;
    END
  END DIG_MON_HV[37]
  PIN DIG_MON_HV[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15334.265 187.44 15334.545 188.44 ;
    END
  END DIG_MON_HV[36]
  PIN DIG_MON_HV[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15329.785 187.44 15330.065 188.44 ;
    END
  END DIG_MON_HV[35]
  PIN DIG_MON_HV[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15268.745 187.44 15269.025 188.44 ;
    END
  END DIG_MON_HV[34]
  PIN DIG_MON_HV[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15251.385 187.44 15251.665 188.44 ;
    END
  END DIG_MON_HV[33]
  PIN DIG_MON_HV[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15178.585 187.44 15178.865 188.44 ;
    END
  END DIG_MON_HV[32]
  PIN DIG_MON_HV[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15174.105 187.44 15174.385 188.44 ;
    END
  END DIG_MON_HV[31]
  PIN DIG_MON_HV[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15108.585 187.44 15108.865 188.44 ;
    END
  END DIG_MON_HV[30]
  PIN DIG_MON_HV[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15104.105 187.44 15104.385 188.44 ;
    END
  END DIG_MON_HV[29]
  PIN DIG_MON_HV[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15028.785 187.44 15029.065 188.44 ;
    END
  END DIG_MON_HV[28]
  PIN DIG_MON_HV[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14998.265 187.44 14998.545 188.44 ;
    END
  END DIG_MON_HV[27]
  PIN DIG_MON_HV[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14920.985 187.44 14921.265 188.44 ;
    END
  END DIG_MON_HV[26]
  PIN DIG_MON_HV[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14916.505 187.44 14916.785 188.44 ;
    END
  END DIG_MON_HV[25]
  PIN DIG_MON_HV[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14855.465 187.44 14855.745 188.44 ;
    END
  END DIG_MON_HV[24]
  PIN DIG_MON_HV[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14850.985 187.44 14851.265 188.44 ;
    END
  END DIG_MON_HV[23]
  PIN DIG_MON_HV[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14774.265 187.44 14774.545 188.44 ;
    END
  END DIG_MON_HV[22]
  PIN DIG_MON_HV[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14769.785 187.44 14770.065 188.44 ;
    END
  END DIG_MON_HV[21]
  PIN DIG_MON_HV[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14708.745 187.44 14709.025 188.44 ;
    END
  END DIG_MON_HV[20]
  PIN DIG_MON_HV[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14691.385 187.44 14691.665 188.44 ;
    END
  END DIG_MON_HV[19]
  PIN DIG_MON_HV[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14618.585 187.44 14618.865 188.44 ;
    END
  END DIG_MON_HV[18]
  PIN DIG_MON_HV[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14614.105 187.44 14614.385 188.44 ;
    END
  END DIG_MON_HV[17]
  PIN DIG_MON_HV[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14548.585 187.44 14548.865 188.44 ;
    END
  END DIG_MON_HV[16]
  PIN DIG_MON_HV[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14544.105 187.44 14544.385 188.44 ;
    END
  END DIG_MON_HV[15]
  PIN DIG_MON_HV[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14468.785 187.44 14469.065 188.44 ;
    END
  END DIG_MON_HV[14]
  PIN DIG_MON_HV[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14438.265 187.44 14438.545 188.44 ;
    END
  END DIG_MON_HV[13]
  PIN DIG_MON_HV[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14360.985 187.44 14361.265 188.44 ;
    END
  END DIG_MON_HV[12]
  PIN DIG_MON_HV[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14356.505 187.44 14356.785 188.44 ;
    END
  END DIG_MON_HV[11]
  PIN DIG_MON_HV[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14295.465 187.44 14295.745 188.44 ;
    END
  END DIG_MON_HV[10]
  PIN DIG_MON_HV[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14290.985 187.44 14291.265 188.44 ;
    END
  END DIG_MON_HV[9]
  PIN DIG_MON_HV[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14214.265 187.44 14214.545 188.44 ;
    END
  END DIG_MON_HV[8]
  PIN DIG_MON_HV[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14209.785 187.44 14210.065 188.44 ;
    END
  END DIG_MON_HV[7]
  PIN DIG_MON_HV[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14148.745 187.44 14149.025 188.44 ;
    END
  END DIG_MON_HV[6]
  PIN DIG_MON_HV[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14131.385 187.44 14131.665 188.44 ;
    END
  END DIG_MON_HV[5]
  PIN DIG_MON_HV[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14058.585 187.44 14058.865 188.44 ;
    END
  END DIG_MON_HV[4]
  PIN DIG_MON_HV[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14054.105 187.44 14054.385 188.44 ;
    END
  END DIG_MON_HV[3]
  PIN DIG_MON_HV[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13988.585 187.44 13988.865 188.44 ;
    END
  END DIG_MON_HV[2]
  PIN DIG_MON_HV[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13984.105 187.44 13984.385 188.44 ;
    END
  END DIG_MON_HV[1]
  PIN DIG_MON_HV[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13908.785 187.44 13909.065 188.44 ;
    END
  END DIG_MON_HV[0]
  PIN BiasSF
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 18489.46 508.445 18490.46 509.445 ;
    END
  END BiasSF
  PIN INJ_IN_MON_L
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 466.545 187.44 466.825 188.44 ;
    END
  END INJ_IN_MON_L
  PIN INJ_IN_MON_R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18361.065 187.44 18361.345 188.44 ;
    END
  END INJ_IN_MON_R
  PIN INJ_IN[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13869.865 187.44 13870.145 188.44 ;
    END
  END INJ_IN[335]
  PIN INJ_IN[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13849.145 187.44 13849.425 188.44 ;
    END
  END INJ_IN[334]
  PIN INJ_IN[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13779.705 187.44 13779.985 188.44 ;
    END
  END INJ_IN[333]
  PIN INJ_IN[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13770.465 187.44 13770.745 188.44 ;
    END
  END INJ_IN[332]
  PIN INJ_IN[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13709.705 187.44 13709.985 188.44 ;
    END
  END INJ_IN[331]
  PIN INJ_IN[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13702.425 187.44 13702.705 188.44 ;
    END
  END INJ_IN[330]
  PIN INJ_IN[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13631.025 187.44 13631.305 188.44 ;
    END
  END INJ_IN[329]
  PIN INJ_IN[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13598.265 187.44 13598.545 188.44 ;
    END
  END INJ_IN[328]
  PIN INJ_IN[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13562.985 187.44 13563.265 188.44 ;
    END
  END INJ_IN[327]
  PIN INJ_IN[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13516.505 187.44 13516.785 188.44 ;
    END
  END INJ_IN[326]
  PIN INJ_IN[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13458.265 187.44 13458.545 188.44 ;
    END
  END INJ_IN[325]
  PIN INJ_IN[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13450.985 187.44 13451.265 188.44 ;
    END
  END INJ_IN[324]
  PIN INJ_IN[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13375.945 187.44 13376.225 188.44 ;
    END
  END INJ_IN[323]
  PIN INJ_IN[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13360.265 187.44 13360.545 188.44 ;
    END
  END INJ_IN[322]
  PIN INJ_IN[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13309.865 187.44 13310.145 188.44 ;
    END
  END INJ_IN[321]
  PIN INJ_IN[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13289.145 187.44 13289.425 188.44 ;
    END
  END INJ_IN[320]
  PIN INJ_IN[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13219.705 187.44 13219.985 188.44 ;
    END
  END INJ_IN[319]
  PIN INJ_IN[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13210.465 187.44 13210.745 188.44 ;
    END
  END INJ_IN[318]
  PIN INJ_IN[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13149.705 187.44 13149.985 188.44 ;
    END
  END INJ_IN[317]
  PIN INJ_IN[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13142.425 187.44 13142.705 188.44 ;
    END
  END INJ_IN[316]
  PIN INJ_IN[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13071.025 187.44 13071.305 188.44 ;
    END
  END INJ_IN[315]
  PIN INJ_IN[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13038.265 187.44 13038.545 188.44 ;
    END
  END INJ_IN[314]
  PIN INJ_IN[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13002.985 187.44 13003.265 188.44 ;
    END
  END INJ_IN[313]
  PIN INJ_IN[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12956.505 187.44 12956.785 188.44 ;
    END
  END INJ_IN[312]
  PIN INJ_IN[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12898.265 187.44 12898.545 188.44 ;
    END
  END INJ_IN[311]
  PIN INJ_IN[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12890.985 187.44 12891.265 188.44 ;
    END
  END INJ_IN[310]
  PIN INJ_IN[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12815.945 187.44 12816.225 188.44 ;
    END
  END INJ_IN[309]
  PIN INJ_IN[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12800.265 187.44 12800.545 188.44 ;
    END
  END INJ_IN[308]
  PIN INJ_IN[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12749.865 187.44 12750.145 188.44 ;
    END
  END INJ_IN[307]
  PIN INJ_IN[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12729.145 187.44 12729.425 188.44 ;
    END
  END INJ_IN[306]
  PIN INJ_IN[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12659.705 187.44 12659.985 188.44 ;
    END
  END INJ_IN[305]
  PIN INJ_IN[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12650.465 187.44 12650.745 188.44 ;
    END
  END INJ_IN[304]
  PIN INJ_IN[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12589.705 187.44 12589.985 188.44 ;
    END
  END INJ_IN[303]
  PIN INJ_IN[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12582.425 187.44 12582.705 188.44 ;
    END
  END INJ_IN[302]
  PIN INJ_IN[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12511.025 187.44 12511.305 188.44 ;
    END
  END INJ_IN[301]
  PIN INJ_IN[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12478.265 187.44 12478.545 188.44 ;
    END
  END INJ_IN[300]
  PIN INJ_IN[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12442.985 187.44 12443.265 188.44 ;
    END
  END INJ_IN[299]
  PIN INJ_IN[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12396.505 187.44 12396.785 188.44 ;
    END
  END INJ_IN[298]
  PIN INJ_IN[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12338.265 187.44 12338.545 188.44 ;
    END
  END INJ_IN[297]
  PIN INJ_IN[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12330.985 187.44 12331.265 188.44 ;
    END
  END INJ_IN[296]
  PIN INJ_IN[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12255.945 187.44 12256.225 188.44 ;
    END
  END INJ_IN[295]
  PIN INJ_IN[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12240.265 187.44 12240.545 188.44 ;
    END
  END INJ_IN[294]
  PIN INJ_IN[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12189.865 187.44 12190.145 188.44 ;
    END
  END INJ_IN[293]
  PIN INJ_IN[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12169.145 187.44 12169.425 188.44 ;
    END
  END INJ_IN[292]
  PIN INJ_IN[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12099.705 187.44 12099.985 188.44 ;
    END
  END INJ_IN[291]
  PIN INJ_IN[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12090.465 187.44 12090.745 188.44 ;
    END
  END INJ_IN[290]
  PIN INJ_IN[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12029.705 187.44 12029.985 188.44 ;
    END
  END INJ_IN[289]
  PIN INJ_IN[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12022.425 187.44 12022.705 188.44 ;
    END
  END INJ_IN[288]
  PIN INJ_IN[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11951.025 187.44 11951.305 188.44 ;
    END
  END INJ_IN[287]
  PIN INJ_IN[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11918.265 187.44 11918.545 188.44 ;
    END
  END INJ_IN[286]
  PIN INJ_IN[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11882.985 187.44 11883.265 188.44 ;
    END
  END INJ_IN[285]
  PIN INJ_IN[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11836.505 187.44 11836.785 188.44 ;
    END
  END INJ_IN[284]
  PIN INJ_IN[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11778.265 187.44 11778.545 188.44 ;
    END
  END INJ_IN[283]
  PIN INJ_IN[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11770.985 187.44 11771.265 188.44 ;
    END
  END INJ_IN[282]
  PIN INJ_IN[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11695.945 187.44 11696.225 188.44 ;
    END
  END INJ_IN[281]
  PIN INJ_IN[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11680.265 187.44 11680.545 188.44 ;
    END
  END INJ_IN[280]
  PIN INJ_IN[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11629.865 187.44 11630.145 188.44 ;
    END
  END INJ_IN[279]
  PIN INJ_IN[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11609.145 187.44 11609.425 188.44 ;
    END
  END INJ_IN[278]
  PIN INJ_IN[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11539.705 187.44 11539.985 188.44 ;
    END
  END INJ_IN[277]
  PIN INJ_IN[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11530.465 187.44 11530.745 188.44 ;
    END
  END INJ_IN[276]
  PIN INJ_IN[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11469.705 187.44 11469.985 188.44 ;
    END
  END INJ_IN[275]
  PIN INJ_IN[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11462.425 187.44 11462.705 188.44 ;
    END
  END INJ_IN[274]
  PIN INJ_IN[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11391.025 187.44 11391.305 188.44 ;
    END
  END INJ_IN[273]
  PIN INJ_IN[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11358.265 187.44 11358.545 188.44 ;
    END
  END INJ_IN[272]
  PIN INJ_IN[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11322.985 187.44 11323.265 188.44 ;
    END
  END INJ_IN[271]
  PIN INJ_IN[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11276.505 187.44 11276.785 188.44 ;
    END
  END INJ_IN[270]
  PIN INJ_IN[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11218.265 187.44 11218.545 188.44 ;
    END
  END INJ_IN[269]
  PIN INJ_IN[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11210.985 187.44 11211.265 188.44 ;
    END
  END INJ_IN[268]
  PIN INJ_IN[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11135.945 187.44 11136.225 188.44 ;
    END
  END INJ_IN[267]
  PIN INJ_IN[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11120.265 187.44 11120.545 188.44 ;
    END
  END INJ_IN[266]
  PIN INJ_IN[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11069.865 187.44 11070.145 188.44 ;
    END
  END INJ_IN[265]
  PIN INJ_IN[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11049.145 187.44 11049.425 188.44 ;
    END
  END INJ_IN[264]
  PIN INJ_IN[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10979.705 187.44 10979.985 188.44 ;
    END
  END INJ_IN[263]
  PIN INJ_IN[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10970.465 187.44 10970.745 188.44 ;
    END
  END INJ_IN[262]
  PIN INJ_IN[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10909.705 187.44 10909.985 188.44 ;
    END
  END INJ_IN[261]
  PIN INJ_IN[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10902.425 187.44 10902.705 188.44 ;
    END
  END INJ_IN[260]
  PIN INJ_IN[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10831.025 187.44 10831.305 188.44 ;
    END
  END INJ_IN[259]
  PIN INJ_IN[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10798.265 187.44 10798.545 188.44 ;
    END
  END INJ_IN[258]
  PIN INJ_IN[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10762.985 187.44 10763.265 188.44 ;
    END
  END INJ_IN[257]
  PIN INJ_IN[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10716.505 187.44 10716.785 188.44 ;
    END
  END INJ_IN[256]
  PIN INJ_IN[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10658.265 187.44 10658.545 188.44 ;
    END
  END INJ_IN[255]
  PIN INJ_IN[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10650.985 187.44 10651.265 188.44 ;
    END
  END INJ_IN[254]
  PIN INJ_IN[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10575.945 187.44 10576.225 188.44 ;
    END
  END INJ_IN[253]
  PIN INJ_IN[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10560.265 187.44 10560.545 188.44 ;
    END
  END INJ_IN[252]
  PIN INJ_IN[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10509.865 187.44 10510.145 188.44 ;
    END
  END INJ_IN[251]
  PIN INJ_IN[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10489.145 187.44 10489.425 188.44 ;
    END
  END INJ_IN[250]
  PIN INJ_IN[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10419.705 187.44 10419.985 188.44 ;
    END
  END INJ_IN[249]
  PIN INJ_IN[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10410.465 187.44 10410.745 188.44 ;
    END
  END INJ_IN[248]
  PIN INJ_IN[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10349.705 187.44 10349.985 188.44 ;
    END
  END INJ_IN[247]
  PIN INJ_IN[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10342.425 187.44 10342.705 188.44 ;
    END
  END INJ_IN[246]
  PIN INJ_IN[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10271.025 187.44 10271.305 188.44 ;
    END
  END INJ_IN[245]
  PIN INJ_IN[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10238.265 187.44 10238.545 188.44 ;
    END
  END INJ_IN[244]
  PIN INJ_IN[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10202.985 187.44 10203.265 188.44 ;
    END
  END INJ_IN[243]
  PIN INJ_IN[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10156.505 187.44 10156.785 188.44 ;
    END
  END INJ_IN[242]
  PIN INJ_IN[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10098.265 187.44 10098.545 188.44 ;
    END
  END INJ_IN[241]
  PIN INJ_IN[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10090.985 187.44 10091.265 188.44 ;
    END
  END INJ_IN[240]
  PIN INJ_IN[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10015.945 187.44 10016.225 188.44 ;
    END
  END INJ_IN[239]
  PIN INJ_IN[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10000.265 187.44 10000.545 188.44 ;
    END
  END INJ_IN[238]
  PIN INJ_IN[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9949.865 187.44 9950.145 188.44 ;
    END
  END INJ_IN[237]
  PIN INJ_IN[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9929.145 187.44 9929.425 188.44 ;
    END
  END INJ_IN[236]
  PIN INJ_IN[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9859.705 187.44 9859.985 188.44 ;
    END
  END INJ_IN[235]
  PIN INJ_IN[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9850.465 187.44 9850.745 188.44 ;
    END
  END INJ_IN[234]
  PIN INJ_IN[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9789.705 187.44 9789.985 188.44 ;
    END
  END INJ_IN[233]
  PIN INJ_IN[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9782.425 187.44 9782.705 188.44 ;
    END
  END INJ_IN[232]
  PIN INJ_IN[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9711.025 187.44 9711.305 188.44 ;
    END
  END INJ_IN[231]
  PIN INJ_IN[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9678.265 187.44 9678.545 188.44 ;
    END
  END INJ_IN[230]
  PIN INJ_IN[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9642.985 187.44 9643.265 188.44 ;
    END
  END INJ_IN[229]
  PIN INJ_IN[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9596.505 187.44 9596.785 188.44 ;
    END
  END INJ_IN[228]
  PIN INJ_IN[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9538.265 187.44 9538.545 188.44 ;
    END
  END INJ_IN[227]
  PIN INJ_IN[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9530.985 187.44 9531.265 188.44 ;
    END
  END INJ_IN[226]
  PIN INJ_IN[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9455.945 187.44 9456.225 188.44 ;
    END
  END INJ_IN[225]
  PIN INJ_IN[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9440.265 187.44 9440.545 188.44 ;
    END
  END INJ_IN[224]
  PIN INJ_IN[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9389.865 187.44 9390.145 188.44 ;
    END
  END INJ_IN[223]
  PIN INJ_IN[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9369.145 187.44 9369.425 188.44 ;
    END
  END INJ_IN[222]
  PIN INJ_IN[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9299.705 187.44 9299.985 188.44 ;
    END
  END INJ_IN[221]
  PIN INJ_IN[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9290.465 187.44 9290.745 188.44 ;
    END
  END INJ_IN[220]
  PIN INJ_IN[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9229.705 187.44 9229.985 188.44 ;
    END
  END INJ_IN[219]
  PIN INJ_IN[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9222.425 187.44 9222.705 188.44 ;
    END
  END INJ_IN[218]
  PIN INJ_IN[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9151.025 187.44 9151.305 188.44 ;
    END
  END INJ_IN[217]
  PIN INJ_IN[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9118.265 187.44 9118.545 188.44 ;
    END
  END INJ_IN[216]
  PIN INJ_IN[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9082.985 187.44 9083.265 188.44 ;
    END
  END INJ_IN[215]
  PIN INJ_IN[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9036.505 187.44 9036.785 188.44 ;
    END
  END INJ_IN[214]
  PIN INJ_IN[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8978.265 187.44 8978.545 188.44 ;
    END
  END INJ_IN[213]
  PIN INJ_IN[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8970.985 187.44 8971.265 188.44 ;
    END
  END INJ_IN[212]
  PIN INJ_IN[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8895.945 187.44 8896.225 188.44 ;
    END
  END INJ_IN[211]
  PIN INJ_IN[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8880.265 187.44 8880.545 188.44 ;
    END
  END INJ_IN[210]
  PIN INJ_IN[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8829.865 187.44 8830.145 188.44 ;
    END
  END INJ_IN[209]
  PIN INJ_IN[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8809.145 187.44 8809.425 188.44 ;
    END
  END INJ_IN[208]
  PIN INJ_IN[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8739.705 187.44 8739.985 188.44 ;
    END
  END INJ_IN[207]
  PIN INJ_IN[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8730.465 187.44 8730.745 188.44 ;
    END
  END INJ_IN[206]
  PIN INJ_IN[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8669.705 187.44 8669.985 188.44 ;
    END
  END INJ_IN[205]
  PIN INJ_IN[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8662.425 187.44 8662.705 188.44 ;
    END
  END INJ_IN[204]
  PIN INJ_IN[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8591.025 187.44 8591.305 188.44 ;
    END
  END INJ_IN[203]
  PIN INJ_IN[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8558.265 187.44 8558.545 188.44 ;
    END
  END INJ_IN[202]
  PIN INJ_IN[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8522.985 187.44 8523.265 188.44 ;
    END
  END INJ_IN[201]
  PIN INJ_IN[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8476.505 187.44 8476.785 188.44 ;
    END
  END INJ_IN[200]
  PIN INJ_IN[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8418.265 187.44 8418.545 188.44 ;
    END
  END INJ_IN[199]
  PIN INJ_IN[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8410.985 187.44 8411.265 188.44 ;
    END
  END INJ_IN[198]
  PIN INJ_IN[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8335.945 187.44 8336.225 188.44 ;
    END
  END INJ_IN[197]
  PIN INJ_IN[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8320.265 187.44 8320.545 188.44 ;
    END
  END INJ_IN[196]
  PIN INJ_IN[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8269.865 187.44 8270.145 188.44 ;
    END
  END INJ_IN[195]
  PIN INJ_IN[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8249.145 187.44 8249.425 188.44 ;
    END
  END INJ_IN[194]
  PIN INJ_IN[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8179.705 187.44 8179.985 188.44 ;
    END
  END INJ_IN[193]
  PIN INJ_IN[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8170.465 187.44 8170.745 188.44 ;
    END
  END INJ_IN[192]
  PIN INJ_IN[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8109.705 187.44 8109.985 188.44 ;
    END
  END INJ_IN[191]
  PIN INJ_IN[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8102.425 187.44 8102.705 188.44 ;
    END
  END INJ_IN[190]
  PIN INJ_IN[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8031.025 187.44 8031.305 188.44 ;
    END
  END INJ_IN[189]
  PIN INJ_IN[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7998.265 187.44 7998.545 188.44 ;
    END
  END INJ_IN[188]
  PIN INJ_IN[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7962.985 187.44 7963.265 188.44 ;
    END
  END INJ_IN[187]
  PIN INJ_IN[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7916.505 187.44 7916.785 188.44 ;
    END
  END INJ_IN[186]
  PIN INJ_IN[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7858.265 187.44 7858.545 188.44 ;
    END
  END INJ_IN[185]
  PIN INJ_IN[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7850.985 187.44 7851.265 188.44 ;
    END
  END INJ_IN[184]
  PIN INJ_IN[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7775.945 187.44 7776.225 188.44 ;
    END
  END INJ_IN[183]
  PIN INJ_IN[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7760.265 187.44 7760.545 188.44 ;
    END
  END INJ_IN[182]
  PIN INJ_IN[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7709.865 187.44 7710.145 188.44 ;
    END
  END INJ_IN[181]
  PIN INJ_IN[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7689.145 187.44 7689.425 188.44 ;
    END
  END INJ_IN[180]
  PIN INJ_IN[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7619.705 187.44 7619.985 188.44 ;
    END
  END INJ_IN[179]
  PIN INJ_IN[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7610.465 187.44 7610.745 188.44 ;
    END
  END INJ_IN[178]
  PIN INJ_IN[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7549.705 187.44 7549.985 188.44 ;
    END
  END INJ_IN[177]
  PIN INJ_IN[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7542.425 187.44 7542.705 188.44 ;
    END
  END INJ_IN[176]
  PIN INJ_IN[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7471.025 187.44 7471.305 188.44 ;
    END
  END INJ_IN[175]
  PIN INJ_IN[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7438.265 187.44 7438.545 188.44 ;
    END
  END INJ_IN[174]
  PIN INJ_IN[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7402.985 187.44 7403.265 188.44 ;
    END
  END INJ_IN[173]
  PIN INJ_IN[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7356.505 187.44 7356.785 188.44 ;
    END
  END INJ_IN[172]
  PIN INJ_IN[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7298.265 187.44 7298.545 188.44 ;
    END
  END INJ_IN[171]
  PIN INJ_IN[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7290.985 187.44 7291.265 188.44 ;
    END
  END INJ_IN[170]
  PIN INJ_IN[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7215.945 187.44 7216.225 188.44 ;
    END
  END INJ_IN[169]
  PIN INJ_IN[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7200.265 187.44 7200.545 188.44 ;
    END
  END INJ_IN[168]
  PIN INJ_IN[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7149.865 187.44 7150.145 188.44 ;
    END
  END INJ_IN[167]
  PIN INJ_IN[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7129.145 187.44 7129.425 188.44 ;
    END
  END INJ_IN[166]
  PIN INJ_IN[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7059.705 187.44 7059.985 188.44 ;
    END
  END INJ_IN[165]
  PIN INJ_IN[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7050.465 187.44 7050.745 188.44 ;
    END
  END INJ_IN[164]
  PIN INJ_IN[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6989.705 187.44 6989.985 188.44 ;
    END
  END INJ_IN[163]
  PIN INJ_IN[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6982.425 187.44 6982.705 188.44 ;
    END
  END INJ_IN[162]
  PIN INJ_IN[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6911.025 187.44 6911.305 188.44 ;
    END
  END INJ_IN[161]
  PIN INJ_IN[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6878.265 187.44 6878.545 188.44 ;
    END
  END INJ_IN[160]
  PIN INJ_IN[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6842.985 187.44 6843.265 188.44 ;
    END
  END INJ_IN[159]
  PIN INJ_IN[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6796.505 187.44 6796.785 188.44 ;
    END
  END INJ_IN[158]
  PIN INJ_IN[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6738.265 187.44 6738.545 188.44 ;
    END
  END INJ_IN[157]
  PIN INJ_IN[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6730.985 187.44 6731.265 188.44 ;
    END
  END INJ_IN[156]
  PIN INJ_IN[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6655.945 187.44 6656.225 188.44 ;
    END
  END INJ_IN[155]
  PIN INJ_IN[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6640.265 187.44 6640.545 188.44 ;
    END
  END INJ_IN[154]
  PIN INJ_IN[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6589.865 187.44 6590.145 188.44 ;
    END
  END INJ_IN[153]
  PIN INJ_IN[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6569.145 187.44 6569.425 188.44 ;
    END
  END INJ_IN[152]
  PIN INJ_IN[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6499.705 187.44 6499.985 188.44 ;
    END
  END INJ_IN[151]
  PIN INJ_IN[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6490.465 187.44 6490.745 188.44 ;
    END
  END INJ_IN[150]
  PIN INJ_IN[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6429.705 187.44 6429.985 188.44 ;
    END
  END INJ_IN[149]
  PIN INJ_IN[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6422.425 187.44 6422.705 188.44 ;
    END
  END INJ_IN[148]
  PIN INJ_IN[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6351.025 187.44 6351.305 188.44 ;
    END
  END INJ_IN[147]
  PIN INJ_IN[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6318.265 187.44 6318.545 188.44 ;
    END
  END INJ_IN[146]
  PIN INJ_IN[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6282.985 187.44 6283.265 188.44 ;
    END
  END INJ_IN[145]
  PIN INJ_IN[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6236.505 187.44 6236.785 188.44 ;
    END
  END INJ_IN[144]
  PIN INJ_IN[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6178.265 187.44 6178.545 188.44 ;
    END
  END INJ_IN[143]
  PIN INJ_IN[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6170.985 187.44 6171.265 188.44 ;
    END
  END INJ_IN[142]
  PIN INJ_IN[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6095.945 187.44 6096.225 188.44 ;
    END
  END INJ_IN[141]
  PIN INJ_IN[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6080.265 187.44 6080.545 188.44 ;
    END
  END INJ_IN[140]
  PIN INJ_IN[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6029.865 187.44 6030.145 188.44 ;
    END
  END INJ_IN[139]
  PIN INJ_IN[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6009.145 187.44 6009.425 188.44 ;
    END
  END INJ_IN[138]
  PIN INJ_IN[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5939.705 187.44 5939.985 188.44 ;
    END
  END INJ_IN[137]
  PIN INJ_IN[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5930.465 187.44 5930.745 188.44 ;
    END
  END INJ_IN[136]
  PIN INJ_IN[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5869.705 187.44 5869.985 188.44 ;
    END
  END INJ_IN[135]
  PIN INJ_IN[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5862.425 187.44 5862.705 188.44 ;
    END
  END INJ_IN[134]
  PIN INJ_IN[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5791.025 187.44 5791.305 188.44 ;
    END
  END INJ_IN[133]
  PIN INJ_IN[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5758.265 187.44 5758.545 188.44 ;
    END
  END INJ_IN[132]
  PIN INJ_IN[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5722.985 187.44 5723.265 188.44 ;
    END
  END INJ_IN[131]
  PIN INJ_IN[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5676.505 187.44 5676.785 188.44 ;
    END
  END INJ_IN[130]
  PIN INJ_IN[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5618.265 187.44 5618.545 188.44 ;
    END
  END INJ_IN[129]
  PIN INJ_IN[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5610.985 187.44 5611.265 188.44 ;
    END
  END INJ_IN[128]
  PIN INJ_IN[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5535.945 187.44 5536.225 188.44 ;
    END
  END INJ_IN[127]
  PIN INJ_IN[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5520.265 187.44 5520.545 188.44 ;
    END
  END INJ_IN[126]
  PIN INJ_IN[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5469.865 187.44 5470.145 188.44 ;
    END
  END INJ_IN[125]
  PIN INJ_IN[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5449.145 187.44 5449.425 188.44 ;
    END
  END INJ_IN[124]
  PIN INJ_IN[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5379.705 187.44 5379.985 188.44 ;
    END
  END INJ_IN[123]
  PIN INJ_IN[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5370.465 187.44 5370.745 188.44 ;
    END
  END INJ_IN[122]
  PIN INJ_IN[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5309.705 187.44 5309.985 188.44 ;
    END
  END INJ_IN[121]
  PIN INJ_IN[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5302.425 187.44 5302.705 188.44 ;
    END
  END INJ_IN[120]
  PIN INJ_IN[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5231.025 187.44 5231.305 188.44 ;
    END
  END INJ_IN[119]
  PIN INJ_IN[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5198.265 187.44 5198.545 188.44 ;
    END
  END INJ_IN[118]
  PIN INJ_IN[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5162.985 187.44 5163.265 188.44 ;
    END
  END INJ_IN[117]
  PIN INJ_IN[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5116.505 187.44 5116.785 188.44 ;
    END
  END INJ_IN[116]
  PIN INJ_IN[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5058.265 187.44 5058.545 188.44 ;
    END
  END INJ_IN[115]
  PIN INJ_IN[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5050.985 187.44 5051.265 188.44 ;
    END
  END INJ_IN[114]
  PIN INJ_IN[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4975.945 187.44 4976.225 188.44 ;
    END
  END INJ_IN[113]
  PIN INJ_IN[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4960.265 187.44 4960.545 188.44 ;
    END
  END INJ_IN[112]
  PIN INJ_IN[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4909.865 187.44 4910.145 188.44 ;
    END
  END INJ_IN[111]
  PIN INJ_IN[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4889.145 187.44 4889.425 188.44 ;
    END
  END INJ_IN[110]
  PIN INJ_IN[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4819.705 187.44 4819.985 188.44 ;
    END
  END INJ_IN[109]
  PIN INJ_IN[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4810.465 187.44 4810.745 188.44 ;
    END
  END INJ_IN[108]
  PIN INJ_IN[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4749.705 187.44 4749.985 188.44 ;
    END
  END INJ_IN[107]
  PIN INJ_IN[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4742.425 187.44 4742.705 188.44 ;
    END
  END INJ_IN[106]
  PIN INJ_IN[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4671.025 187.44 4671.305 188.44 ;
    END
  END INJ_IN[105]
  PIN INJ_IN[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4638.265 187.44 4638.545 188.44 ;
    END
  END INJ_IN[104]
  PIN INJ_IN[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4602.985 187.44 4603.265 188.44 ;
    END
  END INJ_IN[103]
  PIN INJ_IN[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4556.505 187.44 4556.785 188.44 ;
    END
  END INJ_IN[102]
  PIN INJ_IN[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4498.265 187.44 4498.545 188.44 ;
    END
  END INJ_IN[101]
  PIN INJ_IN[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4490.985 187.44 4491.265 188.44 ;
    END
  END INJ_IN[100]
  PIN INJ_IN[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4415.945 187.44 4416.225 188.44 ;
    END
  END INJ_IN[99]
  PIN INJ_IN[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4400.265 187.44 4400.545 188.44 ;
    END
  END INJ_IN[98]
  PIN INJ_IN[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4349.865 187.44 4350.145 188.44 ;
    END
  END INJ_IN[97]
  PIN INJ_IN[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4329.145 187.44 4329.425 188.44 ;
    END
  END INJ_IN[96]
  PIN INJ_IN[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4259.705 187.44 4259.985 188.44 ;
    END
  END INJ_IN[95]
  PIN INJ_IN[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4250.465 187.44 4250.745 188.44 ;
    END
  END INJ_IN[94]
  PIN INJ_IN[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4189.705 187.44 4189.985 188.44 ;
    END
  END INJ_IN[93]
  PIN INJ_IN[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4182.425 187.44 4182.705 188.44 ;
    END
  END INJ_IN[92]
  PIN INJ_IN[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4111.025 187.44 4111.305 188.44 ;
    END
  END INJ_IN[91]
  PIN INJ_IN[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4078.265 187.44 4078.545 188.44 ;
    END
  END INJ_IN[90]
  PIN INJ_IN[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4042.985 187.44 4043.265 188.44 ;
    END
  END INJ_IN[89]
  PIN INJ_IN[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3996.505 187.44 3996.785 188.44 ;
    END
  END INJ_IN[88]
  PIN INJ_IN[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3938.265 187.44 3938.545 188.44 ;
    END
  END INJ_IN[87]
  PIN INJ_IN[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3930.985 187.44 3931.265 188.44 ;
    END
  END INJ_IN[86]
  PIN INJ_IN[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3855.945 187.44 3856.225 188.44 ;
    END
  END INJ_IN[85]
  PIN INJ_IN[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3840.265 187.44 3840.545 188.44 ;
    END
  END INJ_IN[84]
  PIN INJ_IN[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3789.865 187.44 3790.145 188.44 ;
    END
  END INJ_IN[83]
  PIN INJ_IN[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3769.145 187.44 3769.425 188.44 ;
    END
  END INJ_IN[82]
  PIN INJ_IN[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3699.705 187.44 3699.985 188.44 ;
    END
  END INJ_IN[81]
  PIN INJ_IN[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3690.465 187.44 3690.745 188.44 ;
    END
  END INJ_IN[80]
  PIN INJ_IN[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3629.705 187.44 3629.985 188.44 ;
    END
  END INJ_IN[79]
  PIN INJ_IN[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3622.425 187.44 3622.705 188.44 ;
    END
  END INJ_IN[78]
  PIN INJ_IN[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3551.025 187.44 3551.305 188.44 ;
    END
  END INJ_IN[77]
  PIN INJ_IN[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3518.265 187.44 3518.545 188.44 ;
    END
  END INJ_IN[76]
  PIN INJ_IN[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3482.985 187.44 3483.265 188.44 ;
    END
  END INJ_IN[75]
  PIN INJ_IN[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3436.505 187.44 3436.785 188.44 ;
    END
  END INJ_IN[74]
  PIN INJ_IN[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3378.265 187.44 3378.545 188.44 ;
    END
  END INJ_IN[73]
  PIN INJ_IN[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3370.985 187.44 3371.265 188.44 ;
    END
  END INJ_IN[72]
  PIN INJ_IN[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3295.945 187.44 3296.225 188.44 ;
    END
  END INJ_IN[71]
  PIN INJ_IN[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3280.265 187.44 3280.545 188.44 ;
    END
  END INJ_IN[70]
  PIN INJ_IN[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3229.865 187.44 3230.145 188.44 ;
    END
  END INJ_IN[69]
  PIN INJ_IN[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3209.145 187.44 3209.425 188.44 ;
    END
  END INJ_IN[68]
  PIN INJ_IN[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3139.705 187.44 3139.985 188.44 ;
    END
  END INJ_IN[67]
  PIN INJ_IN[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3130.465 187.44 3130.745 188.44 ;
    END
  END INJ_IN[66]
  PIN INJ_IN[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3069.705 187.44 3069.985 188.44 ;
    END
  END INJ_IN[65]
  PIN INJ_IN[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3062.425 187.44 3062.705 188.44 ;
    END
  END INJ_IN[64]
  PIN INJ_IN[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2991.025 187.44 2991.305 188.44 ;
    END
  END INJ_IN[63]
  PIN INJ_IN[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2958.265 187.44 2958.545 188.44 ;
    END
  END INJ_IN[62]
  PIN INJ_IN[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2922.985 187.44 2923.265 188.44 ;
    END
  END INJ_IN[61]
  PIN INJ_IN[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2876.505 187.44 2876.785 188.44 ;
    END
  END INJ_IN[60]
  PIN INJ_IN[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2818.265 187.44 2818.545 188.44 ;
    END
  END INJ_IN[59]
  PIN INJ_IN[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2810.985 187.44 2811.265 188.44 ;
    END
  END INJ_IN[58]
  PIN INJ_IN[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2735.945 187.44 2736.225 188.44 ;
    END
  END INJ_IN[57]
  PIN INJ_IN[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2720.265 187.44 2720.545 188.44 ;
    END
  END INJ_IN[56]
  PIN INJ_IN[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2669.865 187.44 2670.145 188.44 ;
    END
  END INJ_IN[55]
  PIN INJ_IN[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2649.145 187.44 2649.425 188.44 ;
    END
  END INJ_IN[54]
  PIN INJ_IN[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2579.705 187.44 2579.985 188.44 ;
    END
  END INJ_IN[53]
  PIN INJ_IN[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2570.465 187.44 2570.745 188.44 ;
    END
  END INJ_IN[52]
  PIN INJ_IN[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2509.705 187.44 2509.985 188.44 ;
    END
  END INJ_IN[51]
  PIN INJ_IN[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2502.425 187.44 2502.705 188.44 ;
    END
  END INJ_IN[50]
  PIN INJ_IN[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2431.025 187.44 2431.305 188.44 ;
    END
  END INJ_IN[49]
  PIN INJ_IN[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2398.265 187.44 2398.545 188.44 ;
    END
  END INJ_IN[48]
  PIN INJ_IN[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2362.985 187.44 2363.265 188.44 ;
    END
  END INJ_IN[47]
  PIN INJ_IN[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2316.505 187.44 2316.785 188.44 ;
    END
  END INJ_IN[46]
  PIN INJ_IN[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2258.265 187.44 2258.545 188.44 ;
    END
  END INJ_IN[45]
  PIN INJ_IN[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2250.985 187.44 2251.265 188.44 ;
    END
  END INJ_IN[44]
  PIN INJ_IN[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2175.945 187.44 2176.225 188.44 ;
    END
  END INJ_IN[43]
  PIN INJ_IN[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2160.265 187.44 2160.545 188.44 ;
    END
  END INJ_IN[42]
  PIN INJ_IN[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2109.865 187.44 2110.145 188.44 ;
    END
  END INJ_IN[41]
  PIN INJ_IN[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2089.145 187.44 2089.425 188.44 ;
    END
  END INJ_IN[40]
  PIN INJ_IN[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2019.705 187.44 2019.985 188.44 ;
    END
  END INJ_IN[39]
  PIN INJ_IN[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2010.465 187.44 2010.745 188.44 ;
    END
  END INJ_IN[38]
  PIN INJ_IN[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1949.705 187.44 1949.985 188.44 ;
    END
  END INJ_IN[37]
  PIN INJ_IN[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1942.425 187.44 1942.705 188.44 ;
    END
  END INJ_IN[36]
  PIN INJ_IN[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1871.025 187.44 1871.305 188.44 ;
    END
  END INJ_IN[35]
  PIN INJ_IN[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1838.265 187.44 1838.545 188.44 ;
    END
  END INJ_IN[34]
  PIN INJ_IN[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1802.985 187.44 1803.265 188.44 ;
    END
  END INJ_IN[33]
  PIN INJ_IN[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1756.505 187.44 1756.785 188.44 ;
    END
  END INJ_IN[32]
  PIN INJ_IN[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1698.265 187.44 1698.545 188.44 ;
    END
  END INJ_IN[31]
  PIN INJ_IN[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1690.985 187.44 1691.265 188.44 ;
    END
  END INJ_IN[30]
  PIN INJ_IN[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1615.945 187.44 1616.225 188.44 ;
    END
  END INJ_IN[29]
  PIN INJ_IN[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1600.265 187.44 1600.545 188.44 ;
    END
  END INJ_IN[28]
  PIN INJ_IN[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1549.865 187.44 1550.145 188.44 ;
    END
  END INJ_IN[27]
  PIN INJ_IN[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1529.145 187.44 1529.425 188.44 ;
    END
  END INJ_IN[26]
  PIN INJ_IN[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1459.705 187.44 1459.985 188.44 ;
    END
  END INJ_IN[25]
  PIN INJ_IN[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1450.465 187.44 1450.745 188.44 ;
    END
  END INJ_IN[24]
  PIN INJ_IN[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1389.705 187.44 1389.985 188.44 ;
    END
  END INJ_IN[23]
  PIN INJ_IN[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1382.425 187.44 1382.705 188.44 ;
    END
  END INJ_IN[22]
  PIN INJ_IN[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1311.025 187.44 1311.305 188.44 ;
    END
  END INJ_IN[21]
  PIN INJ_IN[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1278.265 187.44 1278.545 188.44 ;
    END
  END INJ_IN[20]
  PIN INJ_IN[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1242.985 187.44 1243.265 188.44 ;
    END
  END INJ_IN[19]
  PIN INJ_IN[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1196.505 187.44 1196.785 188.44 ;
    END
  END INJ_IN[18]
  PIN INJ_IN[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1138.265 187.44 1138.545 188.44 ;
    END
  END INJ_IN[17]
  PIN INJ_IN[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1130.985 187.44 1131.265 188.44 ;
    END
  END INJ_IN[16]
  PIN INJ_IN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1055.945 187.44 1056.225 188.44 ;
    END
  END INJ_IN[15]
  PIN INJ_IN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1040.265 187.44 1040.545 188.44 ;
    END
  END INJ_IN[14]
  PIN INJ_IN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 989.865 187.44 990.145 188.44 ;
    END
  END INJ_IN[13]
  PIN INJ_IN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 969.145 187.44 969.425 188.44 ;
    END
  END INJ_IN[12]
  PIN INJ_IN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 899.705 187.44 899.985 188.44 ;
    END
  END INJ_IN[11]
  PIN INJ_IN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 890.465 187.44 890.745 188.44 ;
    END
  END INJ_IN[10]
  PIN INJ_IN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 829.705 187.44 829.985 188.44 ;
    END
  END INJ_IN[9]
  PIN INJ_IN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 822.425 187.44 822.705 188.44 ;
    END
  END INJ_IN[8]
  PIN INJ_IN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 751.025 187.44 751.305 188.44 ;
    END
  END INJ_IN[7]
  PIN INJ_IN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 718.265 187.44 718.545 188.44 ;
    END
  END INJ_IN[6]
  PIN INJ_IN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 682.985 187.44 683.265 188.44 ;
    END
  END INJ_IN[5]
  PIN INJ_IN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 636.505 187.44 636.785 188.44 ;
    END
  END INJ_IN[4]
  PIN INJ_IN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 578.265 187.44 578.545 188.44 ;
    END
  END INJ_IN[3]
  PIN INJ_IN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 570.985 187.44 571.265 188.44 ;
    END
  END INJ_IN[2]
  PIN INJ_IN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 495.945 187.44 496.225 188.44 ;
    END
  END INJ_IN[1]
  PIN INJ_IN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 480.265 187.44 480.545 188.44 ;
    END
  END INJ_IN[0]
  PIN MASKV[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18356.585 187.44 18356.865 188.44 ;
    END
  END MASKV[447]
  PIN MASKV[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18283.225 187.44 18283.505 188.44 ;
    END
  END MASKV[446]
  PIN MASKV[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18274.825 187.44 18275.105 188.44 ;
    END
  END MASKV[445]
  PIN MASKV[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18217.705 187.44 18217.985 188.44 ;
    END
  END MASKV[444]
  PIN MASKV[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18209.305 187.44 18209.585 188.44 ;
    END
  END MASKV[443]
  PIN MASKV[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18136.505 187.44 18136.785 188.44 ;
    END
  END MASKV[442]
  PIN MASKV[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18119.705 187.44 18119.985 188.44 ;
    END
  END MASKV[441]
  PIN MASKV[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18070.985 187.44 18071.265 188.44 ;
    END
  END MASKV[440]
  PIN MASKV[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18049.705 187.44 18049.985 188.44 ;
    END
  END MASKV[439]
  PIN MASKV[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17980.825 187.44 17981.105 188.44 ;
    END
  END MASKV[438]
  PIN MASKV[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17970.465 187.44 17970.745 188.44 ;
    END
  END MASKV[437]
  PIN MASKV[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17910.825 187.44 17911.105 188.44 ;
    END
  END MASKV[436]
  PIN MASKV[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17902.425 187.44 17902.705 188.44 ;
    END
  END MASKV[435]
  PIN MASKV[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17831.025 187.44 17831.305 188.44 ;
    END
  END MASKV[434]
  PIN MASKV[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17796.585 187.44 17796.865 188.44 ;
    END
  END MASKV[433]
  PIN MASKV[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17723.225 187.44 17723.505 188.44 ;
    END
  END MASKV[432]
  PIN MASKV[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17714.825 187.44 17715.105 188.44 ;
    END
  END MASKV[431]
  PIN MASKV[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17657.705 187.44 17657.985 188.44 ;
    END
  END MASKV[430]
  PIN MASKV[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17649.305 187.44 17649.585 188.44 ;
    END
  END MASKV[429]
  PIN MASKV[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17576.505 187.44 17576.785 188.44 ;
    END
  END MASKV[428]
  PIN MASKV[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17559.705 187.44 17559.985 188.44 ;
    END
  END MASKV[427]
  PIN MASKV[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17510.985 187.44 17511.265 188.44 ;
    END
  END MASKV[426]
  PIN MASKV[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17489.705 187.44 17489.985 188.44 ;
    END
  END MASKV[425]
  PIN MASKV[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17420.825 187.44 17421.105 188.44 ;
    END
  END MASKV[424]
  PIN MASKV[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17410.465 187.44 17410.745 188.44 ;
    END
  END MASKV[423]
  PIN MASKV[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17350.825 187.44 17351.105 188.44 ;
    END
  END MASKV[422]
  PIN MASKV[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17342.425 187.44 17342.705 188.44 ;
    END
  END MASKV[421]
  PIN MASKV[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17271.025 187.44 17271.305 188.44 ;
    END
  END MASKV[420]
  PIN MASKV[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17236.585 187.44 17236.865 188.44 ;
    END
  END MASKV[419]
  PIN MASKV[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17163.225 187.44 17163.505 188.44 ;
    END
  END MASKV[418]
  PIN MASKV[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17154.825 187.44 17155.105 188.44 ;
    END
  END MASKV[417]
  PIN MASKV[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17097.705 187.44 17097.985 188.44 ;
    END
  END MASKV[416]
  PIN MASKV[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17089.305 187.44 17089.585 188.44 ;
    END
  END MASKV[415]
  PIN MASKV[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17016.505 187.44 17016.785 188.44 ;
    END
  END MASKV[414]
  PIN MASKV[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16999.705 187.44 16999.985 188.44 ;
    END
  END MASKV[413]
  PIN MASKV[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16950.985 187.44 16951.265 188.44 ;
    END
  END MASKV[412]
  PIN MASKV[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16929.705 187.44 16929.985 188.44 ;
    END
  END MASKV[411]
  PIN MASKV[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16860.825 187.44 16861.105 188.44 ;
    END
  END MASKV[410]
  PIN MASKV[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16850.465 187.44 16850.745 188.44 ;
    END
  END MASKV[409]
  PIN MASKV[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16790.825 187.44 16791.105 188.44 ;
    END
  END MASKV[408]
  PIN MASKV[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16782.425 187.44 16782.705 188.44 ;
    END
  END MASKV[407]
  PIN MASKV[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16711.025 187.44 16711.305 188.44 ;
    END
  END MASKV[406]
  PIN MASKV[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16676.585 187.44 16676.865 188.44 ;
    END
  END MASKV[405]
  PIN MASKV[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16603.225 187.44 16603.505 188.44 ;
    END
  END MASKV[404]
  PIN MASKV[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16594.825 187.44 16595.105 188.44 ;
    END
  END MASKV[403]
  PIN MASKV[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16537.705 187.44 16537.985 188.44 ;
    END
  END MASKV[402]
  PIN MASKV[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16529.305 187.44 16529.585 188.44 ;
    END
  END MASKV[401]
  PIN MASKV[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16456.505 187.44 16456.785 188.44 ;
    END
  END MASKV[400]
  PIN MASKV[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16439.705 187.44 16439.985 188.44 ;
    END
  END MASKV[399]
  PIN MASKV[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16390.985 187.44 16391.265 188.44 ;
    END
  END MASKV[398]
  PIN MASKV[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16369.705 187.44 16369.985 188.44 ;
    END
  END MASKV[397]
  PIN MASKV[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16300.825 187.44 16301.105 188.44 ;
    END
  END MASKV[396]
  PIN MASKV[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16290.465 187.44 16290.745 188.44 ;
    END
  END MASKV[395]
  PIN MASKV[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16230.825 187.44 16231.105 188.44 ;
    END
  END MASKV[394]
  PIN MASKV[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16222.425 187.44 16222.705 188.44 ;
    END
  END MASKV[393]
  PIN MASKV[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16151.025 187.44 16151.305 188.44 ;
    END
  END MASKV[392]
  PIN MASKV[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16116.585 187.44 16116.865 188.44 ;
    END
  END MASKV[391]
  PIN MASKV[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16043.225 187.44 16043.505 188.44 ;
    END
  END MASKV[390]
  PIN MASKV[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16034.825 187.44 16035.105 188.44 ;
    END
  END MASKV[389]
  PIN MASKV[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15977.705 187.44 15977.985 188.44 ;
    END
  END MASKV[388]
  PIN MASKV[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15969.305 187.44 15969.585 188.44 ;
    END
  END MASKV[387]
  PIN MASKV[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15896.505 187.44 15896.785 188.44 ;
    END
  END MASKV[386]
  PIN MASKV[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15879.705 187.44 15879.985 188.44 ;
    END
  END MASKV[385]
  PIN MASKV[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15830.985 187.44 15831.265 188.44 ;
    END
  END MASKV[384]
  PIN MASKV[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15809.705 187.44 15809.985 188.44 ;
    END
  END MASKV[383]
  PIN MASKV[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15740.825 187.44 15741.105 188.44 ;
    END
  END MASKV[382]
  PIN MASKV[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15730.465 187.44 15730.745 188.44 ;
    END
  END MASKV[381]
  PIN MASKV[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15670.825 187.44 15671.105 188.44 ;
    END
  END MASKV[380]
  PIN MASKV[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15662.425 187.44 15662.705 188.44 ;
    END
  END MASKV[379]
  PIN MASKV[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15591.025 187.44 15591.305 188.44 ;
    END
  END MASKV[378]
  PIN MASKV[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15556.585 187.44 15556.865 188.44 ;
    END
  END MASKV[377]
  PIN MASKV[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15483.225 187.44 15483.505 188.44 ;
    END
  END MASKV[376]
  PIN MASKV[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15474.825 187.44 15475.105 188.44 ;
    END
  END MASKV[375]
  PIN MASKV[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15417.705 187.44 15417.985 188.44 ;
    END
  END MASKV[374]
  PIN MASKV[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15409.305 187.44 15409.585 188.44 ;
    END
  END MASKV[373]
  PIN MASKV[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15336.505 187.44 15336.785 188.44 ;
    END
  END MASKV[372]
  PIN MASKV[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15319.705 187.44 15319.985 188.44 ;
    END
  END MASKV[371]
  PIN MASKV[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15270.985 187.44 15271.265 188.44 ;
    END
  END MASKV[370]
  PIN MASKV[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15249.705 187.44 15249.985 188.44 ;
    END
  END MASKV[369]
  PIN MASKV[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15180.825 187.44 15181.105 188.44 ;
    END
  END MASKV[368]
  PIN MASKV[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15170.465 187.44 15170.745 188.44 ;
    END
  END MASKV[367]
  PIN MASKV[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15110.825 187.44 15111.105 188.44 ;
    END
  END MASKV[366]
  PIN MASKV[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15102.425 187.44 15102.705 188.44 ;
    END
  END MASKV[365]
  PIN MASKV[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15031.025 187.44 15031.305 188.44 ;
    END
  END MASKV[364]
  PIN MASKV[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14996.585 187.44 14996.865 188.44 ;
    END
  END MASKV[363]
  PIN MASKV[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14923.225 187.44 14923.505 188.44 ;
    END
  END MASKV[362]
  PIN MASKV[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14914.825 187.44 14915.105 188.44 ;
    END
  END MASKV[361]
  PIN MASKV[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14857.705 187.44 14857.985 188.44 ;
    END
  END MASKV[360]
  PIN MASKV[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14849.305 187.44 14849.585 188.44 ;
    END
  END MASKV[359]
  PIN MASKV[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14776.505 187.44 14776.785 188.44 ;
    END
  END MASKV[358]
  PIN MASKV[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14759.705 187.44 14759.985 188.44 ;
    END
  END MASKV[357]
  PIN MASKV[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14710.985 187.44 14711.265 188.44 ;
    END
  END MASKV[356]
  PIN MASKV[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14689.705 187.44 14689.985 188.44 ;
    END
  END MASKV[355]
  PIN MASKV[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14620.825 187.44 14621.105 188.44 ;
    END
  END MASKV[354]
  PIN MASKV[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14610.465 187.44 14610.745 188.44 ;
    END
  END MASKV[353]
  PIN MASKV[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14550.825 187.44 14551.105 188.44 ;
    END
  END MASKV[352]
  PIN MASKV[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14542.425 187.44 14542.705 188.44 ;
    END
  END MASKV[351]
  PIN MASKV[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14471.025 187.44 14471.305 188.44 ;
    END
  END MASKV[350]
  PIN MASKV[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14436.585 187.44 14436.865 188.44 ;
    END
  END MASKV[349]
  PIN MASKV[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14363.225 187.44 14363.505 188.44 ;
    END
  END MASKV[348]
  PIN MASKV[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14354.825 187.44 14355.105 188.44 ;
    END
  END MASKV[347]
  PIN MASKV[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14297.705 187.44 14297.985 188.44 ;
    END
  END MASKV[346]
  PIN MASKV[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14289.305 187.44 14289.585 188.44 ;
    END
  END MASKV[345]
  PIN MASKV[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14216.505 187.44 14216.785 188.44 ;
    END
  END MASKV[344]
  PIN MASKV[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14199.705 187.44 14199.985 188.44 ;
    END
  END MASKV[343]
  PIN MASKV[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14150.985 187.44 14151.265 188.44 ;
    END
  END MASKV[342]
  PIN MASKV[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14129.705 187.44 14129.985 188.44 ;
    END
  END MASKV[341]
  PIN MASKV[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14060.825 187.44 14061.105 188.44 ;
    END
  END MASKV[340]
  PIN MASKV[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14050.465 187.44 14050.745 188.44 ;
    END
  END MASKV[339]
  PIN MASKV[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13990.825 187.44 13991.105 188.44 ;
    END
  END MASKV[338]
  PIN MASKV[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13982.425 187.44 13982.705 188.44 ;
    END
  END MASKV[337]
  PIN MASKV[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13911.025 187.44 13911.305 188.44 ;
    END
  END MASKV[336]
  PIN MASKV[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13876.585 187.44 13876.865 188.44 ;
    END
  END MASKV[335]
  PIN MASKV[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13803.225 187.44 13803.505 188.44 ;
    END
  END MASKV[334]
  PIN MASKV[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13794.825 187.44 13795.105 188.44 ;
    END
  END MASKV[333]
  PIN MASKV[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13737.705 187.44 13737.985 188.44 ;
    END
  END MASKV[332]
  PIN MASKV[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13729.305 187.44 13729.585 188.44 ;
    END
  END MASKV[331]
  PIN MASKV[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13656.505 187.44 13656.785 188.44 ;
    END
  END MASKV[330]
  PIN MASKV[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13639.705 187.44 13639.985 188.44 ;
    END
  END MASKV[329]
  PIN MASKV[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13590.985 187.44 13591.265 188.44 ;
    END
  END MASKV[328]
  PIN MASKV[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13569.705 187.44 13569.985 188.44 ;
    END
  END MASKV[327]
  PIN MASKV[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13500.825 187.44 13501.105 188.44 ;
    END
  END MASKV[326]
  PIN MASKV[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13490.465 187.44 13490.745 188.44 ;
    END
  END MASKV[325]
  PIN MASKV[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13430.825 187.44 13431.105 188.44 ;
    END
  END MASKV[324]
  PIN MASKV[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13422.425 187.44 13422.705 188.44 ;
    END
  END MASKV[323]
  PIN MASKV[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13351.025 187.44 13351.305 188.44 ;
    END
  END MASKV[322]
  PIN MASKV[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13316.585 187.44 13316.865 188.44 ;
    END
  END MASKV[321]
  PIN MASKV[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13243.225 187.44 13243.505 188.44 ;
    END
  END MASKV[320]
  PIN MASKV[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13234.825 187.44 13235.105 188.44 ;
    END
  END MASKV[319]
  PIN MASKV[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13177.705 187.44 13177.985 188.44 ;
    END
  END MASKV[318]
  PIN MASKV[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13169.305 187.44 13169.585 188.44 ;
    END
  END MASKV[317]
  PIN MASKV[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13096.505 187.44 13096.785 188.44 ;
    END
  END MASKV[316]
  PIN MASKV[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13079.705 187.44 13079.985 188.44 ;
    END
  END MASKV[315]
  PIN MASKV[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13030.985 187.44 13031.265 188.44 ;
    END
  END MASKV[314]
  PIN MASKV[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13009.705 187.44 13009.985 188.44 ;
    END
  END MASKV[313]
  PIN MASKV[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12940.825 187.44 12941.105 188.44 ;
    END
  END MASKV[312]
  PIN MASKV[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12930.465 187.44 12930.745 188.44 ;
    END
  END MASKV[311]
  PIN MASKV[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12870.825 187.44 12871.105 188.44 ;
    END
  END MASKV[310]
  PIN MASKV[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12862.425 187.44 12862.705 188.44 ;
    END
  END MASKV[309]
  PIN MASKV[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12791.025 187.44 12791.305 188.44 ;
    END
  END MASKV[308]
  PIN MASKV[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12756.585 187.44 12756.865 188.44 ;
    END
  END MASKV[307]
  PIN MASKV[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12683.225 187.44 12683.505 188.44 ;
    END
  END MASKV[306]
  PIN MASKV[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12674.825 187.44 12675.105 188.44 ;
    END
  END MASKV[305]
  PIN MASKV[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12617.705 187.44 12617.985 188.44 ;
    END
  END MASKV[304]
  PIN MASKV[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12609.305 187.44 12609.585 188.44 ;
    END
  END MASKV[303]
  PIN MASKV[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12536.505 187.44 12536.785 188.44 ;
    END
  END MASKV[302]
  PIN MASKV[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12519.705 187.44 12519.985 188.44 ;
    END
  END MASKV[301]
  PIN MASKV[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12470.985 187.44 12471.265 188.44 ;
    END
  END MASKV[300]
  PIN MASKV[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12449.705 187.44 12449.985 188.44 ;
    END
  END MASKV[299]
  PIN MASKV[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12380.825 187.44 12381.105 188.44 ;
    END
  END MASKV[298]
  PIN MASKV[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12370.465 187.44 12370.745 188.44 ;
    END
  END MASKV[297]
  PIN MASKV[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12310.825 187.44 12311.105 188.44 ;
    END
  END MASKV[296]
  PIN MASKV[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12302.425 187.44 12302.705 188.44 ;
    END
  END MASKV[295]
  PIN MASKV[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12231.025 187.44 12231.305 188.44 ;
    END
  END MASKV[294]
  PIN MASKV[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12196.585 187.44 12196.865 188.44 ;
    END
  END MASKV[293]
  PIN MASKV[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12123.225 187.44 12123.505 188.44 ;
    END
  END MASKV[292]
  PIN MASKV[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12114.825 187.44 12115.105 188.44 ;
    END
  END MASKV[291]
  PIN MASKV[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12057.705 187.44 12057.985 188.44 ;
    END
  END MASKV[290]
  PIN MASKV[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12049.305 187.44 12049.585 188.44 ;
    END
  END MASKV[289]
  PIN MASKV[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11976.505 187.44 11976.785 188.44 ;
    END
  END MASKV[288]
  PIN MASKV[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11959.705 187.44 11959.985 188.44 ;
    END
  END MASKV[287]
  PIN MASKV[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11910.985 187.44 11911.265 188.44 ;
    END
  END MASKV[286]
  PIN MASKV[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11889.705 187.44 11889.985 188.44 ;
    END
  END MASKV[285]
  PIN MASKV[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11820.825 187.44 11821.105 188.44 ;
    END
  END MASKV[284]
  PIN MASKV[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11810.465 187.44 11810.745 188.44 ;
    END
  END MASKV[283]
  PIN MASKV[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11750.825 187.44 11751.105 188.44 ;
    END
  END MASKV[282]
  PIN MASKV[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11742.425 187.44 11742.705 188.44 ;
    END
  END MASKV[281]
  PIN MASKV[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11671.025 187.44 11671.305 188.44 ;
    END
  END MASKV[280]
  PIN MASKV[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11636.585 187.44 11636.865 188.44 ;
    END
  END MASKV[279]
  PIN MASKV[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11563.225 187.44 11563.505 188.44 ;
    END
  END MASKV[278]
  PIN MASKV[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11554.825 187.44 11555.105 188.44 ;
    END
  END MASKV[277]
  PIN MASKV[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11497.705 187.44 11497.985 188.44 ;
    END
  END MASKV[276]
  PIN MASKV[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11489.305 187.44 11489.585 188.44 ;
    END
  END MASKV[275]
  PIN MASKV[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11416.505 187.44 11416.785 188.44 ;
    END
  END MASKV[274]
  PIN MASKV[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11399.705 187.44 11399.985 188.44 ;
    END
  END MASKV[273]
  PIN MASKV[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11350.985 187.44 11351.265 188.44 ;
    END
  END MASKV[272]
  PIN MASKV[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11329.705 187.44 11329.985 188.44 ;
    END
  END MASKV[271]
  PIN MASKV[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11260.825 187.44 11261.105 188.44 ;
    END
  END MASKV[270]
  PIN MASKV[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11250.465 187.44 11250.745 188.44 ;
    END
  END MASKV[269]
  PIN MASKV[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11190.825 187.44 11191.105 188.44 ;
    END
  END MASKV[268]
  PIN MASKV[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11182.425 187.44 11182.705 188.44 ;
    END
  END MASKV[267]
  PIN MASKV[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11111.025 187.44 11111.305 188.44 ;
    END
  END MASKV[266]
  PIN MASKV[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11076.585 187.44 11076.865 188.44 ;
    END
  END MASKV[265]
  PIN MASKV[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11003.225 187.44 11003.505 188.44 ;
    END
  END MASKV[264]
  PIN MASKV[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10994.825 187.44 10995.105 188.44 ;
    END
  END MASKV[263]
  PIN MASKV[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10937.705 187.44 10937.985 188.44 ;
    END
  END MASKV[262]
  PIN MASKV[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10929.305 187.44 10929.585 188.44 ;
    END
  END MASKV[261]
  PIN MASKV[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10856.505 187.44 10856.785 188.44 ;
    END
  END MASKV[260]
  PIN MASKV[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10839.705 187.44 10839.985 188.44 ;
    END
  END MASKV[259]
  PIN MASKV[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10790.985 187.44 10791.265 188.44 ;
    END
  END MASKV[258]
  PIN MASKV[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10769.705 187.44 10769.985 188.44 ;
    END
  END MASKV[257]
  PIN MASKV[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10700.825 187.44 10701.105 188.44 ;
    END
  END MASKV[256]
  PIN MASKV[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10690.465 187.44 10690.745 188.44 ;
    END
  END MASKV[255]
  PIN MASKV[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10630.825 187.44 10631.105 188.44 ;
    END
  END MASKV[254]
  PIN MASKV[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10622.425 187.44 10622.705 188.44 ;
    END
  END MASKV[253]
  PIN MASKV[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10551.025 187.44 10551.305 188.44 ;
    END
  END MASKV[252]
  PIN MASKV[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10516.585 187.44 10516.865 188.44 ;
    END
  END MASKV[251]
  PIN MASKV[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10443.225 187.44 10443.505 188.44 ;
    END
  END MASKV[250]
  PIN MASKV[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10434.825 187.44 10435.105 188.44 ;
    END
  END MASKV[249]
  PIN MASKV[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10377.705 187.44 10377.985 188.44 ;
    END
  END MASKV[248]
  PIN MASKV[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10369.305 187.44 10369.585 188.44 ;
    END
  END MASKV[247]
  PIN MASKV[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10296.505 187.44 10296.785 188.44 ;
    END
  END MASKV[246]
  PIN MASKV[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10279.705 187.44 10279.985 188.44 ;
    END
  END MASKV[245]
  PIN MASKV[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10230.985 187.44 10231.265 188.44 ;
    END
  END MASKV[244]
  PIN MASKV[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10209.705 187.44 10209.985 188.44 ;
    END
  END MASKV[243]
  PIN MASKV[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10140.825 187.44 10141.105 188.44 ;
    END
  END MASKV[242]
  PIN MASKV[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10130.465 187.44 10130.745 188.44 ;
    END
  END MASKV[241]
  PIN MASKV[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10070.825 187.44 10071.105 188.44 ;
    END
  END MASKV[240]
  PIN MASKV[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10062.425 187.44 10062.705 188.44 ;
    END
  END MASKV[239]
  PIN MASKV[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9991.025 187.44 9991.305 188.44 ;
    END
  END MASKV[238]
  PIN MASKV[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9956.585 187.44 9956.865 188.44 ;
    END
  END MASKV[237]
  PIN MASKV[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9883.225 187.44 9883.505 188.44 ;
    END
  END MASKV[236]
  PIN MASKV[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9874.825 187.44 9875.105 188.44 ;
    END
  END MASKV[235]
  PIN MASKV[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9817.705 187.44 9817.985 188.44 ;
    END
  END MASKV[234]
  PIN MASKV[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9809.305 187.44 9809.585 188.44 ;
    END
  END MASKV[233]
  PIN MASKV[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9736.505 187.44 9736.785 188.44 ;
    END
  END MASKV[232]
  PIN MASKV[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9719.705 187.44 9719.985 188.44 ;
    END
  END MASKV[231]
  PIN MASKV[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9670.985 187.44 9671.265 188.44 ;
    END
  END MASKV[230]
  PIN MASKV[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9649.705 187.44 9649.985 188.44 ;
    END
  END MASKV[229]
  PIN MASKV[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9580.825 187.44 9581.105 188.44 ;
    END
  END MASKV[228]
  PIN MASKV[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9570.465 187.44 9570.745 188.44 ;
    END
  END MASKV[227]
  PIN MASKV[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9510.825 187.44 9511.105 188.44 ;
    END
  END MASKV[226]
  PIN MASKV[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9502.425 187.44 9502.705 188.44 ;
    END
  END MASKV[225]
  PIN MASKV[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9431.025 187.44 9431.305 188.44 ;
    END
  END MASKV[224]
  PIN MASKV[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9396.585 187.44 9396.865 188.44 ;
    END
  END MASKV[223]
  PIN MASKV[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9323.225 187.44 9323.505 188.44 ;
    END
  END MASKV[222]
  PIN MASKV[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9314.825 187.44 9315.105 188.44 ;
    END
  END MASKV[221]
  PIN MASKV[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9257.705 187.44 9257.985 188.44 ;
    END
  END MASKV[220]
  PIN MASKV[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9249.305 187.44 9249.585 188.44 ;
    END
  END MASKV[219]
  PIN MASKV[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9176.505 187.44 9176.785 188.44 ;
    END
  END MASKV[218]
  PIN MASKV[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9159.705 187.44 9159.985 188.44 ;
    END
  END MASKV[217]
  PIN MASKV[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9110.985 187.44 9111.265 188.44 ;
    END
  END MASKV[216]
  PIN MASKV[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9089.705 187.44 9089.985 188.44 ;
    END
  END MASKV[215]
  PIN MASKV[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9020.825 187.44 9021.105 188.44 ;
    END
  END MASKV[214]
  PIN MASKV[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9010.465 187.44 9010.745 188.44 ;
    END
  END MASKV[213]
  PIN MASKV[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8950.825 187.44 8951.105 188.44 ;
    END
  END MASKV[212]
  PIN MASKV[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8942.425 187.44 8942.705 188.44 ;
    END
  END MASKV[211]
  PIN MASKV[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8871.025 187.44 8871.305 188.44 ;
    END
  END MASKV[210]
  PIN MASKV[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8836.585 187.44 8836.865 188.44 ;
    END
  END MASKV[209]
  PIN MASKV[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8763.225 187.44 8763.505 188.44 ;
    END
  END MASKV[208]
  PIN MASKV[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8754.825 187.44 8755.105 188.44 ;
    END
  END MASKV[207]
  PIN MASKV[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8697.705 187.44 8697.985 188.44 ;
    END
  END MASKV[206]
  PIN MASKV[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8689.305 187.44 8689.585 188.44 ;
    END
  END MASKV[205]
  PIN MASKV[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8616.505 187.44 8616.785 188.44 ;
    END
  END MASKV[204]
  PIN MASKV[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8599.705 187.44 8599.985 188.44 ;
    END
  END MASKV[203]
  PIN MASKV[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8550.985 187.44 8551.265 188.44 ;
    END
  END MASKV[202]
  PIN MASKV[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8529.705 187.44 8529.985 188.44 ;
    END
  END MASKV[201]
  PIN MASKV[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8460.825 187.44 8461.105 188.44 ;
    END
  END MASKV[200]
  PIN MASKV[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8450.465 187.44 8450.745 188.44 ;
    END
  END MASKV[199]
  PIN MASKV[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8390.825 187.44 8391.105 188.44 ;
    END
  END MASKV[198]
  PIN MASKV[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8382.425 187.44 8382.705 188.44 ;
    END
  END MASKV[197]
  PIN MASKV[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8311.025 187.44 8311.305 188.44 ;
    END
  END MASKV[196]
  PIN MASKV[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8276.585 187.44 8276.865 188.44 ;
    END
  END MASKV[195]
  PIN MASKV[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8203.225 187.44 8203.505 188.44 ;
    END
  END MASKV[194]
  PIN MASKV[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8194.825 187.44 8195.105 188.44 ;
    END
  END MASKV[193]
  PIN MASKV[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8137.705 187.44 8137.985 188.44 ;
    END
  END MASKV[192]
  PIN MASKV[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8129.305 187.44 8129.585 188.44 ;
    END
  END MASKV[191]
  PIN MASKV[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8056.505 187.44 8056.785 188.44 ;
    END
  END MASKV[190]
  PIN MASKV[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8039.705 187.44 8039.985 188.44 ;
    END
  END MASKV[189]
  PIN MASKV[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7990.985 187.44 7991.265 188.44 ;
    END
  END MASKV[188]
  PIN MASKV[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7969.705 187.44 7969.985 188.44 ;
    END
  END MASKV[187]
  PIN MASKV[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7900.825 187.44 7901.105 188.44 ;
    END
  END MASKV[186]
  PIN MASKV[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7890.465 187.44 7890.745 188.44 ;
    END
  END MASKV[185]
  PIN MASKV[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7830.825 187.44 7831.105 188.44 ;
    END
  END MASKV[184]
  PIN MASKV[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7822.425 187.44 7822.705 188.44 ;
    END
  END MASKV[183]
  PIN MASKV[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7751.025 187.44 7751.305 188.44 ;
    END
  END MASKV[182]
  PIN MASKV[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7716.585 187.44 7716.865 188.44 ;
    END
  END MASKV[181]
  PIN MASKV[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7643.225 187.44 7643.505 188.44 ;
    END
  END MASKV[180]
  PIN MASKV[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7634.825 187.44 7635.105 188.44 ;
    END
  END MASKV[179]
  PIN MASKV[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7577.705 187.44 7577.985 188.44 ;
    END
  END MASKV[178]
  PIN MASKV[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7569.305 187.44 7569.585 188.44 ;
    END
  END MASKV[177]
  PIN MASKV[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7496.505 187.44 7496.785 188.44 ;
    END
  END MASKV[176]
  PIN MASKV[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7479.705 187.44 7479.985 188.44 ;
    END
  END MASKV[175]
  PIN MASKV[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7430.985 187.44 7431.265 188.44 ;
    END
  END MASKV[174]
  PIN MASKV[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7409.705 187.44 7409.985 188.44 ;
    END
  END MASKV[173]
  PIN MASKV[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7340.825 187.44 7341.105 188.44 ;
    END
  END MASKV[172]
  PIN MASKV[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7330.465 187.44 7330.745 188.44 ;
    END
  END MASKV[171]
  PIN MASKV[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7270.825 187.44 7271.105 188.44 ;
    END
  END MASKV[170]
  PIN MASKV[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7262.425 187.44 7262.705 188.44 ;
    END
  END MASKV[169]
  PIN MASKV[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7191.025 187.44 7191.305 188.44 ;
    END
  END MASKV[168]
  PIN MASKV[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7156.585 187.44 7156.865 188.44 ;
    END
  END MASKV[167]
  PIN MASKV[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7083.225 187.44 7083.505 188.44 ;
    END
  END MASKV[166]
  PIN MASKV[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7074.825 187.44 7075.105 188.44 ;
    END
  END MASKV[165]
  PIN MASKV[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7017.705 187.44 7017.985 188.44 ;
    END
  END MASKV[164]
  PIN MASKV[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7009.305 187.44 7009.585 188.44 ;
    END
  END MASKV[163]
  PIN MASKV[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6936.505 187.44 6936.785 188.44 ;
    END
  END MASKV[162]
  PIN MASKV[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6919.705 187.44 6919.985 188.44 ;
    END
  END MASKV[161]
  PIN MASKV[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6870.985 187.44 6871.265 188.44 ;
    END
  END MASKV[160]
  PIN MASKV[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6849.705 187.44 6849.985 188.44 ;
    END
  END MASKV[159]
  PIN MASKV[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6780.825 187.44 6781.105 188.44 ;
    END
  END MASKV[158]
  PIN MASKV[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6770.465 187.44 6770.745 188.44 ;
    END
  END MASKV[157]
  PIN MASKV[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6710.825 187.44 6711.105 188.44 ;
    END
  END MASKV[156]
  PIN MASKV[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6702.425 187.44 6702.705 188.44 ;
    END
  END MASKV[155]
  PIN MASKV[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6631.025 187.44 6631.305 188.44 ;
    END
  END MASKV[154]
  PIN MASKV[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6596.585 187.44 6596.865 188.44 ;
    END
  END MASKV[153]
  PIN MASKV[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6523.225 187.44 6523.505 188.44 ;
    END
  END MASKV[152]
  PIN MASKV[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6514.825 187.44 6515.105 188.44 ;
    END
  END MASKV[151]
  PIN MASKV[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6457.705 187.44 6457.985 188.44 ;
    END
  END MASKV[150]
  PIN MASKV[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6449.305 187.44 6449.585 188.44 ;
    END
  END MASKV[149]
  PIN MASKV[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6376.505 187.44 6376.785 188.44 ;
    END
  END MASKV[148]
  PIN MASKV[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6359.705 187.44 6359.985 188.44 ;
    END
  END MASKV[147]
  PIN MASKV[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6310.985 187.44 6311.265 188.44 ;
    END
  END MASKV[146]
  PIN MASKV[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6289.705 187.44 6289.985 188.44 ;
    END
  END MASKV[145]
  PIN MASKV[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6220.825 187.44 6221.105 188.44 ;
    END
  END MASKV[144]
  PIN MASKV[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6210.465 187.44 6210.745 188.44 ;
    END
  END MASKV[143]
  PIN MASKV[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6150.825 187.44 6151.105 188.44 ;
    END
  END MASKV[142]
  PIN MASKV[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6142.425 187.44 6142.705 188.44 ;
    END
  END MASKV[141]
  PIN MASKV[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6071.025 187.44 6071.305 188.44 ;
    END
  END MASKV[140]
  PIN MASKV[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6036.585 187.44 6036.865 188.44 ;
    END
  END MASKV[139]
  PIN MASKV[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5963.225 187.44 5963.505 188.44 ;
    END
  END MASKV[138]
  PIN MASKV[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5954.825 187.44 5955.105 188.44 ;
    END
  END MASKV[137]
  PIN MASKV[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5897.705 187.44 5897.985 188.44 ;
    END
  END MASKV[136]
  PIN MASKV[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5889.305 187.44 5889.585 188.44 ;
    END
  END MASKV[135]
  PIN MASKV[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5816.505 187.44 5816.785 188.44 ;
    END
  END MASKV[134]
  PIN MASKV[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5799.705 187.44 5799.985 188.44 ;
    END
  END MASKV[133]
  PIN MASKV[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5750.985 187.44 5751.265 188.44 ;
    END
  END MASKV[132]
  PIN MASKV[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5729.705 187.44 5729.985 188.44 ;
    END
  END MASKV[131]
  PIN MASKV[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5660.825 187.44 5661.105 188.44 ;
    END
  END MASKV[130]
  PIN MASKV[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5650.465 187.44 5650.745 188.44 ;
    END
  END MASKV[129]
  PIN MASKV[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5590.825 187.44 5591.105 188.44 ;
    END
  END MASKV[128]
  PIN MASKV[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5582.425 187.44 5582.705 188.44 ;
    END
  END MASKV[127]
  PIN MASKV[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5511.025 187.44 5511.305 188.44 ;
    END
  END MASKV[126]
  PIN MASKV[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5476.585 187.44 5476.865 188.44 ;
    END
  END MASKV[125]
  PIN MASKV[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5403.225 187.44 5403.505 188.44 ;
    END
  END MASKV[124]
  PIN MASKV[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5394.825 187.44 5395.105 188.44 ;
    END
  END MASKV[123]
  PIN MASKV[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5337.705 187.44 5337.985 188.44 ;
    END
  END MASKV[122]
  PIN MASKV[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5329.305 187.44 5329.585 188.44 ;
    END
  END MASKV[121]
  PIN MASKV[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5256.505 187.44 5256.785 188.44 ;
    END
  END MASKV[120]
  PIN MASKV[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5239.705 187.44 5239.985 188.44 ;
    END
  END MASKV[119]
  PIN MASKV[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5190.985 187.44 5191.265 188.44 ;
    END
  END MASKV[118]
  PIN MASKV[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5169.705 187.44 5169.985 188.44 ;
    END
  END MASKV[117]
  PIN MASKV[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5100.825 187.44 5101.105 188.44 ;
    END
  END MASKV[116]
  PIN MASKV[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5090.465 187.44 5090.745 188.44 ;
    END
  END MASKV[115]
  PIN MASKV[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5030.825 187.44 5031.105 188.44 ;
    END
  END MASKV[114]
  PIN MASKV[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5022.425 187.44 5022.705 188.44 ;
    END
  END MASKV[113]
  PIN MASKV[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4951.025 187.44 4951.305 188.44 ;
    END
  END MASKV[112]
  PIN MASKV[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4916.585 187.44 4916.865 188.44 ;
    END
  END MASKV[111]
  PIN MASKV[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4843.225 187.44 4843.505 188.44 ;
    END
  END MASKV[110]
  PIN MASKV[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4834.825 187.44 4835.105 188.44 ;
    END
  END MASKV[109]
  PIN MASKV[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4777.705 187.44 4777.985 188.44 ;
    END
  END MASKV[108]
  PIN MASKV[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4769.305 187.44 4769.585 188.44 ;
    END
  END MASKV[107]
  PIN MASKV[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4696.505 187.44 4696.785 188.44 ;
    END
  END MASKV[106]
  PIN MASKV[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4679.705 187.44 4679.985 188.44 ;
    END
  END MASKV[105]
  PIN MASKV[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4630.985 187.44 4631.265 188.44 ;
    END
  END MASKV[104]
  PIN MASKV[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4609.705 187.44 4609.985 188.44 ;
    END
  END MASKV[103]
  PIN MASKV[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4540.825 187.44 4541.105 188.44 ;
    END
  END MASKV[102]
  PIN MASKV[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4530.465 187.44 4530.745 188.44 ;
    END
  END MASKV[101]
  PIN MASKV[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4470.825 187.44 4471.105 188.44 ;
    END
  END MASKV[100]
  PIN MASKV[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4462.425 187.44 4462.705 188.44 ;
    END
  END MASKV[99]
  PIN MASKV[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4391.025 187.44 4391.305 188.44 ;
    END
  END MASKV[98]
  PIN MASKV[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4356.585 187.44 4356.865 188.44 ;
    END
  END MASKV[97]
  PIN MASKV[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4283.225 187.44 4283.505 188.44 ;
    END
  END MASKV[96]
  PIN MASKV[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4274.825 187.44 4275.105 188.44 ;
    END
  END MASKV[95]
  PIN MASKV[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4217.705 187.44 4217.985 188.44 ;
    END
  END MASKV[94]
  PIN MASKV[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4209.305 187.44 4209.585 188.44 ;
    END
  END MASKV[93]
  PIN MASKV[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4136.505 187.44 4136.785 188.44 ;
    END
  END MASKV[92]
  PIN MASKV[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4119.705 187.44 4119.985 188.44 ;
    END
  END MASKV[91]
  PIN MASKV[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4070.985 187.44 4071.265 188.44 ;
    END
  END MASKV[90]
  PIN MASKV[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4049.705 187.44 4049.985 188.44 ;
    END
  END MASKV[89]
  PIN MASKV[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3980.825 187.44 3981.105 188.44 ;
    END
  END MASKV[88]
  PIN MASKV[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3970.465 187.44 3970.745 188.44 ;
    END
  END MASKV[87]
  PIN MASKV[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3910.825 187.44 3911.105 188.44 ;
    END
  END MASKV[86]
  PIN MASKV[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3902.425 187.44 3902.705 188.44 ;
    END
  END MASKV[85]
  PIN MASKV[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3831.025 187.44 3831.305 188.44 ;
    END
  END MASKV[84]
  PIN MASKV[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3796.585 187.44 3796.865 188.44 ;
    END
  END MASKV[83]
  PIN MASKV[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3723.225 187.44 3723.505 188.44 ;
    END
  END MASKV[82]
  PIN MASKV[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3714.825 187.44 3715.105 188.44 ;
    END
  END MASKV[81]
  PIN MASKV[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3657.705 187.44 3657.985 188.44 ;
    END
  END MASKV[80]
  PIN MASKV[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3649.305 187.44 3649.585 188.44 ;
    END
  END MASKV[79]
  PIN MASKV[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3576.505 187.44 3576.785 188.44 ;
    END
  END MASKV[78]
  PIN MASKV[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3559.705 187.44 3559.985 188.44 ;
    END
  END MASKV[77]
  PIN MASKV[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3510.985 187.44 3511.265 188.44 ;
    END
  END MASKV[76]
  PIN MASKV[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3489.705 187.44 3489.985 188.44 ;
    END
  END MASKV[75]
  PIN MASKV[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3420.825 187.44 3421.105 188.44 ;
    END
  END MASKV[74]
  PIN MASKV[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3410.465 187.44 3410.745 188.44 ;
    END
  END MASKV[73]
  PIN MASKV[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3350.825 187.44 3351.105 188.44 ;
    END
  END MASKV[72]
  PIN MASKV[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3342.425 187.44 3342.705 188.44 ;
    END
  END MASKV[71]
  PIN MASKV[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3271.025 187.44 3271.305 188.44 ;
    END
  END MASKV[70]
  PIN MASKV[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3236.585 187.44 3236.865 188.44 ;
    END
  END MASKV[69]
  PIN MASKV[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3163.225 187.44 3163.505 188.44 ;
    END
  END MASKV[68]
  PIN MASKV[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3154.825 187.44 3155.105 188.44 ;
    END
  END MASKV[67]
  PIN MASKV[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3097.705 187.44 3097.985 188.44 ;
    END
  END MASKV[66]
  PIN MASKV[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3089.305 187.44 3089.585 188.44 ;
    END
  END MASKV[65]
  PIN MASKV[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3016.505 187.44 3016.785 188.44 ;
    END
  END MASKV[64]
  PIN MASKV[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2999.705 187.44 2999.985 188.44 ;
    END
  END MASKV[63]
  PIN MASKV[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2950.985 187.44 2951.265 188.44 ;
    END
  END MASKV[62]
  PIN MASKV[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2929.705 187.44 2929.985 188.44 ;
    END
  END MASKV[61]
  PIN MASKV[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2860.825 187.44 2861.105 188.44 ;
    END
  END MASKV[60]
  PIN MASKV[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2850.465 187.44 2850.745 188.44 ;
    END
  END MASKV[59]
  PIN MASKV[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2790.825 187.44 2791.105 188.44 ;
    END
  END MASKV[58]
  PIN MASKV[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2782.425 187.44 2782.705 188.44 ;
    END
  END MASKV[57]
  PIN MASKV[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2711.025 187.44 2711.305 188.44 ;
    END
  END MASKV[56]
  PIN MASKV[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2676.585 187.44 2676.865 188.44 ;
    END
  END MASKV[55]
  PIN MASKV[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2603.225 187.44 2603.505 188.44 ;
    END
  END MASKV[54]
  PIN MASKV[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2594.825 187.44 2595.105 188.44 ;
    END
  END MASKV[53]
  PIN MASKV[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2537.705 187.44 2537.985 188.44 ;
    END
  END MASKV[52]
  PIN MASKV[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2529.305 187.44 2529.585 188.44 ;
    END
  END MASKV[51]
  PIN MASKV[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2456.505 187.44 2456.785 188.44 ;
    END
  END MASKV[50]
  PIN MASKV[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2439.705 187.44 2439.985 188.44 ;
    END
  END MASKV[49]
  PIN MASKV[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2390.985 187.44 2391.265 188.44 ;
    END
  END MASKV[48]
  PIN MASKV[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2369.705 187.44 2369.985 188.44 ;
    END
  END MASKV[47]
  PIN MASKV[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2300.825 187.44 2301.105 188.44 ;
    END
  END MASKV[46]
  PIN MASKV[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2290.465 187.44 2290.745 188.44 ;
    END
  END MASKV[45]
  PIN MASKV[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2230.825 187.44 2231.105 188.44 ;
    END
  END MASKV[44]
  PIN MASKV[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2222.425 187.44 2222.705 188.44 ;
    END
  END MASKV[43]
  PIN MASKV[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2151.025 187.44 2151.305 188.44 ;
    END
  END MASKV[42]
  PIN MASKV[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2116.585 187.44 2116.865 188.44 ;
    END
  END MASKV[41]
  PIN MASKV[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2043.225 187.44 2043.505 188.44 ;
    END
  END MASKV[40]
  PIN MASKV[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2034.825 187.44 2035.105 188.44 ;
    END
  END MASKV[39]
  PIN MASKV[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1977.705 187.44 1977.985 188.44 ;
    END
  END MASKV[38]
  PIN MASKV[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1969.305 187.44 1969.585 188.44 ;
    END
  END MASKV[37]
  PIN MASKV[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1896.505 187.44 1896.785 188.44 ;
    END
  END MASKV[36]
  PIN MASKV[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1879.705 187.44 1879.985 188.44 ;
    END
  END MASKV[35]
  PIN MASKV[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1830.985 187.44 1831.265 188.44 ;
    END
  END MASKV[34]
  PIN MASKV[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1809.705 187.44 1809.985 188.44 ;
    END
  END MASKV[33]
  PIN MASKV[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1740.825 187.44 1741.105 188.44 ;
    END
  END MASKV[32]
  PIN MASKV[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1730.465 187.44 1730.745 188.44 ;
    END
  END MASKV[31]
  PIN MASKV[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1670.825 187.44 1671.105 188.44 ;
    END
  END MASKV[30]
  PIN MASKV[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1662.425 187.44 1662.705 188.44 ;
    END
  END MASKV[29]
  PIN MASKV[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1591.025 187.44 1591.305 188.44 ;
    END
  END MASKV[28]
  PIN MASKV[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1556.585 187.44 1556.865 188.44 ;
    END
  END MASKV[27]
  PIN MASKV[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1483.225 187.44 1483.505 188.44 ;
    END
  END MASKV[26]
  PIN MASKV[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1474.825 187.44 1475.105 188.44 ;
    END
  END MASKV[25]
  PIN MASKV[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1417.705 187.44 1417.985 188.44 ;
    END
  END MASKV[24]
  PIN MASKV[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1409.305 187.44 1409.585 188.44 ;
    END
  END MASKV[23]
  PIN MASKV[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1336.505 187.44 1336.785 188.44 ;
    END
  END MASKV[22]
  PIN MASKV[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1319.705 187.44 1319.985 188.44 ;
    END
  END MASKV[21]
  PIN MASKV[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1270.985 187.44 1271.265 188.44 ;
    END
  END MASKV[20]
  PIN MASKV[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1249.705 187.44 1249.985 188.44 ;
    END
  END MASKV[19]
  PIN MASKV[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1180.825 187.44 1181.105 188.44 ;
    END
  END MASKV[18]
  PIN MASKV[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1170.465 187.44 1170.745 188.44 ;
    END
  END MASKV[17]
  PIN MASKV[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1110.825 187.44 1111.105 188.44 ;
    END
  END MASKV[16]
  PIN MASKV[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1102.425 187.44 1102.705 188.44 ;
    END
  END MASKV[15]
  PIN MASKV[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1031.025 187.44 1031.305 188.44 ;
    END
  END MASKV[14]
  PIN MASKV[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 996.585 187.44 996.865 188.44 ;
    END
  END MASKV[13]
  PIN MASKV[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 923.225 187.44 923.505 188.44 ;
    END
  END MASKV[12]
  PIN MASKV[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 914.825 187.44 915.105 188.44 ;
    END
  END MASKV[11]
  PIN MASKV[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 857.705 187.44 857.985 188.44 ;
    END
  END MASKV[10]
  PIN MASKV[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 849.305 187.44 849.585 188.44 ;
    END
  END MASKV[9]
  PIN MASKV[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 776.505 187.44 776.785 188.44 ;
    END
  END MASKV[8]
  PIN MASKV[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 759.705 187.44 759.985 188.44 ;
    END
  END MASKV[7]
  PIN MASKV[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 710.985 187.44 711.265 188.44 ;
    END
  END MASKV[6]
  PIN MASKV[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 689.705 187.44 689.985 188.44 ;
    END
  END MASKV[5]
  PIN MASKV[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 620.825 187.44 621.105 188.44 ;
    END
  END MASKV[4]
  PIN MASKV[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 610.465 187.44 610.745 188.44 ;
    END
  END MASKV[3]
  PIN MASKV[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 550.825 187.44 551.105 188.44 ;
    END
  END MASKV[2]
  PIN MASKV[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 542.425 187.44 542.705 188.44 ;
    END
  END MASKV[1]
  PIN MASKV[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 471.025 187.44 471.305 188.44 ;
    END
  END MASKV[0]
  PIN INJ_ROW[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18357.145 187.44 18357.425 188.44 ;
    END
  END INJ_ROW[223]
  PIN INJ_ROW[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18275.385 187.44 18275.665 188.44 ;
    END
  END INJ_ROW[222]
  PIN INJ_ROW[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18209.865 187.44 18210.145 188.44 ;
    END
  END INJ_ROW[221]
  PIN INJ_ROW[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18120.265 187.44 18120.545 188.44 ;
    END
  END INJ_ROW[220]
  PIN INJ_ROW[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18050.265 187.44 18050.545 188.44 ;
    END
  END INJ_ROW[219]
  PIN INJ_ROW[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17971.025 187.44 17971.305 188.44 ;
    END
  END INJ_ROW[218]
  PIN INJ_ROW[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17902.985 187.44 17903.265 188.44 ;
    END
  END INJ_ROW[217]
  PIN INJ_ROW[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17797.145 187.44 17797.425 188.44 ;
    END
  END INJ_ROW[216]
  PIN INJ_ROW[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17715.385 187.44 17715.665 188.44 ;
    END
  END INJ_ROW[215]
  PIN INJ_ROW[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17649.865 187.44 17650.145 188.44 ;
    END
  END INJ_ROW[214]
  PIN INJ_ROW[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17560.265 187.44 17560.545 188.44 ;
    END
  END INJ_ROW[213]
  PIN INJ_ROW[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17490.265 187.44 17490.545 188.44 ;
    END
  END INJ_ROW[212]
  PIN INJ_ROW[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17411.025 187.44 17411.305 188.44 ;
    END
  END INJ_ROW[211]
  PIN INJ_ROW[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17342.985 187.44 17343.265 188.44 ;
    END
  END INJ_ROW[210]
  PIN INJ_ROW[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17237.145 187.44 17237.425 188.44 ;
    END
  END INJ_ROW[209]
  PIN INJ_ROW[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17155.385 187.44 17155.665 188.44 ;
    END
  END INJ_ROW[208]
  PIN INJ_ROW[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17089.865 187.44 17090.145 188.44 ;
    END
  END INJ_ROW[207]
  PIN INJ_ROW[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17000.265 187.44 17000.545 188.44 ;
    END
  END INJ_ROW[206]
  PIN INJ_ROW[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16930.265 187.44 16930.545 188.44 ;
    END
  END INJ_ROW[205]
  PIN INJ_ROW[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16851.025 187.44 16851.305 188.44 ;
    END
  END INJ_ROW[204]
  PIN INJ_ROW[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16782.985 187.44 16783.265 188.44 ;
    END
  END INJ_ROW[203]
  PIN INJ_ROW[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16677.145 187.44 16677.425 188.44 ;
    END
  END INJ_ROW[202]
  PIN INJ_ROW[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16595.385 187.44 16595.665 188.44 ;
    END
  END INJ_ROW[201]
  PIN INJ_ROW[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16529.865 187.44 16530.145 188.44 ;
    END
  END INJ_ROW[200]
  PIN INJ_ROW[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16440.265 187.44 16440.545 188.44 ;
    END
  END INJ_ROW[199]
  PIN INJ_ROW[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16370.265 187.44 16370.545 188.44 ;
    END
  END INJ_ROW[198]
  PIN INJ_ROW[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16291.025 187.44 16291.305 188.44 ;
    END
  END INJ_ROW[197]
  PIN INJ_ROW[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16222.985 187.44 16223.265 188.44 ;
    END
  END INJ_ROW[196]
  PIN INJ_ROW[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16117.145 187.44 16117.425 188.44 ;
    END
  END INJ_ROW[195]
  PIN INJ_ROW[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16035.385 187.44 16035.665 188.44 ;
    END
  END INJ_ROW[194]
  PIN INJ_ROW[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15969.865 187.44 15970.145 188.44 ;
    END
  END INJ_ROW[193]
  PIN INJ_ROW[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15880.265 187.44 15880.545 188.44 ;
    END
  END INJ_ROW[192]
  PIN INJ_ROW[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15810.265 187.44 15810.545 188.44 ;
    END
  END INJ_ROW[191]
  PIN INJ_ROW[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15731.025 187.44 15731.305 188.44 ;
    END
  END INJ_ROW[190]
  PIN INJ_ROW[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15662.985 187.44 15663.265 188.44 ;
    END
  END INJ_ROW[189]
  PIN INJ_ROW[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15557.145 187.44 15557.425 188.44 ;
    END
  END INJ_ROW[188]
  PIN INJ_ROW[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15475.385 187.44 15475.665 188.44 ;
    END
  END INJ_ROW[187]
  PIN INJ_ROW[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15409.865 187.44 15410.145 188.44 ;
    END
  END INJ_ROW[186]
  PIN INJ_ROW[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15320.265 187.44 15320.545 188.44 ;
    END
  END INJ_ROW[185]
  PIN INJ_ROW[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15250.265 187.44 15250.545 188.44 ;
    END
  END INJ_ROW[184]
  PIN INJ_ROW[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15171.025 187.44 15171.305 188.44 ;
    END
  END INJ_ROW[183]
  PIN INJ_ROW[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15102.985 187.44 15103.265 188.44 ;
    END
  END INJ_ROW[182]
  PIN INJ_ROW[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14997.145 187.44 14997.425 188.44 ;
    END
  END INJ_ROW[181]
  PIN INJ_ROW[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14915.385 187.44 14915.665 188.44 ;
    END
  END INJ_ROW[180]
  PIN INJ_ROW[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14849.865 187.44 14850.145 188.44 ;
    END
  END INJ_ROW[179]
  PIN INJ_ROW[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14760.265 187.44 14760.545 188.44 ;
    END
  END INJ_ROW[178]
  PIN INJ_ROW[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14690.265 187.44 14690.545 188.44 ;
    END
  END INJ_ROW[177]
  PIN INJ_ROW[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14611.025 187.44 14611.305 188.44 ;
    END
  END INJ_ROW[176]
  PIN INJ_ROW[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14542.985 187.44 14543.265 188.44 ;
    END
  END INJ_ROW[175]
  PIN INJ_ROW[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14437.145 187.44 14437.425 188.44 ;
    END
  END INJ_ROW[174]
  PIN INJ_ROW[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14355.385 187.44 14355.665 188.44 ;
    END
  END INJ_ROW[173]
  PIN INJ_ROW[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14289.865 187.44 14290.145 188.44 ;
    END
  END INJ_ROW[172]
  PIN INJ_ROW[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14200.265 187.44 14200.545 188.44 ;
    END
  END INJ_ROW[171]
  PIN INJ_ROW[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14130.265 187.44 14130.545 188.44 ;
    END
  END INJ_ROW[170]
  PIN INJ_ROW[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14051.025 187.44 14051.305 188.44 ;
    END
  END INJ_ROW[169]
  PIN INJ_ROW[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13982.985 187.44 13983.265 188.44 ;
    END
  END INJ_ROW[168]
  PIN INJ_ROW[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13877.145 187.44 13877.425 188.44 ;
    END
  END INJ_ROW[167]
  PIN INJ_ROW[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13795.385 187.44 13795.665 188.44 ;
    END
  END INJ_ROW[166]
  PIN INJ_ROW[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13729.865 187.44 13730.145 188.44 ;
    END
  END INJ_ROW[165]
  PIN INJ_ROW[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13640.265 187.44 13640.545 188.44 ;
    END
  END INJ_ROW[164]
  PIN INJ_ROW[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13570.265 187.44 13570.545 188.44 ;
    END
  END INJ_ROW[163]
  PIN INJ_ROW[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13491.025 187.44 13491.305 188.44 ;
    END
  END INJ_ROW[162]
  PIN INJ_ROW[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13422.985 187.44 13423.265 188.44 ;
    END
  END INJ_ROW[161]
  PIN INJ_ROW[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13317.145 187.44 13317.425 188.44 ;
    END
  END INJ_ROW[160]
  PIN INJ_ROW[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13235.385 187.44 13235.665 188.44 ;
    END
  END INJ_ROW[159]
  PIN INJ_ROW[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13169.865 187.44 13170.145 188.44 ;
    END
  END INJ_ROW[158]
  PIN INJ_ROW[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13080.265 187.44 13080.545 188.44 ;
    END
  END INJ_ROW[157]
  PIN INJ_ROW[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13010.265 187.44 13010.545 188.44 ;
    END
  END INJ_ROW[156]
  PIN INJ_ROW[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12931.025 187.44 12931.305 188.44 ;
    END
  END INJ_ROW[155]
  PIN INJ_ROW[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12862.985 187.44 12863.265 188.44 ;
    END
  END INJ_ROW[154]
  PIN INJ_ROW[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12757.145 187.44 12757.425 188.44 ;
    END
  END INJ_ROW[153]
  PIN INJ_ROW[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12675.385 187.44 12675.665 188.44 ;
    END
  END INJ_ROW[152]
  PIN INJ_ROW[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12609.865 187.44 12610.145 188.44 ;
    END
  END INJ_ROW[151]
  PIN INJ_ROW[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12520.265 187.44 12520.545 188.44 ;
    END
  END INJ_ROW[150]
  PIN INJ_ROW[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12450.265 187.44 12450.545 188.44 ;
    END
  END INJ_ROW[149]
  PIN INJ_ROW[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12371.025 187.44 12371.305 188.44 ;
    END
  END INJ_ROW[148]
  PIN INJ_ROW[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12302.985 187.44 12303.265 188.44 ;
    END
  END INJ_ROW[147]
  PIN INJ_ROW[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12197.145 187.44 12197.425 188.44 ;
    END
  END INJ_ROW[146]
  PIN INJ_ROW[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12115.385 187.44 12115.665 188.44 ;
    END
  END INJ_ROW[145]
  PIN INJ_ROW[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12049.865 187.44 12050.145 188.44 ;
    END
  END INJ_ROW[144]
  PIN INJ_ROW[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11960.265 187.44 11960.545 188.44 ;
    END
  END INJ_ROW[143]
  PIN INJ_ROW[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11890.265 187.44 11890.545 188.44 ;
    END
  END INJ_ROW[142]
  PIN INJ_ROW[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11811.025 187.44 11811.305 188.44 ;
    END
  END INJ_ROW[141]
  PIN INJ_ROW[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11742.985 187.44 11743.265 188.44 ;
    END
  END INJ_ROW[140]
  PIN INJ_ROW[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11637.145 187.44 11637.425 188.44 ;
    END
  END INJ_ROW[139]
  PIN INJ_ROW[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11555.385 187.44 11555.665 188.44 ;
    END
  END INJ_ROW[138]
  PIN INJ_ROW[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11489.865 187.44 11490.145 188.44 ;
    END
  END INJ_ROW[137]
  PIN INJ_ROW[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11400.265 187.44 11400.545 188.44 ;
    END
  END INJ_ROW[136]
  PIN INJ_ROW[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11330.265 187.44 11330.545 188.44 ;
    END
  END INJ_ROW[135]
  PIN INJ_ROW[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11251.025 187.44 11251.305 188.44 ;
    END
  END INJ_ROW[134]
  PIN INJ_ROW[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11182.985 187.44 11183.265 188.44 ;
    END
  END INJ_ROW[133]
  PIN INJ_ROW[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11077.145 187.44 11077.425 188.44 ;
    END
  END INJ_ROW[132]
  PIN INJ_ROW[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10995.385 187.44 10995.665 188.44 ;
    END
  END INJ_ROW[131]
  PIN INJ_ROW[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10929.865 187.44 10930.145 188.44 ;
    END
  END INJ_ROW[130]
  PIN INJ_ROW[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10840.265 187.44 10840.545 188.44 ;
    END
  END INJ_ROW[129]
  PIN INJ_ROW[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10770.265 187.44 10770.545 188.44 ;
    END
  END INJ_ROW[128]
  PIN INJ_ROW[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10691.025 187.44 10691.305 188.44 ;
    END
  END INJ_ROW[127]
  PIN INJ_ROW[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10622.985 187.44 10623.265 188.44 ;
    END
  END INJ_ROW[126]
  PIN INJ_ROW[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10517.145 187.44 10517.425 188.44 ;
    END
  END INJ_ROW[125]
  PIN INJ_ROW[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10435.385 187.44 10435.665 188.44 ;
    END
  END INJ_ROW[124]
  PIN INJ_ROW[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10369.865 187.44 10370.145 188.44 ;
    END
  END INJ_ROW[123]
  PIN INJ_ROW[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10280.265 187.44 10280.545 188.44 ;
    END
  END INJ_ROW[122]
  PIN INJ_ROW[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10210.265 187.44 10210.545 188.44 ;
    END
  END INJ_ROW[121]
  PIN INJ_ROW[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10131.025 187.44 10131.305 188.44 ;
    END
  END INJ_ROW[120]
  PIN INJ_ROW[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10062.985 187.44 10063.265 188.44 ;
    END
  END INJ_ROW[119]
  PIN INJ_ROW[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9957.145 187.44 9957.425 188.44 ;
    END
  END INJ_ROW[118]
  PIN INJ_ROW[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9875.385 187.44 9875.665 188.44 ;
    END
  END INJ_ROW[117]
  PIN INJ_ROW[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9809.865 187.44 9810.145 188.44 ;
    END
  END INJ_ROW[116]
  PIN INJ_ROW[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9720.265 187.44 9720.545 188.44 ;
    END
  END INJ_ROW[115]
  PIN INJ_ROW[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9650.265 187.44 9650.545 188.44 ;
    END
  END INJ_ROW[114]
  PIN INJ_ROW[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9571.025 187.44 9571.305 188.44 ;
    END
  END INJ_ROW[113]
  PIN INJ_ROW[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9502.985 187.44 9503.265 188.44 ;
    END
  END INJ_ROW[112]
  PIN INJ_ROW[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9397.145 187.44 9397.425 188.44 ;
    END
  END INJ_ROW[111]
  PIN INJ_ROW[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9315.385 187.44 9315.665 188.44 ;
    END
  END INJ_ROW[110]
  PIN INJ_ROW[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9249.865 187.44 9250.145 188.44 ;
    END
  END INJ_ROW[109]
  PIN INJ_ROW[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9160.265 187.44 9160.545 188.44 ;
    END
  END INJ_ROW[108]
  PIN INJ_ROW[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9090.265 187.44 9090.545 188.44 ;
    END
  END INJ_ROW[107]
  PIN INJ_ROW[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9011.025 187.44 9011.305 188.44 ;
    END
  END INJ_ROW[106]
  PIN INJ_ROW[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8942.985 187.44 8943.265 188.44 ;
    END
  END INJ_ROW[105]
  PIN INJ_ROW[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8837.145 187.44 8837.425 188.44 ;
    END
  END INJ_ROW[104]
  PIN INJ_ROW[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8755.385 187.44 8755.665 188.44 ;
    END
  END INJ_ROW[103]
  PIN INJ_ROW[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8689.865 187.44 8690.145 188.44 ;
    END
  END INJ_ROW[102]
  PIN INJ_ROW[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8600.265 187.44 8600.545 188.44 ;
    END
  END INJ_ROW[101]
  PIN INJ_ROW[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8530.265 187.44 8530.545 188.44 ;
    END
  END INJ_ROW[100]
  PIN INJ_ROW[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8451.025 187.44 8451.305 188.44 ;
    END
  END INJ_ROW[99]
  PIN INJ_ROW[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8382.985 187.44 8383.265 188.44 ;
    END
  END INJ_ROW[98]
  PIN INJ_ROW[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8277.145 187.44 8277.425 188.44 ;
    END
  END INJ_ROW[97]
  PIN INJ_ROW[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8195.385 187.44 8195.665 188.44 ;
    END
  END INJ_ROW[96]
  PIN INJ_ROW[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8129.865 187.44 8130.145 188.44 ;
    END
  END INJ_ROW[95]
  PIN INJ_ROW[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8040.265 187.44 8040.545 188.44 ;
    END
  END INJ_ROW[94]
  PIN INJ_ROW[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7970.265 187.44 7970.545 188.44 ;
    END
  END INJ_ROW[93]
  PIN INJ_ROW[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7891.025 187.44 7891.305 188.44 ;
    END
  END INJ_ROW[92]
  PIN INJ_ROW[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7822.985 187.44 7823.265 188.44 ;
    END
  END INJ_ROW[91]
  PIN INJ_ROW[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7717.145 187.44 7717.425 188.44 ;
    END
  END INJ_ROW[90]
  PIN INJ_ROW[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7635.385 187.44 7635.665 188.44 ;
    END
  END INJ_ROW[89]
  PIN INJ_ROW[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7569.865 187.44 7570.145 188.44 ;
    END
  END INJ_ROW[88]
  PIN INJ_ROW[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7480.265 187.44 7480.545 188.44 ;
    END
  END INJ_ROW[87]
  PIN INJ_ROW[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7410.265 187.44 7410.545 188.44 ;
    END
  END INJ_ROW[86]
  PIN INJ_ROW[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7331.025 187.44 7331.305 188.44 ;
    END
  END INJ_ROW[85]
  PIN INJ_ROW[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7262.985 187.44 7263.265 188.44 ;
    END
  END INJ_ROW[84]
  PIN INJ_ROW[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7157.145 187.44 7157.425 188.44 ;
    END
  END INJ_ROW[83]
  PIN INJ_ROW[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7075.385 187.44 7075.665 188.44 ;
    END
  END INJ_ROW[82]
  PIN INJ_ROW[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7009.865 187.44 7010.145 188.44 ;
    END
  END INJ_ROW[81]
  PIN INJ_ROW[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6920.265 187.44 6920.545 188.44 ;
    END
  END INJ_ROW[80]
  PIN INJ_ROW[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6850.265 187.44 6850.545 188.44 ;
    END
  END INJ_ROW[79]
  PIN INJ_ROW[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6771.025 187.44 6771.305 188.44 ;
    END
  END INJ_ROW[78]
  PIN INJ_ROW[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6702.985 187.44 6703.265 188.44 ;
    END
  END INJ_ROW[77]
  PIN INJ_ROW[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6597.145 187.44 6597.425 188.44 ;
    END
  END INJ_ROW[76]
  PIN INJ_ROW[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6515.385 187.44 6515.665 188.44 ;
    END
  END INJ_ROW[75]
  PIN INJ_ROW[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6449.865 187.44 6450.145 188.44 ;
    END
  END INJ_ROW[74]
  PIN INJ_ROW[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6360.265 187.44 6360.545 188.44 ;
    END
  END INJ_ROW[73]
  PIN INJ_ROW[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6290.265 187.44 6290.545 188.44 ;
    END
  END INJ_ROW[72]
  PIN INJ_ROW[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6211.025 187.44 6211.305 188.44 ;
    END
  END INJ_ROW[71]
  PIN INJ_ROW[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6142.985 187.44 6143.265 188.44 ;
    END
  END INJ_ROW[70]
  PIN INJ_ROW[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6037.145 187.44 6037.425 188.44 ;
    END
  END INJ_ROW[69]
  PIN INJ_ROW[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5955.385 187.44 5955.665 188.44 ;
    END
  END INJ_ROW[68]
  PIN INJ_ROW[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5889.865 187.44 5890.145 188.44 ;
    END
  END INJ_ROW[67]
  PIN INJ_ROW[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5800.265 187.44 5800.545 188.44 ;
    END
  END INJ_ROW[66]
  PIN INJ_ROW[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5730.265 187.44 5730.545 188.44 ;
    END
  END INJ_ROW[65]
  PIN INJ_ROW[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5651.025 187.44 5651.305 188.44 ;
    END
  END INJ_ROW[64]
  PIN INJ_ROW[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5582.985 187.44 5583.265 188.44 ;
    END
  END INJ_ROW[63]
  PIN INJ_ROW[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5477.145 187.44 5477.425 188.44 ;
    END
  END INJ_ROW[62]
  PIN INJ_ROW[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5395.385 187.44 5395.665 188.44 ;
    END
  END INJ_ROW[61]
  PIN INJ_ROW[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5329.865 187.44 5330.145 188.44 ;
    END
  END INJ_ROW[60]
  PIN INJ_ROW[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5240.265 187.44 5240.545 188.44 ;
    END
  END INJ_ROW[59]
  PIN INJ_ROW[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5170.265 187.44 5170.545 188.44 ;
    END
  END INJ_ROW[58]
  PIN INJ_ROW[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5091.025 187.44 5091.305 188.44 ;
    END
  END INJ_ROW[57]
  PIN INJ_ROW[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5022.985 187.44 5023.265 188.44 ;
    END
  END INJ_ROW[56]
  PIN INJ_ROW[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4917.145 187.44 4917.425 188.44 ;
    END
  END INJ_ROW[55]
  PIN INJ_ROW[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4835.385 187.44 4835.665 188.44 ;
    END
  END INJ_ROW[54]
  PIN INJ_ROW[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4769.865 187.44 4770.145 188.44 ;
    END
  END INJ_ROW[53]
  PIN INJ_ROW[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4680.265 187.44 4680.545 188.44 ;
    END
  END INJ_ROW[52]
  PIN INJ_ROW[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4610.265 187.44 4610.545 188.44 ;
    END
  END INJ_ROW[51]
  PIN INJ_ROW[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4531.025 187.44 4531.305 188.44 ;
    END
  END INJ_ROW[50]
  PIN INJ_ROW[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4462.985 187.44 4463.265 188.44 ;
    END
  END INJ_ROW[49]
  PIN INJ_ROW[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4357.145 187.44 4357.425 188.44 ;
    END
  END INJ_ROW[48]
  PIN INJ_ROW[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4275.385 187.44 4275.665 188.44 ;
    END
  END INJ_ROW[47]
  PIN INJ_ROW[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4209.865 187.44 4210.145 188.44 ;
    END
  END INJ_ROW[46]
  PIN INJ_ROW[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4120.265 187.44 4120.545 188.44 ;
    END
  END INJ_ROW[45]
  PIN INJ_ROW[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4050.265 187.44 4050.545 188.44 ;
    END
  END INJ_ROW[44]
  PIN INJ_ROW[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3971.025 187.44 3971.305 188.44 ;
    END
  END INJ_ROW[43]
  PIN INJ_ROW[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3902.985 187.44 3903.265 188.44 ;
    END
  END INJ_ROW[42]
  PIN INJ_ROW[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3797.145 187.44 3797.425 188.44 ;
    END
  END INJ_ROW[41]
  PIN INJ_ROW[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3715.385 187.44 3715.665 188.44 ;
    END
  END INJ_ROW[40]
  PIN INJ_ROW[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3649.865 187.44 3650.145 188.44 ;
    END
  END INJ_ROW[39]
  PIN INJ_ROW[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3560.265 187.44 3560.545 188.44 ;
    END
  END INJ_ROW[38]
  PIN INJ_ROW[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3490.265 187.44 3490.545 188.44 ;
    END
  END INJ_ROW[37]
  PIN INJ_ROW[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3411.025 187.44 3411.305 188.44 ;
    END
  END INJ_ROW[36]
  PIN INJ_ROW[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3342.985 187.44 3343.265 188.44 ;
    END
  END INJ_ROW[35]
  PIN INJ_ROW[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3237.145 187.44 3237.425 188.44 ;
    END
  END INJ_ROW[34]
  PIN INJ_ROW[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3155.385 187.44 3155.665 188.44 ;
    END
  END INJ_ROW[33]
  PIN INJ_ROW[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3089.865 187.44 3090.145 188.44 ;
    END
  END INJ_ROW[32]
  PIN INJ_ROW[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3000.265 187.44 3000.545 188.44 ;
    END
  END INJ_ROW[31]
  PIN INJ_ROW[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2930.265 187.44 2930.545 188.44 ;
    END
  END INJ_ROW[30]
  PIN INJ_ROW[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2851.025 187.44 2851.305 188.44 ;
    END
  END INJ_ROW[29]
  PIN INJ_ROW[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2782.985 187.44 2783.265 188.44 ;
    END
  END INJ_ROW[28]
  PIN INJ_ROW[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2677.145 187.44 2677.425 188.44 ;
    END
  END INJ_ROW[27]
  PIN INJ_ROW[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2595.385 187.44 2595.665 188.44 ;
    END
  END INJ_ROW[26]
  PIN INJ_ROW[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2529.865 187.44 2530.145 188.44 ;
    END
  END INJ_ROW[25]
  PIN INJ_ROW[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2440.265 187.44 2440.545 188.44 ;
    END
  END INJ_ROW[24]
  PIN INJ_ROW[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2370.265 187.44 2370.545 188.44 ;
    END
  END INJ_ROW[23]
  PIN INJ_ROW[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2291.025 187.44 2291.305 188.44 ;
    END
  END INJ_ROW[22]
  PIN INJ_ROW[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2222.985 187.44 2223.265 188.44 ;
    END
  END INJ_ROW[21]
  PIN INJ_ROW[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2117.145 187.44 2117.425 188.44 ;
    END
  END INJ_ROW[20]
  PIN INJ_ROW[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2035.385 187.44 2035.665 188.44 ;
    END
  END INJ_ROW[19]
  PIN INJ_ROW[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1969.865 187.44 1970.145 188.44 ;
    END
  END INJ_ROW[18]
  PIN INJ_ROW[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1880.265 187.44 1880.545 188.44 ;
    END
  END INJ_ROW[17]
  PIN INJ_ROW[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1810.265 187.44 1810.545 188.44 ;
    END
  END INJ_ROW[16]
  PIN INJ_ROW[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1731.025 187.44 1731.305 188.44 ;
    END
  END INJ_ROW[15]
  PIN INJ_ROW[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1662.985 187.44 1663.265 188.44 ;
    END
  END INJ_ROW[14]
  PIN INJ_ROW[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1557.145 187.44 1557.425 188.44 ;
    END
  END INJ_ROW[13]
  PIN INJ_ROW[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1475.385 187.44 1475.665 188.44 ;
    END
  END INJ_ROW[12]
  PIN INJ_ROW[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1409.865 187.44 1410.145 188.44 ;
    END
  END INJ_ROW[11]
  PIN INJ_ROW[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1320.265 187.44 1320.545 188.44 ;
    END
  END INJ_ROW[10]
  PIN INJ_ROW[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1250.265 187.44 1250.545 188.44 ;
    END
  END INJ_ROW[9]
  PIN INJ_ROW[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1171.025 187.44 1171.305 188.44 ;
    END
  END INJ_ROW[8]
  PIN INJ_ROW[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1102.985 187.44 1103.265 188.44 ;
    END
  END INJ_ROW[7]
  PIN INJ_ROW[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 997.145 187.44 997.425 188.44 ;
    END
  END INJ_ROW[6]
  PIN INJ_ROW[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 915.385 187.44 915.665 188.44 ;
    END
  END INJ_ROW[5]
  PIN INJ_ROW[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 849.865 187.44 850.145 188.44 ;
    END
  END INJ_ROW[4]
  PIN INJ_ROW[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 760.265 187.44 760.545 188.44 ;
    END
  END INJ_ROW[3]
  PIN INJ_ROW[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 690.265 187.44 690.545 188.44 ;
    END
  END INJ_ROW[2]
  PIN INJ_ROW[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 611.025 187.44 611.305 188.44 ;
    END
  END INJ_ROW[1]
  PIN INJ_ROW[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 542.985 187.44 543.265 188.44 ;
    END
  END INJ_ROW[0]
  PIN MASKH[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18282.665 187.44 18282.945 188.44 ;
    END
  END MASKH[223]
  PIN MASKH[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18217.145 187.44 18217.425 188.44 ;
    END
  END MASKH[222]
  PIN MASKH[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18135.945 187.44 18136.225 188.44 ;
    END
  END MASKH[221]
  PIN MASKH[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18070.425 187.44 18070.705 188.44 ;
    END
  END MASKH[220]
  PIN MASKH[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17980.265 187.44 17980.545 188.44 ;
    END
  END MASKH[219]
  PIN MASKH[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17910.265 187.44 17910.545 188.44 ;
    END
  END MASKH[218]
  PIN MASKH[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17830.465 187.44 17830.745 188.44 ;
    END
  END MASKH[217]
  PIN MASKH[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17722.665 187.44 17722.945 188.44 ;
    END
  END MASKH[216]
  PIN MASKH[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17657.145 187.44 17657.425 188.44 ;
    END
  END MASKH[215]
  PIN MASKH[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17575.945 187.44 17576.225 188.44 ;
    END
  END MASKH[214]
  PIN MASKH[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17510.425 187.44 17510.705 188.44 ;
    END
  END MASKH[213]
  PIN MASKH[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17420.265 187.44 17420.545 188.44 ;
    END
  END MASKH[212]
  PIN MASKH[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17350.265 187.44 17350.545 188.44 ;
    END
  END MASKH[211]
  PIN MASKH[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17270.465 187.44 17270.745 188.44 ;
    END
  END MASKH[210]
  PIN MASKH[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17162.665 187.44 17162.945 188.44 ;
    END
  END MASKH[209]
  PIN MASKH[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17097.145 187.44 17097.425 188.44 ;
    END
  END MASKH[208]
  PIN MASKH[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17015.945 187.44 17016.225 188.44 ;
    END
  END MASKH[207]
  PIN MASKH[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16950.425 187.44 16950.705 188.44 ;
    END
  END MASKH[206]
  PIN MASKH[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16860.265 187.44 16860.545 188.44 ;
    END
  END MASKH[205]
  PIN MASKH[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16790.265 187.44 16790.545 188.44 ;
    END
  END MASKH[204]
  PIN MASKH[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16710.465 187.44 16710.745 188.44 ;
    END
  END MASKH[203]
  PIN MASKH[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16602.665 187.44 16602.945 188.44 ;
    END
  END MASKH[202]
  PIN MASKH[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16537.145 187.44 16537.425 188.44 ;
    END
  END MASKH[201]
  PIN MASKH[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16455.945 187.44 16456.225 188.44 ;
    END
  END MASKH[200]
  PIN MASKH[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16390.425 187.44 16390.705 188.44 ;
    END
  END MASKH[199]
  PIN MASKH[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16300.265 187.44 16300.545 188.44 ;
    END
  END MASKH[198]
  PIN MASKH[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16230.265 187.44 16230.545 188.44 ;
    END
  END MASKH[197]
  PIN MASKH[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16150.465 187.44 16150.745 188.44 ;
    END
  END MASKH[196]
  PIN MASKH[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16042.665 187.44 16042.945 188.44 ;
    END
  END MASKH[195]
  PIN MASKH[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15977.145 187.44 15977.425 188.44 ;
    END
  END MASKH[194]
  PIN MASKH[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15895.945 187.44 15896.225 188.44 ;
    END
  END MASKH[193]
  PIN MASKH[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15830.425 187.44 15830.705 188.44 ;
    END
  END MASKH[192]
  PIN MASKH[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15740.265 187.44 15740.545 188.44 ;
    END
  END MASKH[191]
  PIN MASKH[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15670.265 187.44 15670.545 188.44 ;
    END
  END MASKH[190]
  PIN MASKH[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15590.465 187.44 15590.745 188.44 ;
    END
  END MASKH[189]
  PIN MASKH[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15482.665 187.44 15482.945 188.44 ;
    END
  END MASKH[188]
  PIN MASKH[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15417.145 187.44 15417.425 188.44 ;
    END
  END MASKH[187]
  PIN MASKH[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15335.945 187.44 15336.225 188.44 ;
    END
  END MASKH[186]
  PIN MASKH[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15270.425 187.44 15270.705 188.44 ;
    END
  END MASKH[185]
  PIN MASKH[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15180.265 187.44 15180.545 188.44 ;
    END
  END MASKH[184]
  PIN MASKH[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15110.265 187.44 15110.545 188.44 ;
    END
  END MASKH[183]
  PIN MASKH[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15030.465 187.44 15030.745 188.44 ;
    END
  END MASKH[182]
  PIN MASKH[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14922.665 187.44 14922.945 188.44 ;
    END
  END MASKH[181]
  PIN MASKH[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14857.145 187.44 14857.425 188.44 ;
    END
  END MASKH[180]
  PIN MASKH[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14775.945 187.44 14776.225 188.44 ;
    END
  END MASKH[179]
  PIN MASKH[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14710.425 187.44 14710.705 188.44 ;
    END
  END MASKH[178]
  PIN MASKH[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14620.265 187.44 14620.545 188.44 ;
    END
  END MASKH[177]
  PIN MASKH[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14550.265 187.44 14550.545 188.44 ;
    END
  END MASKH[176]
  PIN MASKH[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14470.465 187.44 14470.745 188.44 ;
    END
  END MASKH[175]
  PIN MASKH[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14362.665 187.44 14362.945 188.44 ;
    END
  END MASKH[174]
  PIN MASKH[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14297.145 187.44 14297.425 188.44 ;
    END
  END MASKH[173]
  PIN MASKH[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14215.945 187.44 14216.225 188.44 ;
    END
  END MASKH[172]
  PIN MASKH[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14150.425 187.44 14150.705 188.44 ;
    END
  END MASKH[171]
  PIN MASKH[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14060.265 187.44 14060.545 188.44 ;
    END
  END MASKH[170]
  PIN MASKH[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13990.265 187.44 13990.545 188.44 ;
    END
  END MASKH[169]
  PIN MASKH[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13910.465 187.44 13910.745 188.44 ;
    END
  END MASKH[168]
  PIN MASKH[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13802.665 187.44 13802.945 188.44 ;
    END
  END MASKH[167]
  PIN MASKH[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13737.145 187.44 13737.425 188.44 ;
    END
  END MASKH[166]
  PIN MASKH[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13655.945 187.44 13656.225 188.44 ;
    END
  END MASKH[165]
  PIN MASKH[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13590.425 187.44 13590.705 188.44 ;
    END
  END MASKH[164]
  PIN MASKH[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13500.265 187.44 13500.545 188.44 ;
    END
  END MASKH[163]
  PIN MASKH[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13430.265 187.44 13430.545 188.44 ;
    END
  END MASKH[162]
  PIN MASKH[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13350.465 187.44 13350.745 188.44 ;
    END
  END MASKH[161]
  PIN MASKH[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13242.665 187.44 13242.945 188.44 ;
    END
  END MASKH[160]
  PIN MASKH[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13177.145 187.44 13177.425 188.44 ;
    END
  END MASKH[159]
  PIN MASKH[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13095.945 187.44 13096.225 188.44 ;
    END
  END MASKH[158]
  PIN MASKH[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13030.425 187.44 13030.705 188.44 ;
    END
  END MASKH[157]
  PIN MASKH[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12940.265 187.44 12940.545 188.44 ;
    END
  END MASKH[156]
  PIN MASKH[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12870.265 187.44 12870.545 188.44 ;
    END
  END MASKH[155]
  PIN MASKH[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12790.465 187.44 12790.745 188.44 ;
    END
  END MASKH[154]
  PIN MASKH[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12682.665 187.44 12682.945 188.44 ;
    END
  END MASKH[153]
  PIN MASKH[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12617.145 187.44 12617.425 188.44 ;
    END
  END MASKH[152]
  PIN MASKH[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12535.945 187.44 12536.225 188.44 ;
    END
  END MASKH[151]
  PIN MASKH[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12470.425 187.44 12470.705 188.44 ;
    END
  END MASKH[150]
  PIN MASKH[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12380.265 187.44 12380.545 188.44 ;
    END
  END MASKH[149]
  PIN MASKH[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12310.265 187.44 12310.545 188.44 ;
    END
  END MASKH[148]
  PIN MASKH[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12230.465 187.44 12230.745 188.44 ;
    END
  END MASKH[147]
  PIN MASKH[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12122.665 187.44 12122.945 188.44 ;
    END
  END MASKH[146]
  PIN MASKH[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12057.145 187.44 12057.425 188.44 ;
    END
  END MASKH[145]
  PIN MASKH[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11975.945 187.44 11976.225 188.44 ;
    END
  END MASKH[144]
  PIN MASKH[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11910.425 187.44 11910.705 188.44 ;
    END
  END MASKH[143]
  PIN MASKH[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11820.265 187.44 11820.545 188.44 ;
    END
  END MASKH[142]
  PIN MASKH[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11750.265 187.44 11750.545 188.44 ;
    END
  END MASKH[141]
  PIN MASKH[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11670.465 187.44 11670.745 188.44 ;
    END
  END MASKH[140]
  PIN MASKH[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11562.665 187.44 11562.945 188.44 ;
    END
  END MASKH[139]
  PIN MASKH[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11497.145 187.44 11497.425 188.44 ;
    END
  END MASKH[138]
  PIN MASKH[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11415.945 187.44 11416.225 188.44 ;
    END
  END MASKH[137]
  PIN MASKH[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11350.425 187.44 11350.705 188.44 ;
    END
  END MASKH[136]
  PIN MASKH[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11260.265 187.44 11260.545 188.44 ;
    END
  END MASKH[135]
  PIN MASKH[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11190.265 187.44 11190.545 188.44 ;
    END
  END MASKH[134]
  PIN MASKH[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11110.465 187.44 11110.745 188.44 ;
    END
  END MASKH[133]
  PIN MASKH[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11002.665 187.44 11002.945 188.44 ;
    END
  END MASKH[132]
  PIN MASKH[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10937.145 187.44 10937.425 188.44 ;
    END
  END MASKH[131]
  PIN MASKH[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10855.945 187.44 10856.225 188.44 ;
    END
  END MASKH[130]
  PIN MASKH[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10790.425 187.44 10790.705 188.44 ;
    END
  END MASKH[129]
  PIN MASKH[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10700.265 187.44 10700.545 188.44 ;
    END
  END MASKH[128]
  PIN MASKH[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10630.265 187.44 10630.545 188.44 ;
    END
  END MASKH[127]
  PIN MASKH[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10550.465 187.44 10550.745 188.44 ;
    END
  END MASKH[126]
  PIN MASKH[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10442.665 187.44 10442.945 188.44 ;
    END
  END MASKH[125]
  PIN MASKH[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10377.145 187.44 10377.425 188.44 ;
    END
  END MASKH[124]
  PIN MASKH[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10295.945 187.44 10296.225 188.44 ;
    END
  END MASKH[123]
  PIN MASKH[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10230.425 187.44 10230.705 188.44 ;
    END
  END MASKH[122]
  PIN MASKH[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10140.265 187.44 10140.545 188.44 ;
    END
  END MASKH[121]
  PIN MASKH[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10070.265 187.44 10070.545 188.44 ;
    END
  END MASKH[120]
  PIN MASKH[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9990.465 187.44 9990.745 188.44 ;
    END
  END MASKH[119]
  PIN MASKH[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9882.665 187.44 9882.945 188.44 ;
    END
  END MASKH[118]
  PIN MASKH[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9817.145 187.44 9817.425 188.44 ;
    END
  END MASKH[117]
  PIN MASKH[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9735.945 187.44 9736.225 188.44 ;
    END
  END MASKH[116]
  PIN MASKH[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9670.425 187.44 9670.705 188.44 ;
    END
  END MASKH[115]
  PIN MASKH[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9580.265 187.44 9580.545 188.44 ;
    END
  END MASKH[114]
  PIN MASKH[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9510.265 187.44 9510.545 188.44 ;
    END
  END MASKH[113]
  PIN MASKH[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9430.465 187.44 9430.745 188.44 ;
    END
  END MASKH[112]
  PIN MASKH[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9322.665 187.44 9322.945 188.44 ;
    END
  END MASKH[111]
  PIN MASKH[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9257.145 187.44 9257.425 188.44 ;
    END
  END MASKH[110]
  PIN MASKH[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9175.945 187.44 9176.225 188.44 ;
    END
  END MASKH[109]
  PIN MASKH[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9110.425 187.44 9110.705 188.44 ;
    END
  END MASKH[108]
  PIN MASKH[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9020.265 187.44 9020.545 188.44 ;
    END
  END MASKH[107]
  PIN MASKH[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8950.265 187.44 8950.545 188.44 ;
    END
  END MASKH[106]
  PIN MASKH[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8870.465 187.44 8870.745 188.44 ;
    END
  END MASKH[105]
  PIN MASKH[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8762.665 187.44 8762.945 188.44 ;
    END
  END MASKH[104]
  PIN MASKH[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8697.145 187.44 8697.425 188.44 ;
    END
  END MASKH[103]
  PIN MASKH[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8615.945 187.44 8616.225 188.44 ;
    END
  END MASKH[102]
  PIN MASKH[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8550.425 187.44 8550.705 188.44 ;
    END
  END MASKH[101]
  PIN MASKH[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8460.265 187.44 8460.545 188.44 ;
    END
  END MASKH[100]
  PIN MASKH[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8390.265 187.44 8390.545 188.44 ;
    END
  END MASKH[99]
  PIN MASKH[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8310.465 187.44 8310.745 188.44 ;
    END
  END MASKH[98]
  PIN MASKH[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8202.665 187.44 8202.945 188.44 ;
    END
  END MASKH[97]
  PIN MASKH[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8137.145 187.44 8137.425 188.44 ;
    END
  END MASKH[96]
  PIN MASKH[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8055.945 187.44 8056.225 188.44 ;
    END
  END MASKH[95]
  PIN MASKH[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7990.425 187.44 7990.705 188.44 ;
    END
  END MASKH[94]
  PIN MASKH[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7900.265 187.44 7900.545 188.44 ;
    END
  END MASKH[93]
  PIN MASKH[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7830.265 187.44 7830.545 188.44 ;
    END
  END MASKH[92]
  PIN MASKH[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7750.465 187.44 7750.745 188.44 ;
    END
  END MASKH[91]
  PIN MASKH[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7642.665 187.44 7642.945 188.44 ;
    END
  END MASKH[90]
  PIN MASKH[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7577.145 187.44 7577.425 188.44 ;
    END
  END MASKH[89]
  PIN MASKH[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7495.945 187.44 7496.225 188.44 ;
    END
  END MASKH[88]
  PIN MASKH[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7430.425 187.44 7430.705 188.44 ;
    END
  END MASKH[87]
  PIN MASKH[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7340.265 187.44 7340.545 188.44 ;
    END
  END MASKH[86]
  PIN MASKH[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7270.265 187.44 7270.545 188.44 ;
    END
  END MASKH[85]
  PIN MASKH[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7190.465 187.44 7190.745 188.44 ;
    END
  END MASKH[84]
  PIN MASKH[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7082.665 187.44 7082.945 188.44 ;
    END
  END MASKH[83]
  PIN MASKH[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7017.145 187.44 7017.425 188.44 ;
    END
  END MASKH[82]
  PIN MASKH[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6935.945 187.44 6936.225 188.44 ;
    END
  END MASKH[81]
  PIN MASKH[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6870.425 187.44 6870.705 188.44 ;
    END
  END MASKH[80]
  PIN MASKH[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6780.265 187.44 6780.545 188.44 ;
    END
  END MASKH[79]
  PIN MASKH[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6710.265 187.44 6710.545 188.44 ;
    END
  END MASKH[78]
  PIN MASKH[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6630.465 187.44 6630.745 188.44 ;
    END
  END MASKH[77]
  PIN MASKH[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6522.665 187.44 6522.945 188.44 ;
    END
  END MASKH[76]
  PIN MASKH[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6457.145 187.44 6457.425 188.44 ;
    END
  END MASKH[75]
  PIN MASKH[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6375.945 187.44 6376.225 188.44 ;
    END
  END MASKH[74]
  PIN MASKH[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6310.425 187.44 6310.705 188.44 ;
    END
  END MASKH[73]
  PIN MASKH[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6220.265 187.44 6220.545 188.44 ;
    END
  END MASKH[72]
  PIN MASKH[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6150.265 187.44 6150.545 188.44 ;
    END
  END MASKH[71]
  PIN MASKH[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6070.465 187.44 6070.745 188.44 ;
    END
  END MASKH[70]
  PIN MASKH[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5962.665 187.44 5962.945 188.44 ;
    END
  END MASKH[69]
  PIN MASKH[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5897.145 187.44 5897.425 188.44 ;
    END
  END MASKH[68]
  PIN MASKH[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5815.945 187.44 5816.225 188.44 ;
    END
  END MASKH[67]
  PIN MASKH[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5750.425 187.44 5750.705 188.44 ;
    END
  END MASKH[66]
  PIN MASKH[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5660.265 187.44 5660.545 188.44 ;
    END
  END MASKH[65]
  PIN MASKH[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5590.265 187.44 5590.545 188.44 ;
    END
  END MASKH[64]
  PIN MASKH[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5510.465 187.44 5510.745 188.44 ;
    END
  END MASKH[63]
  PIN MASKH[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5402.665 187.44 5402.945 188.44 ;
    END
  END MASKH[62]
  PIN MASKH[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5337.145 187.44 5337.425 188.44 ;
    END
  END MASKH[61]
  PIN MASKH[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5255.945 187.44 5256.225 188.44 ;
    END
  END MASKH[60]
  PIN MASKH[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5190.425 187.44 5190.705 188.44 ;
    END
  END MASKH[59]
  PIN MASKH[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5100.265 187.44 5100.545 188.44 ;
    END
  END MASKH[58]
  PIN MASKH[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5030.265 187.44 5030.545 188.44 ;
    END
  END MASKH[57]
  PIN MASKH[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4950.465 187.44 4950.745 188.44 ;
    END
  END MASKH[56]
  PIN MASKH[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4842.665 187.44 4842.945 188.44 ;
    END
  END MASKH[55]
  PIN MASKH[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4777.145 187.44 4777.425 188.44 ;
    END
  END MASKH[54]
  PIN MASKH[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4695.945 187.44 4696.225 188.44 ;
    END
  END MASKH[53]
  PIN MASKH[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4630.425 187.44 4630.705 188.44 ;
    END
  END MASKH[52]
  PIN MASKH[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4540.265 187.44 4540.545 188.44 ;
    END
  END MASKH[51]
  PIN MASKH[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4470.265 187.44 4470.545 188.44 ;
    END
  END MASKH[50]
  PIN MASKH[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4390.465 187.44 4390.745 188.44 ;
    END
  END MASKH[49]
  PIN MASKH[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4282.665 187.44 4282.945 188.44 ;
    END
  END MASKH[48]
  PIN MASKH[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4217.145 187.44 4217.425 188.44 ;
    END
  END MASKH[47]
  PIN MASKH[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4135.945 187.44 4136.225 188.44 ;
    END
  END MASKH[46]
  PIN MASKH[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4070.425 187.44 4070.705 188.44 ;
    END
  END MASKH[45]
  PIN MASKH[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3980.265 187.44 3980.545 188.44 ;
    END
  END MASKH[44]
  PIN MASKH[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3910.265 187.44 3910.545 188.44 ;
    END
  END MASKH[43]
  PIN MASKH[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3830.465 187.44 3830.745 188.44 ;
    END
  END MASKH[42]
  PIN MASKH[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3722.665 187.44 3722.945 188.44 ;
    END
  END MASKH[41]
  PIN MASKH[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3657.145 187.44 3657.425 188.44 ;
    END
  END MASKH[40]
  PIN MASKH[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3575.945 187.44 3576.225 188.44 ;
    END
  END MASKH[39]
  PIN MASKH[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3510.425 187.44 3510.705 188.44 ;
    END
  END MASKH[38]
  PIN MASKH[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3420.265 187.44 3420.545 188.44 ;
    END
  END MASKH[37]
  PIN MASKH[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3350.265 187.44 3350.545 188.44 ;
    END
  END MASKH[36]
  PIN MASKH[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3270.465 187.44 3270.745 188.44 ;
    END
  END MASKH[35]
  PIN MASKH[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3162.665 187.44 3162.945 188.44 ;
    END
  END MASKH[34]
  PIN MASKH[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3097.145 187.44 3097.425 188.44 ;
    END
  END MASKH[33]
  PIN MASKH[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3015.945 187.44 3016.225 188.44 ;
    END
  END MASKH[32]
  PIN MASKH[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2950.425 187.44 2950.705 188.44 ;
    END
  END MASKH[31]
  PIN MASKH[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2860.265 187.44 2860.545 188.44 ;
    END
  END MASKH[30]
  PIN MASKH[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2790.265 187.44 2790.545 188.44 ;
    END
  END MASKH[29]
  PIN MASKH[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2710.465 187.44 2710.745 188.44 ;
    END
  END MASKH[28]
  PIN MASKH[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2602.665 187.44 2602.945 188.44 ;
    END
  END MASKH[27]
  PIN MASKH[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2537.145 187.44 2537.425 188.44 ;
    END
  END MASKH[26]
  PIN MASKH[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2455.945 187.44 2456.225 188.44 ;
    END
  END MASKH[25]
  PIN MASKH[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2390.425 187.44 2390.705 188.44 ;
    END
  END MASKH[24]
  PIN MASKH[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2300.265 187.44 2300.545 188.44 ;
    END
  END MASKH[23]
  PIN MASKH[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2230.265 187.44 2230.545 188.44 ;
    END
  END MASKH[22]
  PIN MASKH[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2150.465 187.44 2150.745 188.44 ;
    END
  END MASKH[21]
  PIN MASKH[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2042.665 187.44 2042.945 188.44 ;
    END
  END MASKH[20]
  PIN MASKH[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1977.145 187.44 1977.425 188.44 ;
    END
  END MASKH[19]
  PIN MASKH[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1895.945 187.44 1896.225 188.44 ;
    END
  END MASKH[18]
  PIN MASKH[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1830.425 187.44 1830.705 188.44 ;
    END
  END MASKH[17]
  PIN MASKH[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1740.265 187.44 1740.545 188.44 ;
    END
  END MASKH[16]
  PIN MASKH[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1670.265 187.44 1670.545 188.44 ;
    END
  END MASKH[15]
  PIN MASKH[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1590.465 187.44 1590.745 188.44 ;
    END
  END MASKH[14]
  PIN MASKH[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1482.665 187.44 1482.945 188.44 ;
    END
  END MASKH[13]
  PIN MASKH[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1417.145 187.44 1417.425 188.44 ;
    END
  END MASKH[12]
  PIN MASKH[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1335.945 187.44 1336.225 188.44 ;
    END
  END MASKH[11]
  PIN MASKH[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1270.425 187.44 1270.705 188.44 ;
    END
  END MASKH[10]
  PIN MASKH[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1180.265 187.44 1180.545 188.44 ;
    END
  END MASKH[9]
  PIN MASKH[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1110.265 187.44 1110.545 188.44 ;
    END
  END MASKH[8]
  PIN MASKH[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1030.465 187.44 1030.745 188.44 ;
    END
  END MASKH[7]
  PIN MASKH[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 922.665 187.44 922.945 188.44 ;
    END
  END MASKH[6]
  PIN MASKH[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 857.145 187.44 857.425 188.44 ;
    END
  END MASKH[5]
  PIN MASKH[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 775.945 187.44 776.225 188.44 ;
    END
  END MASKH[4]
  PIN MASKH[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 710.425 187.44 710.705 188.44 ;
    END
  END MASKH[3]
  PIN MASKH[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 620.265 187.44 620.545 188.44 ;
    END
  END MASKH[2]
  PIN MASKH[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 550.265 187.44 550.545 188.44 ;
    END
  END MASKH[1]
  PIN MASKH[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 470.465 187.44 470.745 188.44 ;
    END
  END MASKH[0]
  PIN MASKD[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18359.385 187.44 18359.665 188.44 ;
    END
  END MASKD[447]
  PIN MASKD[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18282.105 187.44 18282.385 188.44 ;
    END
  END MASKD[446]
  PIN MASKD[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18277.625 187.44 18277.905 188.44 ;
    END
  END MASKD[445]
  PIN MASKD[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18216.585 187.44 18216.865 188.44 ;
    END
  END MASKD[444]
  PIN MASKD[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18212.105 187.44 18212.385 188.44 ;
    END
  END MASKD[443]
  PIN MASKD[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18135.385 187.44 18135.665 188.44 ;
    END
  END MASKD[442]
  PIN MASKD[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18130.905 187.44 18131.185 188.44 ;
    END
  END MASKD[441]
  PIN MASKD[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18069.865 187.44 18070.145 188.44 ;
    END
  END MASKD[440]
  PIN MASKD[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18052.505 187.44 18052.785 188.44 ;
    END
  END MASKD[439]
  PIN MASKD[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17979.705 187.44 17979.985 188.44 ;
    END
  END MASKD[438]
  PIN MASKD[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17975.225 187.44 17975.505 188.44 ;
    END
  END MASKD[437]
  PIN MASKD[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17909.705 187.44 17909.985 188.44 ;
    END
  END MASKD[436]
  PIN MASKD[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17905.225 187.44 17905.505 188.44 ;
    END
  END MASKD[435]
  PIN MASKD[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17829.905 187.44 17830.185 188.44 ;
    END
  END MASKD[434]
  PIN MASKD[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17799.385 187.44 17799.665 188.44 ;
    END
  END MASKD[433]
  PIN MASKD[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17722.105 187.44 17722.385 188.44 ;
    END
  END MASKD[432]
  PIN MASKD[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17717.625 187.44 17717.905 188.44 ;
    END
  END MASKD[431]
  PIN MASKD[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17656.585 187.44 17656.865 188.44 ;
    END
  END MASKD[430]
  PIN MASKD[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17652.105 187.44 17652.385 188.44 ;
    END
  END MASKD[429]
  PIN MASKD[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17575.385 187.44 17575.665 188.44 ;
    END
  END MASKD[428]
  PIN MASKD[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17570.905 187.44 17571.185 188.44 ;
    END
  END MASKD[427]
  PIN MASKD[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17509.865 187.44 17510.145 188.44 ;
    END
  END MASKD[426]
  PIN MASKD[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17492.505 187.44 17492.785 188.44 ;
    END
  END MASKD[425]
  PIN MASKD[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17419.705 187.44 17419.985 188.44 ;
    END
  END MASKD[424]
  PIN MASKD[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17415.225 187.44 17415.505 188.44 ;
    END
  END MASKD[423]
  PIN MASKD[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17349.705 187.44 17349.985 188.44 ;
    END
  END MASKD[422]
  PIN MASKD[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17345.225 187.44 17345.505 188.44 ;
    END
  END MASKD[421]
  PIN MASKD[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17269.905 187.44 17270.185 188.44 ;
    END
  END MASKD[420]
  PIN MASKD[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17239.385 187.44 17239.665 188.44 ;
    END
  END MASKD[419]
  PIN MASKD[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17162.105 187.44 17162.385 188.44 ;
    END
  END MASKD[418]
  PIN MASKD[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17157.625 187.44 17157.905 188.44 ;
    END
  END MASKD[417]
  PIN MASKD[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17096.585 187.44 17096.865 188.44 ;
    END
  END MASKD[416]
  PIN MASKD[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17092.105 187.44 17092.385 188.44 ;
    END
  END MASKD[415]
  PIN MASKD[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17015.385 187.44 17015.665 188.44 ;
    END
  END MASKD[414]
  PIN MASKD[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17010.905 187.44 17011.185 188.44 ;
    END
  END MASKD[413]
  PIN MASKD[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16949.865 187.44 16950.145 188.44 ;
    END
  END MASKD[412]
  PIN MASKD[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16932.505 187.44 16932.785 188.44 ;
    END
  END MASKD[411]
  PIN MASKD[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16859.705 187.44 16859.985 188.44 ;
    END
  END MASKD[410]
  PIN MASKD[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16855.225 187.44 16855.505 188.44 ;
    END
  END MASKD[409]
  PIN MASKD[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16789.705 187.44 16789.985 188.44 ;
    END
  END MASKD[408]
  PIN MASKD[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16785.225 187.44 16785.505 188.44 ;
    END
  END MASKD[407]
  PIN MASKD[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16709.905 187.44 16710.185 188.44 ;
    END
  END MASKD[406]
  PIN MASKD[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16679.385 187.44 16679.665 188.44 ;
    END
  END MASKD[405]
  PIN MASKD[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16602.105 187.44 16602.385 188.44 ;
    END
  END MASKD[404]
  PIN MASKD[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16597.625 187.44 16597.905 188.44 ;
    END
  END MASKD[403]
  PIN MASKD[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16536.585 187.44 16536.865 188.44 ;
    END
  END MASKD[402]
  PIN MASKD[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16532.105 187.44 16532.385 188.44 ;
    END
  END MASKD[401]
  PIN MASKD[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16455.385 187.44 16455.665 188.44 ;
    END
  END MASKD[400]
  PIN MASKD[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16450.905 187.44 16451.185 188.44 ;
    END
  END MASKD[399]
  PIN MASKD[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16389.865 187.44 16390.145 188.44 ;
    END
  END MASKD[398]
  PIN MASKD[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16372.505 187.44 16372.785 188.44 ;
    END
  END MASKD[397]
  PIN MASKD[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16299.705 187.44 16299.985 188.44 ;
    END
  END MASKD[396]
  PIN MASKD[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16295.225 187.44 16295.505 188.44 ;
    END
  END MASKD[395]
  PIN MASKD[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16229.705 187.44 16229.985 188.44 ;
    END
  END MASKD[394]
  PIN MASKD[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16225.225 187.44 16225.505 188.44 ;
    END
  END MASKD[393]
  PIN MASKD[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16149.905 187.44 16150.185 188.44 ;
    END
  END MASKD[392]
  PIN MASKD[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16119.385 187.44 16119.665 188.44 ;
    END
  END MASKD[391]
  PIN MASKD[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16042.105 187.44 16042.385 188.44 ;
    END
  END MASKD[390]
  PIN MASKD[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16037.625 187.44 16037.905 188.44 ;
    END
  END MASKD[389]
  PIN MASKD[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15976.585 187.44 15976.865 188.44 ;
    END
  END MASKD[388]
  PIN MASKD[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15972.105 187.44 15972.385 188.44 ;
    END
  END MASKD[387]
  PIN MASKD[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15895.385 187.44 15895.665 188.44 ;
    END
  END MASKD[386]
  PIN MASKD[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15890.905 187.44 15891.185 188.44 ;
    END
  END MASKD[385]
  PIN MASKD[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15829.865 187.44 15830.145 188.44 ;
    END
  END MASKD[384]
  PIN MASKD[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15812.505 187.44 15812.785 188.44 ;
    END
  END MASKD[383]
  PIN MASKD[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15739.705 187.44 15739.985 188.44 ;
    END
  END MASKD[382]
  PIN MASKD[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15735.225 187.44 15735.505 188.44 ;
    END
  END MASKD[381]
  PIN MASKD[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15669.705 187.44 15669.985 188.44 ;
    END
  END MASKD[380]
  PIN MASKD[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15665.225 187.44 15665.505 188.44 ;
    END
  END MASKD[379]
  PIN MASKD[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15589.905 187.44 15590.185 188.44 ;
    END
  END MASKD[378]
  PIN MASKD[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15559.385 187.44 15559.665 188.44 ;
    END
  END MASKD[377]
  PIN MASKD[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15482.105 187.44 15482.385 188.44 ;
    END
  END MASKD[376]
  PIN MASKD[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15477.625 187.44 15477.905 188.44 ;
    END
  END MASKD[375]
  PIN MASKD[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15416.585 187.44 15416.865 188.44 ;
    END
  END MASKD[374]
  PIN MASKD[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15412.105 187.44 15412.385 188.44 ;
    END
  END MASKD[373]
  PIN MASKD[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15335.385 187.44 15335.665 188.44 ;
    END
  END MASKD[372]
  PIN MASKD[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15330.905 187.44 15331.185 188.44 ;
    END
  END MASKD[371]
  PIN MASKD[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15269.865 187.44 15270.145 188.44 ;
    END
  END MASKD[370]
  PIN MASKD[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15252.505 187.44 15252.785 188.44 ;
    END
  END MASKD[369]
  PIN MASKD[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15179.705 187.44 15179.985 188.44 ;
    END
  END MASKD[368]
  PIN MASKD[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15175.225 187.44 15175.505 188.44 ;
    END
  END MASKD[367]
  PIN MASKD[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15109.705 187.44 15109.985 188.44 ;
    END
  END MASKD[366]
  PIN MASKD[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15105.225 187.44 15105.505 188.44 ;
    END
  END MASKD[365]
  PIN MASKD[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15029.905 187.44 15030.185 188.44 ;
    END
  END MASKD[364]
  PIN MASKD[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14999.385 187.44 14999.665 188.44 ;
    END
  END MASKD[363]
  PIN MASKD[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14922.105 187.44 14922.385 188.44 ;
    END
  END MASKD[362]
  PIN MASKD[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14917.625 187.44 14917.905 188.44 ;
    END
  END MASKD[361]
  PIN MASKD[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14856.585 187.44 14856.865 188.44 ;
    END
  END MASKD[360]
  PIN MASKD[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14852.105 187.44 14852.385 188.44 ;
    END
  END MASKD[359]
  PIN MASKD[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14775.385 187.44 14775.665 188.44 ;
    END
  END MASKD[358]
  PIN MASKD[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14770.905 187.44 14771.185 188.44 ;
    END
  END MASKD[357]
  PIN MASKD[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14709.865 187.44 14710.145 188.44 ;
    END
  END MASKD[356]
  PIN MASKD[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14692.505 187.44 14692.785 188.44 ;
    END
  END MASKD[355]
  PIN MASKD[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14619.705 187.44 14619.985 188.44 ;
    END
  END MASKD[354]
  PIN MASKD[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14615.225 187.44 14615.505 188.44 ;
    END
  END MASKD[353]
  PIN MASKD[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14549.705 187.44 14549.985 188.44 ;
    END
  END MASKD[352]
  PIN MASKD[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14545.225 187.44 14545.505 188.44 ;
    END
  END MASKD[351]
  PIN MASKD[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14469.905 187.44 14470.185 188.44 ;
    END
  END MASKD[350]
  PIN MASKD[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14439.385 187.44 14439.665 188.44 ;
    END
  END MASKD[349]
  PIN MASKD[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14362.105 187.44 14362.385 188.44 ;
    END
  END MASKD[348]
  PIN MASKD[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14357.625 187.44 14357.905 188.44 ;
    END
  END MASKD[347]
  PIN MASKD[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14296.585 187.44 14296.865 188.44 ;
    END
  END MASKD[346]
  PIN MASKD[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14292.105 187.44 14292.385 188.44 ;
    END
  END MASKD[345]
  PIN MASKD[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14215.385 187.44 14215.665 188.44 ;
    END
  END MASKD[344]
  PIN MASKD[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14210.905 187.44 14211.185 188.44 ;
    END
  END MASKD[343]
  PIN MASKD[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14149.865 187.44 14150.145 188.44 ;
    END
  END MASKD[342]
  PIN MASKD[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14132.505 187.44 14132.785 188.44 ;
    END
  END MASKD[341]
  PIN MASKD[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14059.705 187.44 14059.985 188.44 ;
    END
  END MASKD[340]
  PIN MASKD[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14055.225 187.44 14055.505 188.44 ;
    END
  END MASKD[339]
  PIN MASKD[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13989.705 187.44 13989.985 188.44 ;
    END
  END MASKD[338]
  PIN MASKD[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13985.225 187.44 13985.505 188.44 ;
    END
  END MASKD[337]
  PIN MASKD[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13909.905 187.44 13910.185 188.44 ;
    END
  END MASKD[336]
  PIN MASKD[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13879.385 187.44 13879.665 188.44 ;
    END
  END MASKD[335]
  PIN MASKD[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13802.105 187.44 13802.385 188.44 ;
    END
  END MASKD[334]
  PIN MASKD[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13797.625 187.44 13797.905 188.44 ;
    END
  END MASKD[333]
  PIN MASKD[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13736.585 187.44 13736.865 188.44 ;
    END
  END MASKD[332]
  PIN MASKD[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13732.105 187.44 13732.385 188.44 ;
    END
  END MASKD[331]
  PIN MASKD[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13655.385 187.44 13655.665 188.44 ;
    END
  END MASKD[330]
  PIN MASKD[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13650.905 187.44 13651.185 188.44 ;
    END
  END MASKD[329]
  PIN MASKD[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13589.865 187.44 13590.145 188.44 ;
    END
  END MASKD[328]
  PIN MASKD[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13572.505 187.44 13572.785 188.44 ;
    END
  END MASKD[327]
  PIN MASKD[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13499.705 187.44 13499.985 188.44 ;
    END
  END MASKD[326]
  PIN MASKD[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13495.225 187.44 13495.505 188.44 ;
    END
  END MASKD[325]
  PIN MASKD[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13429.705 187.44 13429.985 188.44 ;
    END
  END MASKD[324]
  PIN MASKD[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13425.225 187.44 13425.505 188.44 ;
    END
  END MASKD[323]
  PIN MASKD[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13349.905 187.44 13350.185 188.44 ;
    END
  END MASKD[322]
  PIN MASKD[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13319.385 187.44 13319.665 188.44 ;
    END
  END MASKD[321]
  PIN MASKD[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13242.105 187.44 13242.385 188.44 ;
    END
  END MASKD[320]
  PIN MASKD[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13237.625 187.44 13237.905 188.44 ;
    END
  END MASKD[319]
  PIN MASKD[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13176.585 187.44 13176.865 188.44 ;
    END
  END MASKD[318]
  PIN MASKD[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13172.105 187.44 13172.385 188.44 ;
    END
  END MASKD[317]
  PIN MASKD[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13095.385 187.44 13095.665 188.44 ;
    END
  END MASKD[316]
  PIN MASKD[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13090.905 187.44 13091.185 188.44 ;
    END
  END MASKD[315]
  PIN MASKD[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13029.865 187.44 13030.145 188.44 ;
    END
  END MASKD[314]
  PIN MASKD[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13012.505 187.44 13012.785 188.44 ;
    END
  END MASKD[313]
  PIN MASKD[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12939.705 187.44 12939.985 188.44 ;
    END
  END MASKD[312]
  PIN MASKD[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12935.225 187.44 12935.505 188.44 ;
    END
  END MASKD[311]
  PIN MASKD[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12869.705 187.44 12869.985 188.44 ;
    END
  END MASKD[310]
  PIN MASKD[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12865.225 187.44 12865.505 188.44 ;
    END
  END MASKD[309]
  PIN MASKD[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12789.905 187.44 12790.185 188.44 ;
    END
  END MASKD[308]
  PIN MASKD[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12759.385 187.44 12759.665 188.44 ;
    END
  END MASKD[307]
  PIN MASKD[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12682.105 187.44 12682.385 188.44 ;
    END
  END MASKD[306]
  PIN MASKD[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12677.625 187.44 12677.905 188.44 ;
    END
  END MASKD[305]
  PIN MASKD[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12616.585 187.44 12616.865 188.44 ;
    END
  END MASKD[304]
  PIN MASKD[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12612.105 187.44 12612.385 188.44 ;
    END
  END MASKD[303]
  PIN MASKD[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12535.385 187.44 12535.665 188.44 ;
    END
  END MASKD[302]
  PIN MASKD[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12530.905 187.44 12531.185 188.44 ;
    END
  END MASKD[301]
  PIN MASKD[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12469.865 187.44 12470.145 188.44 ;
    END
  END MASKD[300]
  PIN MASKD[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12452.505 187.44 12452.785 188.44 ;
    END
  END MASKD[299]
  PIN MASKD[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12379.705 187.44 12379.985 188.44 ;
    END
  END MASKD[298]
  PIN MASKD[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12375.225 187.44 12375.505 188.44 ;
    END
  END MASKD[297]
  PIN MASKD[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12309.705 187.44 12309.985 188.44 ;
    END
  END MASKD[296]
  PIN MASKD[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12305.225 187.44 12305.505 188.44 ;
    END
  END MASKD[295]
  PIN MASKD[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12229.905 187.44 12230.185 188.44 ;
    END
  END MASKD[294]
  PIN MASKD[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12199.385 187.44 12199.665 188.44 ;
    END
  END MASKD[293]
  PIN MASKD[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12122.105 187.44 12122.385 188.44 ;
    END
  END MASKD[292]
  PIN MASKD[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12117.625 187.44 12117.905 188.44 ;
    END
  END MASKD[291]
  PIN MASKD[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12056.585 187.44 12056.865 188.44 ;
    END
  END MASKD[290]
  PIN MASKD[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12052.105 187.44 12052.385 188.44 ;
    END
  END MASKD[289]
  PIN MASKD[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11975.385 187.44 11975.665 188.44 ;
    END
  END MASKD[288]
  PIN MASKD[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11970.905 187.44 11971.185 188.44 ;
    END
  END MASKD[287]
  PIN MASKD[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11909.865 187.44 11910.145 188.44 ;
    END
  END MASKD[286]
  PIN MASKD[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11892.505 187.44 11892.785 188.44 ;
    END
  END MASKD[285]
  PIN MASKD[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11819.705 187.44 11819.985 188.44 ;
    END
  END MASKD[284]
  PIN MASKD[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11815.225 187.44 11815.505 188.44 ;
    END
  END MASKD[283]
  PIN MASKD[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11749.705 187.44 11749.985 188.44 ;
    END
  END MASKD[282]
  PIN MASKD[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11745.225 187.44 11745.505 188.44 ;
    END
  END MASKD[281]
  PIN MASKD[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11669.905 187.44 11670.185 188.44 ;
    END
  END MASKD[280]
  PIN MASKD[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11639.385 187.44 11639.665 188.44 ;
    END
  END MASKD[279]
  PIN MASKD[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11562.105 187.44 11562.385 188.44 ;
    END
  END MASKD[278]
  PIN MASKD[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11557.625 187.44 11557.905 188.44 ;
    END
  END MASKD[277]
  PIN MASKD[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11496.585 187.44 11496.865 188.44 ;
    END
  END MASKD[276]
  PIN MASKD[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11492.105 187.44 11492.385 188.44 ;
    END
  END MASKD[275]
  PIN MASKD[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11415.385 187.44 11415.665 188.44 ;
    END
  END MASKD[274]
  PIN MASKD[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11410.905 187.44 11411.185 188.44 ;
    END
  END MASKD[273]
  PIN MASKD[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11349.865 187.44 11350.145 188.44 ;
    END
  END MASKD[272]
  PIN MASKD[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11332.505 187.44 11332.785 188.44 ;
    END
  END MASKD[271]
  PIN MASKD[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11259.705 187.44 11259.985 188.44 ;
    END
  END MASKD[270]
  PIN MASKD[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11255.225 187.44 11255.505 188.44 ;
    END
  END MASKD[269]
  PIN MASKD[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11189.705 187.44 11189.985 188.44 ;
    END
  END MASKD[268]
  PIN MASKD[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11185.225 187.44 11185.505 188.44 ;
    END
  END MASKD[267]
  PIN MASKD[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11109.905 187.44 11110.185 188.44 ;
    END
  END MASKD[266]
  PIN MASKD[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11079.385 187.44 11079.665 188.44 ;
    END
  END MASKD[265]
  PIN MASKD[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11002.105 187.44 11002.385 188.44 ;
    END
  END MASKD[264]
  PIN MASKD[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10997.625 187.44 10997.905 188.44 ;
    END
  END MASKD[263]
  PIN MASKD[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10936.585 187.44 10936.865 188.44 ;
    END
  END MASKD[262]
  PIN MASKD[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10932.105 187.44 10932.385 188.44 ;
    END
  END MASKD[261]
  PIN MASKD[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10855.385 187.44 10855.665 188.44 ;
    END
  END MASKD[260]
  PIN MASKD[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10850.905 187.44 10851.185 188.44 ;
    END
  END MASKD[259]
  PIN MASKD[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10789.865 187.44 10790.145 188.44 ;
    END
  END MASKD[258]
  PIN MASKD[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10772.505 187.44 10772.785 188.44 ;
    END
  END MASKD[257]
  PIN MASKD[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10699.705 187.44 10699.985 188.44 ;
    END
  END MASKD[256]
  PIN MASKD[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10695.225 187.44 10695.505 188.44 ;
    END
  END MASKD[255]
  PIN MASKD[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10629.705 187.44 10629.985 188.44 ;
    END
  END MASKD[254]
  PIN MASKD[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10625.225 187.44 10625.505 188.44 ;
    END
  END MASKD[253]
  PIN MASKD[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10549.905 187.44 10550.185 188.44 ;
    END
  END MASKD[252]
  PIN MASKD[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10519.385 187.44 10519.665 188.44 ;
    END
  END MASKD[251]
  PIN MASKD[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10442.105 187.44 10442.385 188.44 ;
    END
  END MASKD[250]
  PIN MASKD[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10437.625 187.44 10437.905 188.44 ;
    END
  END MASKD[249]
  PIN MASKD[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10376.585 187.44 10376.865 188.44 ;
    END
  END MASKD[248]
  PIN MASKD[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10372.105 187.44 10372.385 188.44 ;
    END
  END MASKD[247]
  PIN MASKD[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10295.385 187.44 10295.665 188.44 ;
    END
  END MASKD[246]
  PIN MASKD[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10290.905 187.44 10291.185 188.44 ;
    END
  END MASKD[245]
  PIN MASKD[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10229.865 187.44 10230.145 188.44 ;
    END
  END MASKD[244]
  PIN MASKD[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10212.505 187.44 10212.785 188.44 ;
    END
  END MASKD[243]
  PIN MASKD[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10139.705 187.44 10139.985 188.44 ;
    END
  END MASKD[242]
  PIN MASKD[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10135.225 187.44 10135.505 188.44 ;
    END
  END MASKD[241]
  PIN MASKD[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10069.705 187.44 10069.985 188.44 ;
    END
  END MASKD[240]
  PIN MASKD[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10065.225 187.44 10065.505 188.44 ;
    END
  END MASKD[239]
  PIN MASKD[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9989.905 187.44 9990.185 188.44 ;
    END
  END MASKD[238]
  PIN MASKD[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9959.385 187.44 9959.665 188.44 ;
    END
  END MASKD[237]
  PIN MASKD[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9882.105 187.44 9882.385 188.44 ;
    END
  END MASKD[236]
  PIN MASKD[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9877.625 187.44 9877.905 188.44 ;
    END
  END MASKD[235]
  PIN MASKD[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9816.585 187.44 9816.865 188.44 ;
    END
  END MASKD[234]
  PIN MASKD[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9812.105 187.44 9812.385 188.44 ;
    END
  END MASKD[233]
  PIN MASKD[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9735.385 187.44 9735.665 188.44 ;
    END
  END MASKD[232]
  PIN MASKD[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9730.905 187.44 9731.185 188.44 ;
    END
  END MASKD[231]
  PIN MASKD[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9669.865 187.44 9670.145 188.44 ;
    END
  END MASKD[230]
  PIN MASKD[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9652.505 187.44 9652.785 188.44 ;
    END
  END MASKD[229]
  PIN MASKD[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9579.705 187.44 9579.985 188.44 ;
    END
  END MASKD[228]
  PIN MASKD[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9575.225 187.44 9575.505 188.44 ;
    END
  END MASKD[227]
  PIN MASKD[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9509.705 187.44 9509.985 188.44 ;
    END
  END MASKD[226]
  PIN MASKD[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9505.225 187.44 9505.505 188.44 ;
    END
  END MASKD[225]
  PIN MASKD[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9429.905 187.44 9430.185 188.44 ;
    END
  END MASKD[224]
  PIN MASKD[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9399.385 187.44 9399.665 188.44 ;
    END
  END MASKD[223]
  PIN MASKD[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9322.105 187.44 9322.385 188.44 ;
    END
  END MASKD[222]
  PIN MASKD[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9317.625 187.44 9317.905 188.44 ;
    END
  END MASKD[221]
  PIN MASKD[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9256.585 187.44 9256.865 188.44 ;
    END
  END MASKD[220]
  PIN MASKD[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9252.105 187.44 9252.385 188.44 ;
    END
  END MASKD[219]
  PIN MASKD[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9175.385 187.44 9175.665 188.44 ;
    END
  END MASKD[218]
  PIN MASKD[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9170.905 187.44 9171.185 188.44 ;
    END
  END MASKD[217]
  PIN MASKD[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9109.865 187.44 9110.145 188.44 ;
    END
  END MASKD[216]
  PIN MASKD[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9092.505 187.44 9092.785 188.44 ;
    END
  END MASKD[215]
  PIN MASKD[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9019.705 187.44 9019.985 188.44 ;
    END
  END MASKD[214]
  PIN MASKD[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9015.225 187.44 9015.505 188.44 ;
    END
  END MASKD[213]
  PIN MASKD[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8949.705 187.44 8949.985 188.44 ;
    END
  END MASKD[212]
  PIN MASKD[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8945.225 187.44 8945.505 188.44 ;
    END
  END MASKD[211]
  PIN MASKD[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8869.905 187.44 8870.185 188.44 ;
    END
  END MASKD[210]
  PIN MASKD[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8839.385 187.44 8839.665 188.44 ;
    END
  END MASKD[209]
  PIN MASKD[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8762.105 187.44 8762.385 188.44 ;
    END
  END MASKD[208]
  PIN MASKD[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8757.625 187.44 8757.905 188.44 ;
    END
  END MASKD[207]
  PIN MASKD[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8696.585 187.44 8696.865 188.44 ;
    END
  END MASKD[206]
  PIN MASKD[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8692.105 187.44 8692.385 188.44 ;
    END
  END MASKD[205]
  PIN MASKD[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8615.385 187.44 8615.665 188.44 ;
    END
  END MASKD[204]
  PIN MASKD[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8610.905 187.44 8611.185 188.44 ;
    END
  END MASKD[203]
  PIN MASKD[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8549.865 187.44 8550.145 188.44 ;
    END
  END MASKD[202]
  PIN MASKD[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8532.505 187.44 8532.785 188.44 ;
    END
  END MASKD[201]
  PIN MASKD[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8459.705 187.44 8459.985 188.44 ;
    END
  END MASKD[200]
  PIN MASKD[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8455.225 187.44 8455.505 188.44 ;
    END
  END MASKD[199]
  PIN MASKD[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8389.705 187.44 8389.985 188.44 ;
    END
  END MASKD[198]
  PIN MASKD[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8385.225 187.44 8385.505 188.44 ;
    END
  END MASKD[197]
  PIN MASKD[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8309.905 187.44 8310.185 188.44 ;
    END
  END MASKD[196]
  PIN MASKD[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8279.385 187.44 8279.665 188.44 ;
    END
  END MASKD[195]
  PIN MASKD[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8202.105 187.44 8202.385 188.44 ;
    END
  END MASKD[194]
  PIN MASKD[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8197.625 187.44 8197.905 188.44 ;
    END
  END MASKD[193]
  PIN MASKD[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8136.585 187.44 8136.865 188.44 ;
    END
  END MASKD[192]
  PIN MASKD[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8132.105 187.44 8132.385 188.44 ;
    END
  END MASKD[191]
  PIN MASKD[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8055.385 187.44 8055.665 188.44 ;
    END
  END MASKD[190]
  PIN MASKD[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8050.905 187.44 8051.185 188.44 ;
    END
  END MASKD[189]
  PIN MASKD[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7989.865 187.44 7990.145 188.44 ;
    END
  END MASKD[188]
  PIN MASKD[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7972.505 187.44 7972.785 188.44 ;
    END
  END MASKD[187]
  PIN MASKD[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7899.705 187.44 7899.985 188.44 ;
    END
  END MASKD[186]
  PIN MASKD[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7895.225 187.44 7895.505 188.44 ;
    END
  END MASKD[185]
  PIN MASKD[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7829.705 187.44 7829.985 188.44 ;
    END
  END MASKD[184]
  PIN MASKD[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7825.225 187.44 7825.505 188.44 ;
    END
  END MASKD[183]
  PIN MASKD[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7749.905 187.44 7750.185 188.44 ;
    END
  END MASKD[182]
  PIN MASKD[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7719.385 187.44 7719.665 188.44 ;
    END
  END MASKD[181]
  PIN MASKD[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7642.105 187.44 7642.385 188.44 ;
    END
  END MASKD[180]
  PIN MASKD[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7637.625 187.44 7637.905 188.44 ;
    END
  END MASKD[179]
  PIN MASKD[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7576.585 187.44 7576.865 188.44 ;
    END
  END MASKD[178]
  PIN MASKD[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7572.105 187.44 7572.385 188.44 ;
    END
  END MASKD[177]
  PIN MASKD[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7495.385 187.44 7495.665 188.44 ;
    END
  END MASKD[176]
  PIN MASKD[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7490.905 187.44 7491.185 188.44 ;
    END
  END MASKD[175]
  PIN MASKD[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7429.865 187.44 7430.145 188.44 ;
    END
  END MASKD[174]
  PIN MASKD[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7412.505 187.44 7412.785 188.44 ;
    END
  END MASKD[173]
  PIN MASKD[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7339.705 187.44 7339.985 188.44 ;
    END
  END MASKD[172]
  PIN MASKD[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7335.225 187.44 7335.505 188.44 ;
    END
  END MASKD[171]
  PIN MASKD[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7269.705 187.44 7269.985 188.44 ;
    END
  END MASKD[170]
  PIN MASKD[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7265.225 187.44 7265.505 188.44 ;
    END
  END MASKD[169]
  PIN MASKD[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7189.905 187.44 7190.185 188.44 ;
    END
  END MASKD[168]
  PIN MASKD[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7159.385 187.44 7159.665 188.44 ;
    END
  END MASKD[167]
  PIN MASKD[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7082.105 187.44 7082.385 188.44 ;
    END
  END MASKD[166]
  PIN MASKD[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7077.625 187.44 7077.905 188.44 ;
    END
  END MASKD[165]
  PIN MASKD[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7016.585 187.44 7016.865 188.44 ;
    END
  END MASKD[164]
  PIN MASKD[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7012.105 187.44 7012.385 188.44 ;
    END
  END MASKD[163]
  PIN MASKD[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6935.385 187.44 6935.665 188.44 ;
    END
  END MASKD[162]
  PIN MASKD[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6930.905 187.44 6931.185 188.44 ;
    END
  END MASKD[161]
  PIN MASKD[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6869.865 187.44 6870.145 188.44 ;
    END
  END MASKD[160]
  PIN MASKD[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6852.505 187.44 6852.785 188.44 ;
    END
  END MASKD[159]
  PIN MASKD[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6779.705 187.44 6779.985 188.44 ;
    END
  END MASKD[158]
  PIN MASKD[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6775.225 187.44 6775.505 188.44 ;
    END
  END MASKD[157]
  PIN MASKD[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6709.705 187.44 6709.985 188.44 ;
    END
  END MASKD[156]
  PIN MASKD[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6705.225 187.44 6705.505 188.44 ;
    END
  END MASKD[155]
  PIN MASKD[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6629.905 187.44 6630.185 188.44 ;
    END
  END MASKD[154]
  PIN MASKD[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6599.385 187.44 6599.665 188.44 ;
    END
  END MASKD[153]
  PIN MASKD[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6522.105 187.44 6522.385 188.44 ;
    END
  END MASKD[152]
  PIN MASKD[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6517.625 187.44 6517.905 188.44 ;
    END
  END MASKD[151]
  PIN MASKD[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6456.585 187.44 6456.865 188.44 ;
    END
  END MASKD[150]
  PIN MASKD[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6452.105 187.44 6452.385 188.44 ;
    END
  END MASKD[149]
  PIN MASKD[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6375.385 187.44 6375.665 188.44 ;
    END
  END MASKD[148]
  PIN MASKD[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6370.905 187.44 6371.185 188.44 ;
    END
  END MASKD[147]
  PIN MASKD[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6309.865 187.44 6310.145 188.44 ;
    END
  END MASKD[146]
  PIN MASKD[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6292.505 187.44 6292.785 188.44 ;
    END
  END MASKD[145]
  PIN MASKD[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6219.705 187.44 6219.985 188.44 ;
    END
  END MASKD[144]
  PIN MASKD[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6215.225 187.44 6215.505 188.44 ;
    END
  END MASKD[143]
  PIN MASKD[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6149.705 187.44 6149.985 188.44 ;
    END
  END MASKD[142]
  PIN MASKD[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6145.225 187.44 6145.505 188.44 ;
    END
  END MASKD[141]
  PIN MASKD[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6069.905 187.44 6070.185 188.44 ;
    END
  END MASKD[140]
  PIN MASKD[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6039.385 187.44 6039.665 188.44 ;
    END
  END MASKD[139]
  PIN MASKD[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5962.105 187.44 5962.385 188.44 ;
    END
  END MASKD[138]
  PIN MASKD[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5957.625 187.44 5957.905 188.44 ;
    END
  END MASKD[137]
  PIN MASKD[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5896.585 187.44 5896.865 188.44 ;
    END
  END MASKD[136]
  PIN MASKD[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5892.105 187.44 5892.385 188.44 ;
    END
  END MASKD[135]
  PIN MASKD[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5815.385 187.44 5815.665 188.44 ;
    END
  END MASKD[134]
  PIN MASKD[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5810.905 187.44 5811.185 188.44 ;
    END
  END MASKD[133]
  PIN MASKD[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5749.865 187.44 5750.145 188.44 ;
    END
  END MASKD[132]
  PIN MASKD[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5732.505 187.44 5732.785 188.44 ;
    END
  END MASKD[131]
  PIN MASKD[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5659.705 187.44 5659.985 188.44 ;
    END
  END MASKD[130]
  PIN MASKD[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5655.225 187.44 5655.505 188.44 ;
    END
  END MASKD[129]
  PIN MASKD[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5589.705 187.44 5589.985 188.44 ;
    END
  END MASKD[128]
  PIN MASKD[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5585.225 187.44 5585.505 188.44 ;
    END
  END MASKD[127]
  PIN MASKD[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5509.905 187.44 5510.185 188.44 ;
    END
  END MASKD[126]
  PIN MASKD[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5479.385 187.44 5479.665 188.44 ;
    END
  END MASKD[125]
  PIN MASKD[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5402.105 187.44 5402.385 188.44 ;
    END
  END MASKD[124]
  PIN MASKD[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5397.625 187.44 5397.905 188.44 ;
    END
  END MASKD[123]
  PIN MASKD[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5336.585 187.44 5336.865 188.44 ;
    END
  END MASKD[122]
  PIN MASKD[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5332.105 187.44 5332.385 188.44 ;
    END
  END MASKD[121]
  PIN MASKD[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5255.385 187.44 5255.665 188.44 ;
    END
  END MASKD[120]
  PIN MASKD[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5250.905 187.44 5251.185 188.44 ;
    END
  END MASKD[119]
  PIN MASKD[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5189.865 187.44 5190.145 188.44 ;
    END
  END MASKD[118]
  PIN MASKD[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5172.505 187.44 5172.785 188.44 ;
    END
  END MASKD[117]
  PIN MASKD[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5099.705 187.44 5099.985 188.44 ;
    END
  END MASKD[116]
  PIN MASKD[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5095.225 187.44 5095.505 188.44 ;
    END
  END MASKD[115]
  PIN MASKD[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5029.705 187.44 5029.985 188.44 ;
    END
  END MASKD[114]
  PIN MASKD[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5025.225 187.44 5025.505 188.44 ;
    END
  END MASKD[113]
  PIN MASKD[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4949.905 187.44 4950.185 188.44 ;
    END
  END MASKD[112]
  PIN MASKD[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4919.385 187.44 4919.665 188.44 ;
    END
  END MASKD[111]
  PIN MASKD[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4842.105 187.44 4842.385 188.44 ;
    END
  END MASKD[110]
  PIN MASKD[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4837.625 187.44 4837.905 188.44 ;
    END
  END MASKD[109]
  PIN MASKD[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4776.585 187.44 4776.865 188.44 ;
    END
  END MASKD[108]
  PIN MASKD[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4772.105 187.44 4772.385 188.44 ;
    END
  END MASKD[107]
  PIN MASKD[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4695.385 187.44 4695.665 188.44 ;
    END
  END MASKD[106]
  PIN MASKD[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4690.905 187.44 4691.185 188.44 ;
    END
  END MASKD[105]
  PIN MASKD[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4629.865 187.44 4630.145 188.44 ;
    END
  END MASKD[104]
  PIN MASKD[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4612.505 187.44 4612.785 188.44 ;
    END
  END MASKD[103]
  PIN MASKD[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4539.705 187.44 4539.985 188.44 ;
    END
  END MASKD[102]
  PIN MASKD[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4535.225 187.44 4535.505 188.44 ;
    END
  END MASKD[101]
  PIN MASKD[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4469.705 187.44 4469.985 188.44 ;
    END
  END MASKD[100]
  PIN MASKD[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4465.225 187.44 4465.505 188.44 ;
    END
  END MASKD[99]
  PIN MASKD[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4389.905 187.44 4390.185 188.44 ;
    END
  END MASKD[98]
  PIN MASKD[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4359.385 187.44 4359.665 188.44 ;
    END
  END MASKD[97]
  PIN MASKD[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4282.105 187.44 4282.385 188.44 ;
    END
  END MASKD[96]
  PIN MASKD[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4277.625 187.44 4277.905 188.44 ;
    END
  END MASKD[95]
  PIN MASKD[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4216.585 187.44 4216.865 188.44 ;
    END
  END MASKD[94]
  PIN MASKD[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4212.105 187.44 4212.385 188.44 ;
    END
  END MASKD[93]
  PIN MASKD[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4135.385 187.44 4135.665 188.44 ;
    END
  END MASKD[92]
  PIN MASKD[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4130.905 187.44 4131.185 188.44 ;
    END
  END MASKD[91]
  PIN MASKD[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4069.865 187.44 4070.145 188.44 ;
    END
  END MASKD[90]
  PIN MASKD[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4052.505 187.44 4052.785 188.44 ;
    END
  END MASKD[89]
  PIN MASKD[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3979.705 187.44 3979.985 188.44 ;
    END
  END MASKD[88]
  PIN MASKD[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3975.225 187.44 3975.505 188.44 ;
    END
  END MASKD[87]
  PIN MASKD[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3909.705 187.44 3909.985 188.44 ;
    END
  END MASKD[86]
  PIN MASKD[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3905.225 187.44 3905.505 188.44 ;
    END
  END MASKD[85]
  PIN MASKD[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3829.905 187.44 3830.185 188.44 ;
    END
  END MASKD[84]
  PIN MASKD[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3799.385 187.44 3799.665 188.44 ;
    END
  END MASKD[83]
  PIN MASKD[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3722.105 187.44 3722.385 188.44 ;
    END
  END MASKD[82]
  PIN MASKD[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3717.625 187.44 3717.905 188.44 ;
    END
  END MASKD[81]
  PIN MASKD[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3656.585 187.44 3656.865 188.44 ;
    END
  END MASKD[80]
  PIN MASKD[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3652.105 187.44 3652.385 188.44 ;
    END
  END MASKD[79]
  PIN MASKD[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3575.385 187.44 3575.665 188.44 ;
    END
  END MASKD[78]
  PIN MASKD[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3570.905 187.44 3571.185 188.44 ;
    END
  END MASKD[77]
  PIN MASKD[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3509.865 187.44 3510.145 188.44 ;
    END
  END MASKD[76]
  PIN MASKD[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3492.505 187.44 3492.785 188.44 ;
    END
  END MASKD[75]
  PIN MASKD[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3419.705 187.44 3419.985 188.44 ;
    END
  END MASKD[74]
  PIN MASKD[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3415.225 187.44 3415.505 188.44 ;
    END
  END MASKD[73]
  PIN MASKD[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3349.705 187.44 3349.985 188.44 ;
    END
  END MASKD[72]
  PIN MASKD[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3345.225 187.44 3345.505 188.44 ;
    END
  END MASKD[71]
  PIN MASKD[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3269.905 187.44 3270.185 188.44 ;
    END
  END MASKD[70]
  PIN MASKD[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3239.385 187.44 3239.665 188.44 ;
    END
  END MASKD[69]
  PIN MASKD[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3162.105 187.44 3162.385 188.44 ;
    END
  END MASKD[68]
  PIN MASKD[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3157.625 187.44 3157.905 188.44 ;
    END
  END MASKD[67]
  PIN MASKD[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3096.585 187.44 3096.865 188.44 ;
    END
  END MASKD[66]
  PIN MASKD[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3092.105 187.44 3092.385 188.44 ;
    END
  END MASKD[65]
  PIN MASKD[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3015.385 187.44 3015.665 188.44 ;
    END
  END MASKD[64]
  PIN MASKD[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3010.905 187.44 3011.185 188.44 ;
    END
  END MASKD[63]
  PIN MASKD[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2949.865 187.44 2950.145 188.44 ;
    END
  END MASKD[62]
  PIN MASKD[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2932.505 187.44 2932.785 188.44 ;
    END
  END MASKD[61]
  PIN MASKD[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2859.705 187.44 2859.985 188.44 ;
    END
  END MASKD[60]
  PIN MASKD[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2855.225 187.44 2855.505 188.44 ;
    END
  END MASKD[59]
  PIN MASKD[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2789.705 187.44 2789.985 188.44 ;
    END
  END MASKD[58]
  PIN MASKD[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2785.225 187.44 2785.505 188.44 ;
    END
  END MASKD[57]
  PIN MASKD[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2709.905 187.44 2710.185 188.44 ;
    END
  END MASKD[56]
  PIN MASKD[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2679.385 187.44 2679.665 188.44 ;
    END
  END MASKD[55]
  PIN MASKD[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2602.105 187.44 2602.385 188.44 ;
    END
  END MASKD[54]
  PIN MASKD[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2597.625 187.44 2597.905 188.44 ;
    END
  END MASKD[53]
  PIN MASKD[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2536.585 187.44 2536.865 188.44 ;
    END
  END MASKD[52]
  PIN MASKD[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2532.105 187.44 2532.385 188.44 ;
    END
  END MASKD[51]
  PIN MASKD[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2455.385 187.44 2455.665 188.44 ;
    END
  END MASKD[50]
  PIN MASKD[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2450.905 187.44 2451.185 188.44 ;
    END
  END MASKD[49]
  PIN MASKD[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2389.865 187.44 2390.145 188.44 ;
    END
  END MASKD[48]
  PIN MASKD[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2372.505 187.44 2372.785 188.44 ;
    END
  END MASKD[47]
  PIN MASKD[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2299.705 187.44 2299.985 188.44 ;
    END
  END MASKD[46]
  PIN MASKD[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2295.225 187.44 2295.505 188.44 ;
    END
  END MASKD[45]
  PIN MASKD[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2229.705 187.44 2229.985 188.44 ;
    END
  END MASKD[44]
  PIN MASKD[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2225.225 187.44 2225.505 188.44 ;
    END
  END MASKD[43]
  PIN MASKD[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2149.905 187.44 2150.185 188.44 ;
    END
  END MASKD[42]
  PIN MASKD[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2119.385 187.44 2119.665 188.44 ;
    END
  END MASKD[41]
  PIN MASKD[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2042.105 187.44 2042.385 188.44 ;
    END
  END MASKD[40]
  PIN MASKD[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2037.625 187.44 2037.905 188.44 ;
    END
  END MASKD[39]
  PIN MASKD[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1976.585 187.44 1976.865 188.44 ;
    END
  END MASKD[38]
  PIN MASKD[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1972.105 187.44 1972.385 188.44 ;
    END
  END MASKD[37]
  PIN MASKD[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1895.385 187.44 1895.665 188.44 ;
    END
  END MASKD[36]
  PIN MASKD[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1890.905 187.44 1891.185 188.44 ;
    END
  END MASKD[35]
  PIN MASKD[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1829.865 187.44 1830.145 188.44 ;
    END
  END MASKD[34]
  PIN MASKD[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1812.505 187.44 1812.785 188.44 ;
    END
  END MASKD[33]
  PIN MASKD[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1739.705 187.44 1739.985 188.44 ;
    END
  END MASKD[32]
  PIN MASKD[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1735.225 187.44 1735.505 188.44 ;
    END
  END MASKD[31]
  PIN MASKD[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1669.705 187.44 1669.985 188.44 ;
    END
  END MASKD[30]
  PIN MASKD[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1665.225 187.44 1665.505 188.44 ;
    END
  END MASKD[29]
  PIN MASKD[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1589.905 187.44 1590.185 188.44 ;
    END
  END MASKD[28]
  PIN MASKD[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1559.385 187.44 1559.665 188.44 ;
    END
  END MASKD[27]
  PIN MASKD[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1482.105 187.44 1482.385 188.44 ;
    END
  END MASKD[26]
  PIN MASKD[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1477.625 187.44 1477.905 188.44 ;
    END
  END MASKD[25]
  PIN MASKD[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1416.585 187.44 1416.865 188.44 ;
    END
  END MASKD[24]
  PIN MASKD[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1412.105 187.44 1412.385 188.44 ;
    END
  END MASKD[23]
  PIN MASKD[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1335.385 187.44 1335.665 188.44 ;
    END
  END MASKD[22]
  PIN MASKD[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1330.905 187.44 1331.185 188.44 ;
    END
  END MASKD[21]
  PIN MASKD[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1269.865 187.44 1270.145 188.44 ;
    END
  END MASKD[20]
  PIN MASKD[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1252.505 187.44 1252.785 188.44 ;
    END
  END MASKD[19]
  PIN MASKD[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1179.705 187.44 1179.985 188.44 ;
    END
  END MASKD[18]
  PIN MASKD[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1175.225 187.44 1175.505 188.44 ;
    END
  END MASKD[17]
  PIN MASKD[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1109.705 187.44 1109.985 188.44 ;
    END
  END MASKD[16]
  PIN MASKD[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1105.225 187.44 1105.505 188.44 ;
    END
  END MASKD[15]
  PIN MASKD[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1029.905 187.44 1030.185 188.44 ;
    END
  END MASKD[14]
  PIN MASKD[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 999.385 187.44 999.665 188.44 ;
    END
  END MASKD[13]
  PIN MASKD[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 922.105 187.44 922.385 188.44 ;
    END
  END MASKD[12]
  PIN MASKD[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 917.625 187.44 917.905 188.44 ;
    END
  END MASKD[11]
  PIN MASKD[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 856.585 187.44 856.865 188.44 ;
    END
  END MASKD[10]
  PIN MASKD[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 852.105 187.44 852.385 188.44 ;
    END
  END MASKD[9]
  PIN MASKD[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 775.385 187.44 775.665 188.44 ;
    END
  END MASKD[8]
  PIN MASKD[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 770.905 187.44 771.185 188.44 ;
    END
  END MASKD[7]
  PIN MASKD[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 709.865 187.44 710.145 188.44 ;
    END
  END MASKD[6]
  PIN MASKD[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 692.505 187.44 692.785 188.44 ;
    END
  END MASKD[5]
  PIN MASKD[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 619.705 187.44 619.985 188.44 ;
    END
  END MASKD[4]
  PIN MASKD[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 615.225 187.44 615.505 188.44 ;
    END
  END MASKD[3]
  PIN MASKD[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 549.705 187.44 549.985 188.44 ;
    END
  END MASKD[2]
  PIN MASKD[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 545.225 187.44 545.505 188.44 ;
    END
  END MASKD[1]
  PIN MASKD[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 469.905 187.44 470.185 188.44 ;
    END
  END MASKD[0]
  PIN nRST
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 467.665 187.44 467.945 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 547.465 187.44 547.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 617.465 187.44 617.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 694.745 187.44 695.025 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 773.145 187.44 773.425 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 854.345 187.44 854.625 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 919.865 187.44 920.145 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 1027.665 187.44 1027.945 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 1107.465 187.44 1107.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 1177.465 187.44 1177.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 1254.745 187.44 1255.025 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 1333.145 187.44 1333.425 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 1414.345 187.44 1414.625 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 1479.865 187.44 1480.145 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 1587.665 187.44 1587.945 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 1667.465 187.44 1667.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 1737.465 187.44 1737.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 1814.745 187.44 1815.025 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 1893.145 187.44 1893.425 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 1974.345 187.44 1974.625 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 2039.865 187.44 2040.145 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 2147.665 187.44 2147.945 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 2227.465 187.44 2227.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 2297.465 187.44 2297.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 2374.745 187.44 2375.025 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 2453.145 187.44 2453.425 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 2534.345 187.44 2534.625 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 2599.865 187.44 2600.145 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 2707.665 187.44 2707.945 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 2787.465 187.44 2787.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 2857.465 187.44 2857.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 2934.745 187.44 2935.025 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 3013.145 187.44 3013.425 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 3094.345 187.44 3094.625 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 3159.865 187.44 3160.145 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 3267.665 187.44 3267.945 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 3347.465 187.44 3347.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 3417.465 187.44 3417.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 3494.745 187.44 3495.025 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 3573.145 187.44 3573.425 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 3654.345 187.44 3654.625 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 3719.865 187.44 3720.145 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 3827.665 187.44 3827.945 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 3907.465 187.44 3907.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 3977.465 187.44 3977.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 4054.745 187.44 4055.025 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 4133.145 187.44 4133.425 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 4214.345 187.44 4214.625 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 4279.865 187.44 4280.145 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 4387.665 187.44 4387.945 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 4467.465 187.44 4467.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 4537.465 187.44 4537.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 4614.745 187.44 4615.025 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 4693.145 187.44 4693.425 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 4774.345 187.44 4774.625 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 4839.865 187.44 4840.145 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 4947.665 187.44 4947.945 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 5027.465 187.44 5027.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 5097.465 187.44 5097.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 5174.745 187.44 5175.025 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 5253.145 187.44 5253.425 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 5334.345 187.44 5334.625 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 5399.865 187.44 5400.145 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 5507.665 187.44 5507.945 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 5587.465 187.44 5587.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 5657.465 187.44 5657.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 5734.745 187.44 5735.025 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 5813.145 187.44 5813.425 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 5894.345 187.44 5894.625 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 5959.865 187.44 5960.145 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 6067.665 187.44 6067.945 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 6147.465 187.44 6147.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 6217.465 187.44 6217.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 6294.745 187.44 6295.025 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 6373.145 187.44 6373.425 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 6454.345 187.44 6454.625 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 6519.865 187.44 6520.145 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 6627.665 187.44 6627.945 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 6707.465 187.44 6707.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 6777.465 187.44 6777.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 6854.745 187.44 6855.025 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 6933.145 187.44 6933.425 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 7014.345 187.44 7014.625 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 7079.865 187.44 7080.145 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 7187.665 187.44 7187.945 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 7267.465 187.44 7267.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 7337.465 187.44 7337.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 7414.745 187.44 7415.025 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 7493.145 187.44 7493.425 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 7574.345 187.44 7574.625 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 7639.865 187.44 7640.145 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 7747.665 187.44 7747.945 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 7827.465 187.44 7827.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 7897.465 187.44 7897.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 7974.745 187.44 7975.025 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 8053.145 187.44 8053.425 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 8134.345 187.44 8134.625 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 8199.865 187.44 8200.145 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 8307.665 187.44 8307.945 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 8387.465 187.44 8387.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 8457.465 187.44 8457.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 8534.745 187.44 8535.025 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 8613.145 187.44 8613.425 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 8694.345 187.44 8694.625 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 8759.865 187.44 8760.145 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 8867.665 187.44 8867.945 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 8947.465 187.44 8947.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 9017.465 187.44 9017.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 9094.745 187.44 9095.025 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 9173.145 187.44 9173.425 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 9254.345 187.44 9254.625 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 9319.865 187.44 9320.145 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 9427.665 187.44 9427.945 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 9507.465 187.44 9507.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 9577.465 187.44 9577.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 9654.745 187.44 9655.025 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 9733.145 187.44 9733.425 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 9814.345 187.44 9814.625 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 9879.865 187.44 9880.145 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 9987.665 187.44 9987.945 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 10067.465 187.44 10067.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 10137.465 187.44 10137.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 10214.745 187.44 10215.025 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 10293.145 187.44 10293.425 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 10374.345 187.44 10374.625 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 10439.865 187.44 10440.145 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 10547.665 187.44 10547.945 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 10627.465 187.44 10627.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 10697.465 187.44 10697.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 10774.745 187.44 10775.025 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 10853.145 187.44 10853.425 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 10934.345 187.44 10934.625 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 10999.865 187.44 11000.145 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 11107.665 187.44 11107.945 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 11187.465 187.44 11187.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 11257.465 187.44 11257.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 11334.745 187.44 11335.025 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 11413.145 187.44 11413.425 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 11494.345 187.44 11494.625 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 11559.865 187.44 11560.145 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 11667.665 187.44 11667.945 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 11747.465 187.44 11747.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 11817.465 187.44 11817.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 11894.745 187.44 11895.025 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 11973.145 187.44 11973.425 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 12054.345 187.44 12054.625 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 12119.865 187.44 12120.145 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 12227.665 187.44 12227.945 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 12307.465 187.44 12307.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 12377.465 187.44 12377.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 12454.745 187.44 12455.025 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 12533.145 187.44 12533.425 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 12614.345 187.44 12614.625 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 12679.865 187.44 12680.145 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 12787.665 187.44 12787.945 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 12867.465 187.44 12867.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 12937.465 187.44 12937.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 13014.745 187.44 13015.025 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 13093.145 187.44 13093.425 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 13174.345 187.44 13174.625 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 13239.865 187.44 13240.145 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 13347.665 187.44 13347.945 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 13427.465 187.44 13427.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 13497.465 187.44 13497.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 13574.745 187.44 13575.025 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 13653.145 187.44 13653.425 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 13734.345 187.44 13734.625 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 13799.865 187.44 13800.145 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 13907.665 187.44 13907.945 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 13987.465 187.44 13987.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 14057.465 187.44 14057.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 14134.745 187.44 14135.025 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 14213.145 187.44 14213.425 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 14294.345 187.44 14294.625 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 14359.865 187.44 14360.145 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 14467.665 187.44 14467.945 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 14547.465 187.44 14547.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 14617.465 187.44 14617.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 14694.745 187.44 14695.025 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 14773.145 187.44 14773.425 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 14854.345 187.44 14854.625 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 14919.865 187.44 14920.145 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 15027.665 187.44 15027.945 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 15107.465 187.44 15107.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 15177.465 187.44 15177.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 15254.745 187.44 15255.025 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 15333.145 187.44 15333.425 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 15414.345 187.44 15414.625 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 15479.865 187.44 15480.145 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 15587.665 187.44 15587.945 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 15667.465 187.44 15667.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 15737.465 187.44 15737.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 15814.745 187.44 15815.025 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 15893.145 187.44 15893.425 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 15974.345 187.44 15974.625 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 16039.865 187.44 16040.145 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 16147.665 187.44 16147.945 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 16227.465 187.44 16227.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 16297.465 187.44 16297.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 16374.745 187.44 16375.025 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 16453.145 187.44 16453.425 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 16534.345 187.44 16534.625 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 16599.865 187.44 16600.145 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 16707.665 187.44 16707.945 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 16787.465 187.44 16787.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 16857.465 187.44 16857.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 16934.745 187.44 16935.025 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 17013.145 187.44 17013.425 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 17094.345 187.44 17094.625 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 17159.865 187.44 17160.145 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 17267.665 187.44 17267.945 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 17347.465 187.44 17347.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 17417.465 187.44 17417.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 17494.745 187.44 17495.025 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 17573.145 187.44 17573.425 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 17654.345 187.44 17654.625 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 17719.865 187.44 17720.145 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 17827.665 187.44 17827.945 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 17907.465 187.44 17907.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 17977.465 187.44 17977.745 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 18054.745 187.44 18055.025 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 18133.145 187.44 18133.425 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 18214.345 187.44 18214.625 188.44 ;
    END
    PORT
      LAYER M4 ;
        RECT 18279.865 187.44 18280.145 188.44 ;
    END
  END nRST
  PIN Read_PMOS[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9371.945 187.44 9372.225 188.44 ;
    END
  END Read_PMOS[55]
  PIN Read_PMOS[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9295.225 187.44 9295.505 188.44 ;
    END
  END Read_PMOS[54]
  PIN Read_PMOS[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9225.225 187.44 9225.505 188.44 ;
    END
  END Read_PMOS[53]
  PIN Read_PMOS[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9121.065 187.44 9121.345 188.44 ;
    END
  END Read_PMOS[52]
  PIN Read_PMOS[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9039.305 187.44 9039.585 188.44 ;
    END
  END Read_PMOS[51]
  PIN Read_PMOS[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8973.785 187.44 8974.065 188.44 ;
    END
  END Read_PMOS[50]
  PIN Read_PMOS[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8891.465 187.44 8891.745 188.44 ;
    END
  END Read_PMOS[49]
  PIN Read_PMOS[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8811.945 187.44 8812.225 188.44 ;
    END
  END Read_PMOS[48]
  PIN Read_PMOS[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8735.225 187.44 8735.505 188.44 ;
    END
  END Read_PMOS[47]
  PIN Read_PMOS[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8665.225 187.44 8665.505 188.44 ;
    END
  END Read_PMOS[46]
  PIN Read_PMOS[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8561.065 187.44 8561.345 188.44 ;
    END
  END Read_PMOS[45]
  PIN Read_PMOS[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8479.305 187.44 8479.585 188.44 ;
    END
  END Read_PMOS[44]
  PIN Read_PMOS[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8413.785 187.44 8414.065 188.44 ;
    END
  END Read_PMOS[43]
  PIN Read_PMOS[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8331.465 187.44 8331.745 188.44 ;
    END
  END Read_PMOS[42]
  PIN Read_PMOS[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8251.945 187.44 8252.225 188.44 ;
    END
  END Read_PMOS[41]
  PIN Read_PMOS[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8175.225 187.44 8175.505 188.44 ;
    END
  END Read_PMOS[40]
  PIN Read_PMOS[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8105.225 187.44 8105.505 188.44 ;
    END
  END Read_PMOS[39]
  PIN Read_PMOS[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8001.065 187.44 8001.345 188.44 ;
    END
  END Read_PMOS[38]
  PIN Read_PMOS[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7919.305 187.44 7919.585 188.44 ;
    END
  END Read_PMOS[37]
  PIN Read_PMOS[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7853.785 187.44 7854.065 188.44 ;
    END
  END Read_PMOS[36]
  PIN Read_PMOS[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7771.465 187.44 7771.745 188.44 ;
    END
  END Read_PMOS[35]
  PIN Read_PMOS[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7691.945 187.44 7692.225 188.44 ;
    END
  END Read_PMOS[34]
  PIN Read_PMOS[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7615.225 187.44 7615.505 188.44 ;
    END
  END Read_PMOS[33]
  PIN Read_PMOS[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7545.225 187.44 7545.505 188.44 ;
    END
  END Read_PMOS[32]
  PIN Read_PMOS[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7441.065 187.44 7441.345 188.44 ;
    END
  END Read_PMOS[31]
  PIN Read_PMOS[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7359.305 187.44 7359.585 188.44 ;
    END
  END Read_PMOS[30]
  PIN Read_PMOS[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7293.785 187.44 7294.065 188.44 ;
    END
  END Read_PMOS[29]
  PIN Read_PMOS[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7211.465 187.44 7211.745 188.44 ;
    END
  END Read_PMOS[28]
  PIN Read_PMOS[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7131.945 187.44 7132.225 188.44 ;
    END
  END Read_PMOS[27]
  PIN Read_PMOS[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7055.225 187.44 7055.505 188.44 ;
    END
  END Read_PMOS[26]
  PIN Read_PMOS[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6985.225 187.44 6985.505 188.44 ;
    END
  END Read_PMOS[25]
  PIN Read_PMOS[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6881.065 187.44 6881.345 188.44 ;
    END
  END Read_PMOS[24]
  PIN Read_PMOS[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6799.305 187.44 6799.585 188.44 ;
    END
  END Read_PMOS[23]
  PIN Read_PMOS[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6733.785 187.44 6734.065 188.44 ;
    END
  END Read_PMOS[22]
  PIN Read_PMOS[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6651.465 187.44 6651.745 188.44 ;
    END
  END Read_PMOS[21]
  PIN Read_PMOS[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6571.945 187.44 6572.225 188.44 ;
    END
  END Read_PMOS[20]
  PIN Read_PMOS[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6495.225 187.44 6495.505 188.44 ;
    END
  END Read_PMOS[19]
  PIN Read_PMOS[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6425.225 187.44 6425.505 188.44 ;
    END
  END Read_PMOS[18]
  PIN Read_PMOS[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6321.065 187.44 6321.345 188.44 ;
    END
  END Read_PMOS[17]
  PIN Read_PMOS[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6239.305 187.44 6239.585 188.44 ;
    END
  END Read_PMOS[16]
  PIN Read_PMOS[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6173.785 187.44 6174.065 188.44 ;
    END
  END Read_PMOS[15]
  PIN Read_PMOS[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6091.465 187.44 6091.745 188.44 ;
    END
  END Read_PMOS[14]
  PIN Read_PMOS[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6011.945 187.44 6012.225 188.44 ;
    END
  END Read_PMOS[13]
  PIN Read_PMOS[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5935.225 187.44 5935.505 188.44 ;
    END
  END Read_PMOS[12]
  PIN Read_PMOS[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5865.225 187.44 5865.505 188.44 ;
    END
  END Read_PMOS[11]
  PIN Read_PMOS[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5761.065 187.44 5761.345 188.44 ;
    END
  END Read_PMOS[10]
  PIN Read_PMOS[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5679.305 187.44 5679.585 188.44 ;
    END
  END Read_PMOS[9]
  PIN Read_PMOS[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5613.785 187.44 5614.065 188.44 ;
    END
  END Read_PMOS[8]
  PIN Read_PMOS[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5531.465 187.44 5531.745 188.44 ;
    END
  END Read_PMOS[7]
  PIN Read_PMOS[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5451.945 187.44 5452.225 188.44 ;
    END
  END Read_PMOS[6]
  PIN Read_PMOS[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5375.225 187.44 5375.505 188.44 ;
    END
  END Read_PMOS[5]
  PIN Read_PMOS[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5305.225 187.44 5305.505 188.44 ;
    END
  END Read_PMOS[4]
  PIN Read_PMOS[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5201.065 187.44 5201.345 188.44 ;
    END
  END Read_PMOS[3]
  PIN Read_PMOS[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5119.305 187.44 5119.585 188.44 ;
    END
  END Read_PMOS[2]
  PIN Read_PMOS[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5053.785 187.44 5054.065 188.44 ;
    END
  END Read_PMOS[1]
  PIN Read_PMOS[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4971.465 187.44 4971.745 188.44 ;
    END
  END Read_PMOS[0]
  PIN FREEZE_PMOS[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9372.505 187.44 9372.785 188.44 ;
    END
  END FREEZE_PMOS[55]
  PIN FREEZE_PMOS[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9295.785 187.44 9296.065 188.44 ;
    END
  END FREEZE_PMOS[54]
  PIN FREEZE_PMOS[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9225.785 187.44 9226.065 188.44 ;
    END
  END FREEZE_PMOS[53]
  PIN FREEZE_PMOS[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9121.625 187.44 9121.905 188.44 ;
    END
  END FREEZE_PMOS[52]
  PIN FREEZE_PMOS[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9039.865 187.44 9040.145 188.44 ;
    END
  END FREEZE_PMOS[51]
  PIN FREEZE_PMOS[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8974.345 187.44 8974.625 188.44 ;
    END
  END FREEZE_PMOS[50]
  PIN FREEZE_PMOS[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8892.025 187.44 8892.305 188.44 ;
    END
  END FREEZE_PMOS[49]
  PIN FREEZE_PMOS[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8812.505 187.44 8812.785 188.44 ;
    END
  END FREEZE_PMOS[48]
  PIN FREEZE_PMOS[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8735.785 187.44 8736.065 188.44 ;
    END
  END FREEZE_PMOS[47]
  PIN FREEZE_PMOS[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8665.785 187.44 8666.065 188.44 ;
    END
  END FREEZE_PMOS[46]
  PIN FREEZE_PMOS[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8561.625 187.44 8561.905 188.44 ;
    END
  END FREEZE_PMOS[45]
  PIN FREEZE_PMOS[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8479.865 187.44 8480.145 188.44 ;
    END
  END FREEZE_PMOS[44]
  PIN FREEZE_PMOS[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8414.345 187.44 8414.625 188.44 ;
    END
  END FREEZE_PMOS[43]
  PIN FREEZE_PMOS[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8332.025 187.44 8332.305 188.44 ;
    END
  END FREEZE_PMOS[42]
  PIN FREEZE_PMOS[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8252.505 187.44 8252.785 188.44 ;
    END
  END FREEZE_PMOS[41]
  PIN FREEZE_PMOS[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8175.785 187.44 8176.065 188.44 ;
    END
  END FREEZE_PMOS[40]
  PIN FREEZE_PMOS[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8105.785 187.44 8106.065 188.44 ;
    END
  END FREEZE_PMOS[39]
  PIN FREEZE_PMOS[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8001.625 187.44 8001.905 188.44 ;
    END
  END FREEZE_PMOS[38]
  PIN FREEZE_PMOS[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7919.865 187.44 7920.145 188.44 ;
    END
  END FREEZE_PMOS[37]
  PIN FREEZE_PMOS[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7854.345 187.44 7854.625 188.44 ;
    END
  END FREEZE_PMOS[36]
  PIN FREEZE_PMOS[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7772.025 187.44 7772.305 188.44 ;
    END
  END FREEZE_PMOS[35]
  PIN FREEZE_PMOS[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7692.505 187.44 7692.785 188.44 ;
    END
  END FREEZE_PMOS[34]
  PIN FREEZE_PMOS[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7615.785 187.44 7616.065 188.44 ;
    END
  END FREEZE_PMOS[33]
  PIN FREEZE_PMOS[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7545.785 187.44 7546.065 188.44 ;
    END
  END FREEZE_PMOS[32]
  PIN FREEZE_PMOS[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7441.625 187.44 7441.905 188.44 ;
    END
  END FREEZE_PMOS[31]
  PIN FREEZE_PMOS[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7359.865 187.44 7360.145 188.44 ;
    END
  END FREEZE_PMOS[30]
  PIN FREEZE_PMOS[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7294.345 187.44 7294.625 188.44 ;
    END
  END FREEZE_PMOS[29]
  PIN FREEZE_PMOS[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7212.025 187.44 7212.305 188.44 ;
    END
  END FREEZE_PMOS[28]
  PIN FREEZE_PMOS[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7132.505 187.44 7132.785 188.44 ;
    END
  END FREEZE_PMOS[27]
  PIN FREEZE_PMOS[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7055.785 187.44 7056.065 188.44 ;
    END
  END FREEZE_PMOS[26]
  PIN FREEZE_PMOS[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6985.785 187.44 6986.065 188.44 ;
    END
  END FREEZE_PMOS[25]
  PIN FREEZE_PMOS[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6881.625 187.44 6881.905 188.44 ;
    END
  END FREEZE_PMOS[24]
  PIN FREEZE_PMOS[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6799.865 187.44 6800.145 188.44 ;
    END
  END FREEZE_PMOS[23]
  PIN FREEZE_PMOS[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6734.345 187.44 6734.625 188.44 ;
    END
  END FREEZE_PMOS[22]
  PIN FREEZE_PMOS[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6652.025 187.44 6652.305 188.44 ;
    END
  END FREEZE_PMOS[21]
  PIN FREEZE_PMOS[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6572.505 187.44 6572.785 188.44 ;
    END
  END FREEZE_PMOS[20]
  PIN FREEZE_PMOS[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6495.785 187.44 6496.065 188.44 ;
    END
  END FREEZE_PMOS[19]
  PIN FREEZE_PMOS[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6425.785 187.44 6426.065 188.44 ;
    END
  END FREEZE_PMOS[18]
  PIN FREEZE_PMOS[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6321.625 187.44 6321.905 188.44 ;
    END
  END FREEZE_PMOS[17]
  PIN FREEZE_PMOS[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6239.865 187.44 6240.145 188.44 ;
    END
  END FREEZE_PMOS[16]
  PIN FREEZE_PMOS[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6174.345 187.44 6174.625 188.44 ;
    END
  END FREEZE_PMOS[15]
  PIN FREEZE_PMOS[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6092.025 187.44 6092.305 188.44 ;
    END
  END FREEZE_PMOS[14]
  PIN FREEZE_PMOS[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6012.505 187.44 6012.785 188.44 ;
    END
  END FREEZE_PMOS[13]
  PIN FREEZE_PMOS[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5935.785 187.44 5936.065 188.44 ;
    END
  END FREEZE_PMOS[12]
  PIN FREEZE_PMOS[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5865.785 187.44 5866.065 188.44 ;
    END
  END FREEZE_PMOS[11]
  PIN FREEZE_PMOS[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5761.625 187.44 5761.905 188.44 ;
    END
  END FREEZE_PMOS[10]
  PIN FREEZE_PMOS[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5679.865 187.44 5680.145 188.44 ;
    END
  END FREEZE_PMOS[9]
  PIN FREEZE_PMOS[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5614.345 187.44 5614.625 188.44 ;
    END
  END FREEZE_PMOS[8]
  PIN FREEZE_PMOS[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5532.025 187.44 5532.305 188.44 ;
    END
  END FREEZE_PMOS[7]
  PIN FREEZE_PMOS[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5452.505 187.44 5452.785 188.44 ;
    END
  END FREEZE_PMOS[6]
  PIN FREEZE_PMOS[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5375.785 187.44 5376.065 188.44 ;
    END
  END FREEZE_PMOS[5]
  PIN FREEZE_PMOS[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5305.785 187.44 5306.065 188.44 ;
    END
  END FREEZE_PMOS[4]
  PIN FREEZE_PMOS[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5201.625 187.44 5201.905 188.44 ;
    END
  END FREEZE_PMOS[3]
  PIN FREEZE_PMOS[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5119.865 187.44 5120.145 188.44 ;
    END
  END FREEZE_PMOS[2]
  PIN FREEZE_PMOS[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5054.345 187.44 5054.625 188.44 ;
    END
  END FREEZE_PMOS[1]
  PIN FREEZE_PMOS[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4972.025 187.44 4972.305 188.44 ;
    END
  END FREEZE_PMOS[0]
  PIN INJ_IN[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13920.265 187.44 13920.545 188.44 ;
    END
  END INJ_IN[336]
  PIN INJ_IN[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13935.945 187.44 13936.225 188.44 ;
    END
  END INJ_IN[337]
  PIN INJ_IN[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14010.985 187.44 14011.265 188.44 ;
    END
  END INJ_IN[338]
  PIN INJ_IN[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14018.265 187.44 14018.545 188.44 ;
    END
  END INJ_IN[339]
  PIN INJ_IN[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14076.505 187.44 14076.785 188.44 ;
    END
  END INJ_IN[340]
  PIN INJ_IN[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14122.985 187.44 14123.265 188.44 ;
    END
  END INJ_IN[341]
  PIN INJ_IN[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14158.265 187.44 14158.545 188.44 ;
    END
  END INJ_IN[342]
  PIN INJ_IN[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14191.025 187.44 14191.305 188.44 ;
    END
  END INJ_IN[343]
  PIN INJ_IN[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14262.425 187.44 14262.705 188.44 ;
    END
  END INJ_IN[344]
  PIN INJ_IN[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14269.705 187.44 14269.985 188.44 ;
    END
  END INJ_IN[345]
  PIN INJ_IN[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14330.465 187.44 14330.745 188.44 ;
    END
  END INJ_IN[346]
  PIN Read_COMP[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13851.945 187.44 13852.225 188.44 ;
    END
  END Read_COMP[55]
  PIN Read_COMP[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13775.225 187.44 13775.505 188.44 ;
    END
  END Read_COMP[54]
  PIN Read_COMP[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13705.225 187.44 13705.505 188.44 ;
    END
  END Read_COMP[53]
  PIN Read_COMP[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13601.065 187.44 13601.345 188.44 ;
    END
  END Read_COMP[52]
  PIN Read_COMP[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13519.305 187.44 13519.585 188.44 ;
    END
  END Read_COMP[51]
  PIN Read_COMP[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13453.785 187.44 13454.065 188.44 ;
    END
  END Read_COMP[50]
  PIN Read_COMP[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13371.465 187.44 13371.745 188.44 ;
    END
  END Read_COMP[49]
  PIN Read_COMP[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13291.945 187.44 13292.225 188.44 ;
    END
  END Read_COMP[48]
  PIN Read_COMP[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13215.225 187.44 13215.505 188.44 ;
    END
  END Read_COMP[47]
  PIN Read_COMP[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13145.225 187.44 13145.505 188.44 ;
    END
  END Read_COMP[46]
  PIN Read_COMP[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13041.065 187.44 13041.345 188.44 ;
    END
  END Read_COMP[45]
  PIN Read_COMP[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12959.305 187.44 12959.585 188.44 ;
    END
  END Read_COMP[44]
  PIN Read_COMP[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12893.785 187.44 12894.065 188.44 ;
    END
  END Read_COMP[43]
  PIN Read_COMP[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12811.465 187.44 12811.745 188.44 ;
    END
  END Read_COMP[42]
  PIN Read_COMP[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12731.945 187.44 12732.225 188.44 ;
    END
  END Read_COMP[41]
  PIN Read_COMP[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12655.225 187.44 12655.505 188.44 ;
    END
  END Read_COMP[40]
  PIN Read_COMP[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12585.225 187.44 12585.505 188.44 ;
    END
  END Read_COMP[39]
  PIN Read_COMP[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12481.065 187.44 12481.345 188.44 ;
    END
  END Read_COMP[38]
  PIN Read_COMP[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12399.305 187.44 12399.585 188.44 ;
    END
  END Read_COMP[37]
  PIN Read_COMP[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12333.785 187.44 12334.065 188.44 ;
    END
  END Read_COMP[36]
  PIN Read_COMP[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12251.465 187.44 12251.745 188.44 ;
    END
  END Read_COMP[35]
  PIN Read_COMP[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12171.945 187.44 12172.225 188.44 ;
    END
  END Read_COMP[34]
  PIN Read_COMP[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12095.225 187.44 12095.505 188.44 ;
    END
  END Read_COMP[33]
  PIN Read_COMP[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12025.225 187.44 12025.505 188.44 ;
    END
  END Read_COMP[32]
  PIN Read_COMP[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11921.065 187.44 11921.345 188.44 ;
    END
  END Read_COMP[31]
  PIN Read_COMP[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11839.305 187.44 11839.585 188.44 ;
    END
  END Read_COMP[30]
  PIN Read_COMP[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11773.785 187.44 11774.065 188.44 ;
    END
  END Read_COMP[29]
  PIN Read_COMP[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11691.465 187.44 11691.745 188.44 ;
    END
  END Read_COMP[28]
  PIN Read_COMP[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11611.945 187.44 11612.225 188.44 ;
    END
  END Read_COMP[27]
  PIN Read_COMP[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11535.225 187.44 11535.505 188.44 ;
    END
  END Read_COMP[26]
  PIN Read_COMP[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11465.225 187.44 11465.505 188.44 ;
    END
  END Read_COMP[25]
  PIN Read_COMP[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11361.065 187.44 11361.345 188.44 ;
    END
  END Read_COMP[24]
  PIN Read_COMP[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11279.305 187.44 11279.585 188.44 ;
    END
  END Read_COMP[23]
  PIN Read_COMP[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11213.785 187.44 11214.065 188.44 ;
    END
  END Read_COMP[22]
  PIN Read_COMP[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11131.465 187.44 11131.745 188.44 ;
    END
  END Read_COMP[21]
  PIN Read_COMP[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11051.945 187.44 11052.225 188.44 ;
    END
  END Read_COMP[20]
  PIN Read_COMP[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10975.225 187.44 10975.505 188.44 ;
    END
  END Read_COMP[19]
  PIN Read_COMP[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10905.225 187.44 10905.505 188.44 ;
    END
  END Read_COMP[18]
  PIN Read_COMP[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10801.065 187.44 10801.345 188.44 ;
    END
  END Read_COMP[17]
  PIN Read_COMP[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10719.305 187.44 10719.585 188.44 ;
    END
  END Read_COMP[16]
  PIN Read_COMP[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10653.785 187.44 10654.065 188.44 ;
    END
  END Read_COMP[15]
  PIN Read_COMP[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10571.465 187.44 10571.745 188.44 ;
    END
  END Read_COMP[14]
  PIN Read_COMP[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10491.945 187.44 10492.225 188.44 ;
    END
  END Read_COMP[13]
  PIN Read_COMP[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10415.225 187.44 10415.505 188.44 ;
    END
  END Read_COMP[12]
  PIN Read_COMP[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10345.225 187.44 10345.505 188.44 ;
    END
  END Read_COMP[11]
  PIN Read_COMP[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10241.065 187.44 10241.345 188.44 ;
    END
  END Read_COMP[10]
  PIN Read_COMP[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10159.305 187.44 10159.585 188.44 ;
    END
  END Read_COMP[9]
  PIN Read_COMP[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10093.785 187.44 10094.065 188.44 ;
    END
  END Read_COMP[8]
  PIN Read_COMP[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10011.465 187.44 10011.745 188.44 ;
    END
  END Read_COMP[7]
  PIN Read_COMP[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9931.945 187.44 9932.225 188.44 ;
    END
  END Read_COMP[6]
  PIN Read_COMP[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9855.225 187.44 9855.505 188.44 ;
    END
  END Read_COMP[5]
  PIN Read_COMP[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9785.225 187.44 9785.505 188.44 ;
    END
  END Read_COMP[4]
  PIN Read_COMP[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9681.065 187.44 9681.345 188.44 ;
    END
  END Read_COMP[3]
  PIN Read_COMP[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9599.305 187.44 9599.585 188.44 ;
    END
  END Read_COMP[2]
  PIN Read_COMP[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9533.785 187.44 9534.065 188.44 ;
    END
  END Read_COMP[1]
  PIN Read_COMP[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9451.465 187.44 9451.745 188.44 ;
    END
  END Read_COMP[0]
  PIN INJ_IN[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14339.705 187.44 14339.985 188.44 ;
    END
  END INJ_IN[347]
  PIN INJ_IN[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14409.145 187.44 14409.425 188.44 ;
    END
  END INJ_IN[348]
  PIN INJ_IN[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14429.865 187.44 14430.145 188.44 ;
    END
  END INJ_IN[349]
  PIN INJ_IN[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14480.265 187.44 14480.545 188.44 ;
    END
  END INJ_IN[350]
  PIN INJ_IN[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14495.945 187.44 14496.225 188.44 ;
    END
  END INJ_IN[351]
  PIN INJ_IN[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14570.985 187.44 14571.265 188.44 ;
    END
  END INJ_IN[352]
  PIN INJ_IN[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14578.265 187.44 14578.545 188.44 ;
    END
  END INJ_IN[353]
  PIN INJ_IN[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14636.505 187.44 14636.785 188.44 ;
    END
  END INJ_IN[354]
  PIN INJ_IN[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14682.985 187.44 14683.265 188.44 ;
    END
  END INJ_IN[355]
  PIN INJ_IN[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14718.265 187.44 14718.545 188.44 ;
    END
  END INJ_IN[356]
  PIN INJ_IN[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14751.025 187.44 14751.305 188.44 ;
    END
  END INJ_IN[357]
  PIN INJ_IN[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14822.425 187.44 14822.705 188.44 ;
    END
  END INJ_IN[358]
  PIN INJ_IN[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14829.705 187.44 14829.985 188.44 ;
    END
  END INJ_IN[359]
  PIN INJ_IN[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14890.465 187.44 14890.745 188.44 ;
    END
  END INJ_IN[360]
  PIN INJ_IN[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14899.705 187.44 14899.985 188.44 ;
    END
  END INJ_IN[361]
  PIN INJ_IN[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14969.145 187.44 14969.425 188.44 ;
    END
  END INJ_IN[362]
  PIN INJ_IN[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14989.865 187.44 14990.145 188.44 ;
    END
  END INJ_IN[363]
  PIN INJ_IN[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15040.265 187.44 15040.545 188.44 ;
    END
  END INJ_IN[364]
  PIN INJ_IN[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15055.945 187.44 15056.225 188.44 ;
    END
  END INJ_IN[365]
  PIN INJ_IN[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15130.985 187.44 15131.265 188.44 ;
    END
  END INJ_IN[366]
  PIN INJ_IN[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15138.265 187.44 15138.545 188.44 ;
    END
  END INJ_IN[367]
  PIN INJ_IN[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15196.505 187.44 15196.785 188.44 ;
    END
  END INJ_IN[368]
  PIN INJ_IN[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15242.985 187.44 15243.265 188.44 ;
    END
  END INJ_IN[369]
  PIN INJ_IN[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15278.265 187.44 15278.545 188.44 ;
    END
  END INJ_IN[370]
  PIN INJ_IN[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15311.025 187.44 15311.305 188.44 ;
    END
  END INJ_IN[371]
  PIN INJ_IN[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15382.425 187.44 15382.705 188.44 ;
    END
  END INJ_IN[372]
  PIN INJ_IN[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15389.705 187.44 15389.985 188.44 ;
    END
  END INJ_IN[373]
  PIN INJ_IN[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15450.465 187.44 15450.745 188.44 ;
    END
  END INJ_IN[374]
  PIN INJ_IN[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15459.705 187.44 15459.985 188.44 ;
    END
  END INJ_IN[375]
  PIN INJ_IN[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15529.145 187.44 15529.425 188.44 ;
    END
  END INJ_IN[376]
  PIN INJ_IN[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15549.865 187.44 15550.145 188.44 ;
    END
  END INJ_IN[377]
  PIN INJ_IN[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15600.265 187.44 15600.545 188.44 ;
    END
  END INJ_IN[378]
  PIN INJ_IN[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15615.945 187.44 15616.225 188.44 ;
    END
  END INJ_IN[379]
  PIN INJ_IN[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15690.985 187.44 15691.265 188.44 ;
    END
  END INJ_IN[380]
  PIN INJ_IN[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15698.265 187.44 15698.545 188.44 ;
    END
  END INJ_IN[381]
  PIN INJ_IN[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15756.505 187.44 15756.785 188.44 ;
    END
  END INJ_IN[382]
  PIN INJ_IN[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15802.985 187.44 15803.265 188.44 ;
    END
  END INJ_IN[383]
  PIN INJ_IN[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15838.265 187.44 15838.545 188.44 ;
    END
  END INJ_IN[384]
  PIN INJ_IN[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15871.025 187.44 15871.305 188.44 ;
    END
  END INJ_IN[385]
  PIN INJ_IN[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15942.425 187.44 15942.705 188.44 ;
    END
  END INJ_IN[386]
  PIN INJ_IN[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15949.705 187.44 15949.985 188.44 ;
    END
  END INJ_IN[387]
  PIN INJ_IN[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16010.465 187.44 16010.745 188.44 ;
    END
  END INJ_IN[388]
  PIN INJ_IN[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16019.705 187.44 16019.985 188.44 ;
    END
  END INJ_IN[389]
  PIN INJ_IN[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16089.145 187.44 16089.425 188.44 ;
    END
  END INJ_IN[390]
  PIN INJ_IN[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16109.865 187.44 16110.145 188.44 ;
    END
  END INJ_IN[391]
  PIN INJ_IN[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16160.265 187.44 16160.545 188.44 ;
    END
  END INJ_IN[392]
  PIN INJ_IN[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16175.945 187.44 16176.225 188.44 ;
    END
  END INJ_IN[393]
  PIN INJ_IN[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16250.985 187.44 16251.265 188.44 ;
    END
  END INJ_IN[394]
  PIN INJ_IN[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16258.265 187.44 16258.545 188.44 ;
    END
  END INJ_IN[395]
  PIN INJ_IN[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16316.505 187.44 16316.785 188.44 ;
    END
  END INJ_IN[396]
  PIN INJ_IN[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16362.985 187.44 16363.265 188.44 ;
    END
  END INJ_IN[397]
  PIN INJ_IN[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16398.265 187.44 16398.545 188.44 ;
    END
  END INJ_IN[398]
  PIN INJ_IN[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16431.025 187.44 16431.305 188.44 ;
    END
  END INJ_IN[399]
  PIN INJ_IN[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16502.425 187.44 16502.705 188.44 ;
    END
  END INJ_IN[400]
  PIN INJ_IN[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16509.705 187.44 16509.985 188.44 ;
    END
  END INJ_IN[401]
  PIN INJ_IN[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16570.465 187.44 16570.745 188.44 ;
    END
  END INJ_IN[402]
  PIN INJ_IN[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16579.705 187.44 16579.985 188.44 ;
    END
  END INJ_IN[403]
  PIN FREEZE_COMP[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13852.505 187.44 13852.785 188.44 ;
    END
  END FREEZE_COMP[55]
  PIN FREEZE_COMP[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13775.785 187.44 13776.065 188.44 ;
    END
  END FREEZE_COMP[54]
  PIN FREEZE_COMP[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13705.785 187.44 13706.065 188.44 ;
    END
  END FREEZE_COMP[53]
  PIN FREEZE_COMP[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13601.625 187.44 13601.905 188.44 ;
    END
  END FREEZE_COMP[52]
  PIN FREEZE_COMP[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13519.865 187.44 13520.145 188.44 ;
    END
  END FREEZE_COMP[51]
  PIN FREEZE_COMP[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13454.345 187.44 13454.625 188.44 ;
    END
  END FREEZE_COMP[50]
  PIN FREEZE_COMP[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13372.025 187.44 13372.305 188.44 ;
    END
  END FREEZE_COMP[49]
  PIN FREEZE_COMP[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13292.505 187.44 13292.785 188.44 ;
    END
  END FREEZE_COMP[48]
  PIN FREEZE_COMP[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13215.785 187.44 13216.065 188.44 ;
    END
  END FREEZE_COMP[47]
  PIN FREEZE_COMP[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13145.785 187.44 13146.065 188.44 ;
    END
  END FREEZE_COMP[46]
  PIN FREEZE_COMP[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13041.625 187.44 13041.905 188.44 ;
    END
  END FREEZE_COMP[45]
  PIN FREEZE_COMP[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12959.865 187.44 12960.145 188.44 ;
    END
  END FREEZE_COMP[44]
  PIN FREEZE_COMP[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12894.345 187.44 12894.625 188.44 ;
    END
  END FREEZE_COMP[43]
  PIN FREEZE_COMP[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12812.025 187.44 12812.305 188.44 ;
    END
  END FREEZE_COMP[42]
  PIN FREEZE_COMP[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12732.505 187.44 12732.785 188.44 ;
    END
  END FREEZE_COMP[41]
  PIN FREEZE_COMP[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12655.785 187.44 12656.065 188.44 ;
    END
  END FREEZE_COMP[40]
  PIN FREEZE_COMP[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12585.785 187.44 12586.065 188.44 ;
    END
  END FREEZE_COMP[39]
  PIN FREEZE_COMP[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12481.625 187.44 12481.905 188.44 ;
    END
  END FREEZE_COMP[38]
  PIN FREEZE_COMP[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12399.865 187.44 12400.145 188.44 ;
    END
  END FREEZE_COMP[37]
  PIN FREEZE_COMP[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12334.345 187.44 12334.625 188.44 ;
    END
  END FREEZE_COMP[36]
  PIN FREEZE_COMP[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12252.025 187.44 12252.305 188.44 ;
    END
  END FREEZE_COMP[35]
  PIN FREEZE_COMP[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12172.505 187.44 12172.785 188.44 ;
    END
  END FREEZE_COMP[34]
  PIN FREEZE_COMP[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12095.785 187.44 12096.065 188.44 ;
    END
  END FREEZE_COMP[33]
  PIN FREEZE_COMP[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12025.785 187.44 12026.065 188.44 ;
    END
  END FREEZE_COMP[32]
  PIN FREEZE_COMP[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11921.625 187.44 11921.905 188.44 ;
    END
  END FREEZE_COMP[31]
  PIN FREEZE_COMP[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11839.865 187.44 11840.145 188.44 ;
    END
  END FREEZE_COMP[30]
  PIN FREEZE_COMP[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11774.345 187.44 11774.625 188.44 ;
    END
  END FREEZE_COMP[29]
  PIN FREEZE_COMP[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11692.025 187.44 11692.305 188.44 ;
    END
  END FREEZE_COMP[28]
  PIN FREEZE_COMP[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11612.505 187.44 11612.785 188.44 ;
    END
  END FREEZE_COMP[27]
  PIN FREEZE_COMP[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11535.785 187.44 11536.065 188.44 ;
    END
  END FREEZE_COMP[26]
  PIN FREEZE_COMP[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11465.785 187.44 11466.065 188.44 ;
    END
  END FREEZE_COMP[25]
  PIN FREEZE_COMP[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11361.625 187.44 11361.905 188.44 ;
    END
  END FREEZE_COMP[24]
  PIN FREEZE_COMP[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11279.865 187.44 11280.145 188.44 ;
    END
  END FREEZE_COMP[23]
  PIN FREEZE_COMP[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11214.345 187.44 11214.625 188.44 ;
    END
  END FREEZE_COMP[22]
  PIN FREEZE_COMP[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11132.025 187.44 11132.305 188.44 ;
    END
  END FREEZE_COMP[21]
  PIN FREEZE_COMP[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11052.505 187.44 11052.785 188.44 ;
    END
  END FREEZE_COMP[20]
  PIN FREEZE_COMP[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10975.785 187.44 10976.065 188.44 ;
    END
  END FREEZE_COMP[19]
  PIN FREEZE_COMP[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10905.785 187.44 10906.065 188.44 ;
    END
  END FREEZE_COMP[18]
  PIN FREEZE_COMP[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10801.625 187.44 10801.905 188.44 ;
    END
  END FREEZE_COMP[17]
  PIN FREEZE_COMP[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10719.865 187.44 10720.145 188.44 ;
    END
  END FREEZE_COMP[16]
  PIN FREEZE_COMP[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10654.345 187.44 10654.625 188.44 ;
    END
  END FREEZE_COMP[15]
  PIN FREEZE_COMP[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10572.025 187.44 10572.305 188.44 ;
    END
  END FREEZE_COMP[14]
  PIN FREEZE_COMP[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10492.505 187.44 10492.785 188.44 ;
    END
  END FREEZE_COMP[13]
  PIN FREEZE_COMP[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10415.785 187.44 10416.065 188.44 ;
    END
  END FREEZE_COMP[12]
  PIN FREEZE_COMP[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10345.785 187.44 10346.065 188.44 ;
    END
  END FREEZE_COMP[11]
  PIN FREEZE_COMP[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10241.625 187.44 10241.905 188.44 ;
    END
  END FREEZE_COMP[10]
  PIN FREEZE_COMP[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10159.865 187.44 10160.145 188.44 ;
    END
  END FREEZE_COMP[9]
  PIN FREEZE_COMP[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10094.345 187.44 10094.625 188.44 ;
    END
  END FREEZE_COMP[8]
  PIN FREEZE_COMP[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10012.025 187.44 10012.305 188.44 ;
    END
  END FREEZE_COMP[7]
  PIN FREEZE_COMP[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9932.505 187.44 9932.785 188.44 ;
    END
  END FREEZE_COMP[6]
  PIN FREEZE_COMP[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9855.785 187.44 9856.065 188.44 ;
    END
  END FREEZE_COMP[5]
  PIN FREEZE_COMP[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9785.785 187.44 9786.065 188.44 ;
    END
  END FREEZE_COMP[4]
  PIN FREEZE_COMP[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9681.625 187.44 9681.905 188.44 ;
    END
  END FREEZE_COMP[3]
  PIN FREEZE_COMP[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9599.865 187.44 9600.145 188.44 ;
    END
  END FREEZE_COMP[2]
  PIN FREEZE_COMP[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9534.345 187.44 9534.625 188.44 ;
    END
  END FREEZE_COMP[1]
  PIN FREEZE_COMP[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9452.025 187.44 9452.305 188.44 ;
    END
  END FREEZE_COMP[0]
  PIN INJ_IN[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16649.145 187.44 16649.425 188.44 ;
    END
  END INJ_IN[404]
  PIN INJ_IN[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16669.865 187.44 16670.145 188.44 ;
    END
  END INJ_IN[405]
  PIN INJ_IN[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16720.265 187.44 16720.545 188.44 ;
    END
  END INJ_IN[406]
  PIN INJ_IN[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16735.945 187.44 16736.225 188.44 ;
    END
  END INJ_IN[407]
  PIN INJ_IN[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16810.985 187.44 16811.265 188.44 ;
    END
  END INJ_IN[408]
  PIN INJ_IN[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16818.265 187.44 16818.545 188.44 ;
    END
  END INJ_IN[409]
  PIN INJ_IN[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16876.505 187.44 16876.785 188.44 ;
    END
  END INJ_IN[410]
  PIN INJ_IN[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16922.985 187.44 16923.265 188.44 ;
    END
  END INJ_IN[411]
  PIN INJ_IN[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16958.265 187.44 16958.545 188.44 ;
    END
  END INJ_IN[412]
  PIN INJ_IN[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16991.025 187.44 16991.305 188.44 ;
    END
  END INJ_IN[413]
  PIN INJ_IN[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17062.425 187.44 17062.705 188.44 ;
    END
  END INJ_IN[414]
  PIN INJ_IN[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17069.705 187.44 17069.985 188.44 ;
    END
  END INJ_IN[415]
  PIN INJ_IN[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17130.465 187.44 17130.745 188.44 ;
    END
  END INJ_IN[416]
  PIN INJ_IN[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17139.705 187.44 17139.985 188.44 ;
    END
  END INJ_IN[417]
  PIN INJ_IN[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17209.145 187.44 17209.425 188.44 ;
    END
  END INJ_IN[418]
  PIN INJ_IN[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17229.865 187.44 17230.145 188.44 ;
    END
  END INJ_IN[419]
  PIN INJ_IN[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17280.265 187.44 17280.545 188.44 ;
    END
  END INJ_IN[420]
  PIN INJ_IN[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17295.945 187.44 17296.225 188.44 ;
    END
  END INJ_IN[421]
  PIN INJ_IN[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17370.985 187.44 17371.265 188.44 ;
    END
  END INJ_IN[422]
  PIN INJ_IN[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17378.265 187.44 17378.545 188.44 ;
    END
  END INJ_IN[423]
  PIN INJ_IN[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17436.505 187.44 17436.785 188.44 ;
    END
  END INJ_IN[424]
  PIN INJ_IN[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17482.985 187.44 17483.265 188.44 ;
    END
  END INJ_IN[425]
  PIN INJ_IN[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17518.265 187.44 17518.545 188.44 ;
    END
  END INJ_IN[426]
  PIN INJ_IN[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17551.025 187.44 17551.305 188.44 ;
    END
  END INJ_IN[427]
  PIN INJ_IN[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17622.425 187.44 17622.705 188.44 ;
    END
  END INJ_IN[428]
  PIN INJ_IN[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17629.705 187.44 17629.985 188.44 ;
    END
  END INJ_IN[429]
  PIN INJ_IN[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17690.465 187.44 17690.745 188.44 ;
    END
  END INJ_IN[430]
  PIN INJ_IN[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17699.705 187.44 17699.985 188.44 ;
    END
  END INJ_IN[431]
  PIN INJ_IN[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17769.145 187.44 17769.425 188.44 ;
    END
  END INJ_IN[432]
  PIN INJ_IN[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17789.865 187.44 17790.145 188.44 ;
    END
  END INJ_IN[433]
  PIN INJ_IN[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17840.265 187.44 17840.545 188.44 ;
    END
  END INJ_IN[434]
  PIN INJ_IN[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17855.945 187.44 17856.225 188.44 ;
    END
  END INJ_IN[435]
  PIN INJ_IN[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17930.985 187.44 17931.265 188.44 ;
    END
  END INJ_IN[436]
  PIN INJ_IN[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17938.265 187.44 17938.545 188.44 ;
    END
  END INJ_IN[437]
  PIN INJ_IN[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17996.505 187.44 17996.785 188.44 ;
    END
  END INJ_IN[438]
  PIN INJ_IN[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18042.985 187.44 18043.265 188.44 ;
    END
  END INJ_IN[439]
  PIN INJ_IN[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18078.265 187.44 18078.545 188.44 ;
    END
  END INJ_IN[440]
  PIN INJ_IN[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18111.025 187.44 18111.305 188.44 ;
    END
  END INJ_IN[441]
  PIN INJ_IN[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18182.425 187.44 18182.705 188.44 ;
    END
  END INJ_IN[442]
  PIN INJ_IN[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18189.705 187.44 18189.985 188.44 ;
    END
  END INJ_IN[443]
  PIN INJ_IN[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18250.465 187.44 18250.745 188.44 ;
    END
  END INJ_IN[444]
  PIN INJ_IN[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18259.705 187.44 18259.985 188.44 ;
    END
  END INJ_IN[445]
  PIN INJ_IN[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18329.145 187.44 18329.425 188.44 ;
    END
  END INJ_IN[446]
  PIN INJ_IN[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18349.865 187.44 18350.145 188.44 ;
    END
  END INJ_IN[447]
  PIN Read_HV[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18331.945 187.44 18332.225 188.44 ;
    END
  END Read_HV[55]
  PIN Read_HV[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18255.225 187.44 18255.505 188.44 ;
    END
  END Read_HV[54]
  PIN Read_HV[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18185.225 187.44 18185.505 188.44 ;
    END
  END Read_HV[53]
  PIN Read_HV[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18081.065 187.44 18081.345 188.44 ;
    END
  END Read_HV[52]
  PIN Read_HV[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17999.305 187.44 17999.585 188.44 ;
    END
  END Read_HV[51]
  PIN Read_HV[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17933.785 187.44 17934.065 188.44 ;
    END
  END Read_HV[50]
  PIN Read_HV[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17851.465 187.44 17851.745 188.44 ;
    END
  END Read_HV[49]
  PIN Read_HV[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17771.945 187.44 17772.225 188.44 ;
    END
  END Read_HV[48]
  PIN Read_HV[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17695.225 187.44 17695.505 188.44 ;
    END
  END Read_HV[47]
  PIN Read_HV[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17625.225 187.44 17625.505 188.44 ;
    END
  END Read_HV[46]
  PIN Read_HV[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17521.065 187.44 17521.345 188.44 ;
    END
  END Read_HV[45]
  PIN Read_HV[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17439.305 187.44 17439.585 188.44 ;
    END
  END Read_HV[44]
  PIN Read_HV[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17373.785 187.44 17374.065 188.44 ;
    END
  END Read_HV[43]
  PIN Read_HV[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17291.465 187.44 17291.745 188.44 ;
    END
  END Read_HV[42]
  PIN Read_HV[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17211.945 187.44 17212.225 188.44 ;
    END
  END Read_HV[41]
  PIN Read_HV[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17135.225 187.44 17135.505 188.44 ;
    END
  END Read_HV[40]
  PIN Read_HV[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17065.225 187.44 17065.505 188.44 ;
    END
  END Read_HV[39]
  PIN Read_HV[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16961.065 187.44 16961.345 188.44 ;
    END
  END Read_HV[38]
  PIN Read_HV[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16879.305 187.44 16879.585 188.44 ;
    END
  END Read_HV[37]
  PIN Read_HV[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16813.785 187.44 16814.065 188.44 ;
    END
  END Read_HV[36]
  PIN Read_HV[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16731.465 187.44 16731.745 188.44 ;
    END
  END Read_HV[35]
  PIN Read_HV[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16651.945 187.44 16652.225 188.44 ;
    END
  END Read_HV[34]
  PIN Read_HV[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16575.225 187.44 16575.505 188.44 ;
    END
  END Read_HV[33]
  PIN Read_HV[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16505.225 187.44 16505.505 188.44 ;
    END
  END Read_HV[32]
  PIN Read_HV[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16401.065 187.44 16401.345 188.44 ;
    END
  END Read_HV[31]
  PIN Read_HV[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16319.305 187.44 16319.585 188.44 ;
    END
  END Read_HV[30]
  PIN Read_HV[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16253.785 187.44 16254.065 188.44 ;
    END
  END Read_HV[29]
  PIN Read_HV[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16171.465 187.44 16171.745 188.44 ;
    END
  END Read_HV[28]
  PIN Read_HV[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16091.945 187.44 16092.225 188.44 ;
    END
  END Read_HV[27]
  PIN Read_HV[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16015.225 187.44 16015.505 188.44 ;
    END
  END Read_HV[26]
  PIN Read_HV[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15945.225 187.44 15945.505 188.44 ;
    END
  END Read_HV[25]
  PIN Read_HV[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15841.065 187.44 15841.345 188.44 ;
    END
  END Read_HV[24]
  PIN Read_HV[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15759.305 187.44 15759.585 188.44 ;
    END
  END Read_HV[23]
  PIN Read_HV[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15693.785 187.44 15694.065 188.44 ;
    END
  END Read_HV[22]
  PIN Read_HV[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15611.465 187.44 15611.745 188.44 ;
    END
  END Read_HV[21]
  PIN Read_HV[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15531.945 187.44 15532.225 188.44 ;
    END
  END Read_HV[20]
  PIN Read_HV[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15455.225 187.44 15455.505 188.44 ;
    END
  END Read_HV[19]
  PIN Read_HV[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15385.225 187.44 15385.505 188.44 ;
    END
  END Read_HV[18]
  PIN Read_HV[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15281.065 187.44 15281.345 188.44 ;
    END
  END Read_HV[17]
  PIN Read_HV[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15199.305 187.44 15199.585 188.44 ;
    END
  END Read_HV[16]
  PIN Read_HV[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15133.785 187.44 15134.065 188.44 ;
    END
  END Read_HV[15]
  PIN Read_HV[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15051.465 187.44 15051.745 188.44 ;
    END
  END Read_HV[14]
  PIN Read_HV[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14971.945 187.44 14972.225 188.44 ;
    END
  END Read_HV[13]
  PIN Read_HV[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14895.225 187.44 14895.505 188.44 ;
    END
  END Read_HV[12]
  PIN Read_HV[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14825.225 187.44 14825.505 188.44 ;
    END
  END Read_HV[11]
  PIN Read_HV[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14721.065 187.44 14721.345 188.44 ;
    END
  END Read_HV[10]
  PIN Read_HV[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14639.305 187.44 14639.585 188.44 ;
    END
  END Read_HV[9]
  PIN Read_HV[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14573.785 187.44 14574.065 188.44 ;
    END
  END Read_HV[8]
  PIN Read_HV[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14491.465 187.44 14491.745 188.44 ;
    END
  END Read_HV[7]
  PIN Read_HV[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14411.945 187.44 14412.225 188.44 ;
    END
  END Read_HV[6]
  PIN Read_HV[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14335.225 187.44 14335.505 188.44 ;
    END
  END Read_HV[5]
  PIN Read_HV[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14265.225 187.44 14265.505 188.44 ;
    END
  END Read_HV[4]
  PIN Read_HV[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14161.065 187.44 14161.345 188.44 ;
    END
  END Read_HV[3]
  PIN Read_HV[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14079.305 187.44 14079.585 188.44 ;
    END
  END Read_HV[2]
  PIN Read_HV[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14013.785 187.44 14014.065 188.44 ;
    END
  END Read_HV[1]
  PIN Read_HV[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13931.465 187.44 13931.745 188.44 ;
    END
  END Read_HV[0]
  PIN FREEZE_HV[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18332.505 187.44 18332.785 188.44 ;
    END
  END FREEZE_HV[55]
  PIN FREEZE_HV[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18255.785 187.44 18256.065 188.44 ;
    END
  END FREEZE_HV[54]
  PIN FREEZE_HV[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18185.785 187.44 18186.065 188.44 ;
    END
  END FREEZE_HV[53]
  PIN FREEZE_HV[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18081.625 187.44 18081.905 188.44 ;
    END
  END FREEZE_HV[52]
  PIN FREEZE_HV[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17999.865 187.44 18000.145 188.44 ;
    END
  END FREEZE_HV[51]
  PIN FREEZE_HV[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17934.345 187.44 17934.625 188.44 ;
    END
  END FREEZE_HV[50]
  PIN FREEZE_HV[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17852.025 187.44 17852.305 188.44 ;
    END
  END FREEZE_HV[49]
  PIN FREEZE_HV[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17772.505 187.44 17772.785 188.44 ;
    END
  END FREEZE_HV[48]
  PIN FREEZE_HV[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17695.785 187.44 17696.065 188.44 ;
    END
  END FREEZE_HV[47]
  PIN FREEZE_HV[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17625.785 187.44 17626.065 188.44 ;
    END
  END FREEZE_HV[46]
  PIN FREEZE_HV[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17521.625 187.44 17521.905 188.44 ;
    END
  END FREEZE_HV[45]
  PIN FREEZE_HV[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17439.865 187.44 17440.145 188.44 ;
    END
  END FREEZE_HV[44]
  PIN FREEZE_HV[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17374.345 187.44 17374.625 188.44 ;
    END
  END FREEZE_HV[43]
  PIN FREEZE_HV[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17292.025 187.44 17292.305 188.44 ;
    END
  END FREEZE_HV[42]
  PIN FREEZE_HV[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17212.505 187.44 17212.785 188.44 ;
    END
  END FREEZE_HV[41]
  PIN FREEZE_HV[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17135.785 187.44 17136.065 188.44 ;
    END
  END FREEZE_HV[40]
  PIN FREEZE_HV[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17065.785 187.44 17066.065 188.44 ;
    END
  END FREEZE_HV[39]
  PIN FREEZE_HV[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16961.625 187.44 16961.905 188.44 ;
    END
  END FREEZE_HV[38]
  PIN FREEZE_HV[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16879.865 187.44 16880.145 188.44 ;
    END
  END FREEZE_HV[37]
  PIN FREEZE_HV[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16814.345 187.44 16814.625 188.44 ;
    END
  END FREEZE_HV[36]
  PIN FREEZE_HV[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16732.025 187.44 16732.305 188.44 ;
    END
  END FREEZE_HV[35]
  PIN FREEZE_HV[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16652.505 187.44 16652.785 188.44 ;
    END
  END FREEZE_HV[34]
  PIN FREEZE_HV[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16575.785 187.44 16576.065 188.44 ;
    END
  END FREEZE_HV[33]
  PIN FREEZE_HV[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16505.785 187.44 16506.065 188.44 ;
    END
  END FREEZE_HV[32]
  PIN FREEZE_HV[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16401.625 187.44 16401.905 188.44 ;
    END
  END FREEZE_HV[31]
  PIN FREEZE_HV[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16319.865 187.44 16320.145 188.44 ;
    END
  END FREEZE_HV[30]
  PIN FREEZE_HV[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16254.345 187.44 16254.625 188.44 ;
    END
  END FREEZE_HV[29]
  PIN FREEZE_HV[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16172.025 187.44 16172.305 188.44 ;
    END
  END FREEZE_HV[28]
  PIN FREEZE_HV[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16092.505 187.44 16092.785 188.44 ;
    END
  END FREEZE_HV[27]
  PIN FREEZE_HV[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16015.785 187.44 16016.065 188.44 ;
    END
  END FREEZE_HV[26]
  PIN FREEZE_HV[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15945.785 187.44 15946.065 188.44 ;
    END
  END FREEZE_HV[25]
  PIN FREEZE_HV[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15841.625 187.44 15841.905 188.44 ;
    END
  END FREEZE_HV[24]
  PIN FREEZE_HV[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15759.865 187.44 15760.145 188.44 ;
    END
  END FREEZE_HV[23]
  PIN FREEZE_HV[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15694.345 187.44 15694.625 188.44 ;
    END
  END FREEZE_HV[22]
  PIN FREEZE_HV[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15612.025 187.44 15612.305 188.44 ;
    END
  END FREEZE_HV[21]
  PIN FREEZE_HV[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15532.505 187.44 15532.785 188.44 ;
    END
  END FREEZE_HV[20]
  PIN FREEZE_HV[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15455.785 187.44 15456.065 188.44 ;
    END
  END FREEZE_HV[19]
  PIN FREEZE_HV[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15385.785 187.44 15386.065 188.44 ;
    END
  END FREEZE_HV[18]
  PIN FREEZE_HV[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15281.625 187.44 15281.905 188.44 ;
    END
  END FREEZE_HV[17]
  PIN FREEZE_HV[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15199.865 187.44 15200.145 188.44 ;
    END
  END FREEZE_HV[16]
  PIN FREEZE_HV[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15134.345 187.44 15134.625 188.44 ;
    END
  END FREEZE_HV[15]
  PIN FREEZE_HV[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15052.025 187.44 15052.305 188.44 ;
    END
  END FREEZE_HV[14]
  PIN FREEZE_HV[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14972.505 187.44 14972.785 188.44 ;
    END
  END FREEZE_HV[13]
  PIN FREEZE_HV[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14895.785 187.44 14896.065 188.44 ;
    END
  END FREEZE_HV[12]
  PIN FREEZE_HV[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14825.785 187.44 14826.065 188.44 ;
    END
  END FREEZE_HV[11]
  PIN FREEZE_HV[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14721.625 187.44 14721.905 188.44 ;
    END
  END FREEZE_HV[10]
  PIN FREEZE_HV[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14639.865 187.44 14640.145 188.44 ;
    END
  END FREEZE_HV[9]
  PIN FREEZE_HV[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14574.345 187.44 14574.625 188.44 ;
    END
  END FREEZE_HV[8]
  PIN FREEZE_HV[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14492.025 187.44 14492.305 188.44 ;
    END
  END FREEZE_HV[7]
  PIN FREEZE_HV[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14412.505 187.44 14412.785 188.44 ;
    END
  END FREEZE_HV[6]
  PIN FREEZE_HV[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14335.785 187.44 14336.065 188.44 ;
    END
  END FREEZE_HV[5]
  PIN FREEZE_HV[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14265.785 187.44 14266.065 188.44 ;
    END
  END FREEZE_HV[4]
  PIN FREEZE_HV[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14161.625 187.44 14161.905 188.44 ;
    END
  END FREEZE_HV[3]
  PIN FREEZE_HV[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14079.865 187.44 14080.145 188.44 ;
    END
  END FREEZE_HV[2]
  PIN FREEZE_HV[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14014.345 187.44 14014.625 188.44 ;
    END
  END FREEZE_HV[1]
  PIN FREEZE_HV[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13932.025 187.44 13932.305 188.44 ;
    END
  END FREEZE_HV[0]
  PIN DIG_MON_SEL[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18360.505 187.44 18360.785 188.44 ;
    END
  END DIG_MON_SEL[447]
  PIN DIG_MON_SEL[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18279.305 187.44 18279.585 188.44 ;
    END
  END DIG_MON_SEL[446]
  PIN DIG_MON_SEL[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18278.745 187.44 18279.025 188.44 ;
    END
  END DIG_MON_SEL[445]
  PIN DIG_MON_SEL[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18213.785 187.44 18214.065 188.44 ;
    END
  END DIG_MON_SEL[444]
  PIN DIG_MON_SEL[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18213.225 187.44 18213.505 188.44 ;
    END
  END DIG_MON_SEL[443]
  PIN DIG_MON_SEL[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18132.585 187.44 18132.865 188.44 ;
    END
  END DIG_MON_SEL[442]
  PIN DIG_MON_SEL[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18132.025 187.44 18132.305 188.44 ;
    END
  END DIG_MON_SEL[441]
  PIN DIG_MON_SEL[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18054.185 187.44 18054.465 188.44 ;
    END
  END DIG_MON_SEL[440]
  PIN DIG_MON_SEL[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18053.625 187.44 18053.905 188.44 ;
    END
  END DIG_MON_SEL[439]
  PIN DIG_MON_SEL[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17976.905 187.44 17977.185 188.44 ;
    END
  END DIG_MON_SEL[438]
  PIN DIG_MON_SEL[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17976.345 187.44 17976.625 188.44 ;
    END
  END DIG_MON_SEL[437]
  PIN DIG_MON_SEL[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17906.905 187.44 17907.185 188.44 ;
    END
  END DIG_MON_SEL[436]
  PIN DIG_MON_SEL[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17906.345 187.44 17906.625 188.44 ;
    END
  END DIG_MON_SEL[435]
  PIN DIG_MON_SEL[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17827.105 187.44 17827.385 188.44 ;
    END
  END DIG_MON_SEL[434]
  PIN DIG_MON_SEL[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17800.505 187.44 17800.785 188.44 ;
    END
  END DIG_MON_SEL[433]
  PIN DIG_MON_SEL[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17719.305 187.44 17719.585 188.44 ;
    END
  END DIG_MON_SEL[432]
  PIN DIG_MON_SEL[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17718.745 187.44 17719.025 188.44 ;
    END
  END DIG_MON_SEL[431]
  PIN DIG_MON_SEL[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17653.785 187.44 17654.065 188.44 ;
    END
  END DIG_MON_SEL[430]
  PIN DIG_MON_SEL[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17653.225 187.44 17653.505 188.44 ;
    END
  END DIG_MON_SEL[429]
  PIN DIG_MON_SEL[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17572.585 187.44 17572.865 188.44 ;
    END
  END DIG_MON_SEL[428]
  PIN DIG_MON_SEL[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17572.025 187.44 17572.305 188.44 ;
    END
  END DIG_MON_SEL[427]
  PIN DIG_MON_SEL[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17494.185 187.44 17494.465 188.44 ;
    END
  END DIG_MON_SEL[426]
  PIN DIG_MON_SEL[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17493.625 187.44 17493.905 188.44 ;
    END
  END DIG_MON_SEL[425]
  PIN DIG_MON_SEL[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17416.905 187.44 17417.185 188.44 ;
    END
  END DIG_MON_SEL[424]
  PIN DIG_MON_SEL[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17416.345 187.44 17416.625 188.44 ;
    END
  END DIG_MON_SEL[423]
  PIN DIG_MON_SEL[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17346.905 187.44 17347.185 188.44 ;
    END
  END DIG_MON_SEL[422]
  PIN DIG_MON_SEL[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17346.345 187.44 17346.625 188.44 ;
    END
  END DIG_MON_SEL[421]
  PIN DIG_MON_SEL[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17267.105 187.44 17267.385 188.44 ;
    END
  END DIG_MON_SEL[420]
  PIN DIG_MON_SEL[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17240.505 187.44 17240.785 188.44 ;
    END
  END DIG_MON_SEL[419]
  PIN DIG_MON_SEL[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17159.305 187.44 17159.585 188.44 ;
    END
  END DIG_MON_SEL[418]
  PIN DIG_MON_SEL[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17158.745 187.44 17159.025 188.44 ;
    END
  END DIG_MON_SEL[417]
  PIN DIG_MON_SEL[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17093.785 187.44 17094.065 188.44 ;
    END
  END DIG_MON_SEL[416]
  PIN DIG_MON_SEL[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17093.225 187.44 17093.505 188.44 ;
    END
  END DIG_MON_SEL[415]
  PIN DIG_MON_SEL[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17012.585 187.44 17012.865 188.44 ;
    END
  END DIG_MON_SEL[414]
  PIN DIG_MON_SEL[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17012.025 187.44 17012.305 188.44 ;
    END
  END DIG_MON_SEL[413]
  PIN DIG_MON_SEL[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16934.185 187.44 16934.465 188.44 ;
    END
  END DIG_MON_SEL[412]
  PIN DIG_MON_SEL[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16933.625 187.44 16933.905 188.44 ;
    END
  END DIG_MON_SEL[411]
  PIN DIG_MON_SEL[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16856.905 187.44 16857.185 188.44 ;
    END
  END DIG_MON_SEL[410]
  PIN DIG_MON_SEL[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16856.345 187.44 16856.625 188.44 ;
    END
  END DIG_MON_SEL[409]
  PIN DIG_MON_SEL[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16786.905 187.44 16787.185 188.44 ;
    END
  END DIG_MON_SEL[408]
  PIN DIG_MON_SEL[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16786.345 187.44 16786.625 188.44 ;
    END
  END DIG_MON_SEL[407]
  PIN DIG_MON_SEL[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16707.105 187.44 16707.385 188.44 ;
    END
  END DIG_MON_SEL[406]
  PIN DIG_MON_SEL[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16680.505 187.44 16680.785 188.44 ;
    END
  END DIG_MON_SEL[405]
  PIN DIG_MON_SEL[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16599.305 187.44 16599.585 188.44 ;
    END
  END DIG_MON_SEL[404]
  PIN DIG_MON_SEL[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16598.745 187.44 16599.025 188.44 ;
    END
  END DIG_MON_SEL[403]
  PIN DIG_MON_SEL[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16533.785 187.44 16534.065 188.44 ;
    END
  END DIG_MON_SEL[402]
  PIN DIG_MON_SEL[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16533.225 187.44 16533.505 188.44 ;
    END
  END DIG_MON_SEL[401]
  PIN DIG_MON_SEL[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16452.585 187.44 16452.865 188.44 ;
    END
  END DIG_MON_SEL[400]
  PIN DIG_MON_SEL[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16452.025 187.44 16452.305 188.44 ;
    END
  END DIG_MON_SEL[399]
  PIN DIG_MON_SEL[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16374.185 187.44 16374.465 188.44 ;
    END
  END DIG_MON_SEL[398]
  PIN DIG_MON_SEL[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16373.625 187.44 16373.905 188.44 ;
    END
  END DIG_MON_SEL[397]
  PIN DIG_MON_SEL[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16296.905 187.44 16297.185 188.44 ;
    END
  END DIG_MON_SEL[396]
  PIN DIG_MON_SEL[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16296.345 187.44 16296.625 188.44 ;
    END
  END DIG_MON_SEL[395]
  PIN DIG_MON_SEL[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16226.905 187.44 16227.185 188.44 ;
    END
  END DIG_MON_SEL[394]
  PIN DIG_MON_SEL[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16226.345 187.44 16226.625 188.44 ;
    END
  END DIG_MON_SEL[393]
  PIN DIG_MON_SEL[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16147.105 187.44 16147.385 188.44 ;
    END
  END DIG_MON_SEL[392]
  PIN DIG_MON_SEL[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16120.505 187.44 16120.785 188.44 ;
    END
  END DIG_MON_SEL[391]
  PIN DIG_MON_SEL[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16039.305 187.44 16039.585 188.44 ;
    END
  END DIG_MON_SEL[390]
  PIN DIG_MON_SEL[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16038.745 187.44 16039.025 188.44 ;
    END
  END DIG_MON_SEL[389]
  PIN DIG_MON_SEL[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15973.785 187.44 15974.065 188.44 ;
    END
  END DIG_MON_SEL[388]
  PIN DIG_MON_SEL[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15973.225 187.44 15973.505 188.44 ;
    END
  END DIG_MON_SEL[387]
  PIN DIG_MON_SEL[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15892.585 187.44 15892.865 188.44 ;
    END
  END DIG_MON_SEL[386]
  PIN DIG_MON_SEL[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15892.025 187.44 15892.305 188.44 ;
    END
  END DIG_MON_SEL[385]
  PIN DIG_MON_SEL[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15814.185 187.44 15814.465 188.44 ;
    END
  END DIG_MON_SEL[384]
  PIN DIG_MON_SEL[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15813.625 187.44 15813.905 188.44 ;
    END
  END DIG_MON_SEL[383]
  PIN DIG_MON_SEL[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15736.905 187.44 15737.185 188.44 ;
    END
  END DIG_MON_SEL[382]
  PIN DIG_MON_SEL[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15736.345 187.44 15736.625 188.44 ;
    END
  END DIG_MON_SEL[381]
  PIN DIG_MON_SEL[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15666.905 187.44 15667.185 188.44 ;
    END
  END DIG_MON_SEL[380]
  PIN DIG_MON_SEL[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15666.345 187.44 15666.625 188.44 ;
    END
  END DIG_MON_SEL[379]
  PIN DIG_MON_SEL[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15587.105 187.44 15587.385 188.44 ;
    END
  END DIG_MON_SEL[378]
  PIN DIG_MON_SEL[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15560.505 187.44 15560.785 188.44 ;
    END
  END DIG_MON_SEL[377]
  PIN DIG_MON_SEL[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15479.305 187.44 15479.585 188.44 ;
    END
  END DIG_MON_SEL[376]
  PIN DIG_MON_SEL[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15478.745 187.44 15479.025 188.44 ;
    END
  END DIG_MON_SEL[375]
  PIN DIG_MON_SEL[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15413.785 187.44 15414.065 188.44 ;
    END
  END DIG_MON_SEL[374]
  PIN DIG_MON_SEL[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15413.225 187.44 15413.505 188.44 ;
    END
  END DIG_MON_SEL[373]
  PIN DIG_MON_SEL[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15332.585 187.44 15332.865 188.44 ;
    END
  END DIG_MON_SEL[372]
  PIN DIG_MON_SEL[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15332.025 187.44 15332.305 188.44 ;
    END
  END DIG_MON_SEL[371]
  PIN DIG_MON_SEL[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15254.185 187.44 15254.465 188.44 ;
    END
  END DIG_MON_SEL[370]
  PIN DIG_MON_SEL[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15253.625 187.44 15253.905 188.44 ;
    END
  END DIG_MON_SEL[369]
  PIN DIG_MON_SEL[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15176.905 187.44 15177.185 188.44 ;
    END
  END DIG_MON_SEL[368]
  PIN DIG_MON_SEL[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15176.345 187.44 15176.625 188.44 ;
    END
  END DIG_MON_SEL[367]
  PIN DIG_MON_SEL[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15106.905 187.44 15107.185 188.44 ;
    END
  END DIG_MON_SEL[366]
  PIN DIG_MON_SEL[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15106.345 187.44 15106.625 188.44 ;
    END
  END DIG_MON_SEL[365]
  PIN DIG_MON_SEL[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15027.105 187.44 15027.385 188.44 ;
    END
  END DIG_MON_SEL[364]
  PIN DIG_MON_SEL[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15000.505 187.44 15000.785 188.44 ;
    END
  END DIG_MON_SEL[363]
  PIN DIG_MON_SEL[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14919.305 187.44 14919.585 188.44 ;
    END
  END DIG_MON_SEL[362]
  PIN DIG_MON_SEL[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14918.745 187.44 14919.025 188.44 ;
    END
  END DIG_MON_SEL[361]
  PIN DIG_MON_SEL[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14853.785 187.44 14854.065 188.44 ;
    END
  END DIG_MON_SEL[360]
  PIN DIG_MON_SEL[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14853.225 187.44 14853.505 188.44 ;
    END
  END DIG_MON_SEL[359]
  PIN DIG_MON_SEL[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14772.585 187.44 14772.865 188.44 ;
    END
  END DIG_MON_SEL[358]
  PIN DIG_MON_SEL[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14772.025 187.44 14772.305 188.44 ;
    END
  END DIG_MON_SEL[357]
  PIN DIG_MON_SEL[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14694.185 187.44 14694.465 188.44 ;
    END
  END DIG_MON_SEL[356]
  PIN DIG_MON_SEL[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14693.625 187.44 14693.905 188.44 ;
    END
  END DIG_MON_SEL[355]
  PIN DIG_MON_SEL[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14616.905 187.44 14617.185 188.44 ;
    END
  END DIG_MON_SEL[354]
  PIN DIG_MON_SEL[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14616.345 187.44 14616.625 188.44 ;
    END
  END DIG_MON_SEL[353]
  PIN DIG_MON_SEL[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14546.905 187.44 14547.185 188.44 ;
    END
  END DIG_MON_SEL[352]
  PIN DIG_MON_SEL[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14546.345 187.44 14546.625 188.44 ;
    END
  END DIG_MON_SEL[351]
  PIN DIG_MON_SEL[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14467.105 187.44 14467.385 188.44 ;
    END
  END DIG_MON_SEL[350]
  PIN DIG_MON_SEL[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14440.505 187.44 14440.785 188.44 ;
    END
  END DIG_MON_SEL[349]
  PIN DIG_MON_SEL[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14359.305 187.44 14359.585 188.44 ;
    END
  END DIG_MON_SEL[348]
  PIN DIG_MON_SEL[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14358.745 187.44 14359.025 188.44 ;
    END
  END DIG_MON_SEL[347]
  PIN DIG_MON_SEL[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14293.785 187.44 14294.065 188.44 ;
    END
  END DIG_MON_SEL[346]
  PIN DIG_MON_SEL[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14293.225 187.44 14293.505 188.44 ;
    END
  END DIG_MON_SEL[345]
  PIN DIG_MON_SEL[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14212.585 187.44 14212.865 188.44 ;
    END
  END DIG_MON_SEL[344]
  PIN DIG_MON_SEL[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14212.025 187.44 14212.305 188.44 ;
    END
  END DIG_MON_SEL[343]
  PIN DIG_MON_SEL[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14134.185 187.44 14134.465 188.44 ;
    END
  END DIG_MON_SEL[342]
  PIN DIG_MON_SEL[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14133.625 187.44 14133.905 188.44 ;
    END
  END DIG_MON_SEL[341]
  PIN DIG_MON_SEL[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14056.905 187.44 14057.185 188.44 ;
    END
  END DIG_MON_SEL[340]
  PIN DIG_MON_SEL[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14056.345 187.44 14056.625 188.44 ;
    END
  END DIG_MON_SEL[339]
  PIN DIG_MON_SEL[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13986.905 187.44 13987.185 188.44 ;
    END
  END DIG_MON_SEL[338]
  PIN DIG_MON_SEL[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13986.345 187.44 13986.625 188.44 ;
    END
  END DIG_MON_SEL[337]
  PIN DIG_MON_SEL[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13907.105 187.44 13907.385 188.44 ;
    END
  END DIG_MON_SEL[336]
  PIN DIG_MON_SEL[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13880.505 187.44 13880.785 188.44 ;
    END
  END DIG_MON_SEL[335]
  PIN DIG_MON_SEL[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13799.305 187.44 13799.585 188.44 ;
    END
  END DIG_MON_SEL[334]
  PIN DIG_MON_SEL[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13798.745 187.44 13799.025 188.44 ;
    END
  END DIG_MON_SEL[333]
  PIN DIG_MON_SEL[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13733.785 187.44 13734.065 188.44 ;
    END
  END DIG_MON_SEL[332]
  PIN DIG_MON_SEL[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13733.225 187.44 13733.505 188.44 ;
    END
  END DIG_MON_SEL[331]
  PIN DIG_MON_SEL[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13652.585 187.44 13652.865 188.44 ;
    END
  END DIG_MON_SEL[330]
  PIN DIG_MON_SEL[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13652.025 187.44 13652.305 188.44 ;
    END
  END DIG_MON_SEL[329]
  PIN DIG_MON_SEL[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13574.185 187.44 13574.465 188.44 ;
    END
  END DIG_MON_SEL[328]
  PIN DIG_MON_SEL[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13573.625 187.44 13573.905 188.44 ;
    END
  END DIG_MON_SEL[327]
  PIN DIG_MON_SEL[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13496.905 187.44 13497.185 188.44 ;
    END
  END DIG_MON_SEL[326]
  PIN DIG_MON_SEL[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13496.345 187.44 13496.625 188.44 ;
    END
  END DIG_MON_SEL[325]
  PIN DIG_MON_SEL[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13426.905 187.44 13427.185 188.44 ;
    END
  END DIG_MON_SEL[324]
  PIN DIG_MON_SEL[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13426.345 187.44 13426.625 188.44 ;
    END
  END DIG_MON_SEL[323]
  PIN DIG_MON_SEL[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13347.105 187.44 13347.385 188.44 ;
    END
  END DIG_MON_SEL[322]
  PIN DIG_MON_SEL[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13320.505 187.44 13320.785 188.44 ;
    END
  END DIG_MON_SEL[321]
  PIN DIG_MON_SEL[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13239.305 187.44 13239.585 188.44 ;
    END
  END DIG_MON_SEL[320]
  PIN DIG_MON_SEL[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13238.745 187.44 13239.025 188.44 ;
    END
  END DIG_MON_SEL[319]
  PIN DIG_MON_SEL[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13173.785 187.44 13174.065 188.44 ;
    END
  END DIG_MON_SEL[318]
  PIN DIG_MON_SEL[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13173.225 187.44 13173.505 188.44 ;
    END
  END DIG_MON_SEL[317]
  PIN DIG_MON_SEL[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13092.585 187.44 13092.865 188.44 ;
    END
  END DIG_MON_SEL[316]
  PIN DIG_MON_SEL[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13092.025 187.44 13092.305 188.44 ;
    END
  END DIG_MON_SEL[315]
  PIN DIG_MON_SEL[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13014.185 187.44 13014.465 188.44 ;
    END
  END DIG_MON_SEL[314]
  PIN DIG_MON_SEL[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13013.625 187.44 13013.905 188.44 ;
    END
  END DIG_MON_SEL[313]
  PIN DIG_MON_SEL[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12936.905 187.44 12937.185 188.44 ;
    END
  END DIG_MON_SEL[312]
  PIN DIG_MON_SEL[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12936.345 187.44 12936.625 188.44 ;
    END
  END DIG_MON_SEL[311]
  PIN DIG_MON_SEL[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12866.905 187.44 12867.185 188.44 ;
    END
  END DIG_MON_SEL[310]
  PIN DIG_MON_SEL[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12866.345 187.44 12866.625 188.44 ;
    END
  END DIG_MON_SEL[309]
  PIN DIG_MON_SEL[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12787.105 187.44 12787.385 188.44 ;
    END
  END DIG_MON_SEL[308]
  PIN DIG_MON_SEL[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12760.505 187.44 12760.785 188.44 ;
    END
  END DIG_MON_SEL[307]
  PIN DIG_MON_SEL[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12679.305 187.44 12679.585 188.44 ;
    END
  END DIG_MON_SEL[306]
  PIN DIG_MON_SEL[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12678.745 187.44 12679.025 188.44 ;
    END
  END DIG_MON_SEL[305]
  PIN DIG_MON_SEL[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12613.785 187.44 12614.065 188.44 ;
    END
  END DIG_MON_SEL[304]
  PIN DIG_MON_SEL[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12613.225 187.44 12613.505 188.44 ;
    END
  END DIG_MON_SEL[303]
  PIN DIG_MON_SEL[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12532.585 187.44 12532.865 188.44 ;
    END
  END DIG_MON_SEL[302]
  PIN DIG_MON_SEL[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12532.025 187.44 12532.305 188.44 ;
    END
  END DIG_MON_SEL[301]
  PIN DIG_MON_SEL[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12454.185 187.44 12454.465 188.44 ;
    END
  END DIG_MON_SEL[300]
  PIN DIG_MON_SEL[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12453.625 187.44 12453.905 188.44 ;
    END
  END DIG_MON_SEL[299]
  PIN DIG_MON_SEL[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12376.905 187.44 12377.185 188.44 ;
    END
  END DIG_MON_SEL[298]
  PIN DIG_MON_SEL[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12376.345 187.44 12376.625 188.44 ;
    END
  END DIG_MON_SEL[297]
  PIN DIG_MON_SEL[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12306.905 187.44 12307.185 188.44 ;
    END
  END DIG_MON_SEL[296]
  PIN DIG_MON_SEL[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12306.345 187.44 12306.625 188.44 ;
    END
  END DIG_MON_SEL[295]
  PIN DIG_MON_SEL[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12227.105 187.44 12227.385 188.44 ;
    END
  END DIG_MON_SEL[294]
  PIN DIG_MON_SEL[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12200.505 187.44 12200.785 188.44 ;
    END
  END DIG_MON_SEL[293]
  PIN DIG_MON_SEL[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12119.305 187.44 12119.585 188.44 ;
    END
  END DIG_MON_SEL[292]
  PIN DIG_MON_SEL[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12118.745 187.44 12119.025 188.44 ;
    END
  END DIG_MON_SEL[291]
  PIN DIG_MON_SEL[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12053.785 187.44 12054.065 188.44 ;
    END
  END DIG_MON_SEL[290]
  PIN DIG_MON_SEL[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12053.225 187.44 12053.505 188.44 ;
    END
  END DIG_MON_SEL[289]
  PIN DIG_MON_SEL[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11972.585 187.44 11972.865 188.44 ;
    END
  END DIG_MON_SEL[288]
  PIN DIG_MON_SEL[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11972.025 187.44 11972.305 188.44 ;
    END
  END DIG_MON_SEL[287]
  PIN DIG_MON_SEL[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11894.185 187.44 11894.465 188.44 ;
    END
  END DIG_MON_SEL[286]
  PIN DIG_MON_SEL[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11893.625 187.44 11893.905 188.44 ;
    END
  END DIG_MON_SEL[285]
  PIN DIG_MON_SEL[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11816.905 187.44 11817.185 188.44 ;
    END
  END DIG_MON_SEL[284]
  PIN DIG_MON_SEL[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11816.345 187.44 11816.625 188.44 ;
    END
  END DIG_MON_SEL[283]
  PIN DIG_MON_SEL[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11746.905 187.44 11747.185 188.44 ;
    END
  END DIG_MON_SEL[282]
  PIN DIG_MON_SEL[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11746.345 187.44 11746.625 188.44 ;
    END
  END DIG_MON_SEL[281]
  PIN DIG_MON_SEL[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11667.105 187.44 11667.385 188.44 ;
    END
  END DIG_MON_SEL[280]
  PIN DIG_MON_SEL[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11640.505 187.44 11640.785 188.44 ;
    END
  END DIG_MON_SEL[279]
  PIN DIG_MON_SEL[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11559.305 187.44 11559.585 188.44 ;
    END
  END DIG_MON_SEL[278]
  PIN DIG_MON_SEL[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11558.745 187.44 11559.025 188.44 ;
    END
  END DIG_MON_SEL[277]
  PIN DIG_MON_SEL[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11493.785 187.44 11494.065 188.44 ;
    END
  END DIG_MON_SEL[276]
  PIN DIG_MON_SEL[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11493.225 187.44 11493.505 188.44 ;
    END
  END DIG_MON_SEL[275]
  PIN DIG_MON_SEL[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11412.585 187.44 11412.865 188.44 ;
    END
  END DIG_MON_SEL[274]
  PIN DIG_MON_SEL[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11412.025 187.44 11412.305 188.44 ;
    END
  END DIG_MON_SEL[273]
  PIN DIG_MON_SEL[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11334.185 187.44 11334.465 188.44 ;
    END
  END DIG_MON_SEL[272]
  PIN DIG_MON_SEL[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11333.625 187.44 11333.905 188.44 ;
    END
  END DIG_MON_SEL[271]
  PIN DIG_MON_SEL[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11256.905 187.44 11257.185 188.44 ;
    END
  END DIG_MON_SEL[270]
  PIN DIG_MON_SEL[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11256.345 187.44 11256.625 188.44 ;
    END
  END DIG_MON_SEL[269]
  PIN DIG_MON_SEL[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11186.905 187.44 11187.185 188.44 ;
    END
  END DIG_MON_SEL[268]
  PIN DIG_MON_SEL[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11186.345 187.44 11186.625 188.44 ;
    END
  END DIG_MON_SEL[267]
  PIN DIG_MON_SEL[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11107.105 187.44 11107.385 188.44 ;
    END
  END DIG_MON_SEL[266]
  PIN DIG_MON_SEL[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11080.505 187.44 11080.785 188.44 ;
    END
  END DIG_MON_SEL[265]
  PIN DIG_MON_SEL[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10999.305 187.44 10999.585 188.44 ;
    END
  END DIG_MON_SEL[264]
  PIN DIG_MON_SEL[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10998.745 187.44 10999.025 188.44 ;
    END
  END DIG_MON_SEL[263]
  PIN DIG_MON_SEL[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10933.785 187.44 10934.065 188.44 ;
    END
  END DIG_MON_SEL[262]
  PIN DIG_MON_SEL[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10933.225 187.44 10933.505 188.44 ;
    END
  END DIG_MON_SEL[261]
  PIN DIG_MON_SEL[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10852.585 187.44 10852.865 188.44 ;
    END
  END DIG_MON_SEL[260]
  PIN DIG_MON_SEL[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10852.025 187.44 10852.305 188.44 ;
    END
  END DIG_MON_SEL[259]
  PIN DIG_MON_SEL[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10774.185 187.44 10774.465 188.44 ;
    END
  END DIG_MON_SEL[258]
  PIN DIG_MON_SEL[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10773.625 187.44 10773.905 188.44 ;
    END
  END DIG_MON_SEL[257]
  PIN DIG_MON_SEL[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10696.905 187.44 10697.185 188.44 ;
    END
  END DIG_MON_SEL[256]
  PIN DIG_MON_SEL[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10696.345 187.44 10696.625 188.44 ;
    END
  END DIG_MON_SEL[255]
  PIN DIG_MON_SEL[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10626.905 187.44 10627.185 188.44 ;
    END
  END DIG_MON_SEL[254]
  PIN DIG_MON_SEL[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10626.345 187.44 10626.625 188.44 ;
    END
  END DIG_MON_SEL[253]
  PIN DIG_MON_SEL[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10547.105 187.44 10547.385 188.44 ;
    END
  END DIG_MON_SEL[252]
  PIN DIG_MON_SEL[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10520.505 187.44 10520.785 188.44 ;
    END
  END DIG_MON_SEL[251]
  PIN DIG_MON_SEL[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10439.305 187.44 10439.585 188.44 ;
    END
  END DIG_MON_SEL[250]
  PIN DIG_MON_SEL[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10438.745 187.44 10439.025 188.44 ;
    END
  END DIG_MON_SEL[249]
  PIN DIG_MON_SEL[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10373.785 187.44 10374.065 188.44 ;
    END
  END DIG_MON_SEL[248]
  PIN DIG_MON_SEL[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10373.225 187.44 10373.505 188.44 ;
    END
  END DIG_MON_SEL[247]
  PIN DIG_MON_SEL[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10292.585 187.44 10292.865 188.44 ;
    END
  END DIG_MON_SEL[246]
  PIN DIG_MON_SEL[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10292.025 187.44 10292.305 188.44 ;
    END
  END DIG_MON_SEL[245]
  PIN DIG_MON_SEL[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10214.185 187.44 10214.465 188.44 ;
    END
  END DIG_MON_SEL[244]
  PIN DIG_MON_SEL[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10213.625 187.44 10213.905 188.44 ;
    END
  END DIG_MON_SEL[243]
  PIN DIG_MON_SEL[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10136.905 187.44 10137.185 188.44 ;
    END
  END DIG_MON_SEL[242]
  PIN DIG_MON_SEL[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10136.345 187.44 10136.625 188.44 ;
    END
  END DIG_MON_SEL[241]
  PIN DIG_MON_SEL[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10066.905 187.44 10067.185 188.44 ;
    END
  END DIG_MON_SEL[240]
  PIN DIG_MON_SEL[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10066.345 187.44 10066.625 188.44 ;
    END
  END DIG_MON_SEL[239]
  PIN DIG_MON_SEL[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9987.105 187.44 9987.385 188.44 ;
    END
  END DIG_MON_SEL[238]
  PIN DIG_MON_SEL[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9960.505 187.44 9960.785 188.44 ;
    END
  END DIG_MON_SEL[237]
  PIN DIG_MON_SEL[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9879.305 187.44 9879.585 188.44 ;
    END
  END DIG_MON_SEL[236]
  PIN DIG_MON_SEL[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9878.745 187.44 9879.025 188.44 ;
    END
  END DIG_MON_SEL[235]
  PIN DIG_MON_SEL[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9813.785 187.44 9814.065 188.44 ;
    END
  END DIG_MON_SEL[234]
  PIN DIG_MON_SEL[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9813.225 187.44 9813.505 188.44 ;
    END
  END DIG_MON_SEL[233]
  PIN DIG_MON_SEL[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9732.585 187.44 9732.865 188.44 ;
    END
  END DIG_MON_SEL[232]
  PIN DIG_MON_SEL[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9732.025 187.44 9732.305 188.44 ;
    END
  END DIG_MON_SEL[231]
  PIN DIG_MON_SEL[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9654.185 187.44 9654.465 188.44 ;
    END
  END DIG_MON_SEL[230]
  PIN DIG_MON_SEL[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9653.625 187.44 9653.905 188.44 ;
    END
  END DIG_MON_SEL[229]
  PIN DIG_MON_SEL[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9576.905 187.44 9577.185 188.44 ;
    END
  END DIG_MON_SEL[228]
  PIN DIG_MON_SEL[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9576.345 187.44 9576.625 188.44 ;
    END
  END DIG_MON_SEL[227]
  PIN DIG_MON_SEL[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9506.905 187.44 9507.185 188.44 ;
    END
  END DIG_MON_SEL[226]
  PIN DIG_MON_SEL[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9506.345 187.44 9506.625 188.44 ;
    END
  END DIG_MON_SEL[225]
  PIN DIG_MON_SEL[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9427.105 187.44 9427.385 188.44 ;
    END
  END DIG_MON_SEL[224]
  PIN DIG_MON_SEL[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9400.505 187.44 9400.785 188.44 ;
    END
  END DIG_MON_SEL[223]
  PIN DIG_MON_SEL[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9319.305 187.44 9319.585 188.44 ;
    END
  END DIG_MON_SEL[222]
  PIN DIG_MON_SEL[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9318.745 187.44 9319.025 188.44 ;
    END
  END DIG_MON_SEL[221]
  PIN DIG_MON_SEL[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9253.785 187.44 9254.065 188.44 ;
    END
  END DIG_MON_SEL[220]
  PIN DIG_MON_SEL[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9253.225 187.44 9253.505 188.44 ;
    END
  END DIG_MON_SEL[219]
  PIN DIG_MON_SEL[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9172.585 187.44 9172.865 188.44 ;
    END
  END DIG_MON_SEL[218]
  PIN DIG_MON_SEL[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9172.025 187.44 9172.305 188.44 ;
    END
  END DIG_MON_SEL[217]
  PIN DIG_MON_SEL[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9094.185 187.44 9094.465 188.44 ;
    END
  END DIG_MON_SEL[216]
  PIN DIG_MON_SEL[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9093.625 187.44 9093.905 188.44 ;
    END
  END DIG_MON_SEL[215]
  PIN DIG_MON_SEL[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9016.905 187.44 9017.185 188.44 ;
    END
  END DIG_MON_SEL[214]
  PIN DIG_MON_SEL[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9016.345 187.44 9016.625 188.44 ;
    END
  END DIG_MON_SEL[213]
  PIN DIG_MON_SEL[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8946.905 187.44 8947.185 188.44 ;
    END
  END DIG_MON_SEL[212]
  PIN DIG_MON_SEL[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8946.345 187.44 8946.625 188.44 ;
    END
  END DIG_MON_SEL[211]
  PIN DIG_MON_SEL[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8867.105 187.44 8867.385 188.44 ;
    END
  END DIG_MON_SEL[210]
  PIN DIG_MON_SEL[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8840.505 187.44 8840.785 188.44 ;
    END
  END DIG_MON_SEL[209]
  PIN DIG_MON_SEL[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8759.305 187.44 8759.585 188.44 ;
    END
  END DIG_MON_SEL[208]
  PIN DIG_MON_SEL[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8758.745 187.44 8759.025 188.44 ;
    END
  END DIG_MON_SEL[207]
  PIN DIG_MON_SEL[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8693.785 187.44 8694.065 188.44 ;
    END
  END DIG_MON_SEL[206]
  PIN DIG_MON_SEL[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8693.225 187.44 8693.505 188.44 ;
    END
  END DIG_MON_SEL[205]
  PIN DIG_MON_SEL[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8612.585 187.44 8612.865 188.44 ;
    END
  END DIG_MON_SEL[204]
  PIN DIG_MON_SEL[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8612.025 187.44 8612.305 188.44 ;
    END
  END DIG_MON_SEL[203]
  PIN DIG_MON_SEL[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8534.185 187.44 8534.465 188.44 ;
    END
  END DIG_MON_SEL[202]
  PIN DIG_MON_SEL[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8533.625 187.44 8533.905 188.44 ;
    END
  END DIG_MON_SEL[201]
  PIN DIG_MON_SEL[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8456.905 187.44 8457.185 188.44 ;
    END
  END DIG_MON_SEL[200]
  PIN DIG_MON_SEL[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8456.345 187.44 8456.625 188.44 ;
    END
  END DIG_MON_SEL[199]
  PIN DIG_MON_SEL[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8386.905 187.44 8387.185 188.44 ;
    END
  END DIG_MON_SEL[198]
  PIN DIG_MON_SEL[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8386.345 187.44 8386.625 188.44 ;
    END
  END DIG_MON_SEL[197]
  PIN DIG_MON_SEL[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8307.105 187.44 8307.385 188.44 ;
    END
  END DIG_MON_SEL[196]
  PIN DIG_MON_SEL[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8280.505 187.44 8280.785 188.44 ;
    END
  END DIG_MON_SEL[195]
  PIN DIG_MON_SEL[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8199.305 187.44 8199.585 188.44 ;
    END
  END DIG_MON_SEL[194]
  PIN DIG_MON_SEL[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8198.745 187.44 8199.025 188.44 ;
    END
  END DIG_MON_SEL[193]
  PIN DIG_MON_SEL[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8133.785 187.44 8134.065 188.44 ;
    END
  END DIG_MON_SEL[192]
  PIN DIG_MON_SEL[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8133.225 187.44 8133.505 188.44 ;
    END
  END DIG_MON_SEL[191]
  PIN DIG_MON_SEL[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8052.585 187.44 8052.865 188.44 ;
    END
  END DIG_MON_SEL[190]
  PIN DIG_MON_SEL[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8052.025 187.44 8052.305 188.44 ;
    END
  END DIG_MON_SEL[189]
  PIN DIG_MON_SEL[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7974.185 187.44 7974.465 188.44 ;
    END
  END DIG_MON_SEL[188]
  PIN DIG_MON_SEL[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7973.625 187.44 7973.905 188.44 ;
    END
  END DIG_MON_SEL[187]
  PIN DIG_MON_SEL[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7896.905 187.44 7897.185 188.44 ;
    END
  END DIG_MON_SEL[186]
  PIN DIG_MON_SEL[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7896.345 187.44 7896.625 188.44 ;
    END
  END DIG_MON_SEL[185]
  PIN DIG_MON_SEL[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7826.905 187.44 7827.185 188.44 ;
    END
  END DIG_MON_SEL[184]
  PIN DIG_MON_SEL[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7826.345 187.44 7826.625 188.44 ;
    END
  END DIG_MON_SEL[183]
  PIN DIG_MON_SEL[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7747.105 187.44 7747.385 188.44 ;
    END
  END DIG_MON_SEL[182]
  PIN DIG_MON_SEL[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7720.505 187.44 7720.785 188.44 ;
    END
  END DIG_MON_SEL[181]
  PIN DIG_MON_SEL[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7639.305 187.44 7639.585 188.44 ;
    END
  END DIG_MON_SEL[180]
  PIN DIG_MON_SEL[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7638.745 187.44 7639.025 188.44 ;
    END
  END DIG_MON_SEL[179]
  PIN DIG_MON_SEL[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7573.785 187.44 7574.065 188.44 ;
    END
  END DIG_MON_SEL[178]
  PIN DIG_MON_SEL[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7573.225 187.44 7573.505 188.44 ;
    END
  END DIG_MON_SEL[177]
  PIN DIG_MON_SEL[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7492.585 187.44 7492.865 188.44 ;
    END
  END DIG_MON_SEL[176]
  PIN DIG_MON_SEL[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7492.025 187.44 7492.305 188.44 ;
    END
  END DIG_MON_SEL[175]
  PIN DIG_MON_SEL[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7414.185 187.44 7414.465 188.44 ;
    END
  END DIG_MON_SEL[174]
  PIN DIG_MON_SEL[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7413.625 187.44 7413.905 188.44 ;
    END
  END DIG_MON_SEL[173]
  PIN DIG_MON_SEL[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7336.905 187.44 7337.185 188.44 ;
    END
  END DIG_MON_SEL[172]
  PIN DIG_MON_SEL[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7336.345 187.44 7336.625 188.44 ;
    END
  END DIG_MON_SEL[171]
  PIN DIG_MON_SEL[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7266.905 187.44 7267.185 188.44 ;
    END
  END DIG_MON_SEL[170]
  PIN DIG_MON_SEL[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7266.345 187.44 7266.625 188.44 ;
    END
  END DIG_MON_SEL[169]
  PIN DIG_MON_SEL[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7187.105 187.44 7187.385 188.44 ;
    END
  END DIG_MON_SEL[168]
  PIN DIG_MON_SEL[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7160.505 187.44 7160.785 188.44 ;
    END
  END DIG_MON_SEL[167]
  PIN DIG_MON_SEL[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7079.305 187.44 7079.585 188.44 ;
    END
  END DIG_MON_SEL[166]
  PIN DIG_MON_SEL[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7078.745 187.44 7079.025 188.44 ;
    END
  END DIG_MON_SEL[165]
  PIN DIG_MON_SEL[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7013.785 187.44 7014.065 188.44 ;
    END
  END DIG_MON_SEL[164]
  PIN DIG_MON_SEL[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7013.225 187.44 7013.505 188.44 ;
    END
  END DIG_MON_SEL[163]
  PIN DIG_MON_SEL[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6932.585 187.44 6932.865 188.44 ;
    END
  END DIG_MON_SEL[162]
  PIN DIG_MON_SEL[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6932.025 187.44 6932.305 188.44 ;
    END
  END DIG_MON_SEL[161]
  PIN DIG_MON_SEL[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6854.185 187.44 6854.465 188.44 ;
    END
  END DIG_MON_SEL[160]
  PIN DIG_MON_SEL[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6853.625 187.44 6853.905 188.44 ;
    END
  END DIG_MON_SEL[159]
  PIN DIG_MON_SEL[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6776.905 187.44 6777.185 188.44 ;
    END
  END DIG_MON_SEL[158]
  PIN DIG_MON_SEL[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6776.345 187.44 6776.625 188.44 ;
    END
  END DIG_MON_SEL[157]
  PIN DIG_MON_SEL[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6706.905 187.44 6707.185 188.44 ;
    END
  END DIG_MON_SEL[156]
  PIN DIG_MON_SEL[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6706.345 187.44 6706.625 188.44 ;
    END
  END DIG_MON_SEL[155]
  PIN DIG_MON_SEL[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6627.105 187.44 6627.385 188.44 ;
    END
  END DIG_MON_SEL[154]
  PIN DIG_MON_SEL[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6600.505 187.44 6600.785 188.44 ;
    END
  END DIG_MON_SEL[153]
  PIN DIG_MON_SEL[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6519.305 187.44 6519.585 188.44 ;
    END
  END DIG_MON_SEL[152]
  PIN DIG_MON_SEL[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6518.745 187.44 6519.025 188.44 ;
    END
  END DIG_MON_SEL[151]
  PIN DIG_MON_SEL[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6453.785 187.44 6454.065 188.44 ;
    END
  END DIG_MON_SEL[150]
  PIN DIG_MON_SEL[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6453.225 187.44 6453.505 188.44 ;
    END
  END DIG_MON_SEL[149]
  PIN DIG_MON_SEL[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6372.585 187.44 6372.865 188.44 ;
    END
  END DIG_MON_SEL[148]
  PIN DIG_MON_SEL[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6372.025 187.44 6372.305 188.44 ;
    END
  END DIG_MON_SEL[147]
  PIN DIG_MON_SEL[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6294.185 187.44 6294.465 188.44 ;
    END
  END DIG_MON_SEL[146]
  PIN DIG_MON_SEL[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6293.625 187.44 6293.905 188.44 ;
    END
  END DIG_MON_SEL[145]
  PIN DIG_MON_SEL[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6216.905 187.44 6217.185 188.44 ;
    END
  END DIG_MON_SEL[144]
  PIN DIG_MON_SEL[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6216.345 187.44 6216.625 188.44 ;
    END
  END DIG_MON_SEL[143]
  PIN DIG_MON_SEL[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6146.905 187.44 6147.185 188.44 ;
    END
  END DIG_MON_SEL[142]
  PIN DIG_MON_SEL[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6146.345 187.44 6146.625 188.44 ;
    END
  END DIG_MON_SEL[141]
  PIN DIG_MON_SEL[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6067.105 187.44 6067.385 188.44 ;
    END
  END DIG_MON_SEL[140]
  PIN DIG_MON_SEL[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6040.505 187.44 6040.785 188.44 ;
    END
  END DIG_MON_SEL[139]
  PIN DIG_MON_SEL[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5959.305 187.44 5959.585 188.44 ;
    END
  END DIG_MON_SEL[138]
  PIN DIG_MON_SEL[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5958.745 187.44 5959.025 188.44 ;
    END
  END DIG_MON_SEL[137]
  PIN DIG_MON_SEL[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5893.785 187.44 5894.065 188.44 ;
    END
  END DIG_MON_SEL[136]
  PIN DIG_MON_SEL[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5893.225 187.44 5893.505 188.44 ;
    END
  END DIG_MON_SEL[135]
  PIN DIG_MON_SEL[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5812.585 187.44 5812.865 188.44 ;
    END
  END DIG_MON_SEL[134]
  PIN DIG_MON_SEL[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5812.025 187.44 5812.305 188.44 ;
    END
  END DIG_MON_SEL[133]
  PIN DIG_MON_SEL[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5734.185 187.44 5734.465 188.44 ;
    END
  END DIG_MON_SEL[132]
  PIN DIG_MON_SEL[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5733.625 187.44 5733.905 188.44 ;
    END
  END DIG_MON_SEL[131]
  PIN DIG_MON_SEL[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5656.905 187.44 5657.185 188.44 ;
    END
  END DIG_MON_SEL[130]
  PIN DIG_MON_SEL[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5656.345 187.44 5656.625 188.44 ;
    END
  END DIG_MON_SEL[129]
  PIN DIG_MON_SEL[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5586.905 187.44 5587.185 188.44 ;
    END
  END DIG_MON_SEL[128]
  PIN DIG_MON_SEL[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5586.345 187.44 5586.625 188.44 ;
    END
  END DIG_MON_SEL[127]
  PIN DIG_MON_SEL[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5507.105 187.44 5507.385 188.44 ;
    END
  END DIG_MON_SEL[126]
  PIN DIG_MON_SEL[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5480.505 187.44 5480.785 188.44 ;
    END
  END DIG_MON_SEL[125]
  PIN DIG_MON_SEL[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5399.305 187.44 5399.585 188.44 ;
    END
  END DIG_MON_SEL[124]
  PIN DIG_MON_SEL[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5398.745 187.44 5399.025 188.44 ;
    END
  END DIG_MON_SEL[123]
  PIN DIG_MON_SEL[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5333.785 187.44 5334.065 188.44 ;
    END
  END DIG_MON_SEL[122]
  PIN DIG_MON_SEL[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5333.225 187.44 5333.505 188.44 ;
    END
  END DIG_MON_SEL[121]
  PIN DIG_MON_SEL[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5252.585 187.44 5252.865 188.44 ;
    END
  END DIG_MON_SEL[120]
  PIN DIG_MON_SEL[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5252.025 187.44 5252.305 188.44 ;
    END
  END DIG_MON_SEL[119]
  PIN DIG_MON_SEL[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5174.185 187.44 5174.465 188.44 ;
    END
  END DIG_MON_SEL[118]
  PIN DIG_MON_SEL[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5173.625 187.44 5173.905 188.44 ;
    END
  END DIG_MON_SEL[117]
  PIN DIG_MON_SEL[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5096.905 187.44 5097.185 188.44 ;
    END
  END DIG_MON_SEL[116]
  PIN DIG_MON_SEL[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5096.345 187.44 5096.625 188.44 ;
    END
  END DIG_MON_SEL[115]
  PIN DIG_MON_SEL[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5026.905 187.44 5027.185 188.44 ;
    END
  END DIG_MON_SEL[114]
  PIN DIG_MON_SEL[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5026.345 187.44 5026.625 188.44 ;
    END
  END DIG_MON_SEL[113]
  PIN DIG_MON_SEL[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4947.105 187.44 4947.385 188.44 ;
    END
  END DIG_MON_SEL[112]
  PIN DIG_MON_SEL[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4920.505 187.44 4920.785 188.44 ;
    END
  END DIG_MON_SEL[111]
  PIN DIG_MON_SEL[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4839.305 187.44 4839.585 188.44 ;
    END
  END DIG_MON_SEL[110]
  PIN DIG_MON_SEL[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4838.745 187.44 4839.025 188.44 ;
    END
  END DIG_MON_SEL[109]
  PIN DIG_MON_SEL[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4773.785 187.44 4774.065 188.44 ;
    END
  END DIG_MON_SEL[108]
  PIN DIG_MON_SEL[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4773.225 187.44 4773.505 188.44 ;
    END
  END DIG_MON_SEL[107]
  PIN DIG_MON_SEL[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4692.585 187.44 4692.865 188.44 ;
    END
  END DIG_MON_SEL[106]
  PIN DIG_MON_SEL[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4692.025 187.44 4692.305 188.44 ;
    END
  END DIG_MON_SEL[105]
  PIN DIG_MON_SEL[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4614.185 187.44 4614.465 188.44 ;
    END
  END DIG_MON_SEL[104]
  PIN DIG_MON_SEL[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4613.625 187.44 4613.905 188.44 ;
    END
  END DIG_MON_SEL[103]
  PIN DIG_MON_SEL[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4536.905 187.44 4537.185 188.44 ;
    END
  END DIG_MON_SEL[102]
  PIN DIG_MON_SEL[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4536.345 187.44 4536.625 188.44 ;
    END
  END DIG_MON_SEL[101]
  PIN DIG_MON_SEL[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4466.905 187.44 4467.185 188.44 ;
    END
  END DIG_MON_SEL[100]
  PIN DIG_MON_SEL[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4466.345 187.44 4466.625 188.44 ;
    END
  END DIG_MON_SEL[99]
  PIN DIG_MON_SEL[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4387.105 187.44 4387.385 188.44 ;
    END
  END DIG_MON_SEL[98]
  PIN DIG_MON_SEL[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4360.505 187.44 4360.785 188.44 ;
    END
  END DIG_MON_SEL[97]
  PIN DIG_MON_SEL[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4279.305 187.44 4279.585 188.44 ;
    END
  END DIG_MON_SEL[96]
  PIN DIG_MON_SEL[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4278.745 187.44 4279.025 188.44 ;
    END
  END DIG_MON_SEL[95]
  PIN DIG_MON_SEL[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4213.785 187.44 4214.065 188.44 ;
    END
  END DIG_MON_SEL[94]
  PIN DIG_MON_SEL[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4213.225 187.44 4213.505 188.44 ;
    END
  END DIG_MON_SEL[93]
  PIN DIG_MON_SEL[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4132.585 187.44 4132.865 188.44 ;
    END
  END DIG_MON_SEL[92]
  PIN DIG_MON_SEL[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4132.025 187.44 4132.305 188.44 ;
    END
  END DIG_MON_SEL[91]
  PIN DIG_MON_SEL[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4054.185 187.44 4054.465 188.44 ;
    END
  END DIG_MON_SEL[90]
  PIN DIG_MON_SEL[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4053.625 187.44 4053.905 188.44 ;
    END
  END DIG_MON_SEL[89]
  PIN DIG_MON_SEL[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3976.905 187.44 3977.185 188.44 ;
    END
  END DIG_MON_SEL[88]
  PIN DIG_MON_SEL[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3976.345 187.44 3976.625 188.44 ;
    END
  END DIG_MON_SEL[87]
  PIN DIG_MON_SEL[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3906.905 187.44 3907.185 188.44 ;
    END
  END DIG_MON_SEL[86]
  PIN DIG_MON_SEL[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3906.345 187.44 3906.625 188.44 ;
    END
  END DIG_MON_SEL[85]
  PIN DIG_MON_SEL[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3827.105 187.44 3827.385 188.44 ;
    END
  END DIG_MON_SEL[84]
  PIN DIG_MON_SEL[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3800.505 187.44 3800.785 188.44 ;
    END
  END DIG_MON_SEL[83]
  PIN DIG_MON_SEL[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3719.305 187.44 3719.585 188.44 ;
    END
  END DIG_MON_SEL[82]
  PIN DIG_MON_SEL[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3718.745 187.44 3719.025 188.44 ;
    END
  END DIG_MON_SEL[81]
  PIN DIG_MON_SEL[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3653.785 187.44 3654.065 188.44 ;
    END
  END DIG_MON_SEL[80]
  PIN DIG_MON_SEL[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3653.225 187.44 3653.505 188.44 ;
    END
  END DIG_MON_SEL[79]
  PIN DIG_MON_SEL[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3572.585 187.44 3572.865 188.44 ;
    END
  END DIG_MON_SEL[78]
  PIN DIG_MON_SEL[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3572.025 187.44 3572.305 188.44 ;
    END
  END DIG_MON_SEL[77]
  PIN DIG_MON_SEL[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3494.185 187.44 3494.465 188.44 ;
    END
  END DIG_MON_SEL[76]
  PIN DIG_MON_SEL[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3493.625 187.44 3493.905 188.44 ;
    END
  END DIG_MON_SEL[75]
  PIN DIG_MON_SEL[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3416.905 187.44 3417.185 188.44 ;
    END
  END DIG_MON_SEL[74]
  PIN DIG_MON_SEL[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3416.345 187.44 3416.625 188.44 ;
    END
  END DIG_MON_SEL[73]
  PIN DIG_MON_SEL[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3346.905 187.44 3347.185 188.44 ;
    END
  END DIG_MON_SEL[72]
  PIN DIG_MON_SEL[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3346.345 187.44 3346.625 188.44 ;
    END
  END DIG_MON_SEL[71]
  PIN DIG_MON_SEL[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3267.105 187.44 3267.385 188.44 ;
    END
  END DIG_MON_SEL[70]
  PIN DIG_MON_SEL[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3240.505 187.44 3240.785 188.44 ;
    END
  END DIG_MON_SEL[69]
  PIN DIG_MON_SEL[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3159.305 187.44 3159.585 188.44 ;
    END
  END DIG_MON_SEL[68]
  PIN DIG_MON_SEL[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3158.745 187.44 3159.025 188.44 ;
    END
  END DIG_MON_SEL[67]
  PIN DIG_MON_SEL[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3093.785 187.44 3094.065 188.44 ;
    END
  END DIG_MON_SEL[66]
  PIN DIG_MON_SEL[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3093.225 187.44 3093.505 188.44 ;
    END
  END DIG_MON_SEL[65]
  PIN DIG_MON_SEL[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3012.585 187.44 3012.865 188.44 ;
    END
  END DIG_MON_SEL[64]
  PIN DIG_MON_SEL[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3012.025 187.44 3012.305 188.44 ;
    END
  END DIG_MON_SEL[63]
  PIN DIG_MON_SEL[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2934.185 187.44 2934.465 188.44 ;
    END
  END DIG_MON_SEL[62]
  PIN DIG_MON_SEL[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2933.625 187.44 2933.905 188.44 ;
    END
  END DIG_MON_SEL[61]
  PIN DIG_MON_SEL[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2856.905 187.44 2857.185 188.44 ;
    END
  END DIG_MON_SEL[60]
  PIN DIG_MON_SEL[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2856.345 187.44 2856.625 188.44 ;
    END
  END DIG_MON_SEL[59]
  PIN DIG_MON_SEL[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2786.905 187.44 2787.185 188.44 ;
    END
  END DIG_MON_SEL[58]
  PIN DIG_MON_SEL[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2786.345 187.44 2786.625 188.44 ;
    END
  END DIG_MON_SEL[57]
  PIN DIG_MON_SEL[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2707.105 187.44 2707.385 188.44 ;
    END
  END DIG_MON_SEL[56]
  PIN DIG_MON_SEL[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2680.505 187.44 2680.785 188.44 ;
    END
  END DIG_MON_SEL[55]
  PIN DIG_MON_SEL[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2599.305 187.44 2599.585 188.44 ;
    END
  END DIG_MON_SEL[54]
  PIN DIG_MON_SEL[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2598.745 187.44 2599.025 188.44 ;
    END
  END DIG_MON_SEL[53]
  PIN DIG_MON_SEL[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2533.785 187.44 2534.065 188.44 ;
    END
  END DIG_MON_SEL[52]
  PIN DIG_MON_SEL[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2533.225 187.44 2533.505 188.44 ;
    END
  END DIG_MON_SEL[51]
  PIN DIG_MON_SEL[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2452.585 187.44 2452.865 188.44 ;
    END
  END DIG_MON_SEL[50]
  PIN DIG_MON_SEL[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2452.025 187.44 2452.305 188.44 ;
    END
  END DIG_MON_SEL[49]
  PIN DIG_MON_SEL[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2374.185 187.44 2374.465 188.44 ;
    END
  END DIG_MON_SEL[48]
  PIN DIG_MON_SEL[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2373.625 187.44 2373.905 188.44 ;
    END
  END DIG_MON_SEL[47]
  PIN DIG_MON_SEL[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2296.905 187.44 2297.185 188.44 ;
    END
  END DIG_MON_SEL[46]
  PIN DIG_MON_SEL[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2296.345 187.44 2296.625 188.44 ;
    END
  END DIG_MON_SEL[45]
  PIN DIG_MON_SEL[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2226.905 187.44 2227.185 188.44 ;
    END
  END DIG_MON_SEL[44]
  PIN DIG_MON_SEL[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2226.345 187.44 2226.625 188.44 ;
    END
  END DIG_MON_SEL[43]
  PIN DIG_MON_SEL[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2147.105 187.44 2147.385 188.44 ;
    END
  END DIG_MON_SEL[42]
  PIN DIG_MON_SEL[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2120.505 187.44 2120.785 188.44 ;
    END
  END DIG_MON_SEL[41]
  PIN DIG_MON_SEL[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2039.305 187.44 2039.585 188.44 ;
    END
  END DIG_MON_SEL[40]
  PIN DIG_MON_SEL[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2038.745 187.44 2039.025 188.44 ;
    END
  END DIG_MON_SEL[39]
  PIN DIG_MON_SEL[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1973.785 187.44 1974.065 188.44 ;
    END
  END DIG_MON_SEL[38]
  PIN DIG_MON_SEL[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1973.225 187.44 1973.505 188.44 ;
    END
  END DIG_MON_SEL[37]
  PIN DIG_MON_SEL[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1892.585 187.44 1892.865 188.44 ;
    END
  END DIG_MON_SEL[36]
  PIN DIG_MON_SEL[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1892.025 187.44 1892.305 188.44 ;
    END
  END DIG_MON_SEL[35]
  PIN DIG_MON_SEL[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1814.185 187.44 1814.465 188.44 ;
    END
  END DIG_MON_SEL[34]
  PIN DIG_MON_SEL[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1813.625 187.44 1813.905 188.44 ;
    END
  END DIG_MON_SEL[33]
  PIN DIG_MON_SEL[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1736.905 187.44 1737.185 188.44 ;
    END
  END DIG_MON_SEL[32]
  PIN DIG_MON_SEL[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1736.345 187.44 1736.625 188.44 ;
    END
  END DIG_MON_SEL[31]
  PIN DIG_MON_SEL[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1666.905 187.44 1667.185 188.44 ;
    END
  END DIG_MON_SEL[30]
  PIN DIG_MON_SEL[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1666.345 187.44 1666.625 188.44 ;
    END
  END DIG_MON_SEL[29]
  PIN DIG_MON_SEL[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1587.105 187.44 1587.385 188.44 ;
    END
  END DIG_MON_SEL[28]
  PIN DIG_MON_SEL[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1560.505 187.44 1560.785 188.44 ;
    END
  END DIG_MON_SEL[27]
  PIN DIG_MON_SEL[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1479.305 187.44 1479.585 188.44 ;
    END
  END DIG_MON_SEL[26]
  PIN DIG_MON_SEL[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1478.745 187.44 1479.025 188.44 ;
    END
  END DIG_MON_SEL[25]
  PIN DIG_MON_SEL[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1413.785 187.44 1414.065 188.44 ;
    END
  END DIG_MON_SEL[24]
  PIN DIG_MON_SEL[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1413.225 187.44 1413.505 188.44 ;
    END
  END DIG_MON_SEL[23]
  PIN DIG_MON_SEL[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1332.585 187.44 1332.865 188.44 ;
    END
  END DIG_MON_SEL[22]
  PIN DIG_MON_SEL[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1332.025 187.44 1332.305 188.44 ;
    END
  END DIG_MON_SEL[21]
  PIN DIG_MON_SEL[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1254.185 187.44 1254.465 188.44 ;
    END
  END DIG_MON_SEL[20]
  PIN DIG_MON_SEL[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1253.625 187.44 1253.905 188.44 ;
    END
  END DIG_MON_SEL[19]
  PIN DIG_MON_SEL[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1176.905 187.44 1177.185 188.44 ;
    END
  END DIG_MON_SEL[18]
  PIN DIG_MON_SEL[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1176.345 187.44 1176.625 188.44 ;
    END
  END DIG_MON_SEL[17]
  PIN DIG_MON_SEL[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1106.905 187.44 1107.185 188.44 ;
    END
  END DIG_MON_SEL[16]
  PIN DIG_MON_SEL[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1106.345 187.44 1106.625 188.44 ;
    END
  END DIG_MON_SEL[15]
  PIN DIG_MON_SEL[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1027.105 187.44 1027.385 188.44 ;
    END
  END DIG_MON_SEL[14]
  PIN DIG_MON_SEL[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1000.505 187.44 1000.785 188.44 ;
    END
  END DIG_MON_SEL[13]
  PIN DIG_MON_SEL[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 919.305 187.44 919.585 188.44 ;
    END
  END DIG_MON_SEL[12]
  PIN DIG_MON_SEL[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 918.745 187.44 919.025 188.44 ;
    END
  END DIG_MON_SEL[11]
  PIN DIG_MON_SEL[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 853.785 187.44 854.065 188.44 ;
    END
  END DIG_MON_SEL[10]
  PIN DIG_MON_SEL[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 853.225 187.44 853.505 188.44 ;
    END
  END DIG_MON_SEL[9]
  PIN DIG_MON_SEL[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 772.585 187.44 772.865 188.44 ;
    END
  END DIG_MON_SEL[8]
  PIN DIG_MON_SEL[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 772.025 187.44 772.305 188.44 ;
    END
  END DIG_MON_SEL[7]
  PIN DIG_MON_SEL[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 694.185 187.44 694.465 188.44 ;
    END
  END DIG_MON_SEL[6]
  PIN DIG_MON_SEL[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 693.625 187.44 693.905 188.44 ;
    END
  END DIG_MON_SEL[5]
  PIN DIG_MON_SEL[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 616.905 187.44 617.185 188.44 ;
    END
  END DIG_MON_SEL[4]
  PIN DIG_MON_SEL[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 616.345 187.44 616.625 188.44 ;
    END
  END DIG_MON_SEL[3]
  PIN DIG_MON_SEL[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 546.905 187.44 547.185 188.44 ;
    END
  END DIG_MON_SEL[2]
  PIN DIG_MON_SEL[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 546.345 187.44 546.625 188.44 ;
    END
  END DIG_MON_SEL[1]
  PIN DIG_MON_SEL[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 467.105 187.44 467.385 188.44 ;
    END
  END DIG_MON_SEL[0]
  PIN VDDA
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 326.66 8595.365 327.66 8599.975 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8523.365 327.66 8532.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8451.365 327.66 8460.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8379.365 327.66 8388.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8307.365 327.66 8316.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8235.365 327.66 8244.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8163.365 327.66 8172.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8091.365 327.66 8100.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8019.365 327.66 8028.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7947.365 327.66 7956.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7875.365 327.66 7884.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7803.365 327.66 7812.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7731.365 327.66 7740.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7659.365 327.66 7668.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7587.365 327.66 7596.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7515.365 327.66 7524.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7443.365 327.66 7452.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7371.365 327.66 7380.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7299.365 327.66 7308.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7227.365 327.66 7236.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7155.365 327.66 7164.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7083.365 327.66 7092.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7011.365 327.66 7020.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6939.365 327.66 6948.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6867.365 327.66 6876.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6795.365 327.66 6804.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6723.365 327.66 6732.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6651.365 327.66 6660.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6579.365 327.66 6588.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6507.365 327.66 6516.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6435.365 327.66 6444.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6363.365 327.66 6372.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6291.365 327.66 6300.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6219.365 327.66 6228.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6147.365 327.66 6156.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6075.365 327.66 6084.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6003.365 327.66 6012.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5931.365 327.66 5940.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5859.365 327.66 5868.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5787.365 327.66 5796.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5715.365 327.66 5724.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5643.365 327.66 5652.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5571.365 327.66 5580.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5499.365 327.66 5508.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5427.365 327.66 5436.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5355.365 327.66 5364.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5283.365 327.66 5292.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5211.365 327.66 5220.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5139.365 327.66 5148.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5067.365 327.66 5076.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4995.365 327.66 5004.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4923.365 327.66 4932.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4851.365 327.66 4860.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4779.365 327.66 4788.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4707.365 327.66 4716.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4635.365 327.66 4644.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4563.365 327.66 4572.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4491.365 327.66 4500.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4419.365 327.66 4428.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4347.365 327.66 4356.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4275.365 327.66 4284.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4203.365 327.66 4212.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4131.365 327.66 4140.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4059.365 327.66 4068.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3987.365 327.66 3996.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3915.365 327.66 3924.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3843.365 327.66 3852.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3771.365 327.66 3780.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3699.365 327.66 3708.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3627.365 327.66 3636.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3555.365 327.66 3564.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3483.365 327.66 3492.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3411.365 327.66 3420.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3339.365 327.66 3348.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3267.365 327.66 3276.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3195.365 327.66 3204.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3123.365 327.66 3132.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3051.365 327.66 3060.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2979.365 327.66 2988.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2907.365 327.66 2916.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2835.365 327.66 2844.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2763.365 327.66 2772.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2691.365 327.66 2700.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2619.365 327.66 2628.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2547.365 327.66 2556.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2475.365 327.66 2484.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2403.365 327.66 2412.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2331.365 327.66 2340.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2259.365 327.66 2268.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2187.365 327.66 2196.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2115.365 327.66 2124.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2043.365 327.66 2052.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1971.365 327.66 1980.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1899.365 327.66 1908.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1827.365 327.66 1836.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1755.365 327.66 1764.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1683.365 327.66 1692.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1611.365 327.66 1620.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1539.365 327.66 1548.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1467.365 327.66 1476.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1395.365 327.66 1404.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1323.365 327.66 1332.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1251.365 327.66 1260.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1179.365 327.66 1188.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1107.365 327.66 1116.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1035.365 327.66 1044.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 963.365 327.66 972.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 891.365 327.66 900.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 819.365 327.66 828.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 747.365 327.66 756.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 675.365 327.66 684.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 603.365 327.66 612.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 535.975 327.66 540.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8595.365 18490.46 8599.975 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8523.365 18490.46 8532.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8451.365 18490.46 8460.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8379.365 18490.46 8388.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8307.365 18490.46 8316.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8235.365 18490.46 8244.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8163.365 18490.46 8172.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8091.365 18490.46 8100.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8019.365 18490.46 8028.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7947.365 18490.46 7956.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7875.365 18490.46 7884.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7803.365 18490.46 7812.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7731.365 18490.46 7740.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7659.365 18490.46 7668.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7587.365 18490.46 7596.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7515.365 18490.46 7524.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7443.365 18490.46 7452.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7371.365 18490.46 7380.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7299.365 18490.46 7308.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7227.365 18490.46 7236.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7155.365 18490.46 7164.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7083.365 18490.46 7092.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7011.365 18490.46 7020.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6939.365 18490.46 6948.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6867.365 18490.46 6876.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6795.365 18490.46 6804.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6723.365 18490.46 6732.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6651.365 18490.46 6660.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6579.365 18490.46 6588.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6507.365 18490.46 6516.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6435.365 18490.46 6444.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6363.365 18490.46 6372.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6291.365 18490.46 6300.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6219.365 18490.46 6228.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6147.365 18490.46 6156.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6075.365 18490.46 6084.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6003.365 18490.46 6012.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5931.365 18490.46 5940.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5859.365 18490.46 5868.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5787.365 18490.46 5796.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5715.365 18490.46 5724.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5643.365 18490.46 5652.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5571.365 18490.46 5580.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5499.365 18490.46 5508.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5427.365 18490.46 5436.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5355.365 18490.46 5364.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5283.365 18490.46 5292.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5211.365 18490.46 5220.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5139.365 18490.46 5148.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5067.365 18490.46 5076.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4995.365 18490.46 5004.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4923.365 18490.46 4932.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4851.365 18490.46 4860.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4779.365 18490.46 4788.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4707.365 18490.46 4716.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4635.365 18490.46 4644.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4563.365 18490.46 4572.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4491.365 18490.46 4500.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4419.365 18490.46 4428.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4347.365 18490.46 4356.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4275.365 18490.46 4284.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4203.365 18490.46 4212.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4131.365 18490.46 4140.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4059.365 18490.46 4068.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3987.365 18490.46 3996.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3915.365 18490.46 3924.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3843.365 18490.46 3852.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3771.365 18490.46 3780.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3699.365 18490.46 3708.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3627.365 18490.46 3636.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3555.365 18490.46 3564.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3483.365 18490.46 3492.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3411.365 18490.46 3420.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3339.365 18490.46 3348.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3267.365 18490.46 3276.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3195.365 18490.46 3204.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3123.365 18490.46 3132.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3051.365 18490.46 3060.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2979.365 18490.46 2988.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2907.365 18490.46 2916.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2835.365 18490.46 2844.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2763.365 18490.46 2772.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2691.365 18490.46 2700.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2619.365 18490.46 2628.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2547.365 18490.46 2556.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2475.365 18490.46 2484.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2403.365 18490.46 2412.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2331.365 18490.46 2340.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2259.365 18490.46 2268.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2187.365 18490.46 2196.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2115.365 18490.46 2124.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2043.365 18490.46 2052.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1971.365 18490.46 1980.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1899.365 18490.46 1908.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1827.365 18490.46 1836.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1755.365 18490.46 1764.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1683.365 18490.46 1692.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1611.365 18490.46 1620.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1539.365 18490.46 1548.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1467.365 18490.46 1476.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1395.365 18490.46 1404.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1323.365 18490.46 1332.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1251.365 18490.46 1260.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1179.365 18490.46 1188.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1107.365 18490.46 1116.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1035.365 18490.46 1044.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 963.365 18490.46 972.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 891.365 18490.46 900.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 819.365 18490.46 828.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 747.365 18490.46 756.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 675.365 18490.46 684.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 603.365 18490.46 612.585 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 535.975 18490.46 540.585 ;
    END
  END VDDA
  PIN VDDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER TOP_M ;
        RECT 326.66 8558.205 327.66 8569.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8486.205 327.66 8497.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8414.205 327.66 8425.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8342.205 327.66 8353.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8270.205 327.66 8281.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8198.205 327.66 8209.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8126.205 327.66 8137.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8054.205 327.66 8065.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7982.205 327.66 7993.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7910.205 327.66 7921.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7838.205 327.66 7849.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7766.205 327.66 7777.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7694.205 327.66 7705.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7622.205 327.66 7633.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7550.205 327.66 7561.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7478.205 327.66 7489.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7406.205 327.66 7417.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7334.205 327.66 7345.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7262.205 327.66 7273.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7190.205 327.66 7201.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7118.205 327.66 7129.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7046.205 327.66 7057.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6974.205 327.66 6985.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6902.205 327.66 6913.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6830.205 327.66 6841.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6758.205 327.66 6769.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6686.205 327.66 6697.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6614.205 327.66 6625.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6542.205 327.66 6553.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6470.205 327.66 6481.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6398.205 327.66 6409.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6326.205 327.66 6337.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6254.205 327.66 6265.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6182.205 327.66 6193.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6110.205 327.66 6121.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6038.205 327.66 6049.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5966.205 327.66 5977.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5894.205 327.66 5905.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5822.205 327.66 5833.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5750.205 327.66 5761.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5678.205 327.66 5689.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5606.205 327.66 5617.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5534.205 327.66 5545.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5462.205 327.66 5473.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5390.205 327.66 5401.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5318.205 327.66 5329.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5246.205 327.66 5257.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5174.205 327.66 5185.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5102.205 327.66 5113.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5030.205 327.66 5041.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4958.205 327.66 4969.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4886.205 327.66 4897.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4814.205 327.66 4825.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4742.205 327.66 4753.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4670.205 327.66 4681.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4598.205 327.66 4609.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4526.205 327.66 4537.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4454.205 327.66 4465.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4382.205 327.66 4393.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4310.205 327.66 4321.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4238.205 327.66 4249.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4166.205 327.66 4177.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4094.205 327.66 4105.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4022.205 327.66 4033.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3950.205 327.66 3961.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3878.205 327.66 3889.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3806.205 327.66 3817.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3734.205 327.66 3745.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3662.205 327.66 3673.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3590.205 327.66 3601.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3518.205 327.66 3529.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3446.205 327.66 3457.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3374.205 327.66 3385.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3302.205 327.66 3313.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3230.205 327.66 3241.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3158.205 327.66 3169.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3086.205 327.66 3097.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3014.205 327.66 3025.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2942.205 327.66 2953.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2870.205 327.66 2881.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2798.205 327.66 2809.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2726.205 327.66 2737.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2654.205 327.66 2665.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2582.205 327.66 2593.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2510.205 327.66 2521.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2438.205 327.66 2449.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2366.205 327.66 2377.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2294.205 327.66 2305.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2222.205 327.66 2233.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2150.205 327.66 2161.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2078.205 327.66 2089.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2006.205 327.66 2017.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1934.205 327.66 1945.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1862.205 327.66 1873.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1790.205 327.66 1801.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1718.205 327.66 1729.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1646.205 327.66 1657.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1574.205 327.66 1585.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1502.205 327.66 1513.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1430.205 327.66 1441.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1358.205 327.66 1369.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1286.205 327.66 1297.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1214.205 327.66 1225.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1142.205 327.66 1153.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1070.205 327.66 1081.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 998.205 327.66 1009.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 926.205 327.66 937.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 854.205 327.66 865.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 782.205 327.66 793.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 710.205 327.66 721.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 638.205 327.66 649.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 566.205 327.66 577.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8558.205 18490.46 8569.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8486.205 18490.46 8497.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8414.205 18490.46 8425.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8342.205 18490.46 8353.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8270.205 18490.46 8281.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8198.205 18490.46 8209.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8126.205 18490.46 8137.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8054.205 18490.46 8065.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7982.205 18490.46 7993.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7910.205 18490.46 7921.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7838.205 18490.46 7849.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7766.205 18490.46 7777.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7694.205 18490.46 7705.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7622.205 18490.46 7633.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7550.205 18490.46 7561.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7478.205 18490.46 7489.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7406.205 18490.46 7417.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7334.205 18490.46 7345.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7262.205 18490.46 7273.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7190.205 18490.46 7201.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7118.205 18490.46 7129.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7046.205 18490.46 7057.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6974.205 18490.46 6985.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6902.205 18490.46 6913.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6830.205 18490.46 6841.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6758.205 18490.46 6769.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6686.205 18490.46 6697.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6614.205 18490.46 6625.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6542.205 18490.46 6553.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6470.205 18490.46 6481.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6398.205 18490.46 6409.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6326.205 18490.46 6337.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6254.205 18490.46 6265.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6182.205 18490.46 6193.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6110.205 18490.46 6121.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6038.205 18490.46 6049.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5966.205 18490.46 5977.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5894.205 18490.46 5905.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5822.205 18490.46 5833.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5750.205 18490.46 5761.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5678.205 18490.46 5689.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5606.205 18490.46 5617.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5534.205 18490.46 5545.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5462.205 18490.46 5473.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5390.205 18490.46 5401.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5318.205 18490.46 5329.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5246.205 18490.46 5257.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5174.205 18490.46 5185.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5102.205 18490.46 5113.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5030.205 18490.46 5041.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4958.205 18490.46 4969.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4886.205 18490.46 4897.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4814.205 18490.46 4825.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4742.205 18490.46 4753.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4670.205 18490.46 4681.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4598.205 18490.46 4609.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4526.205 18490.46 4537.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4454.205 18490.46 4465.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4382.205 18490.46 4393.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4310.205 18490.46 4321.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4238.205 18490.46 4249.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4166.205 18490.46 4177.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4094.205 18490.46 4105.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4022.205 18490.46 4033.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3950.205 18490.46 3961.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3878.205 18490.46 3889.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3806.205 18490.46 3817.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3734.205 18490.46 3745.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3662.205 18490.46 3673.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3590.205 18490.46 3601.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3518.205 18490.46 3529.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3446.205 18490.46 3457.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3374.205 18490.46 3385.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3302.205 18490.46 3313.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3230.205 18490.46 3241.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3158.205 18490.46 3169.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3086.205 18490.46 3097.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3014.205 18490.46 3025.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2942.205 18490.46 2953.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2870.205 18490.46 2881.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2798.205 18490.46 2809.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2726.205 18490.46 2737.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2654.205 18490.46 2665.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2582.205 18490.46 2593.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2510.205 18490.46 2521.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2438.205 18490.46 2449.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2366.205 18490.46 2377.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2294.205 18490.46 2305.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2222.205 18490.46 2233.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2150.205 18490.46 2161.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2078.205 18490.46 2089.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2006.205 18490.46 2017.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1934.205 18490.46 1945.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1862.205 18490.46 1873.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1790.205 18490.46 1801.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1718.205 18490.46 1729.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1646.205 18490.46 1657.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1574.205 18490.46 1585.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1502.205 18490.46 1513.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1430.205 18490.46 1441.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1358.205 18490.46 1369.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1286.205 18490.46 1297.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1214.205 18490.46 1225.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1142.205 18490.46 1153.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1070.205 18490.46 1081.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 998.205 18490.46 1009.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 926.205 18490.46 937.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 854.205 18490.46 865.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 782.205 18490.46 793.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 710.205 18490.46 721.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 638.205 18490.46 649.745 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 566.205 18490.46 577.745 ;
    END
  END VDDD
  PIN GNDA
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 326.66 8588.755 327.66 8593.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8534.585 327.66 8539.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8516.755 327.66 8521.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8462.585 327.66 8467.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8444.755 327.66 8449.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8390.585 327.66 8395.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8372.755 327.66 8377.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8318.585 327.66 8323.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8300.755 327.66 8305.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8246.585 327.66 8251.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8228.755 327.66 8233.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8174.585 327.66 8179.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8156.755 327.66 8161.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8102.585 327.66 8107.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8084.755 327.66 8089.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8030.585 327.66 8035.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8012.755 327.66 8017.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7958.585 327.66 7963.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7940.755 327.66 7945.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7886.585 327.66 7891.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7868.755 327.66 7873.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7814.585 327.66 7819.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7796.755 327.66 7801.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7742.585 327.66 7747.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7724.755 327.66 7729.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7670.585 327.66 7675.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7652.755 327.66 7657.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7598.585 327.66 7603.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7580.755 327.66 7585.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7526.585 327.66 7531.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7508.755 327.66 7513.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7454.585 327.66 7459.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7436.755 327.66 7441.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7382.585 327.66 7387.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7364.755 327.66 7369.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7310.585 327.66 7315.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7292.755 327.66 7297.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7238.585 327.66 7243.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7220.755 327.66 7225.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7166.585 327.66 7171.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7148.755 327.66 7153.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7094.585 327.66 7099.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7076.755 327.66 7081.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7022.585 327.66 7027.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7004.755 327.66 7009.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6950.585 327.66 6955.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6932.755 327.66 6937.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6878.585 327.66 6883.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6860.755 327.66 6865.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6806.585 327.66 6811.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6788.755 327.66 6793.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6734.585 327.66 6739.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6716.755 327.66 6721.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6662.585 327.66 6667.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6644.755 327.66 6649.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6590.585 327.66 6595.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6572.755 327.66 6577.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6518.585 327.66 6523.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6500.755 327.66 6505.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6446.585 327.66 6451.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6428.755 327.66 6433.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6374.585 327.66 6379.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6356.755 327.66 6361.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6302.585 327.66 6307.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6284.755 327.66 6289.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6230.585 327.66 6235.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6212.755 327.66 6217.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6158.585 327.66 6163.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6140.755 327.66 6145.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6086.585 327.66 6091.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6068.755 327.66 6073.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6014.585 327.66 6019.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5996.755 327.66 6001.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5942.585 327.66 5947.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5924.755 327.66 5929.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5870.585 327.66 5875.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5852.755 327.66 5857.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5798.585 327.66 5803.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5780.755 327.66 5785.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5726.585 327.66 5731.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5708.755 327.66 5713.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5654.585 327.66 5659.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5636.755 327.66 5641.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5582.585 327.66 5587.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5564.755 327.66 5569.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5510.585 327.66 5515.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5492.755 327.66 5497.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5438.585 327.66 5443.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5420.755 327.66 5425.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5366.585 327.66 5371.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5348.755 327.66 5353.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5294.585 327.66 5299.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5276.755 327.66 5281.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5222.585 327.66 5227.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5204.755 327.66 5209.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5150.585 327.66 5155.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5132.755 327.66 5137.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5078.585 327.66 5083.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5060.755 327.66 5065.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5006.585 327.66 5011.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4988.755 327.66 4993.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4934.585 327.66 4939.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4916.755 327.66 4921.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4862.585 327.66 4867.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4844.755 327.66 4849.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4790.585 327.66 4795.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4772.755 327.66 4777.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4718.585 327.66 4723.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4700.755 327.66 4705.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4646.585 327.66 4651.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4628.755 327.66 4633.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4574.585 327.66 4579.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4556.755 327.66 4561.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4502.585 327.66 4507.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4484.755 327.66 4489.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4430.585 327.66 4435.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4412.755 327.66 4417.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4358.585 327.66 4363.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4340.755 327.66 4345.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4286.585 327.66 4291.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4268.755 327.66 4273.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4214.585 327.66 4219.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4196.755 327.66 4201.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4142.585 327.66 4147.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4124.755 327.66 4129.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4070.585 327.66 4075.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4052.755 327.66 4057.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3998.585 327.66 4003.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3980.755 327.66 3985.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3926.585 327.66 3931.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3908.755 327.66 3913.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3854.585 327.66 3859.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3836.755 327.66 3841.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3782.585 327.66 3787.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3764.755 327.66 3769.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3710.585 327.66 3715.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3692.755 327.66 3697.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3638.585 327.66 3643.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3620.755 327.66 3625.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3566.585 327.66 3571.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3548.755 327.66 3553.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3494.585 327.66 3499.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3476.755 327.66 3481.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3422.585 327.66 3427.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3404.755 327.66 3409.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3350.585 327.66 3355.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3332.755 327.66 3337.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3278.585 327.66 3283.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3260.755 327.66 3265.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3206.585 327.66 3211.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3188.755 327.66 3193.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3134.585 327.66 3139.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3116.755 327.66 3121.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3062.585 327.66 3067.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3044.755 327.66 3049.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2990.585 327.66 2995.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2972.755 327.66 2977.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2918.585 327.66 2923.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2900.755 327.66 2905.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2846.585 327.66 2851.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2828.755 327.66 2833.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2774.585 327.66 2779.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2756.755 327.66 2761.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2702.585 327.66 2707.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2684.755 327.66 2689.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2630.585 327.66 2635.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2612.755 327.66 2617.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2558.585 327.66 2563.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2540.755 327.66 2545.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2486.585 327.66 2491.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2468.755 327.66 2473.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2414.585 327.66 2419.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2396.755 327.66 2401.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2342.585 327.66 2347.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2324.755 327.66 2329.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2270.585 327.66 2275.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2252.755 327.66 2257.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2198.585 327.66 2203.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2180.755 327.66 2185.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2126.585 327.66 2131.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2108.755 327.66 2113.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2054.585 327.66 2059.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2036.755 327.66 2041.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1982.585 327.66 1987.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1964.755 327.66 1969.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1910.585 327.66 1915.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1892.755 327.66 1897.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1838.585 327.66 1843.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1820.755 327.66 1825.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1766.585 327.66 1771.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1748.755 327.66 1753.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1694.585 327.66 1699.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1676.755 327.66 1681.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1622.585 327.66 1627.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1604.755 327.66 1609.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1550.585 327.66 1555.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1532.755 327.66 1537.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1478.585 327.66 1483.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1460.755 327.66 1465.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1406.585 327.66 1411.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1388.755 327.66 1393.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1334.585 327.66 1339.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1316.755 327.66 1321.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1262.585 327.66 1267.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1244.755 327.66 1249.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1190.585 327.66 1195.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1172.755 327.66 1177.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1118.585 327.66 1123.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1100.755 327.66 1105.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1046.585 327.66 1051.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1028.755 327.66 1033.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 974.585 327.66 979.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 956.755 327.66 961.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 902.585 327.66 907.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 884.755 327.66 889.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 830.585 327.66 835.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 812.755 327.66 817.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 758.585 327.66 763.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 740.755 327.66 745.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 686.585 327.66 691.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 668.755 327.66 673.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 614.585 327.66 619.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 596.755 327.66 601.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 542.585 327.66 547.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8588.755 18490.46 8593.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8534.585 18490.46 8539.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8516.755 18490.46 8521.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8462.585 18490.46 8467.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8444.755 18490.46 8449.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8390.585 18490.46 8395.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8372.755 18490.46 8377.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8318.585 18490.46 8323.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8300.755 18490.46 8305.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8246.585 18490.46 8251.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8228.755 18490.46 8233.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8174.585 18490.46 8179.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8156.755 18490.46 8161.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8102.585 18490.46 8107.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8084.755 18490.46 8089.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8030.585 18490.46 8035.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8012.755 18490.46 8017.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7958.585 18490.46 7963.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7940.755 18490.46 7945.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7886.585 18490.46 7891.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7868.755 18490.46 7873.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7814.585 18490.46 7819.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7796.755 18490.46 7801.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7742.585 18490.46 7747.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7724.755 18490.46 7729.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7670.585 18490.46 7675.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7652.755 18490.46 7657.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7598.585 18490.46 7603.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7580.755 18490.46 7585.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7526.585 18490.46 7531.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7508.755 18490.46 7513.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7454.585 18490.46 7459.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7436.755 18490.46 7441.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7382.585 18490.46 7387.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7364.755 18490.46 7369.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7310.585 18490.46 7315.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7292.755 18490.46 7297.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7238.585 18490.46 7243.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7220.755 18490.46 7225.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7166.585 18490.46 7171.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7148.755 18490.46 7153.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7094.585 18490.46 7099.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7076.755 18490.46 7081.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7022.585 18490.46 7027.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7004.755 18490.46 7009.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6950.585 18490.46 6955.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6932.755 18490.46 6937.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6878.585 18490.46 6883.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6860.755 18490.46 6865.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6806.585 18490.46 6811.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6788.755 18490.46 6793.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6734.585 18490.46 6739.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6716.755 18490.46 6721.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6662.585 18490.46 6667.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6644.755 18490.46 6649.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6590.585 18490.46 6595.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6572.755 18490.46 6577.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6518.585 18490.46 6523.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6500.755 18490.46 6505.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6446.585 18490.46 6451.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6428.755 18490.46 6433.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6374.585 18490.46 6379.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6356.755 18490.46 6361.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6302.585 18490.46 6307.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6284.755 18490.46 6289.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6230.585 18490.46 6235.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6212.755 18490.46 6217.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6158.585 18490.46 6163.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6140.755 18490.46 6145.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6086.585 18490.46 6091.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6068.755 18490.46 6073.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6014.585 18490.46 6019.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5996.755 18490.46 6001.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5942.585 18490.46 5947.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5924.755 18490.46 5929.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5870.585 18490.46 5875.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5852.755 18490.46 5857.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5798.585 18490.46 5803.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5780.755 18490.46 5785.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5726.585 18490.46 5731.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5708.755 18490.46 5713.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5654.585 18490.46 5659.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5636.755 18490.46 5641.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5582.585 18490.46 5587.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5564.755 18490.46 5569.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5510.585 18490.46 5515.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5492.755 18490.46 5497.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5438.585 18490.46 5443.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5420.755 18490.46 5425.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5366.585 18490.46 5371.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5348.755 18490.46 5353.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5294.585 18490.46 5299.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5276.755 18490.46 5281.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5222.585 18490.46 5227.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5204.755 18490.46 5209.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5150.585 18490.46 5155.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5132.755 18490.46 5137.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5078.585 18490.46 5083.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5060.755 18490.46 5065.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5006.585 18490.46 5011.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4988.755 18490.46 4993.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4934.585 18490.46 4939.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4916.755 18490.46 4921.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4862.585 18490.46 4867.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4844.755 18490.46 4849.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4790.585 18490.46 4795.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4772.755 18490.46 4777.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4718.585 18490.46 4723.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4700.755 18490.46 4705.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4646.585 18490.46 4651.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4628.755 18490.46 4633.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4574.585 18490.46 4579.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4556.755 18490.46 4561.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4502.585 18490.46 4507.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4484.755 18490.46 4489.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4430.585 18490.46 4435.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4412.755 18490.46 4417.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4358.585 18490.46 4363.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4340.755 18490.46 4345.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4286.585 18490.46 4291.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4268.755 18490.46 4273.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4214.585 18490.46 4219.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4196.755 18490.46 4201.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4142.585 18490.46 4147.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4124.755 18490.46 4129.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4070.585 18490.46 4075.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4052.755 18490.46 4057.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3998.585 18490.46 4003.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3980.755 18490.46 3985.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3926.585 18490.46 3931.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3908.755 18490.46 3913.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3854.585 18490.46 3859.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3836.755 18490.46 3841.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3782.585 18490.46 3787.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3764.755 18490.46 3769.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3710.585 18490.46 3715.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3692.755 18490.46 3697.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3638.585 18490.46 3643.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3620.755 18490.46 3625.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3566.585 18490.46 3571.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3548.755 18490.46 3553.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3494.585 18490.46 3499.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3476.755 18490.46 3481.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3422.585 18490.46 3427.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3404.755 18490.46 3409.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3350.585 18490.46 3355.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3332.755 18490.46 3337.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3278.585 18490.46 3283.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3260.755 18490.46 3265.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3206.585 18490.46 3211.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3188.755 18490.46 3193.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3134.585 18490.46 3139.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3116.755 18490.46 3121.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3062.585 18490.46 3067.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3044.755 18490.46 3049.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2990.585 18490.46 2995.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2972.755 18490.46 2977.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2918.585 18490.46 2923.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2900.755 18490.46 2905.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2846.585 18490.46 2851.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2828.755 18490.46 2833.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2774.585 18490.46 2779.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2756.755 18490.46 2761.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2702.585 18490.46 2707.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2684.755 18490.46 2689.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2630.585 18490.46 2635.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2612.755 18490.46 2617.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2558.585 18490.46 2563.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2540.755 18490.46 2545.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2486.585 18490.46 2491.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2468.755 18490.46 2473.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2414.585 18490.46 2419.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2396.755 18490.46 2401.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2342.585 18490.46 2347.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2324.755 18490.46 2329.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2270.585 18490.46 2275.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2252.755 18490.46 2257.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2198.585 18490.46 2203.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2180.755 18490.46 2185.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2126.585 18490.46 2131.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2108.755 18490.46 2113.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2054.585 18490.46 2059.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2036.755 18490.46 2041.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1982.585 18490.46 1987.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1964.755 18490.46 1969.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1910.585 18490.46 1915.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1892.755 18490.46 1897.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1838.585 18490.46 1843.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1820.755 18490.46 1825.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1766.585 18490.46 1771.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1748.755 18490.46 1753.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1694.585 18490.46 1699.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1676.755 18490.46 1681.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1622.585 18490.46 1627.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1604.755 18490.46 1609.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1550.585 18490.46 1555.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1532.755 18490.46 1537.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1478.585 18490.46 1483.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1460.755 18490.46 1465.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1406.585 18490.46 1411.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1388.755 18490.46 1393.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1334.585 18490.46 1339.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1316.755 18490.46 1321.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1262.585 18490.46 1267.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1244.755 18490.46 1249.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1190.585 18490.46 1195.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1172.755 18490.46 1177.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1118.585 18490.46 1123.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1100.755 18490.46 1105.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1046.585 18490.46 1051.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1028.755 18490.46 1033.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 974.585 18490.46 979.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 956.755 18490.46 961.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 902.585 18490.46 907.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 884.755 18490.46 889.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 830.585 18490.46 835.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 812.755 18490.46 817.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 758.585 18490.46 763.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 740.755 18490.46 745.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 686.585 18490.46 691.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 668.755 18490.46 673.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 614.585 18490.46 619.195 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 596.755 18490.46 601.365 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 542.585 18490.46 547.195 ;
    END
  END GNDA
  PIN GNDD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER TOP_M ;
        RECT 326.66 8571.745 327.66 8577.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8550.435 327.66 8556.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8499.745 327.66 8505.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8478.435 327.66 8484.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8427.745 327.66 8433.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8406.435 327.66 8412.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8355.745 327.66 8361.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8334.435 327.66 8340.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8283.745 327.66 8289.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8262.435 327.66 8268.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8211.745 327.66 8217.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8190.435 327.66 8196.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8139.745 327.66 8145.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8118.435 327.66 8124.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8067.745 327.66 8073.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8046.435 327.66 8052.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7995.745 327.66 8001.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7974.435 327.66 7980.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7923.745 327.66 7929.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7902.435 327.66 7908.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7851.745 327.66 7857.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7830.435 327.66 7836.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7779.745 327.66 7785.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7758.435 327.66 7764.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7707.745 327.66 7713.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7686.435 327.66 7692.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7635.745 327.66 7641.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7614.435 327.66 7620.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7563.745 327.66 7569.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7542.435 327.66 7548.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7491.745 327.66 7497.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7470.435 327.66 7476.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7419.745 327.66 7425.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7398.435 327.66 7404.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7347.745 327.66 7353.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7326.435 327.66 7332.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7275.745 327.66 7281.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7254.435 327.66 7260.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7203.745 327.66 7209.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7182.435 327.66 7188.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7131.745 327.66 7137.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7110.435 327.66 7116.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7059.745 327.66 7065.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7038.435 327.66 7044.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6987.745 327.66 6993.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6966.435 327.66 6972.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6915.745 327.66 6921.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6894.435 327.66 6900.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6843.745 327.66 6849.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6822.435 327.66 6828.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6771.745 327.66 6777.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6750.435 327.66 6756.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6699.745 327.66 6705.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6678.435 327.66 6684.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6627.745 327.66 6633.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6606.435 327.66 6612.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6555.745 327.66 6561.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6534.435 327.66 6540.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6483.745 327.66 6489.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6462.435 327.66 6468.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6411.745 327.66 6417.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6390.435 327.66 6396.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6339.745 327.66 6345.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6318.435 327.66 6324.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6267.745 327.66 6273.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6246.435 327.66 6252.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6195.745 327.66 6201.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6174.435 327.66 6180.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6123.745 327.66 6129.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6102.435 327.66 6108.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6051.745 327.66 6057.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6030.435 327.66 6036.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5979.745 327.66 5985.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5958.435 327.66 5964.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5907.745 327.66 5913.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5886.435 327.66 5892.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5835.745 327.66 5841.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5814.435 327.66 5820.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5763.745 327.66 5769.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5742.435 327.66 5748.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5691.745 327.66 5697.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5670.435 327.66 5676.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5619.745 327.66 5625.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5598.435 327.66 5604.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5547.745 327.66 5553.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5526.435 327.66 5532.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5475.745 327.66 5481.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5454.435 327.66 5460.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5403.745 327.66 5409.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5382.435 327.66 5388.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5331.745 327.66 5337.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5310.435 327.66 5316.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5259.745 327.66 5265.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5238.435 327.66 5244.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5187.745 327.66 5193.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5166.435 327.66 5172.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5115.745 327.66 5121.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5094.435 327.66 5100.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5043.745 327.66 5049.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5022.435 327.66 5028.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4971.745 327.66 4977.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4950.435 327.66 4956.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4899.745 327.66 4905.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4878.435 327.66 4884.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4827.745 327.66 4833.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4806.435 327.66 4812.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4755.745 327.66 4761.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4734.435 327.66 4740.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4683.745 327.66 4689.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4662.435 327.66 4668.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4611.745 327.66 4617.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4590.435 327.66 4596.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4539.745 327.66 4545.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4518.435 327.66 4524.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4467.745 327.66 4473.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4446.435 327.66 4452.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4395.745 327.66 4401.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4374.435 327.66 4380.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4323.745 327.66 4329.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4302.435 327.66 4308.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4251.745 327.66 4257.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4230.435 327.66 4236.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4179.745 327.66 4185.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4158.435 327.66 4164.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4107.745 327.66 4113.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4086.435 327.66 4092.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4035.745 327.66 4041.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4014.435 327.66 4020.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3963.745 327.66 3969.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3942.435 327.66 3948.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3891.745 327.66 3897.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3870.435 327.66 3876.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3819.745 327.66 3825.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3798.435 327.66 3804.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3747.745 327.66 3753.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3726.435 327.66 3732.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3675.745 327.66 3681.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3654.435 327.66 3660.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3603.745 327.66 3609.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3582.435 327.66 3588.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3531.745 327.66 3537.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3510.435 327.66 3516.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3459.745 327.66 3465.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3438.435 327.66 3444.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3387.745 327.66 3393.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3366.435 327.66 3372.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3315.745 327.66 3321.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3294.435 327.66 3300.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3243.745 327.66 3249.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3222.435 327.66 3228.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3171.745 327.66 3177.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3150.435 327.66 3156.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3099.745 327.66 3105.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3078.435 327.66 3084.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3027.745 327.66 3033.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3006.435 327.66 3012.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2955.745 327.66 2961.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2934.435 327.66 2940.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2883.745 327.66 2889.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2862.435 327.66 2868.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2811.745 327.66 2817.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2790.435 327.66 2796.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2739.745 327.66 2745.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2718.435 327.66 2724.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2667.745 327.66 2673.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2646.435 327.66 2652.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2595.745 327.66 2601.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2574.435 327.66 2580.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2523.745 327.66 2529.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2502.435 327.66 2508.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2451.745 327.66 2457.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2430.435 327.66 2436.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2379.745 327.66 2385.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2358.435 327.66 2364.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2307.745 327.66 2313.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2286.435 327.66 2292.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2235.745 327.66 2241.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2214.435 327.66 2220.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2163.745 327.66 2169.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2142.435 327.66 2148.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2091.745 327.66 2097.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2070.435 327.66 2076.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2019.745 327.66 2025.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1998.435 327.66 2004.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1947.745 327.66 1953.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1926.435 327.66 1932.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1875.745 327.66 1881.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1854.435 327.66 1860.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1803.745 327.66 1809.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1782.435 327.66 1788.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1731.745 327.66 1737.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1710.435 327.66 1716.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1659.745 327.66 1665.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1638.435 327.66 1644.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1587.745 327.66 1593.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1566.435 327.66 1572.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1515.745 327.66 1521.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1494.435 327.66 1500.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1443.745 327.66 1449.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1422.435 327.66 1428.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1371.745 327.66 1377.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1350.435 327.66 1356.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1299.745 327.66 1305.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1278.435 327.66 1284.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1227.745 327.66 1233.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1206.435 327.66 1212.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1155.745 327.66 1161.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1134.435 327.66 1140.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1083.745 327.66 1089.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1062.435 327.66 1068.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1011.745 327.66 1017.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 990.435 327.66 996.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 939.745 327.66 945.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 918.435 327.66 924.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 867.745 327.66 873.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 846.435 327.66 852.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 795.745 327.66 801.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 774.435 327.66 780.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 723.745 327.66 729.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 702.435 327.66 708.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 651.745 327.66 657.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 630.435 327.66 636.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 579.745 327.66 585.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 558.435 327.66 564.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8571.745 18490.46 8577.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8550.435 18490.46 8556.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8499.745 18490.46 8505.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8478.435 18490.46 8484.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8427.745 18490.46 8433.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8406.435 18490.46 8412.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8355.745 18490.46 8361.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8334.435 18490.46 8340.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8283.745 18490.46 8289.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8262.435 18490.46 8268.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8211.745 18490.46 8217.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8190.435 18490.46 8196.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8139.745 18490.46 8145.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8118.435 18490.46 8124.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8067.745 18490.46 8073.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8046.435 18490.46 8052.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7995.745 18490.46 8001.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7974.435 18490.46 7980.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7923.745 18490.46 7929.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7902.435 18490.46 7908.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7851.745 18490.46 7857.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7830.435 18490.46 7836.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7779.745 18490.46 7785.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7758.435 18490.46 7764.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7707.745 18490.46 7713.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7686.435 18490.46 7692.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7635.745 18490.46 7641.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7614.435 18490.46 7620.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7563.745 18490.46 7569.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7542.435 18490.46 7548.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7491.745 18490.46 7497.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7470.435 18490.46 7476.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7419.745 18490.46 7425.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7398.435 18490.46 7404.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7347.745 18490.46 7353.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7326.435 18490.46 7332.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7275.745 18490.46 7281.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7254.435 18490.46 7260.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7203.745 18490.46 7209.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7182.435 18490.46 7188.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7131.745 18490.46 7137.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7110.435 18490.46 7116.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7059.745 18490.46 7065.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7038.435 18490.46 7044.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6987.745 18490.46 6993.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6966.435 18490.46 6972.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6915.745 18490.46 6921.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6894.435 18490.46 6900.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6843.745 18490.46 6849.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6822.435 18490.46 6828.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6771.745 18490.46 6777.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6750.435 18490.46 6756.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6699.745 18490.46 6705.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6678.435 18490.46 6684.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6627.745 18490.46 6633.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6606.435 18490.46 6612.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6555.745 18490.46 6561.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6534.435 18490.46 6540.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6483.745 18490.46 6489.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6462.435 18490.46 6468.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6411.745 18490.46 6417.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6390.435 18490.46 6396.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6339.745 18490.46 6345.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6318.435 18490.46 6324.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6267.745 18490.46 6273.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6246.435 18490.46 6252.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6195.745 18490.46 6201.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6174.435 18490.46 6180.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6123.745 18490.46 6129.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6102.435 18490.46 6108.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6051.745 18490.46 6057.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6030.435 18490.46 6036.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5979.745 18490.46 5985.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5958.435 18490.46 5964.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5907.745 18490.46 5913.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5886.435 18490.46 5892.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5835.745 18490.46 5841.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5814.435 18490.46 5820.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5763.745 18490.46 5769.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5742.435 18490.46 5748.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5691.745 18490.46 5697.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5670.435 18490.46 5676.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5619.745 18490.46 5625.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5598.435 18490.46 5604.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5547.745 18490.46 5553.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5526.435 18490.46 5532.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5475.745 18490.46 5481.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5454.435 18490.46 5460.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5403.745 18490.46 5409.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5382.435 18490.46 5388.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5331.745 18490.46 5337.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5310.435 18490.46 5316.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5259.745 18490.46 5265.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5238.435 18490.46 5244.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5187.745 18490.46 5193.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5166.435 18490.46 5172.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5115.745 18490.46 5121.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5094.435 18490.46 5100.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5043.745 18490.46 5049.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5022.435 18490.46 5028.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4971.745 18490.46 4977.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4950.435 18490.46 4956.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4899.745 18490.46 4905.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4878.435 18490.46 4884.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4827.745 18490.46 4833.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4806.435 18490.46 4812.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4755.745 18490.46 4761.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4734.435 18490.46 4740.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4683.745 18490.46 4689.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4662.435 18490.46 4668.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4611.745 18490.46 4617.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4590.435 18490.46 4596.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4539.745 18490.46 4545.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4518.435 18490.46 4524.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4467.745 18490.46 4473.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4446.435 18490.46 4452.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4395.745 18490.46 4401.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4374.435 18490.46 4380.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4323.745 18490.46 4329.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4302.435 18490.46 4308.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4251.745 18490.46 4257.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4230.435 18490.46 4236.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4179.745 18490.46 4185.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4158.435 18490.46 4164.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4107.745 18490.46 4113.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4086.435 18490.46 4092.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4035.745 18490.46 4041.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4014.435 18490.46 4020.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3963.745 18490.46 3969.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3942.435 18490.46 3948.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3891.745 18490.46 3897.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3870.435 18490.46 3876.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3819.745 18490.46 3825.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3798.435 18490.46 3804.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3747.745 18490.46 3753.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3726.435 18490.46 3732.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3675.745 18490.46 3681.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3654.435 18490.46 3660.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3603.745 18490.46 3609.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3582.435 18490.46 3588.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3531.745 18490.46 3537.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3510.435 18490.46 3516.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3459.745 18490.46 3465.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3438.435 18490.46 3444.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3387.745 18490.46 3393.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3366.435 18490.46 3372.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3315.745 18490.46 3321.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3294.435 18490.46 3300.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3243.745 18490.46 3249.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3222.435 18490.46 3228.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3171.745 18490.46 3177.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3150.435 18490.46 3156.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3099.745 18490.46 3105.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3078.435 18490.46 3084.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3027.745 18490.46 3033.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3006.435 18490.46 3012.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2955.745 18490.46 2961.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2934.435 18490.46 2940.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2883.745 18490.46 2889.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2862.435 18490.46 2868.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2811.745 18490.46 2817.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2790.435 18490.46 2796.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2739.745 18490.46 2745.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2718.435 18490.46 2724.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2667.745 18490.46 2673.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2646.435 18490.46 2652.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2595.745 18490.46 2601.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2574.435 18490.46 2580.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2523.745 18490.46 2529.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2502.435 18490.46 2508.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2451.745 18490.46 2457.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2430.435 18490.46 2436.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2379.745 18490.46 2385.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2358.435 18490.46 2364.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2307.745 18490.46 2313.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2286.435 18490.46 2292.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2235.745 18490.46 2241.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2214.435 18490.46 2220.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2163.745 18490.46 2169.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2142.435 18490.46 2148.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2091.745 18490.46 2097.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2070.435 18490.46 2076.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2019.745 18490.46 2025.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1998.435 18490.46 2004.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1947.745 18490.46 1953.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1926.435 18490.46 1932.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1875.745 18490.46 1881.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1854.435 18490.46 1860.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1803.745 18490.46 1809.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1782.435 18490.46 1788.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1731.745 18490.46 1737.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1710.435 18490.46 1716.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1659.745 18490.46 1665.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1638.435 18490.46 1644.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1587.745 18490.46 1593.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1566.435 18490.46 1572.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1515.745 18490.46 1521.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1494.435 18490.46 1500.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1443.745 18490.46 1449.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1422.435 18490.46 1428.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1371.745 18490.46 1377.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1350.435 18490.46 1356.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1299.745 18490.46 1305.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1278.435 18490.46 1284.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1227.745 18490.46 1233.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1206.435 18490.46 1212.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1155.745 18490.46 1161.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1134.435 18490.46 1140.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1083.745 18490.46 1089.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1062.435 18490.46 1068.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1011.745 18490.46 1017.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 990.435 18490.46 996.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 939.745 18490.46 945.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 918.435 18490.46 924.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 867.745 18490.46 873.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 846.435 18490.46 852.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 795.745 18490.46 801.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 774.435 18490.46 780.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 723.745 18490.46 729.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 702.435 18490.46 708.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 651.745 18490.46 657.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 630.435 18490.46 636.205 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 579.745 18490.46 585.515 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 558.435 18490.46 564.205 ;
    END
  END GNDD
  PIN PWELL
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 326.66 8585.635 327.66 8586.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8541.195 327.66 8542.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8513.635 327.66 8514.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8469.195 327.66 8470.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8441.635 327.66 8442.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8397.195 327.66 8398.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8369.635 327.66 8370.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8325.195 327.66 8326.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8297.635 327.66 8298.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8253.195 327.66 8254.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8225.635 327.66 8226.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8181.195 327.66 8182.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8153.635 327.66 8154.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8109.195 327.66 8110.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8081.635 327.66 8082.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8037.195 327.66 8038.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8009.635 327.66 8010.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7965.195 327.66 7966.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7937.635 327.66 7938.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7893.195 327.66 7894.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7865.635 327.66 7866.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7821.195 327.66 7822.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7793.635 327.66 7794.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7749.195 327.66 7750.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7721.635 327.66 7722.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7677.195 327.66 7678.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7649.635 327.66 7650.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7605.195 327.66 7606.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7577.635 327.66 7578.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7533.195 327.66 7534.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7505.635 327.66 7506.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7461.195 327.66 7462.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7433.635 327.66 7434.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7389.195 327.66 7390.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7361.635 327.66 7362.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7317.195 327.66 7318.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7289.635 327.66 7290.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7245.195 327.66 7246.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7217.635 327.66 7218.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7173.195 327.66 7174.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7145.635 327.66 7146.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7101.195 327.66 7102.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7073.635 327.66 7074.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7029.195 327.66 7030.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 7001.635 327.66 7002.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6957.195 327.66 6958.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6929.635 327.66 6930.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6885.195 327.66 6886.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6857.635 327.66 6858.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6813.195 327.66 6814.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6785.635 327.66 6786.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6741.195 327.66 6742.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6713.635 327.66 6714.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6669.195 327.66 6670.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6641.635 327.66 6642.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6597.195 327.66 6598.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6569.635 327.66 6570.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6525.195 327.66 6526.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6497.635 327.66 6498.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6453.195 327.66 6454.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6425.635 327.66 6426.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6381.195 327.66 6382.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6353.635 327.66 6354.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6309.195 327.66 6310.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6281.635 327.66 6282.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6237.195 327.66 6238.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6209.635 327.66 6210.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6165.195 327.66 6166.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6137.635 327.66 6138.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6093.195 327.66 6094.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6065.635 327.66 6066.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 6021.195 327.66 6022.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5993.635 327.66 5994.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5949.195 327.66 5950.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5921.635 327.66 5922.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5877.195 327.66 5878.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5849.635 327.66 5850.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5805.195 327.66 5806.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5777.635 327.66 5778.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5733.195 327.66 5734.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5705.635 327.66 5706.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5661.195 327.66 5662.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5633.635 327.66 5634.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5589.195 327.66 5590.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5561.635 327.66 5562.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5517.195 327.66 5518.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5489.635 327.66 5490.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5445.195 327.66 5446.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5417.635 327.66 5418.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5373.195 327.66 5374.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5345.635 327.66 5346.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5301.195 327.66 5302.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5273.635 327.66 5274.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5229.195 327.66 5230.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5201.635 327.66 5202.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5157.195 327.66 5158.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5129.635 327.66 5130.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5085.195 327.66 5086.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5057.635 327.66 5058.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 5013.195 327.66 5014.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4985.635 327.66 4986.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4941.195 327.66 4942.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4913.635 327.66 4914.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4869.195 327.66 4870.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4841.635 327.66 4842.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4797.195 327.66 4798.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4769.635 327.66 4770.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4725.195 327.66 4726.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4697.635 327.66 4698.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4653.195 327.66 4654.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4625.635 327.66 4626.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4581.195 327.66 4582.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4553.635 327.66 4554.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4509.195 327.66 4510.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4481.635 327.66 4482.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4437.195 327.66 4438.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4409.635 327.66 4410.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4365.195 327.66 4366.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4337.635 327.66 4338.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4293.195 327.66 4294.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4265.635 327.66 4266.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4221.195 327.66 4222.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4193.635 327.66 4194.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4149.195 327.66 4150.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4121.635 327.66 4122.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4077.195 327.66 4078.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4049.635 327.66 4050.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 4005.195 327.66 4006.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3977.635 327.66 3978.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3933.195 327.66 3934.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3905.635 327.66 3906.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3861.195 327.66 3862.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3833.635 327.66 3834.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3789.195 327.66 3790.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3761.635 327.66 3762.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3717.195 327.66 3718.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3689.635 327.66 3690.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3645.195 327.66 3646.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3617.635 327.66 3618.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3573.195 327.66 3574.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3545.635 327.66 3546.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3501.195 327.66 3502.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3473.635 327.66 3474.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3429.195 327.66 3430.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3401.635 327.66 3402.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3357.195 327.66 3358.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3329.635 327.66 3330.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3285.195 327.66 3286.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3257.635 327.66 3258.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3213.195 327.66 3214.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3185.635 327.66 3186.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3141.195 327.66 3142.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3113.635 327.66 3114.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3069.195 327.66 3070.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 3041.635 327.66 3042.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2997.195 327.66 2998.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2969.635 327.66 2970.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2925.195 327.66 2926.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2897.635 327.66 2898.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2853.195 327.66 2854.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2825.635 327.66 2826.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2781.195 327.66 2782.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2753.635 327.66 2754.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2709.195 327.66 2710.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2681.635 327.66 2682.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2637.195 327.66 2638.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2609.635 327.66 2610.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2565.195 327.66 2566.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2537.635 327.66 2538.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2493.195 327.66 2494.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2465.635 327.66 2466.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2421.195 327.66 2422.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2393.635 327.66 2394.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2349.195 327.66 2350.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2321.635 327.66 2322.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2277.195 327.66 2278.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2249.635 327.66 2250.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2205.195 327.66 2206.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2177.635 327.66 2178.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2133.195 327.66 2134.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2105.635 327.66 2106.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2061.195 327.66 2062.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 2033.635 327.66 2034.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1989.195 327.66 1990.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1961.635 327.66 1962.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1917.195 327.66 1918.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1889.635 327.66 1890.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1845.195 327.66 1846.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1817.635 327.66 1818.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1773.195 327.66 1774.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1745.635 327.66 1746.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1701.195 327.66 1702.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1673.635 327.66 1674.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1629.195 327.66 1630.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1601.635 327.66 1602.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1557.195 327.66 1558.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1529.635 327.66 1530.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1485.195 327.66 1486.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1457.635 327.66 1458.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1413.195 327.66 1414.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1385.635 327.66 1386.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1341.195 327.66 1342.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1313.635 327.66 1314.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1269.195 327.66 1270.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1241.635 327.66 1242.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1197.195 327.66 1198.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1169.635 327.66 1170.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1125.195 327.66 1126.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1097.635 327.66 1098.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1053.195 327.66 1054.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 1025.635 327.66 1026.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 981.195 327.66 982.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 953.635 327.66 954.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 909.195 327.66 910.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 881.635 327.66 882.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 837.195 327.66 838.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 809.635 327.66 810.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 765.195 327.66 766.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 737.635 327.66 738.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 693.195 327.66 694.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 665.635 327.66 666.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 621.195 327.66 622.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 593.635 327.66 594.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 549.195 327.66 550.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 521.56 327.66 522.68 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8585.635 18490.46 8586.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8541.195 18490.46 8542.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8513.635 18490.46 8514.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8469.195 18490.46 8470.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8441.635 18490.46 8442.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8397.195 18490.46 8398.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8369.635 18490.46 8370.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8325.195 18490.46 8326.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8297.635 18490.46 8298.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8253.195 18490.46 8254.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8225.635 18490.46 8226.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8181.195 18490.46 8182.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8153.635 18490.46 8154.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8109.195 18490.46 8110.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8081.635 18490.46 8082.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8037.195 18490.46 8038.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 8009.635 18490.46 8010.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7965.195 18490.46 7966.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7937.635 18490.46 7938.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7893.195 18490.46 7894.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7865.635 18490.46 7866.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7821.195 18490.46 7822.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7793.635 18490.46 7794.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7749.195 18490.46 7750.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7721.635 18490.46 7722.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7677.195 18490.46 7678.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7649.635 18490.46 7650.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7605.195 18490.46 7606.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7577.635 18490.46 7578.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7533.195 18490.46 7534.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7505.635 18490.46 7506.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7461.195 18490.46 7462.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7433.635 18490.46 7434.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7389.195 18490.46 7390.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7361.635 18490.46 7362.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7317.195 18490.46 7318.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7289.635 18490.46 7290.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7245.195 18490.46 7246.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7217.635 18490.46 7218.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7173.195 18490.46 7174.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7145.635 18490.46 7146.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7101.195 18490.46 7102.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7073.635 18490.46 7074.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7029.195 18490.46 7030.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 7001.635 18490.46 7002.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6957.195 18490.46 6958.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6929.635 18490.46 6930.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6885.195 18490.46 6886.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6857.635 18490.46 6858.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6813.195 18490.46 6814.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6785.635 18490.46 6786.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6741.195 18490.46 6742.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6713.635 18490.46 6714.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6669.195 18490.46 6670.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6641.635 18490.46 6642.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6597.195 18490.46 6598.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6569.635 18490.46 6570.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6525.195 18490.46 6526.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6497.635 18490.46 6498.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6453.195 18490.46 6454.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6425.635 18490.46 6426.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6381.195 18490.46 6382.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6353.635 18490.46 6354.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6309.195 18490.46 6310.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6281.635 18490.46 6282.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6237.195 18490.46 6238.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6209.635 18490.46 6210.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6165.195 18490.46 6166.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6137.635 18490.46 6138.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6093.195 18490.46 6094.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6065.635 18490.46 6066.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 6021.195 18490.46 6022.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5993.635 18490.46 5994.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5949.195 18490.46 5950.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5921.635 18490.46 5922.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5877.195 18490.46 5878.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5849.635 18490.46 5850.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5805.195 18490.46 5806.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5777.635 18490.46 5778.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5733.195 18490.46 5734.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5705.635 18490.46 5706.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5661.195 18490.46 5662.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5633.635 18490.46 5634.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5589.195 18490.46 5590.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5561.635 18490.46 5562.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5517.195 18490.46 5518.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5489.635 18490.46 5490.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5445.195 18490.46 5446.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5417.635 18490.46 5418.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5373.195 18490.46 5374.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5345.635 18490.46 5346.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5301.195 18490.46 5302.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5273.635 18490.46 5274.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5229.195 18490.46 5230.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5201.635 18490.46 5202.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5157.195 18490.46 5158.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5129.635 18490.46 5130.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5085.195 18490.46 5086.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5057.635 18490.46 5058.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 5013.195 18490.46 5014.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4985.635 18490.46 4986.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4941.195 18490.46 4942.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4913.635 18490.46 4914.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4869.195 18490.46 4870.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4841.635 18490.46 4842.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4797.195 18490.46 4798.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4769.635 18490.46 4770.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4725.195 18490.46 4726.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4697.635 18490.46 4698.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4653.195 18490.46 4654.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4625.635 18490.46 4626.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4581.195 18490.46 4582.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4553.635 18490.46 4554.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4509.195 18490.46 4510.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4481.635 18490.46 4482.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4437.195 18490.46 4438.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4409.635 18490.46 4410.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4365.195 18490.46 4366.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4337.635 18490.46 4338.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4293.195 18490.46 4294.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4265.635 18490.46 4266.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4221.195 18490.46 4222.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4193.635 18490.46 4194.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4149.195 18490.46 4150.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4121.635 18490.46 4122.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4077.195 18490.46 4078.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4049.635 18490.46 4050.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 4005.195 18490.46 4006.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3977.635 18490.46 3978.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3933.195 18490.46 3934.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3905.635 18490.46 3906.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3861.195 18490.46 3862.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3833.635 18490.46 3834.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3789.195 18490.46 3790.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3761.635 18490.46 3762.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3717.195 18490.46 3718.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3689.635 18490.46 3690.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3645.195 18490.46 3646.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3617.635 18490.46 3618.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3573.195 18490.46 3574.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3545.635 18490.46 3546.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3501.195 18490.46 3502.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3473.635 18490.46 3474.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3429.195 18490.46 3430.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3401.635 18490.46 3402.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3357.195 18490.46 3358.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3329.635 18490.46 3330.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3285.195 18490.46 3286.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3257.635 18490.46 3258.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3213.195 18490.46 3214.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3185.635 18490.46 3186.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3141.195 18490.46 3142.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3113.635 18490.46 3114.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3069.195 18490.46 3070.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 3041.635 18490.46 3042.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2997.195 18490.46 2998.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2969.635 18490.46 2970.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2925.195 18490.46 2926.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2897.635 18490.46 2898.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2853.195 18490.46 2854.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2825.635 18490.46 2826.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2781.195 18490.46 2782.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2753.635 18490.46 2754.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2709.195 18490.46 2710.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2681.635 18490.46 2682.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2637.195 18490.46 2638.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2609.635 18490.46 2610.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2565.195 18490.46 2566.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2537.635 18490.46 2538.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2493.195 18490.46 2494.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2465.635 18490.46 2466.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2421.195 18490.46 2422.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2393.635 18490.46 2394.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2349.195 18490.46 2350.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2321.635 18490.46 2322.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2277.195 18490.46 2278.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2249.635 18490.46 2250.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2205.195 18490.46 2206.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2177.635 18490.46 2178.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2133.195 18490.46 2134.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2105.635 18490.46 2106.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2061.195 18490.46 2062.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 2033.635 18490.46 2034.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1989.195 18490.46 1990.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1961.635 18490.46 1962.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1917.195 18490.46 1918.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1889.635 18490.46 1890.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1845.195 18490.46 1846.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1817.635 18490.46 1818.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1773.195 18490.46 1774.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1745.635 18490.46 1746.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1701.195 18490.46 1702.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1673.635 18490.46 1674.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1629.195 18490.46 1630.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1601.635 18490.46 1602.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1557.195 18490.46 1558.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1529.635 18490.46 1530.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1485.195 18490.46 1486.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1457.635 18490.46 1458.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1413.195 18490.46 1414.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1385.635 18490.46 1386.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1341.195 18490.46 1342.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1313.635 18490.46 1314.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1269.195 18490.46 1270.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1241.635 18490.46 1242.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1197.195 18490.46 1198.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1169.635 18490.46 1170.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1125.195 18490.46 1126.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1097.635 18490.46 1098.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1053.195 18490.46 1054.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 1025.635 18490.46 1026.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 981.195 18490.46 982.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 953.635 18490.46 954.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 909.195 18490.46 910.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 881.635 18490.46 882.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 837.195 18490.46 838.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 809.635 18490.46 810.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 765.195 18490.46 766.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 737.635 18490.46 738.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 693.195 18490.46 694.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 665.635 18490.46 666.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 621.195 18490.46 622.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 593.635 18490.46 594.755 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 549.195 18490.46 550.315 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 521.56 18490.46 522.68 ;
    END
  END PWELL
  PIN PSUB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER TOP_M ;
        RECT 326.66 512.265 327.66 514.265 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 191.275 327.66 193.275 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 8611.565 18490.46 8613.565 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 512.265 18490.46 514.265 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 191.275 18490.46 193.275 ;
    END
  END PSUB
  PIN HV_DIODE
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 18488.96 8583.075 18490.46 8583.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 8544.315 18490.46 8544.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 8511.075 18490.46 8511.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 8472.315 18490.46 8472.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 8439.075 18490.46 8439.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 8400.315 18490.46 8400.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 8367.075 18490.46 8367.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 8328.315 18490.46 8328.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 8295.075 18490.46 8295.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 8256.315 18490.46 8256.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 8223.075 18490.46 8223.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 8184.315 18490.46 8184.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 8151.075 18490.46 8151.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 8112.315 18490.46 8112.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 8079.075 18490.46 8079.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 8040.315 18490.46 8040.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 8007.075 18490.46 8007.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 7968.315 18490.46 7968.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 7935.075 18490.46 7935.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 7896.315 18490.46 7896.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 7863.075 18490.46 7863.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 7824.315 18490.46 7824.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 7791.075 18490.46 7791.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 7752.315 18490.46 7752.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 7719.075 18490.46 7719.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 7680.315 18490.46 7680.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 7647.075 18490.46 7647.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 7608.315 18490.46 7608.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 7575.075 18490.46 7575.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 7536.315 18490.46 7536.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 7503.075 18490.46 7503.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 7464.315 18490.46 7464.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 7431.075 18490.46 7431.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 7392.315 18490.46 7392.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 7359.075 18490.46 7359.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 7320.315 18490.46 7320.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 7287.075 18490.46 7287.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 7248.315 18490.46 7248.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 7215.075 18490.46 7215.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 7176.315 18490.46 7176.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 7143.075 18490.46 7143.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 7104.315 18490.46 7104.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 7071.075 18490.46 7071.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 7032.315 18490.46 7032.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 6999.075 18490.46 6999.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 6960.315 18490.46 6960.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 6927.075 18490.46 6927.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 6888.315 18490.46 6888.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 6855.075 18490.46 6855.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 6816.315 18490.46 6816.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 6783.075 18490.46 6783.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 6744.315 18490.46 6744.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 6711.075 18490.46 6711.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 6672.315 18490.46 6672.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 6639.075 18490.46 6639.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 6600.315 18490.46 6600.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 6567.075 18490.46 6567.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 6528.315 18490.46 6528.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 6495.075 18490.46 6495.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 6456.315 18490.46 6456.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 6423.075 18490.46 6423.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 6384.315 18490.46 6384.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 6351.075 18490.46 6351.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 6312.315 18490.46 6312.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 6279.075 18490.46 6279.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 6240.315 18490.46 6240.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 6207.075 18490.46 6207.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 6168.315 18490.46 6168.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 6135.075 18490.46 6135.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 6096.315 18490.46 6096.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 6063.075 18490.46 6063.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 6024.315 18490.46 6024.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 5991.075 18490.46 5991.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 5952.315 18490.46 5952.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 5919.075 18490.46 5919.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 5880.315 18490.46 5880.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 5847.075 18490.46 5847.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 5808.315 18490.46 5808.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 5775.075 18490.46 5775.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 5736.315 18490.46 5736.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 5703.075 18490.46 5703.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 5664.315 18490.46 5664.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 5631.075 18490.46 5631.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 5592.315 18490.46 5592.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 5559.075 18490.46 5559.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 5520.315 18490.46 5520.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 5487.075 18490.46 5487.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 5448.315 18490.46 5448.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 5415.075 18490.46 5415.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 5376.315 18490.46 5376.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 5343.075 18490.46 5343.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 5304.315 18490.46 5304.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 5271.075 18490.46 5271.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 5232.315 18490.46 5232.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 5199.075 18490.46 5199.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 5160.315 18490.46 5160.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 5127.075 18490.46 5127.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 5088.315 18490.46 5088.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 5055.075 18490.46 5055.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 5016.315 18490.46 5016.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 4983.075 18490.46 4983.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 4944.315 18490.46 4944.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 4911.075 18490.46 4911.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 4872.315 18490.46 4872.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 4839.075 18490.46 4839.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 4800.315 18490.46 4800.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 4767.075 18490.46 4767.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 4728.315 18490.46 4728.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 4695.075 18490.46 4695.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 4656.315 18490.46 4656.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 4623.075 18490.46 4623.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 4584.315 18490.46 4584.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 4551.075 18490.46 4551.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 4512.315 18490.46 4512.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 4479.075 18490.46 4479.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 4440.315 18490.46 4440.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 4407.075 18490.46 4407.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 4368.315 18490.46 4368.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 4335.075 18490.46 4335.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 4296.315 18490.46 4296.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 4263.075 18490.46 4263.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 4224.315 18490.46 4224.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 4191.075 18490.46 4191.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 4152.315 18490.46 4152.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 4119.075 18490.46 4119.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 4080.315 18490.46 4080.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 4047.075 18490.46 4047.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 4008.315 18490.46 4008.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 3975.075 18490.46 3975.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 3936.315 18490.46 3936.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 3903.075 18490.46 3903.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 3864.315 18490.46 3864.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 3831.075 18490.46 3831.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 3792.315 18490.46 3792.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 3759.075 18490.46 3759.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 3720.315 18490.46 3720.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 3687.075 18490.46 3687.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 3648.315 18490.46 3648.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 3615.075 18490.46 3615.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 3576.315 18490.46 3576.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 3543.075 18490.46 3543.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 3504.315 18490.46 3504.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 3471.075 18490.46 3471.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 3432.315 18490.46 3432.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 3399.075 18490.46 3399.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 3360.315 18490.46 3360.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 3327.075 18490.46 3327.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 3288.315 18490.46 3288.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 3255.075 18490.46 3255.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 3216.315 18490.46 3216.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 3183.075 18490.46 3183.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 3144.315 18490.46 3144.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 3111.075 18490.46 3111.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 3072.315 18490.46 3072.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 3039.075 18490.46 3039.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 3000.315 18490.46 3000.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 2967.075 18490.46 2967.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 2928.315 18490.46 2928.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 2895.075 18490.46 2895.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 2856.315 18490.46 2856.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 2823.075 18490.46 2823.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 2784.315 18490.46 2784.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 2751.075 18490.46 2751.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 2712.315 18490.46 2712.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 2679.075 18490.46 2679.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 2640.315 18490.46 2640.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 2607.075 18490.46 2607.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 2568.315 18490.46 2568.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 2535.075 18490.46 2535.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 2496.315 18490.46 2496.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 2463.075 18490.46 2463.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 2424.315 18490.46 2424.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 2391.075 18490.46 2391.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 2352.315 18490.46 2352.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 2319.075 18490.46 2319.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 2280.315 18490.46 2280.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 2247.075 18490.46 2247.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 2208.315 18490.46 2208.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 2175.075 18490.46 2175.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 2136.315 18490.46 2136.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 2103.075 18490.46 2103.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 2064.315 18490.46 2064.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 2031.075 18490.46 2031.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 1992.315 18490.46 1992.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 1959.075 18490.46 1959.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 1920.315 18490.46 1920.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 1887.075 18490.46 1887.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 1848.315 18490.46 1848.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 1815.075 18490.46 1815.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 1776.315 18490.46 1776.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 1743.075 18490.46 1743.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 1704.315 18490.46 1704.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 1671.075 18490.46 1671.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 1632.315 18490.46 1632.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 1599.075 18490.46 1599.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 1560.315 18490.46 1560.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 1527.075 18490.46 1527.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 1488.315 18490.46 1488.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 1455.075 18490.46 1455.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 1416.315 18490.46 1416.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 1383.075 18490.46 1383.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 1344.315 18490.46 1344.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 1311.075 18490.46 1311.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 1272.315 18490.46 1272.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 1239.075 18490.46 1239.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 1200.315 18490.46 1200.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 1167.075 18490.46 1167.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 1128.315 18490.46 1128.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 1095.075 18490.46 1095.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 1056.315 18490.46 1056.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 1023.075 18490.46 1023.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 984.315 18490.46 984.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 951.075 18490.46 951.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 912.315 18490.46 912.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 879.075 18490.46 879.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 840.315 18490.46 840.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 807.075 18490.46 807.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 768.315 18490.46 768.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 735.075 18490.46 735.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 696.315 18490.46 696.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 663.075 18490.46 663.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 624.315 18490.46 624.875 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 591.075 18490.46 591.635 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18488.96 552.315 18490.46 552.875 ;
    END
  END HV_DIODE
  PIN SET_VCLIP[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18352.875 187.44 18353.155 188.44 ;
    END
  END SET_VCLIP[127]
  PIN SET_VCLIP[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18212.875 187.44 18213.155 188.44 ;
    END
  END SET_VCLIP[126]
  PIN SET_VCLIP[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18072.875 187.44 18073.155 188.44 ;
    END
  END SET_VCLIP[125]
  PIN SET_VCLIP[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17932.875 187.44 17933.155 188.44 ;
    END
  END SET_VCLIP[124]
  PIN SET_VCLIP[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17792.875 187.44 17793.155 188.44 ;
    END
  END SET_VCLIP[123]
  PIN SET_VCLIP[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17652.875 187.44 17653.155 188.44 ;
    END
  END SET_VCLIP[122]
  PIN SET_VCLIP[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17512.875 187.44 17513.155 188.44 ;
    END
  END SET_VCLIP[121]
  PIN SET_VCLIP[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17372.875 187.44 17373.155 188.44 ;
    END
  END SET_VCLIP[120]
  PIN SET_VCLIP[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17232.875 187.44 17233.155 188.44 ;
    END
  END SET_VCLIP[119]
  PIN SET_VCLIP[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17092.875 187.44 17093.155 188.44 ;
    END
  END SET_VCLIP[118]
  PIN SET_VCLIP[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16952.875 187.44 16953.155 188.44 ;
    END
  END SET_VCLIP[117]
  PIN SET_VCLIP[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16812.875 187.44 16813.155 188.44 ;
    END
  END SET_VCLIP[116]
  PIN SET_VCLIP[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16672.875 187.44 16673.155 188.44 ;
    END
  END SET_VCLIP[115]
  PIN SET_VCLIP[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16532.875 187.44 16533.155 188.44 ;
    END
  END SET_VCLIP[114]
  PIN SET_VCLIP[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16392.875 187.44 16393.155 188.44 ;
    END
  END SET_VCLIP[113]
  PIN SET_VCLIP[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16252.875 187.44 16253.155 188.44 ;
    END
  END SET_VCLIP[112]
  PIN SET_VCLIP[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16112.875 187.44 16113.155 188.44 ;
    END
  END SET_VCLIP[111]
  PIN SET_VCLIP[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15972.875 187.44 15973.155 188.44 ;
    END
  END SET_VCLIP[110]
  PIN SET_VCLIP[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15832.875 187.44 15833.155 188.44 ;
    END
  END SET_VCLIP[109]
  PIN SET_VCLIP[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15692.875 187.44 15693.155 188.44 ;
    END
  END SET_VCLIP[108]
  PIN SET_VCLIP[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15552.875 187.44 15553.155 188.44 ;
    END
  END SET_VCLIP[107]
  PIN SET_VCLIP[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15412.875 187.44 15413.155 188.44 ;
    END
  END SET_VCLIP[106]
  PIN SET_VCLIP[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15272.875 187.44 15273.155 188.44 ;
    END
  END SET_VCLIP[105]
  PIN SET_VCLIP[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15132.875 187.44 15133.155 188.44 ;
    END
  END SET_VCLIP[104]
  PIN SET_VCLIP[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14992.875 187.44 14993.155 188.44 ;
    END
  END SET_VCLIP[103]
  PIN SET_VCLIP[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14852.875 187.44 14853.155 188.44 ;
    END
  END SET_VCLIP[102]
  PIN SET_VCLIP[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14712.875 187.44 14713.155 188.44 ;
    END
  END SET_VCLIP[101]
  PIN SET_VCLIP[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14572.875 187.44 14573.155 188.44 ;
    END
  END SET_VCLIP[100]
  PIN SET_VCLIP[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14432.875 187.44 14433.155 188.44 ;
    END
  END SET_VCLIP[99]
  PIN SET_VCLIP[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14292.875 187.44 14293.155 188.44 ;
    END
  END SET_VCLIP[98]
  PIN SET_VCLIP[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14152.875 187.44 14153.155 188.44 ;
    END
  END SET_VCLIP[97]
  PIN SET_VCLIP[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14012.875 187.44 14013.155 188.44 ;
    END
  END SET_VCLIP[96]
  PIN SET_VCLIP[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13872.875 187.44 13873.155 188.44 ;
    END
  END SET_VCLIP[95]
  PIN SET_VCLIP[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13732.875 187.44 13733.155 188.44 ;
    END
  END SET_VCLIP[94]
  PIN SET_VCLIP[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13592.875 187.44 13593.155 188.44 ;
    END
  END SET_VCLIP[93]
  PIN SET_VCLIP[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13452.875 187.44 13453.155 188.44 ;
    END
  END SET_VCLIP[92]
  PIN SET_VCLIP[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13312.875 187.44 13313.155 188.44 ;
    END
  END SET_VCLIP[91]
  PIN SET_VCLIP[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13172.875 187.44 13173.155 188.44 ;
    END
  END SET_VCLIP[90]
  PIN SET_VCLIP[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13032.875 187.44 13033.155 188.44 ;
    END
  END SET_VCLIP[89]
  PIN SET_VCLIP[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12892.875 187.44 12893.155 188.44 ;
    END
  END SET_VCLIP[88]
  PIN SET_VCLIP[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12752.875 187.44 12753.155 188.44 ;
    END
  END SET_VCLIP[87]
  PIN SET_VCLIP[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12612.875 187.44 12613.155 188.44 ;
    END
  END SET_VCLIP[86]
  PIN SET_VCLIP[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12472.875 187.44 12473.155 188.44 ;
    END
  END SET_VCLIP[85]
  PIN SET_VCLIP[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12332.875 187.44 12333.155 188.44 ;
    END
  END SET_VCLIP[84]
  PIN SET_VCLIP[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12192.875 187.44 12193.155 188.44 ;
    END
  END SET_VCLIP[83]
  PIN SET_VCLIP[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12052.875 187.44 12053.155 188.44 ;
    END
  END SET_VCLIP[82]
  PIN SET_VCLIP[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11912.875 187.44 11913.155 188.44 ;
    END
  END SET_VCLIP[81]
  PIN SET_VCLIP[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11772.875 187.44 11773.155 188.44 ;
    END
  END SET_VCLIP[80]
  PIN SET_VCLIP[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11632.875 187.44 11633.155 188.44 ;
    END
  END SET_VCLIP[79]
  PIN SET_VCLIP[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11492.875 187.44 11493.155 188.44 ;
    END
  END SET_VCLIP[78]
  PIN SET_VCLIP[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11352.875 187.44 11353.155 188.44 ;
    END
  END SET_VCLIP[77]
  PIN SET_VCLIP[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11212.875 187.44 11213.155 188.44 ;
    END
  END SET_VCLIP[76]
  PIN SET_VCLIP[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11072.875 187.44 11073.155 188.44 ;
    END
  END SET_VCLIP[75]
  PIN SET_VCLIP[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10932.875 187.44 10933.155 188.44 ;
    END
  END SET_VCLIP[74]
  PIN SET_VCLIP[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10792.875 187.44 10793.155 188.44 ;
    END
  END SET_VCLIP[73]
  PIN SET_VCLIP[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10652.875 187.44 10653.155 188.44 ;
    END
  END SET_VCLIP[72]
  PIN SET_VCLIP[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10512.875 187.44 10513.155 188.44 ;
    END
  END SET_VCLIP[71]
  PIN SET_VCLIP[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10372.875 187.44 10373.155 188.44 ;
    END
  END SET_VCLIP[70]
  PIN SET_VCLIP[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10232.875 187.44 10233.155 188.44 ;
    END
  END SET_VCLIP[69]
  PIN SET_VCLIP[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10092.875 187.44 10093.155 188.44 ;
    END
  END SET_VCLIP[68]
  PIN SET_VCLIP[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9952.875 187.44 9953.155 188.44 ;
    END
  END SET_VCLIP[67]
  PIN SET_VCLIP[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9812.875 187.44 9813.155 188.44 ;
    END
  END SET_VCLIP[66]
  PIN SET_VCLIP[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9672.875 187.44 9673.155 188.44 ;
    END
  END SET_VCLIP[65]
  PIN SET_VCLIP[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9532.875 187.44 9533.155 188.44 ;
    END
  END SET_VCLIP[64]
  PIN SET_VCLIP[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9392.875 187.44 9393.155 188.44 ;
    END
  END SET_VCLIP[63]
  PIN SET_VCLIP[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9252.875 187.44 9253.155 188.44 ;
    END
  END SET_VCLIP[62]
  PIN SET_VCLIP[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9112.875 187.44 9113.155 188.44 ;
    END
  END SET_VCLIP[61]
  PIN SET_VCLIP[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8972.875 187.44 8973.155 188.44 ;
    END
  END SET_VCLIP[60]
  PIN SET_VCLIP[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8832.875 187.44 8833.155 188.44 ;
    END
  END SET_VCLIP[59]
  PIN SET_VCLIP[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8692.875 187.44 8693.155 188.44 ;
    END
  END SET_VCLIP[58]
  PIN SET_VCLIP[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8552.875 187.44 8553.155 188.44 ;
    END
  END SET_VCLIP[57]
  PIN SET_VCLIP[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8412.875 187.44 8413.155 188.44 ;
    END
  END SET_VCLIP[56]
  PIN SET_VCLIP[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8272.875 187.44 8273.155 188.44 ;
    END
  END SET_VCLIP[55]
  PIN SET_VCLIP[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8132.875 187.44 8133.155 188.44 ;
    END
  END SET_VCLIP[54]
  PIN SET_VCLIP[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7992.875 187.44 7993.155 188.44 ;
    END
  END SET_VCLIP[53]
  PIN SET_VCLIP[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7852.875 187.44 7853.155 188.44 ;
    END
  END SET_VCLIP[52]
  PIN SET_VCLIP[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7712.875 187.44 7713.155 188.44 ;
    END
  END SET_VCLIP[51]
  PIN SET_VCLIP[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7572.875 187.44 7573.155 188.44 ;
    END
  END SET_VCLIP[50]
  PIN SET_VCLIP[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7432.875 187.44 7433.155 188.44 ;
    END
  END SET_VCLIP[49]
  PIN SET_VCLIP[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7292.875 187.44 7293.155 188.44 ;
    END
  END SET_VCLIP[48]
  PIN SET_VCLIP[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7152.875 187.44 7153.155 188.44 ;
    END
  END SET_VCLIP[47]
  PIN SET_VCLIP[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7012.875 187.44 7013.155 188.44 ;
    END
  END SET_VCLIP[46]
  PIN SET_VCLIP[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6872.875 187.44 6873.155 188.44 ;
    END
  END SET_VCLIP[45]
  PIN SET_VCLIP[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6732.875 187.44 6733.155 188.44 ;
    END
  END SET_VCLIP[44]
  PIN SET_VCLIP[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6592.875 187.44 6593.155 188.44 ;
    END
  END SET_VCLIP[43]
  PIN SET_VCLIP[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6452.875 187.44 6453.155 188.44 ;
    END
  END SET_VCLIP[42]
  PIN SET_VCLIP[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6312.875 187.44 6313.155 188.44 ;
    END
  END SET_VCLIP[41]
  PIN SET_VCLIP[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6172.875 187.44 6173.155 188.44 ;
    END
  END SET_VCLIP[40]
  PIN SET_VCLIP[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6032.875 187.44 6033.155 188.44 ;
    END
  END SET_VCLIP[39]
  PIN SET_VCLIP[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5892.875 187.44 5893.155 188.44 ;
    END
  END SET_VCLIP[38]
  PIN SET_VCLIP[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5752.875 187.44 5753.155 188.44 ;
    END
  END SET_VCLIP[37]
  PIN SET_VCLIP[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5612.875 187.44 5613.155 188.44 ;
    END
  END SET_VCLIP[36]
  PIN SET_VCLIP[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5472.875 187.44 5473.155 188.44 ;
    END
  END SET_VCLIP[35]
  PIN SET_VCLIP[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5332.875 187.44 5333.155 188.44 ;
    END
  END SET_VCLIP[34]
  PIN SET_VCLIP[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5192.875 187.44 5193.155 188.44 ;
    END
  END SET_VCLIP[33]
  PIN SET_VCLIP[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5052.875 187.44 5053.155 188.44 ;
    END
  END SET_VCLIP[32]
  PIN SET_VCLIP[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4912.875 187.44 4913.155 188.44 ;
    END
  END SET_VCLIP[31]
  PIN SET_VCLIP[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4772.875 187.44 4773.155 188.44 ;
    END
  END SET_VCLIP[30]
  PIN SET_VCLIP[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4632.875 187.44 4633.155 188.44 ;
    END
  END SET_VCLIP[29]
  PIN SET_VCLIP[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4492.875 187.44 4493.155 188.44 ;
    END
  END SET_VCLIP[28]
  PIN SET_VCLIP[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4352.875 187.44 4353.155 188.44 ;
    END
  END SET_VCLIP[27]
  PIN SET_VCLIP[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4212.875 187.44 4213.155 188.44 ;
    END
  END SET_VCLIP[26]
  PIN SET_VCLIP[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4072.875 187.44 4073.155 188.44 ;
    END
  END SET_VCLIP[25]
  PIN SET_VCLIP[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3932.875 187.44 3933.155 188.44 ;
    END
  END SET_VCLIP[24]
  PIN SET_VCLIP[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3792.875 187.44 3793.155 188.44 ;
    END
  END SET_VCLIP[23]
  PIN SET_VCLIP[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3652.875 187.44 3653.155 188.44 ;
    END
  END SET_VCLIP[22]
  PIN SET_VCLIP[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3512.875 187.44 3513.155 188.44 ;
    END
  END SET_VCLIP[21]
  PIN SET_VCLIP[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3372.875 187.44 3373.155 188.44 ;
    END
  END SET_VCLIP[20]
  PIN SET_VCLIP[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3232.875 187.44 3233.155 188.44 ;
    END
  END SET_VCLIP[19]
  PIN SET_VCLIP[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3092.875 187.44 3093.155 188.44 ;
    END
  END SET_VCLIP[18]
  PIN SET_VCLIP[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2952.875 187.44 2953.155 188.44 ;
    END
  END SET_VCLIP[17]
  PIN SET_VCLIP[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2812.875 187.44 2813.155 188.44 ;
    END
  END SET_VCLIP[16]
  PIN SET_VCLIP[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2672.875 187.44 2673.155 188.44 ;
    END
  END SET_VCLIP[15]
  PIN SET_VCLIP[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2532.875 187.44 2533.155 188.44 ;
    END
  END SET_VCLIP[14]
  PIN SET_VCLIP[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2392.875 187.44 2393.155 188.44 ;
    END
  END SET_VCLIP[13]
  PIN SET_VCLIP[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2252.875 187.44 2253.155 188.44 ;
    END
  END SET_VCLIP[12]
  PIN SET_VCLIP[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2112.875 187.44 2113.155 188.44 ;
    END
  END SET_VCLIP[11]
  PIN SET_VCLIP[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1972.875 187.44 1973.155 188.44 ;
    END
  END SET_VCLIP[10]
  PIN SET_VCLIP[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1832.875 187.44 1833.155 188.44 ;
    END
  END SET_VCLIP[9]
  PIN SET_VCLIP[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1692.875 187.44 1693.155 188.44 ;
    END
  END SET_VCLIP[8]
  PIN SET_VCLIP[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1552.875 187.44 1553.155 188.44 ;
    END
  END SET_VCLIP[7]
  PIN SET_VCLIP[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1412.875 187.44 1413.155 188.44 ;
    END
  END SET_VCLIP[6]
  PIN SET_VCLIP[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1272.875 187.44 1273.155 188.44 ;
    END
  END SET_VCLIP[5]
  PIN SET_VCLIP[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1132.875 187.44 1133.155 188.44 ;
    END
  END SET_VCLIP[4]
  PIN SET_VCLIP[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 992.875 187.44 993.155 188.44 ;
    END
  END SET_VCLIP[3]
  PIN SET_VCLIP[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 852.875 187.44 853.155 188.44 ;
    END
  END SET_VCLIP[2]
  PIN SET_VCLIP[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 712.875 187.44 713.155 188.44 ;
    END
  END SET_VCLIP[1]
  PIN SET_VCLIP[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 572.875 187.44 573.155 188.44 ;
    END
  END SET_VCLIP[0]
  PIN GNDA_IDAC
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 326.66 261.245 327.66 289.275 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 261.245 18490.46 289.275 ;
    END
  END GNDA_IDAC
  PIN VDDA_IDAC
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 326.66 230.245 327.66 258.275 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 230.245 18490.46 258.275 ;
    END
  END VDDA_IDAC
  PIN VDDA_VDAC
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 326.66 292.245 327.66 306.275 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 213.245 327.66 227.275 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 292.245 18490.46 306.275 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 213.245 18490.46 227.275 ;
    END
  END VDDA_VDAC
  PIN SET_VRESET_P[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18349.235 187.44 18349.515 188.44 ;
    END
  END SET_VRESET_P[127]
  PIN SET_VRESET_P[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18209.235 187.44 18209.515 188.44 ;
    END
  END SET_VRESET_P[126]
  PIN SET_VRESET_P[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18069.235 187.44 18069.515 188.44 ;
    END
  END SET_VRESET_P[125]
  PIN SET_VRESET_P[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17929.235 187.44 17929.515 188.44 ;
    END
  END SET_VRESET_P[124]
  PIN SET_VRESET_P[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17789.235 187.44 17789.515 188.44 ;
    END
  END SET_VRESET_P[123]
  PIN SET_VRESET_P[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17649.235 187.44 17649.515 188.44 ;
    END
  END SET_VRESET_P[122]
  PIN SET_VRESET_P[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17509.235 187.44 17509.515 188.44 ;
    END
  END SET_VRESET_P[121]
  PIN SET_VRESET_P[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17369.235 187.44 17369.515 188.44 ;
    END
  END SET_VRESET_P[120]
  PIN SET_VRESET_P[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17229.235 187.44 17229.515 188.44 ;
    END
  END SET_VRESET_P[119]
  PIN SET_VRESET_P[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17089.235 187.44 17089.515 188.44 ;
    END
  END SET_VRESET_P[118]
  PIN SET_VRESET_P[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16949.235 187.44 16949.515 188.44 ;
    END
  END SET_VRESET_P[117]
  PIN SET_VRESET_P[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16809.235 187.44 16809.515 188.44 ;
    END
  END SET_VRESET_P[116]
  PIN SET_VRESET_P[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16669.235 187.44 16669.515 188.44 ;
    END
  END SET_VRESET_P[115]
  PIN SET_VRESET_P[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16529.235 187.44 16529.515 188.44 ;
    END
  END SET_VRESET_P[114]
  PIN SET_VRESET_P[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16389.235 187.44 16389.515 188.44 ;
    END
  END SET_VRESET_P[113]
  PIN SET_VRESET_P[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16249.235 187.44 16249.515 188.44 ;
    END
  END SET_VRESET_P[112]
  PIN SET_VRESET_P[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16109.235 187.44 16109.515 188.44 ;
    END
  END SET_VRESET_P[111]
  PIN SET_VRESET_P[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15969.235 187.44 15969.515 188.44 ;
    END
  END SET_VRESET_P[110]
  PIN SET_VRESET_P[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15829.235 187.44 15829.515 188.44 ;
    END
  END SET_VRESET_P[109]
  PIN SET_VRESET_P[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15689.235 187.44 15689.515 188.44 ;
    END
  END SET_VRESET_P[108]
  PIN SET_VRESET_P[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15549.235 187.44 15549.515 188.44 ;
    END
  END SET_VRESET_P[107]
  PIN SET_VRESET_P[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15409.235 187.44 15409.515 188.44 ;
    END
  END SET_VRESET_P[106]
  PIN SET_VRESET_P[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15269.235 187.44 15269.515 188.44 ;
    END
  END SET_VRESET_P[105]
  PIN SET_VRESET_P[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15129.235 187.44 15129.515 188.44 ;
    END
  END SET_VRESET_P[104]
  PIN SET_VRESET_P[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14989.235 187.44 14989.515 188.44 ;
    END
  END SET_VRESET_P[103]
  PIN SET_VRESET_P[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14849.235 187.44 14849.515 188.44 ;
    END
  END SET_VRESET_P[102]
  PIN SET_VRESET_P[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14709.235 187.44 14709.515 188.44 ;
    END
  END SET_VRESET_P[101]
  PIN SET_VRESET_P[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14569.235 187.44 14569.515 188.44 ;
    END
  END SET_VRESET_P[100]
  PIN SET_VRESET_P[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14429.235 187.44 14429.515 188.44 ;
    END
  END SET_VRESET_P[99]
  PIN SET_VRESET_P[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14289.235 187.44 14289.515 188.44 ;
    END
  END SET_VRESET_P[98]
  PIN SET_VRESET_P[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14149.235 187.44 14149.515 188.44 ;
    END
  END SET_VRESET_P[97]
  PIN SET_VRESET_P[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14009.235 187.44 14009.515 188.44 ;
    END
  END SET_VRESET_P[96]
  PIN SET_VRESET_P[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13869.235 187.44 13869.515 188.44 ;
    END
  END SET_VRESET_P[95]
  PIN SET_VRESET_P[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13729.235 187.44 13729.515 188.44 ;
    END
  END SET_VRESET_P[94]
  PIN SET_VRESET_P[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13589.235 187.44 13589.515 188.44 ;
    END
  END SET_VRESET_P[93]
  PIN SET_VRESET_P[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13449.235 187.44 13449.515 188.44 ;
    END
  END SET_VRESET_P[92]
  PIN SET_VRESET_P[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13309.235 187.44 13309.515 188.44 ;
    END
  END SET_VRESET_P[91]
  PIN SET_VRESET_P[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13169.235 187.44 13169.515 188.44 ;
    END
  END SET_VRESET_P[90]
  PIN SET_VRESET_P[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13029.235 187.44 13029.515 188.44 ;
    END
  END SET_VRESET_P[89]
  PIN SET_VRESET_P[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12889.235 187.44 12889.515 188.44 ;
    END
  END SET_VRESET_P[88]
  PIN SET_VRESET_P[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12749.235 187.44 12749.515 188.44 ;
    END
  END SET_VRESET_P[87]
  PIN SET_VRESET_P[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12609.235 187.44 12609.515 188.44 ;
    END
  END SET_VRESET_P[86]
  PIN SET_VRESET_P[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12469.235 187.44 12469.515 188.44 ;
    END
  END SET_VRESET_P[85]
  PIN SET_VRESET_P[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12329.235 187.44 12329.515 188.44 ;
    END
  END SET_VRESET_P[84]
  PIN SET_VRESET_P[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12189.235 187.44 12189.515 188.44 ;
    END
  END SET_VRESET_P[83]
  PIN SET_VRESET_P[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12049.235 187.44 12049.515 188.44 ;
    END
  END SET_VRESET_P[82]
  PIN SET_VRESET_P[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11909.235 187.44 11909.515 188.44 ;
    END
  END SET_VRESET_P[81]
  PIN SET_VRESET_P[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11769.235 187.44 11769.515 188.44 ;
    END
  END SET_VRESET_P[80]
  PIN SET_VRESET_P[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11629.235 187.44 11629.515 188.44 ;
    END
  END SET_VRESET_P[79]
  PIN SET_VRESET_P[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11489.235 187.44 11489.515 188.44 ;
    END
  END SET_VRESET_P[78]
  PIN SET_VRESET_P[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11349.235 187.44 11349.515 188.44 ;
    END
  END SET_VRESET_P[77]
  PIN SET_VRESET_P[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11209.235 187.44 11209.515 188.44 ;
    END
  END SET_VRESET_P[76]
  PIN SET_VRESET_P[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11069.235 187.44 11069.515 188.44 ;
    END
  END SET_VRESET_P[75]
  PIN SET_VRESET_P[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10929.235 187.44 10929.515 188.44 ;
    END
  END SET_VRESET_P[74]
  PIN SET_VRESET_P[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10789.235 187.44 10789.515 188.44 ;
    END
  END SET_VRESET_P[73]
  PIN SET_VRESET_P[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10649.235 187.44 10649.515 188.44 ;
    END
  END SET_VRESET_P[72]
  PIN SET_VRESET_P[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10509.235 187.44 10509.515 188.44 ;
    END
  END SET_VRESET_P[71]
  PIN SET_VRESET_P[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10369.235 187.44 10369.515 188.44 ;
    END
  END SET_VRESET_P[70]
  PIN SET_VRESET_P[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10229.235 187.44 10229.515 188.44 ;
    END
  END SET_VRESET_P[69]
  PIN SET_VRESET_P[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10089.235 187.44 10089.515 188.44 ;
    END
  END SET_VRESET_P[68]
  PIN SET_VRESET_P[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9949.235 187.44 9949.515 188.44 ;
    END
  END SET_VRESET_P[67]
  PIN SET_VRESET_P[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9809.235 187.44 9809.515 188.44 ;
    END
  END SET_VRESET_P[66]
  PIN SET_VRESET_P[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9669.235 187.44 9669.515 188.44 ;
    END
  END SET_VRESET_P[65]
  PIN SET_VRESET_P[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9529.235 187.44 9529.515 188.44 ;
    END
  END SET_VRESET_P[64]
  PIN SET_VRESET_P[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9389.235 187.44 9389.515 188.44 ;
    END
  END SET_VRESET_P[63]
  PIN SET_VRESET_P[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9249.235 187.44 9249.515 188.44 ;
    END
  END SET_VRESET_P[62]
  PIN SET_VRESET_P[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9109.235 187.44 9109.515 188.44 ;
    END
  END SET_VRESET_P[61]
  PIN SET_VRESET_P[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8969.235 187.44 8969.515 188.44 ;
    END
  END SET_VRESET_P[60]
  PIN SET_VRESET_P[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8829.235 187.44 8829.515 188.44 ;
    END
  END SET_VRESET_P[59]
  PIN SET_VRESET_P[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8689.235 187.44 8689.515 188.44 ;
    END
  END SET_VRESET_P[58]
  PIN SET_VRESET_P[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8549.235 187.44 8549.515 188.44 ;
    END
  END SET_VRESET_P[57]
  PIN SET_VRESET_P[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8409.235 187.44 8409.515 188.44 ;
    END
  END SET_VRESET_P[56]
  PIN SET_VRESET_P[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8269.235 187.44 8269.515 188.44 ;
    END
  END SET_VRESET_P[55]
  PIN SET_VRESET_P[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8129.235 187.44 8129.515 188.44 ;
    END
  END SET_VRESET_P[54]
  PIN SET_VRESET_P[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7989.235 187.44 7989.515 188.44 ;
    END
  END SET_VRESET_P[53]
  PIN SET_VRESET_P[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7849.235 187.44 7849.515 188.44 ;
    END
  END SET_VRESET_P[52]
  PIN SET_VRESET_P[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7709.235 187.44 7709.515 188.44 ;
    END
  END SET_VRESET_P[51]
  PIN SET_VRESET_P[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7569.235 187.44 7569.515 188.44 ;
    END
  END SET_VRESET_P[50]
  PIN SET_VRESET_P[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7429.235 187.44 7429.515 188.44 ;
    END
  END SET_VRESET_P[49]
  PIN SET_VRESET_P[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7289.235 187.44 7289.515 188.44 ;
    END
  END SET_VRESET_P[48]
  PIN SET_VRESET_P[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7149.235 187.44 7149.515 188.44 ;
    END
  END SET_VRESET_P[47]
  PIN SET_VRESET_P[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7009.235 187.44 7009.515 188.44 ;
    END
  END SET_VRESET_P[46]
  PIN SET_VRESET_P[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6869.235 187.44 6869.515 188.44 ;
    END
  END SET_VRESET_P[45]
  PIN SET_VRESET_P[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6729.235 187.44 6729.515 188.44 ;
    END
  END SET_VRESET_P[44]
  PIN SET_VRESET_P[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6589.235 187.44 6589.515 188.44 ;
    END
  END SET_VRESET_P[43]
  PIN SET_VRESET_P[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6449.235 187.44 6449.515 188.44 ;
    END
  END SET_VRESET_P[42]
  PIN SET_VRESET_P[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6309.235 187.44 6309.515 188.44 ;
    END
  END SET_VRESET_P[41]
  PIN SET_VRESET_P[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6169.235 187.44 6169.515 188.44 ;
    END
  END SET_VRESET_P[40]
  PIN SET_VRESET_P[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6029.235 187.44 6029.515 188.44 ;
    END
  END SET_VRESET_P[39]
  PIN SET_VRESET_P[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5889.235 187.44 5889.515 188.44 ;
    END
  END SET_VRESET_P[38]
  PIN SET_VCASN[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18216.515 187.44 18216.795 188.44 ;
    END
  END SET_VCASN[126]
  PIN SET_VCASN[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18076.515 187.44 18076.795 188.44 ;
    END
  END SET_VCASN[125]
  PIN SET_VCASN[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17936.515 187.44 17936.795 188.44 ;
    END
  END SET_VCASN[124]
  PIN SET_VCASN[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17796.515 187.44 17796.795 188.44 ;
    END
  END SET_VCASN[123]
  PIN SET_VCASN[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17656.515 187.44 17656.795 188.44 ;
    END
  END SET_VCASN[122]
  PIN SET_VCASN[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17516.515 187.44 17516.795 188.44 ;
    END
  END SET_VCASN[121]
  PIN SET_VCASN[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17376.515 187.44 17376.795 188.44 ;
    END
  END SET_VCASN[120]
  PIN SET_VCASN[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17236.515 187.44 17236.795 188.44 ;
    END
  END SET_VCASN[119]
  PIN SET_VCASN[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17096.515 187.44 17096.795 188.44 ;
    END
  END SET_VCASN[118]
  PIN SET_VCASN[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16956.515 187.44 16956.795 188.44 ;
    END
  END SET_VCASN[117]
  PIN SET_VCASN[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16816.515 187.44 16816.795 188.44 ;
    END
  END SET_VCASN[116]
  PIN SET_VCASN[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16676.515 187.44 16676.795 188.44 ;
    END
  END SET_VCASN[115]
  PIN SET_VCASN[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16536.515 187.44 16536.795 188.44 ;
    END
  END SET_VCASN[114]
  PIN SET_VCASN[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16396.515 187.44 16396.795 188.44 ;
    END
  END SET_VCASN[113]
  PIN SET_VCASN[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16256.515 187.44 16256.795 188.44 ;
    END
  END SET_VCASN[112]
  PIN SET_VCASN[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16116.515 187.44 16116.795 188.44 ;
    END
  END SET_VCASN[111]
  PIN SET_VCASN[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15976.515 187.44 15976.795 188.44 ;
    END
  END SET_VCASN[110]
  PIN SET_VCASN[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15836.515 187.44 15836.795 188.44 ;
    END
  END SET_VCASN[109]
  PIN SET_VCASN[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15696.515 187.44 15696.795 188.44 ;
    END
  END SET_VCASN[108]
  PIN SET_VCASN[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15556.515 187.44 15556.795 188.44 ;
    END
  END SET_VCASN[107]
  PIN SET_VCASN[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15416.515 187.44 15416.795 188.44 ;
    END
  END SET_VCASN[106]
  PIN SET_VCASN[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15276.515 187.44 15276.795 188.44 ;
    END
  END SET_VCASN[105]
  PIN SET_VCASN[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15136.515 187.44 15136.795 188.44 ;
    END
  END SET_VCASN[104]
  PIN SET_VCASN[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14996.515 187.44 14996.795 188.44 ;
    END
  END SET_VCASN[103]
  PIN SET_VCASN[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14856.515 187.44 14856.795 188.44 ;
    END
  END SET_VCASN[102]
  PIN SET_VCASN[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14716.515 187.44 14716.795 188.44 ;
    END
  END SET_VCASN[101]
  PIN SET_VCASN[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14576.515 187.44 14576.795 188.44 ;
    END
  END SET_VCASN[100]
  PIN SET_VCASN[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14436.515 187.44 14436.795 188.44 ;
    END
  END SET_VCASN[99]
  PIN SET_VCASN[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14296.515 187.44 14296.795 188.44 ;
    END
  END SET_VCASN[98]
  PIN SET_VCASN[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14156.515 187.44 14156.795 188.44 ;
    END
  END SET_VCASN[97]
  PIN SET_VCASN[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14016.515 187.44 14016.795 188.44 ;
    END
  END SET_VCASN[96]
  PIN SET_VCASN[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13876.515 187.44 13876.795 188.44 ;
    END
  END SET_VCASN[95]
  PIN SET_VCASN[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13736.515 187.44 13736.795 188.44 ;
    END
  END SET_VCASN[94]
  PIN SET_VCASN[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13036.515 187.44 13036.795 188.44 ;
    END
  END SET_VCASN[89]
  PIN SET_VCASN[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13456.515 187.44 13456.795 188.44 ;
    END
  END SET_VCASN[92]
  PIN SET_VCASN[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13316.515 187.44 13316.795 188.44 ;
    END
  END SET_VCASN[91]
  PIN SET_VCASN[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13176.515 187.44 13176.795 188.44 ;
    END
  END SET_VCASN[90]
  PIN SET_VCASN[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12896.515 187.44 12896.795 188.44 ;
    END
  END SET_VCASN[88]
  PIN SET_VCASN[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12756.515 187.44 12756.795 188.44 ;
    END
  END SET_VCASN[87]
  PIN SET_VCASN[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12616.515 187.44 12616.795 188.44 ;
    END
  END SET_VCASN[86]
  PIN SET_VCASN[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12476.515 187.44 12476.795 188.44 ;
    END
  END SET_VCASN[85]
  PIN SET_VCASN[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12336.515 187.44 12336.795 188.44 ;
    END
  END SET_VCASN[84]
  PIN SET_VCASN[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12196.515 187.44 12196.795 188.44 ;
    END
  END SET_VCASN[83]
  PIN SET_VCASN[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12056.515 187.44 12056.795 188.44 ;
    END
  END SET_VCASN[82]
  PIN SET_VCASN[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11916.515 187.44 11916.795 188.44 ;
    END
  END SET_VCASN[81]
  PIN SET_VCASN[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11776.515 187.44 11776.795 188.44 ;
    END
  END SET_VCASN[80]
  PIN SET_VCASN[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11636.515 187.44 11636.795 188.44 ;
    END
  END SET_VCASN[79]
  PIN SET_VCASN[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11496.515 187.44 11496.795 188.44 ;
    END
  END SET_VCASN[78]
  PIN SET_VCASN[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11356.515 187.44 11356.795 188.44 ;
    END
  END SET_VCASN[77]
  PIN SET_VCASN[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11216.515 187.44 11216.795 188.44 ;
    END
  END SET_VCASN[76]
  PIN SET_VCASN[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11076.515 187.44 11076.795 188.44 ;
    END
  END SET_VCASN[75]
  PIN SET_VCASN[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10936.515 187.44 10936.795 188.44 ;
    END
  END SET_VCASN[74]
  PIN SET_VCASN[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10796.515 187.44 10796.795 188.44 ;
    END
  END SET_VCASN[73]
  PIN SET_VCASN[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10656.515 187.44 10656.795 188.44 ;
    END
  END SET_VCASN[72]
  PIN SET_VCASN[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10516.515 187.44 10516.795 188.44 ;
    END
  END SET_VCASN[71]
  PIN SET_VCASN[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10376.515 187.44 10376.795 188.44 ;
    END
  END SET_VCASN[70]
  PIN SET_VCASN[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10236.515 187.44 10236.795 188.44 ;
    END
  END SET_VCASN[69]
  PIN SET_VCASN[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10096.515 187.44 10096.795 188.44 ;
    END
  END SET_VCASN[68]
  PIN SET_VCASN[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9956.515 187.44 9956.795 188.44 ;
    END
  END SET_VCASN[67]
  PIN SET_VCASN[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9816.515 187.44 9816.795 188.44 ;
    END
  END SET_VCASN[66]
  PIN SET_VCASN[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9676.515 187.44 9676.795 188.44 ;
    END
  END SET_VCASN[65]
  PIN SET_VCASN[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9536.515 187.44 9536.795 188.44 ;
    END
  END SET_VCASN[64]
  PIN SET_VCASN[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9396.515 187.44 9396.795 188.44 ;
    END
  END SET_VCASN[63]
  PIN SET_VCASN[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9256.515 187.44 9256.795 188.44 ;
    END
  END SET_VCASN[62]
  PIN SET_VCASN[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9116.515 187.44 9116.795 188.44 ;
    END
  END SET_VCASN[61]
  PIN SET_VCASN[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8976.515 187.44 8976.795 188.44 ;
    END
  END SET_VCASN[60]
  PIN SET_VCASN[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8836.515 187.44 8836.795 188.44 ;
    END
  END SET_VCASN[59]
  PIN SET_VCASN[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8696.515 187.44 8696.795 188.44 ;
    END
  END SET_VCASN[58]
  PIN SET_VCASN[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8556.515 187.44 8556.795 188.44 ;
    END
  END SET_VCASN[57]
  PIN SET_VCASN[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8416.515 187.44 8416.795 188.44 ;
    END
  END SET_VCASN[56]
  PIN SET_VCASN[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8276.515 187.44 8276.795 188.44 ;
    END
  END SET_VCASN[55]
  PIN SET_VCASN[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8136.515 187.44 8136.795 188.44 ;
    END
  END SET_VCASN[54]
  PIN SET_VCASN[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7996.515 187.44 7996.795 188.44 ;
    END
  END SET_VCASN[53]
  PIN SET_VCASN[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7856.515 187.44 7856.795 188.44 ;
    END
  END SET_VCASN[52]
  PIN SET_VCASN[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7716.515 187.44 7716.795 188.44 ;
    END
  END SET_VCASN[51]
  PIN SET_VCASN[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7576.515 187.44 7576.795 188.44 ;
    END
  END SET_VCASN[50]
  PIN SET_VCASN[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7436.515 187.44 7436.795 188.44 ;
    END
  END SET_VCASN[49]
  PIN SET_VCASN[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7296.515 187.44 7296.795 188.44 ;
    END
  END SET_VCASN[48]
  PIN SET_VCASN[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7156.515 187.44 7156.795 188.44 ;
    END
  END SET_VCASN[47]
  PIN SET_VCASN[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7016.515 187.44 7016.795 188.44 ;
    END
  END SET_VCASN[46]
  PIN SET_VCASN[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6876.515 187.44 6876.795 188.44 ;
    END
  END SET_VCASN[45]
  PIN SET_VCASN[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6736.515 187.44 6736.795 188.44 ;
    END
  END SET_VCASN[44]
  PIN SET_VCASN[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6596.515 187.44 6596.795 188.44 ;
    END
  END SET_VCASN[43]
  PIN SET_VCASN[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6456.515 187.44 6456.795 188.44 ;
    END
  END SET_VCASN[42]
  PIN SET_VCASN[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6316.515 187.44 6316.795 188.44 ;
    END
  END SET_VCASN[41]
  PIN SET_VCASN[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6176.515 187.44 6176.795 188.44 ;
    END
  END SET_VCASN[40]
  PIN SET_VCASN[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6036.515 187.44 6036.795 188.44 ;
    END
  END SET_VCASN[39]
  PIN SET_VCASN[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5896.515 187.44 5896.795 188.44 ;
    END
  END SET_VCASN[38]
  PIN SET_VCASN[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5756.515 187.44 5756.795 188.44 ;
    END
  END SET_VCASN[37]
  PIN SET_VCASN[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5616.515 187.44 5616.795 188.44 ;
    END
  END SET_VCASN[36]
  PIN SET_VCASN[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5476.515 187.44 5476.795 188.44 ;
    END
  END SET_VCASN[35]
  PIN SET_VCASN[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5336.515 187.44 5336.795 188.44 ;
    END
  END SET_VCASN[34]
  PIN SET_VCASN[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5196.515 187.44 5196.795 188.44 ;
    END
  END SET_VCASN[33]
  PIN SET_VCASN[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5056.515 187.44 5056.795 188.44 ;
    END
  END SET_VCASN[32]
  PIN SET_VCASN[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4916.515 187.44 4916.795 188.44 ;
    END
  END SET_VCASN[31]
  PIN SET_VCASN[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4776.515 187.44 4776.795 188.44 ;
    END
  END SET_VCASN[30]
  PIN SET_VCASN[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4636.515 187.44 4636.795 188.44 ;
    END
  END SET_VCASN[29]
  PIN SET_VCASN[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4496.515 187.44 4496.795 188.44 ;
    END
  END SET_VCASN[28]
  PIN SET_VCASN[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4356.515 187.44 4356.795 188.44 ;
    END
  END SET_VCASN[27]
  PIN SET_VCASN[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4216.515 187.44 4216.795 188.44 ;
    END
  END SET_VCASN[26]
  PIN SET_VCASN[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4076.515 187.44 4076.795 188.44 ;
    END
  END SET_VCASN[25]
  PIN SET_VCASN[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3936.515 187.44 3936.795 188.44 ;
    END
  END SET_VCASN[24]
  PIN SET_VCASN[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3796.515 187.44 3796.795 188.44 ;
    END
  END SET_VCASN[23]
  PIN SET_VCASN[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3656.515 187.44 3656.795 188.44 ;
    END
  END SET_VCASN[22]
  PIN SET_VCASN[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3516.515 187.44 3516.795 188.44 ;
    END
  END SET_VCASN[21]
  PIN SET_VCASN[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3376.515 187.44 3376.795 188.44 ;
    END
  END SET_VCASN[20]
  PIN SET_VCASN[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3236.515 187.44 3236.795 188.44 ;
    END
  END SET_VCASN[19]
  PIN SET_VCASN[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3096.515 187.44 3096.795 188.44 ;
    END
  END SET_VCASN[18]
  PIN SET_VCASN[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2956.515 187.44 2956.795 188.44 ;
    END
  END SET_VCASN[17]
  PIN SET_VCASN[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2816.515 187.44 2816.795 188.44 ;
    END
  END SET_VCASN[16]
  PIN SET_VCASN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2676.515 187.44 2676.795 188.44 ;
    END
  END SET_VCASN[15]
  PIN SET_VCASN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2536.515 187.44 2536.795 188.44 ;
    END
  END SET_VCASN[14]
  PIN SET_VCASN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2396.515 187.44 2396.795 188.44 ;
    END
  END SET_VCASN[13]
  PIN SET_VCASN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2256.515 187.44 2256.795 188.44 ;
    END
  END SET_VCASN[12]
  PIN SET_VCASN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2116.515 187.44 2116.795 188.44 ;
    END
  END SET_VCASN[11]
  PIN SET_VCASN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1976.515 187.44 1976.795 188.44 ;
    END
  END SET_VCASN[10]
  PIN SET_VCASN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1836.515 187.44 1836.795 188.44 ;
    END
  END SET_VCASN[9]
  PIN SET_VCASN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1696.515 187.44 1696.795 188.44 ;
    END
  END SET_VCASN[8]
  PIN SET_VCASN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1556.515 187.44 1556.795 188.44 ;
    END
  END SET_VCASN[7]
  PIN SET_VCASN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1416.515 187.44 1416.795 188.44 ;
    END
  END SET_VCASN[6]
  PIN SET_VCASN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1276.515 187.44 1276.795 188.44 ;
    END
  END SET_VCASN[5]
  PIN SET_VCASN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1136.515 187.44 1136.795 188.44 ;
    END
  END SET_VCASN[4]
  PIN SET_VCASN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 996.515 187.44 996.795 188.44 ;
    END
  END SET_VCASN[3]
  PIN SET_VCASN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 856.515 187.44 856.795 188.44 ;
    END
  END SET_VCASN[2]
  PIN SET_VCASN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 716.515 187.44 716.795 188.44 ;
    END
  END SET_VCASN[1]
  PIN SET_VCASN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 576.515 187.44 576.795 188.44 ;
    END
  END SET_VCASN[0]
  PIN SET_VCASN[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13596.515 187.44 13596.795 188.44 ;
    END
  END SET_VCASN[93]
  PIN SET_VRESET_P[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5749.235 187.44 5749.515 188.44 ;
    END
  END SET_VRESET_P[37]
  PIN SET_VRESET_P[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5609.235 187.44 5609.515 188.44 ;
    END
  END SET_VRESET_P[36]
  PIN SET_VRESET_P[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5469.235 187.44 5469.515 188.44 ;
    END
  END SET_VRESET_P[35]
  PIN SET_VRESET_P[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5329.235 187.44 5329.515 188.44 ;
    END
  END SET_VRESET_P[34]
  PIN SET_VRESET_P[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5189.235 187.44 5189.515 188.44 ;
    END
  END SET_VRESET_P[33]
  PIN SET_VRESET_P[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5049.235 187.44 5049.515 188.44 ;
    END
  END SET_VRESET_P[32]
  PIN SET_VRESET_P[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4909.235 187.44 4909.515 188.44 ;
    END
  END SET_VRESET_P[31]
  PIN SET_VRESET_P[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4769.235 187.44 4769.515 188.44 ;
    END
  END SET_VRESET_P[30]
  PIN SET_VRESET_P[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4629.235 187.44 4629.515 188.44 ;
    END
  END SET_VRESET_P[29]
  PIN SET_VRESET_P[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4489.235 187.44 4489.515 188.44 ;
    END
  END SET_VRESET_P[28]
  PIN SET_VRESET_P[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4349.235 187.44 4349.515 188.44 ;
    END
  END SET_VRESET_P[27]
  PIN SET_VRESET_P[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4209.235 187.44 4209.515 188.44 ;
    END
  END SET_VRESET_P[26]
  PIN SET_VRESET_P[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4069.235 187.44 4069.515 188.44 ;
    END
  END SET_VRESET_P[25]
  PIN SET_VRESET_P[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3929.235 187.44 3929.515 188.44 ;
    END
  END SET_VRESET_P[24]
  PIN SET_VRESET_P[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3789.235 187.44 3789.515 188.44 ;
    END
  END SET_VRESET_P[23]
  PIN SET_VRESET_P[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3649.235 187.44 3649.515 188.44 ;
    END
  END SET_VRESET_P[22]
  PIN SET_VRESET_P[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3509.235 187.44 3509.515 188.44 ;
    END
  END SET_VRESET_P[21]
  PIN SET_VRESET_P[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3369.235 187.44 3369.515 188.44 ;
    END
  END SET_VRESET_P[20]
  PIN SET_VRESET_P[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3229.235 187.44 3229.515 188.44 ;
    END
  END SET_VRESET_P[19]
  PIN SET_VRESET_P[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3089.235 187.44 3089.515 188.44 ;
    END
  END SET_VRESET_P[18]
  PIN SET_VRESET_P[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2949.235 187.44 2949.515 188.44 ;
    END
  END SET_VRESET_P[17]
  PIN SET_VRESET_P[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2809.235 187.44 2809.515 188.44 ;
    END
  END SET_VRESET_P[16]
  PIN SET_VRESET_P[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2669.235 187.44 2669.515 188.44 ;
    END
  END SET_VRESET_P[15]
  PIN SET_VRESET_P[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2529.235 187.44 2529.515 188.44 ;
    END
  END SET_VRESET_P[14]
  PIN SET_VRESET_P[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2389.235 187.44 2389.515 188.44 ;
    END
  END SET_VRESET_P[13]
  PIN SET_VRESET_P[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2249.235 187.44 2249.515 188.44 ;
    END
  END SET_VRESET_P[12]
  PIN SET_VRESET_P[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2109.235 187.44 2109.515 188.44 ;
    END
  END SET_VRESET_P[11]
  PIN SET_VRESET_P[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1969.235 187.44 1969.515 188.44 ;
    END
  END SET_VRESET_P[10]
  PIN SET_VRESET_P[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1829.235 187.44 1829.515 188.44 ;
    END
  END SET_VRESET_P[9]
  PIN SET_VRESET_P[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1689.235 187.44 1689.515 188.44 ;
    END
  END SET_VRESET_P[8]
  PIN SET_VRESET_P[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1549.235 187.44 1549.515 188.44 ;
    END
  END SET_VRESET_P[7]
  PIN SET_VRESET_P[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1409.235 187.44 1409.515 188.44 ;
    END
  END SET_VRESET_P[6]
  PIN SET_VRESET_P[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1269.235 187.44 1269.515 188.44 ;
    END
  END SET_VRESET_P[5]
  PIN SET_VRESET_P[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1129.235 187.44 1129.515 188.44 ;
    END
  END SET_VRESET_P[4]
  PIN SET_VRESET_P[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 989.235 187.44 989.515 188.44 ;
    END
  END SET_VRESET_P[3]
  PIN SET_VRESET_P[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 849.235 187.44 849.515 188.44 ;
    END
  END SET_VRESET_P[2]
  PIN SET_VRESET_P[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 709.235 187.44 709.515 188.44 ;
    END
  END SET_VRESET_P[1]
  PIN SET_VRESET_P[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 569.235 187.44 569.515 188.44 ;
    END
  END SET_VRESET_P[0]
  PIN SET_VH[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18345.595 187.44 18345.875 188.44 ;
    END
  END SET_VH[127]
  PIN SET_VH[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18205.595 187.44 18205.875 188.44 ;
    END
  END SET_VH[126]
  PIN SWCNTL_IDB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9411.475 187.44 9412.035 188.44 ;
    END
  END SWCNTL_IDB
  PIN SET_VH[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18065.595 187.44 18065.875 188.44 ;
    END
  END SET_VH[125]
  PIN SET_VH[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17925.595 187.44 17925.875 188.44 ;
    END
  END SET_VH[124]
  PIN SET_VH[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17785.595 187.44 17785.875 188.44 ;
    END
  END SET_VH[123]
  PIN SET_VH[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17645.595 187.44 17645.875 188.44 ;
    END
  END SET_VH[122]
  PIN SET_VH[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17505.595 187.44 17505.875 188.44 ;
    END
  END SET_VH[121]
  PIN SET_VH[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17365.595 187.44 17365.875 188.44 ;
    END
  END SET_VH[120]
  PIN SET_VH[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17225.595 187.44 17225.875 188.44 ;
    END
  END SET_VH[119]
  PIN SET_VH[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17085.595 187.44 17085.875 188.44 ;
    END
  END SET_VH[118]
  PIN SET_VH[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16945.595 187.44 16945.875 188.44 ;
    END
  END SET_VH[117]
  PIN SET_VH[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16805.595 187.44 16805.875 188.44 ;
    END
  END SET_VH[116]
  PIN SET_VH[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16665.595 187.44 16665.875 188.44 ;
    END
  END SET_VH[115]
  PIN SET_VH[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16525.595 187.44 16525.875 188.44 ;
    END
  END SET_VH[114]
  PIN SET_VH[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16385.595 187.44 16385.875 188.44 ;
    END
  END SET_VH[113]
  PIN SET_VH[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16245.595 187.44 16245.875 188.44 ;
    END
  END SET_VH[112]
  PIN SET_VH[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16105.595 187.44 16105.875 188.44 ;
    END
  END SET_VH[111]
  PIN SET_VH[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15965.595 187.44 15965.875 188.44 ;
    END
  END SET_VH[110]
  PIN SET_VH[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15825.595 187.44 15825.875 188.44 ;
    END
  END SET_VH[109]
  PIN SET_VH[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15685.595 187.44 15685.875 188.44 ;
    END
  END SET_VH[108]
  PIN SET_VH[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15545.595 187.44 15545.875 188.44 ;
    END
  END SET_VH[107]
  PIN SET_VH[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15405.595 187.44 15405.875 188.44 ;
    END
  END SET_VH[106]
  PIN SET_VH[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15265.595 187.44 15265.875 188.44 ;
    END
  END SET_VH[105]
  PIN SET_VH[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15125.595 187.44 15125.875 188.44 ;
    END
  END SET_VH[104]
  PIN SET_VH[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14985.595 187.44 14985.875 188.44 ;
    END
  END SET_VH[103]
  PIN SET_VH[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14845.595 187.44 14845.875 188.44 ;
    END
  END SET_VH[102]
  PIN SET_VH[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14705.595 187.44 14705.875 188.44 ;
    END
  END SET_VH[101]
  PIN SET_VH[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14565.595 187.44 14565.875 188.44 ;
    END
  END SET_VH[100]
  PIN SET_VH[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14425.595 187.44 14425.875 188.44 ;
    END
  END SET_VH[99]
  PIN SET_VH[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14285.595 187.44 14285.875 188.44 ;
    END
  END SET_VH[98]
  PIN SET_VH[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14145.595 187.44 14145.875 188.44 ;
    END
  END SET_VH[97]
  PIN SET_VH[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14005.595 187.44 14005.875 188.44 ;
    END
  END SET_VH[96]
  PIN SET_VH[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13865.595 187.44 13865.875 188.44 ;
    END
  END SET_VH[95]
  PIN SET_VH[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13725.595 187.44 13725.875 188.44 ;
    END
  END SET_VH[94]
  PIN SET_VH[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13585.595 187.44 13585.875 188.44 ;
    END
  END SET_VH[93]
  PIN SET_VH[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13445.595 187.44 13445.875 188.44 ;
    END
  END SET_VH[92]
  PIN SET_VH[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13305.595 187.44 13305.875 188.44 ;
    END
  END SET_VH[91]
  PIN SET_VH[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13165.595 187.44 13165.875 188.44 ;
    END
  END SET_VH[90]
  PIN SET_VH[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13025.595 187.44 13025.875 188.44 ;
    END
  END SET_VH[89]
  PIN SET_VH[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12885.595 187.44 12885.875 188.44 ;
    END
  END SET_VH[88]
  PIN SET_VH[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12745.595 187.44 12745.875 188.44 ;
    END
  END SET_VH[87]
  PIN SET_VH[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12605.595 187.44 12605.875 188.44 ;
    END
  END SET_VH[86]
  PIN SET_VH[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12465.595 187.44 12465.875 188.44 ;
    END
  END SET_VH[85]
  PIN SET_VH[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12325.595 187.44 12325.875 188.44 ;
    END
  END SET_VH[84]
  PIN SET_VH[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12185.595 187.44 12185.875 188.44 ;
    END
  END SET_VH[83]
  PIN SET_VH[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12045.595 187.44 12045.875 188.44 ;
    END
  END SET_VH[82]
  PIN SET_VH[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11905.595 187.44 11905.875 188.44 ;
    END
  END SET_VH[81]
  PIN SET_VH[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11765.595 187.44 11765.875 188.44 ;
    END
  END SET_VH[80]
  PIN SET_VH[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11625.595 187.44 11625.875 188.44 ;
    END
  END SET_VH[79]
  PIN SET_VH[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11485.595 187.44 11485.875 188.44 ;
    END
  END SET_VH[78]
  PIN SET_VH[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11345.595 187.44 11345.875 188.44 ;
    END
  END SET_VH[77]
  PIN SET_VH[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11205.595 187.44 11205.875 188.44 ;
    END
  END SET_VH[76]
  PIN SET_VH[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11065.595 187.44 11065.875 188.44 ;
    END
  END SET_VH[75]
  PIN SET_VH[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10925.595 187.44 10925.875 188.44 ;
    END
  END SET_VH[74]
  PIN SET_VH[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10785.595 187.44 10785.875 188.44 ;
    END
  END SET_VH[73]
  PIN SET_VH[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10645.595 187.44 10645.875 188.44 ;
    END
  END SET_VH[72]
  PIN SET_VH[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10505.595 187.44 10505.875 188.44 ;
    END
  END SET_VH[71]
  PIN SET_VH[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10365.595 187.44 10365.875 188.44 ;
    END
  END SET_VH[70]
  PIN SET_VH[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10225.595 187.44 10225.875 188.44 ;
    END
  END SET_VH[69]
  PIN SET_VH[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10085.595 187.44 10085.875 188.44 ;
    END
  END SET_VH[68]
  PIN SET_VH[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9945.595 187.44 9945.875 188.44 ;
    END
  END SET_VH[67]
  PIN SET_VH[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9805.595 187.44 9805.875 188.44 ;
    END
  END SET_VH[66]
  PIN SET_VH[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9665.595 187.44 9665.875 188.44 ;
    END
  END SET_VH[65]
  PIN SET_VH[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9525.595 187.44 9525.875 188.44 ;
    END
  END SET_VH[64]
  PIN SET_VH[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9385.595 187.44 9385.875 188.44 ;
    END
  END SET_VH[63]
  PIN SET_VH[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9245.595 187.44 9245.875 188.44 ;
    END
  END SET_VH[62]
  PIN SET_VH[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9105.595 187.44 9105.875 188.44 ;
    END
  END SET_VH[61]
  PIN SET_VH[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8965.595 187.44 8965.875 188.44 ;
    END
  END SET_VH[60]
  PIN SET_VH[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8825.595 187.44 8825.875 188.44 ;
    END
  END SET_VH[59]
  PIN SET_VH[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8685.595 187.44 8685.875 188.44 ;
    END
  END SET_VH[58]
  PIN SET_VH[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8545.595 187.44 8545.875 188.44 ;
    END
  END SET_VH[57]
  PIN SET_VH[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8405.595 187.44 8405.875 188.44 ;
    END
  END SET_VH[56]
  PIN SET_VH[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8265.595 187.44 8265.875 188.44 ;
    END
  END SET_VH[55]
  PIN SET_VH[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8125.595 187.44 8125.875 188.44 ;
    END
  END SET_VH[54]
  PIN SET_VH[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7985.595 187.44 7985.875 188.44 ;
    END
  END SET_VH[53]
  PIN SET_VH[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7845.595 187.44 7845.875 188.44 ;
    END
  END SET_VH[52]
  PIN SET_VH[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7705.595 187.44 7705.875 188.44 ;
    END
  END SET_VH[51]
  PIN SET_VH[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7565.595 187.44 7565.875 188.44 ;
    END
  END SET_VH[50]
  PIN SET_VH[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7425.595 187.44 7425.875 188.44 ;
    END
  END SET_VH[49]
  PIN SET_VH[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7285.595 187.44 7285.875 188.44 ;
    END
  END SET_VH[48]
  PIN SET_VH[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7145.595 187.44 7145.875 188.44 ;
    END
  END SET_VH[47]
  PIN SET_VH[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7005.595 187.44 7005.875 188.44 ;
    END
  END SET_VH[46]
  PIN SET_VH[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6865.595 187.44 6865.875 188.44 ;
    END
  END SET_VH[45]
  PIN SET_VH[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6725.595 187.44 6725.875 188.44 ;
    END
  END SET_VH[44]
  PIN SET_VH[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6585.595 187.44 6585.875 188.44 ;
    END
  END SET_VH[43]
  PIN SET_VH[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6445.595 187.44 6445.875 188.44 ;
    END
  END SET_VH[42]
  PIN SET_VH[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6305.595 187.44 6305.875 188.44 ;
    END
  END SET_VH[41]
  PIN SET_VH[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6165.595 187.44 6165.875 188.44 ;
    END
  END SET_VH[40]
  PIN SET_VH[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6025.595 187.44 6025.875 188.44 ;
    END
  END SET_VH[39]
  PIN SET_VH[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5885.595 187.44 5885.875 188.44 ;
    END
  END SET_VH[38]
  PIN SET_VH[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5745.595 187.44 5745.875 188.44 ;
    END
  END SET_VH[37]
  PIN SET_VH[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5605.595 187.44 5605.875 188.44 ;
    END
  END SET_VH[36]
  PIN SET_VH[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5465.595 187.44 5465.875 188.44 ;
    END
  END SET_VH[35]
  PIN SET_VH[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5325.595 187.44 5325.875 188.44 ;
    END
  END SET_VH[34]
  PIN SET_VH[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5185.595 187.44 5185.875 188.44 ;
    END
  END SET_VH[33]
  PIN SET_VH[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5045.595 187.44 5045.875 188.44 ;
    END
  END SET_VH[32]
  PIN SET_VH[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4905.595 187.44 4905.875 188.44 ;
    END
  END SET_VH[31]
  PIN SET_VH[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4765.595 187.44 4765.875 188.44 ;
    END
  END SET_VH[30]
  PIN SET_VH[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4625.595 187.44 4625.875 188.44 ;
    END
  END SET_VH[29]
  PIN SET_VH[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4485.595 187.44 4485.875 188.44 ;
    END
  END SET_VH[28]
  PIN SET_VH[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4345.595 187.44 4345.875 188.44 ;
    END
  END SET_VH[27]
  PIN SET_VH[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4205.595 187.44 4205.875 188.44 ;
    END
  END SET_VH[26]
  PIN SET_VH[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4065.595 187.44 4065.875 188.44 ;
    END
  END SET_VH[25]
  PIN SET_VH[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3925.595 187.44 3925.875 188.44 ;
    END
  END SET_VH[24]
  PIN SET_VH[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3785.595 187.44 3785.875 188.44 ;
    END
  END SET_VH[23]
  PIN SET_VH[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3645.595 187.44 3645.875 188.44 ;
    END
  END SET_VH[22]
  PIN SET_VH[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3505.595 187.44 3505.875 188.44 ;
    END
  END SET_VH[21]
  PIN SET_VH[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3365.595 187.44 3365.875 188.44 ;
    END
  END SET_VH[20]
  PIN SET_VH[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3225.595 187.44 3225.875 188.44 ;
    END
  END SET_VH[19]
  PIN SET_VH[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3085.595 187.44 3085.875 188.44 ;
    END
  END SET_VH[18]
  PIN SET_VH[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2945.595 187.44 2945.875 188.44 ;
    END
  END SET_VH[17]
  PIN SET_VH[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2805.595 187.44 2805.875 188.44 ;
    END
  END SET_VH[16]
  PIN SET_VH[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2665.595 187.44 2665.875 188.44 ;
    END
  END SET_VH[15]
  PIN SET_VH[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2525.595 187.44 2525.875 188.44 ;
    END
  END SET_VH[14]
  PIN SET_VH[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2385.595 187.44 2385.875 188.44 ;
    END
  END SET_VH[13]
  PIN SET_VH[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2245.595 187.44 2245.875 188.44 ;
    END
  END SET_VH[12]
  PIN SET_VH[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2105.595 187.44 2105.875 188.44 ;
    END
  END SET_VH[11]
  PIN SET_VH[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1965.595 187.44 1965.875 188.44 ;
    END
  END SET_VH[10]
  PIN SET_VH[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1825.595 187.44 1825.875 188.44 ;
    END
  END SET_VH[9]
  PIN SET_VH[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1685.595 187.44 1685.875 188.44 ;
    END
  END SET_VH[8]
  PIN SET_VH[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1545.595 187.44 1545.875 188.44 ;
    END
  END SET_VH[7]
  PIN SET_VH[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1405.595 187.44 1405.875 188.44 ;
    END
  END SET_VH[6]
  PIN SET_VH[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1265.595 187.44 1265.875 188.44 ;
    END
  END SET_VH[5]
  PIN SET_VH[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1125.595 187.44 1125.875 188.44 ;
    END
  END SET_VH[4]
  PIN SET_VH[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 985.595 187.44 985.875 188.44 ;
    END
  END SET_VH[3]
  PIN SET_VH[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 845.595 187.44 845.875 188.44 ;
    END
  END SET_VH[2]
  PIN SET_VH[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 705.595 187.44 705.875 188.44 ;
    END
  END SET_VH[1]
  PIN SET_VH[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 565.595 187.44 565.875 188.44 ;
    END
  END SET_VH[0]
  PIN SET_VL[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18341.955 187.44 18342.235 188.44 ;
    END
  END SET_VL[127]
  PIN SET_VL[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18201.955 187.44 18202.235 188.44 ;
    END
  END SET_VL[126]
  PIN SWCNTL_ICASN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9414.835 187.44 9415.395 188.44 ;
    END
  END SWCNTL_ICASN
  PIN SWCNTL_VRESET_D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9416.515 187.44 9417.075 188.44 ;
    END
  END SWCNTL_VRESET_D
  PIN SWCNTL_VL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9418.195 187.44 9418.755 188.44 ;
    END
  END SWCNTL_VL
  PIN SWCNTL_VH
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9419.875 187.44 9420.435 188.44 ;
    END
  END SWCNTL_VH
  PIN SWCNTL_VRESET_P
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9421.555 187.44 9422.115 188.44 ;
    END
  END SWCNTL_VRESET_P
  PIN SWCNTL_VCLIP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9423.235 187.44 9423.795 188.44 ;
    END
  END SWCNTL_VCLIP
  PIN DACMON_VH
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER M5 ;
        RECT 18489.46 264.79 18490.46 265.99 ;
    END
  END DACMON_VH
  PIN SWCNTL_VCASN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9424.915 187.44 9425.475 188.44 ;
    END
  END SWCNTL_VCASN
  PIN SWCNTL_DACMONI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9426.595 187.44 9427.155 188.44 ;
    END
  END SWCNTL_DACMONI
  PIN SWCNTL_DACMONV
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9428.275 187.44 9428.835 188.44 ;
    END
  END SWCNTL_DACMONV
  PIN SWCNTL_IREF
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9429.955 187.44 9430.515 188.44 ;
    END
  END SWCNTL_IREF
  PIN DACMON_IBIAS
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER M5 ;
        RECT 326.66 267.19 327.66 268.39 ;
    END
  END DACMON_IBIAS
  PIN DACMON_ITHR
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER M5 ;
        RECT 326.66 264.79 327.66 265.99 ;
    END
  END DACMON_ITHR
  PIN DACMON_IDB
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER M5 ;
        RECT 326.66 262.39 327.66 263.59 ;
    END
  END DACMON_IDB
  PIN DACMON_IRESET
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER M5 ;
        RECT 326.66 259.99 327.66 261.19 ;
    END
  END DACMON_IRESET
  PIN DACMON_ICASN
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER M5 ;
        RECT 326.66 257.59 327.66 258.79 ;
    END
  END DACMON_ICASN
  PIN DACMON_VRESET_P
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER M5 ;
        RECT 18489.46 262.39 18490.46 263.59 ;
    END
  END DACMON_VRESET_P
  PIN DACMON_VL
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER M5 ;
        RECT 18489.46 267.19 18490.46 268.39 ;
    END
  END DACMON_VL
  PIN SET_VL[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18061.955 187.44 18062.235 188.44 ;
    END
  END SET_VL[125]
  PIN SET_VL[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17921.955 187.44 17922.235 188.44 ;
    END
  END SET_VL[124]
  PIN SET_VL[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17781.955 187.44 17782.235 188.44 ;
    END
  END SET_VL[123]
  PIN SET_VL[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17641.955 187.44 17642.235 188.44 ;
    END
  END SET_VL[122]
  PIN SET_VL[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17501.955 187.44 17502.235 188.44 ;
    END
  END SET_VL[121]
  PIN SET_VL[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17361.955 187.44 17362.235 188.44 ;
    END
  END SET_VL[120]
  PIN SET_VL[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17221.955 187.44 17222.235 188.44 ;
    END
  END SET_VL[119]
  PIN SET_VL[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17081.955 187.44 17082.235 188.44 ;
    END
  END SET_VL[118]
  PIN SET_VL[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16941.955 187.44 16942.235 188.44 ;
    END
  END SET_VL[117]
  PIN SET_VL[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16801.955 187.44 16802.235 188.44 ;
    END
  END SET_VL[116]
  PIN SET_VL[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16661.955 187.44 16662.235 188.44 ;
    END
  END SET_VL[115]
  PIN SET_VL[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16521.955 187.44 16522.235 188.44 ;
    END
  END SET_VL[114]
  PIN SET_VL[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16381.955 187.44 16382.235 188.44 ;
    END
  END SET_VL[113]
  PIN SET_VL[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16241.955 187.44 16242.235 188.44 ;
    END
  END SET_VL[112]
  PIN SET_VL[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16101.955 187.44 16102.235 188.44 ;
    END
  END SET_VL[111]
  PIN SET_VL[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15961.955 187.44 15962.235 188.44 ;
    END
  END SET_VL[110]
  PIN SET_VL[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15821.955 187.44 15822.235 188.44 ;
    END
  END SET_VL[109]
  PIN SET_VL[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15681.955 187.44 15682.235 188.44 ;
    END
  END SET_VL[108]
  PIN SET_VL[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15541.955 187.44 15542.235 188.44 ;
    END
  END SET_VL[107]
  PIN SET_VL[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15401.955 187.44 15402.235 188.44 ;
    END
  END SET_VL[106]
  PIN SET_VL[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15261.955 187.44 15262.235 188.44 ;
    END
  END SET_VL[105]
  PIN SET_VL[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15121.955 187.44 15122.235 188.44 ;
    END
  END SET_VL[104]
  PIN SET_VL[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14981.955 187.44 14982.235 188.44 ;
    END
  END SET_VL[103]
  PIN SET_VL[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14841.955 187.44 14842.235 188.44 ;
    END
  END SET_VL[102]
  PIN SET_VL[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14701.955 187.44 14702.235 188.44 ;
    END
  END SET_VL[101]
  PIN SET_VL[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14561.955 187.44 14562.235 188.44 ;
    END
  END SET_VL[100]
  PIN SET_VL[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14421.955 187.44 14422.235 188.44 ;
    END
  END SET_VL[99]
  PIN SET_VL[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14281.955 187.44 14282.235 188.44 ;
    END
  END SET_VL[98]
  PIN SET_VL[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14141.955 187.44 14142.235 188.44 ;
    END
  END SET_VL[97]
  PIN SET_VL[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14001.955 187.44 14002.235 188.44 ;
    END
  END SET_VL[96]
  PIN SET_VL[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13861.955 187.44 13862.235 188.44 ;
    END
  END SET_VL[95]
  PIN SET_VL[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13721.955 187.44 13722.235 188.44 ;
    END
  END SET_VL[94]
  PIN SET_VL[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13581.955 187.44 13582.235 188.44 ;
    END
  END SET_VL[93]
  PIN SET_VL[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13441.955 187.44 13442.235 188.44 ;
    END
  END SET_VL[92]
  PIN SET_VL[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13301.955 187.44 13302.235 188.44 ;
    END
  END SET_VL[91]
  PIN SET_VL[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13161.955 187.44 13162.235 188.44 ;
    END
  END SET_VL[90]
  PIN SET_VL[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13021.955 187.44 13022.235 188.44 ;
    END
  END SET_VL[89]
  PIN SET_VL[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12881.955 187.44 12882.235 188.44 ;
    END
  END SET_VL[88]
  PIN SET_VL[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12741.955 187.44 12742.235 188.44 ;
    END
  END SET_VL[87]
  PIN SET_VL[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12601.955 187.44 12602.235 188.44 ;
    END
  END SET_VL[86]
  PIN SET_VL[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12461.955 187.44 12462.235 188.44 ;
    END
  END SET_VL[85]
  PIN SET_VL[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12321.955 187.44 12322.235 188.44 ;
    END
  END SET_VL[84]
  PIN SET_VL[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12181.955 187.44 12182.235 188.44 ;
    END
  END SET_VL[83]
  PIN SET_VL[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12041.955 187.44 12042.235 188.44 ;
    END
  END SET_VL[82]
  PIN SET_VL[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11901.955 187.44 11902.235 188.44 ;
    END
  END SET_VL[81]
  PIN SET_VL[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11761.955 187.44 11762.235 188.44 ;
    END
  END SET_VL[80]
  PIN SET_VL[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11621.955 187.44 11622.235 188.44 ;
    END
  END SET_VL[79]
  PIN SET_VL[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11481.955 187.44 11482.235 188.44 ;
    END
  END SET_VL[78]
  PIN SET_VL[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11341.955 187.44 11342.235 188.44 ;
    END
  END SET_VL[77]
  PIN SET_VL[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11201.955 187.44 11202.235 188.44 ;
    END
  END SET_VL[76]
  PIN SET_VL[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11061.955 187.44 11062.235 188.44 ;
    END
  END SET_VL[75]
  PIN SET_VL[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10921.955 187.44 10922.235 188.44 ;
    END
  END SET_VL[74]
  PIN SET_VL[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10781.955 187.44 10782.235 188.44 ;
    END
  END SET_VL[73]
  PIN SET_VL[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10641.955 187.44 10642.235 188.44 ;
    END
  END SET_VL[72]
  PIN SET_VL[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10501.955 187.44 10502.235 188.44 ;
    END
  END SET_VL[71]
  PIN SET_VL[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10361.955 187.44 10362.235 188.44 ;
    END
  END SET_VL[70]
  PIN SET_VL[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10221.955 187.44 10222.235 188.44 ;
    END
  END SET_VL[69]
  PIN SET_VL[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10081.955 187.44 10082.235 188.44 ;
    END
  END SET_VL[68]
  PIN SET_VL[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9941.955 187.44 9942.235 188.44 ;
    END
  END SET_VL[67]
  PIN SET_VL[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9801.955 187.44 9802.235 188.44 ;
    END
  END SET_VL[66]
  PIN SET_VL[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9661.955 187.44 9662.235 188.44 ;
    END
  END SET_VL[65]
  PIN SET_VL[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9521.955 187.44 9522.235 188.44 ;
    END
  END SET_VL[64]
  PIN SET_VL[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9381.955 187.44 9382.235 188.44 ;
    END
  END SET_VL[63]
  PIN SET_VL[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9241.955 187.44 9242.235 188.44 ;
    END
  END SET_VL[62]
  PIN SET_VL[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9101.955 187.44 9102.235 188.44 ;
    END
  END SET_VL[61]
  PIN SET_VL[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8961.955 187.44 8962.235 188.44 ;
    END
  END SET_VL[60]
  PIN SET_VL[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8821.955 187.44 8822.235 188.44 ;
    END
  END SET_VL[59]
  PIN SET_VL[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8681.955 187.44 8682.235 188.44 ;
    END
  END SET_VL[58]
  PIN SET_VL[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8541.955 187.44 8542.235 188.44 ;
    END
  END SET_VL[57]
  PIN SET_VL[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8401.955 187.44 8402.235 188.44 ;
    END
  END SET_VL[56]
  PIN SET_VL[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8261.955 187.44 8262.235 188.44 ;
    END
  END SET_VL[55]
  PIN SET_VL[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8121.955 187.44 8122.235 188.44 ;
    END
  END SET_VL[54]
  PIN SET_VL[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7981.955 187.44 7982.235 188.44 ;
    END
  END SET_VL[53]
  PIN SET_VL[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7841.955 187.44 7842.235 188.44 ;
    END
  END SET_VL[52]
  PIN SET_VL[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7701.955 187.44 7702.235 188.44 ;
    END
  END SET_VL[51]
  PIN SET_VL[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7561.955 187.44 7562.235 188.44 ;
    END
  END SET_VL[50]
  PIN SET_VL[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7421.955 187.44 7422.235 188.44 ;
    END
  END SET_VL[49]
  PIN SET_VL[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7281.955 187.44 7282.235 188.44 ;
    END
  END SET_VL[48]
  PIN SET_VL[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7141.955 187.44 7142.235 188.44 ;
    END
  END SET_VL[47]
  PIN SET_VL[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7001.955 187.44 7002.235 188.44 ;
    END
  END SET_VL[46]
  PIN SET_VL[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6861.955 187.44 6862.235 188.44 ;
    END
  END SET_VL[45]
  PIN SET_VL[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6721.955 187.44 6722.235 188.44 ;
    END
  END SET_VL[44]
  PIN SET_VL[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6581.955 187.44 6582.235 188.44 ;
    END
  END SET_VL[43]
  PIN SET_VL[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6441.955 187.44 6442.235 188.44 ;
    END
  END SET_VL[42]
  PIN SET_VL[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6301.955 187.44 6302.235 188.44 ;
    END
  END SET_VL[41]
  PIN SET_VL[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6161.955 187.44 6162.235 188.44 ;
    END
  END SET_VL[40]
  PIN SET_VL[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6021.955 187.44 6022.235 188.44 ;
    END
  END SET_VL[39]
  PIN SET_VL[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5881.955 187.44 5882.235 188.44 ;
    END
  END SET_VL[38]
  PIN SET_VL[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5741.955 187.44 5742.235 188.44 ;
    END
  END SET_VL[37]
  PIN SET_VL[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5601.955 187.44 5602.235 188.44 ;
    END
  END SET_VL[36]
  PIN SET_VL[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5461.955 187.44 5462.235 188.44 ;
    END
  END SET_VL[35]
  PIN SET_VL[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5321.955 187.44 5322.235 188.44 ;
    END
  END SET_VL[34]
  PIN SET_VL[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5181.955 187.44 5182.235 188.44 ;
    END
  END SET_VL[33]
  PIN SET_VL[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5041.955 187.44 5042.235 188.44 ;
    END
  END SET_VL[32]
  PIN SET_VL[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4901.955 187.44 4902.235 188.44 ;
    END
  END SET_VL[31]
  PIN SET_VL[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4761.955 187.44 4762.235 188.44 ;
    END
  END SET_VL[30]
  PIN SET_VL[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4621.955 187.44 4622.235 188.44 ;
    END
  END SET_VL[29]
  PIN SET_VL[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4481.955 187.44 4482.235 188.44 ;
    END
  END SET_VL[28]
  PIN SET_VL[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4341.955 187.44 4342.235 188.44 ;
    END
  END SET_VL[27]
  PIN SET_VL[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4201.955 187.44 4202.235 188.44 ;
    END
  END SET_VL[26]
  PIN SET_VL[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4061.955 187.44 4062.235 188.44 ;
    END
  END SET_VL[25]
  PIN SET_VL[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3921.955 187.44 3922.235 188.44 ;
    END
  END SET_VL[24]
  PIN SET_VL[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3781.955 187.44 3782.235 188.44 ;
    END
  END SET_VL[23]
  PIN SET_VL[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3641.955 187.44 3642.235 188.44 ;
    END
  END SET_VL[22]
  PIN SET_VL[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3501.955 187.44 3502.235 188.44 ;
    END
  END SET_VL[21]
  PIN SET_VL[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3361.955 187.44 3362.235 188.44 ;
    END
  END SET_VL[20]
  PIN SET_VL[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3221.955 187.44 3222.235 188.44 ;
    END
  END SET_VL[19]
  PIN SET_VL[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3081.955 187.44 3082.235 188.44 ;
    END
  END SET_VL[18]
  PIN SET_VL[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2941.955 187.44 2942.235 188.44 ;
    END
  END SET_VL[17]
  PIN SET_VL[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2801.955 187.44 2802.235 188.44 ;
    END
  END SET_VL[16]
  PIN SET_VL[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2661.955 187.44 2662.235 188.44 ;
    END
  END SET_VL[15]
  PIN SET_VL[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2521.955 187.44 2522.235 188.44 ;
    END
  END SET_VL[14]
  PIN SET_VL[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2381.955 187.44 2382.235 188.44 ;
    END
  END SET_VL[13]
  PIN SET_VL[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2241.955 187.44 2242.235 188.44 ;
    END
  END SET_VL[12]
  PIN SET_VL[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2101.955 187.44 2102.235 188.44 ;
    END
  END SET_VL[11]
  PIN SET_VL[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1961.955 187.44 1962.235 188.44 ;
    END
  END SET_VL[10]
  PIN SET_VL[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1821.955 187.44 1822.235 188.44 ;
    END
  END SET_VL[9]
  PIN SET_VL[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1681.955 187.44 1682.235 188.44 ;
    END
  END SET_VL[8]
  PIN SET_VL[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1541.955 187.44 1542.235 188.44 ;
    END
  END SET_VL[7]
  PIN SET_VL[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1401.955 187.44 1402.235 188.44 ;
    END
  END SET_VL[6]
  PIN SET_VL[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1261.955 187.44 1262.235 188.44 ;
    END
  END SET_VL[5]
  PIN SET_VL[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1121.955 187.44 1122.235 188.44 ;
    END
  END SET_VL[4]
  PIN SET_VL[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 981.955 187.44 982.235 188.44 ;
    END
  END SET_VL[3]
  PIN SET_VL[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 841.955 187.44 842.235 188.44 ;
    END
  END SET_VL[2]
  PIN SET_VL[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 701.955 187.44 702.235 188.44 ;
    END
  END SET_VL[1]
  PIN SET_VL[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 561.955 187.44 562.235 188.44 ;
    END
  END SET_VL[0]
  PIN SET_VRESET_D[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18338.315 187.44 18338.595 188.44 ;
    END
  END SET_VRESET_D[127]
  PIN SET_VRESET_D[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18198.315 187.44 18198.595 188.44 ;
    END
  END SET_VRESET_D[126]
  PIN VCASN_MON_L
    DIRECTION OUTPUT ;
    USE ANALOG ;
    PORT
      LAYER M4 ;
        RECT 326.66 8438.095 327.66 8439.515 ;
    END
  END VCASN_MON_L
  PIN SWCNTL_IRESET
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9413.155 187.44 9413.715 188.44 ;
    END
  END SWCNTL_IRESET
  PIN SET_VRESET_D[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18058.315 187.44 18058.595 188.44 ;
    END
  END SET_VRESET_D[125]
  PIN SET_VRESET_D[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17918.315 187.44 17918.595 188.44 ;
    END
  END SET_VRESET_D[124]
  PIN SET_VRESET_D[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17778.315 187.44 17778.595 188.44 ;
    END
  END SET_VRESET_D[123]
  PIN SET_VRESET_D[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17638.315 187.44 17638.595 188.44 ;
    END
  END SET_VRESET_D[122]
  PIN SET_VRESET_D[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17498.315 187.44 17498.595 188.44 ;
    END
  END SET_VRESET_D[121]
  PIN SET_VRESET_D[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17358.315 187.44 17358.595 188.44 ;
    END
  END SET_VRESET_D[120]
  PIN SET_VRESET_D[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17218.315 187.44 17218.595 188.44 ;
    END
  END SET_VRESET_D[119]
  PIN SET_VRESET_D[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17078.315 187.44 17078.595 188.44 ;
    END
  END SET_VRESET_D[118]
  PIN SET_VRESET_D[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16938.315 187.44 16938.595 188.44 ;
    END
  END SET_VRESET_D[117]
  PIN SET_VRESET_D[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16798.315 187.44 16798.595 188.44 ;
    END
  END SET_VRESET_D[116]
  PIN SET_VRESET_D[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16658.315 187.44 16658.595 188.44 ;
    END
  END SET_VRESET_D[115]
  PIN SET_VRESET_D[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16518.315 187.44 16518.595 188.44 ;
    END
  END SET_VRESET_D[114]
  PIN SET_VRESET_D[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16378.315 187.44 16378.595 188.44 ;
    END
  END SET_VRESET_D[113]
  PIN SET_VRESET_D[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16238.315 187.44 16238.595 188.44 ;
    END
  END SET_VRESET_D[112]
  PIN SET_VRESET_D[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16098.315 187.44 16098.595 188.44 ;
    END
  END SET_VRESET_D[111]
  PIN SET_VRESET_D[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15958.315 187.44 15958.595 188.44 ;
    END
  END SET_VRESET_D[110]
  PIN SET_VRESET_D[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15818.315 187.44 15818.595 188.44 ;
    END
  END SET_VRESET_D[109]
  PIN SET_VRESET_D[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15678.315 187.44 15678.595 188.44 ;
    END
  END SET_VRESET_D[108]
  PIN SET_VRESET_D[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15538.315 187.44 15538.595 188.44 ;
    END
  END SET_VRESET_D[107]
  PIN SET_VRESET_D[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15398.315 187.44 15398.595 188.44 ;
    END
  END SET_VRESET_D[106]
  PIN SET_VRESET_D[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15258.315 187.44 15258.595 188.44 ;
    END
  END SET_VRESET_D[105]
  PIN SET_VRESET_D[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15118.315 187.44 15118.595 188.44 ;
    END
  END SET_VRESET_D[104]
  PIN SET_VRESET_D[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14978.315 187.44 14978.595 188.44 ;
    END
  END SET_VRESET_D[103]
  PIN SET_VRESET_D[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14838.315 187.44 14838.595 188.44 ;
    END
  END SET_VRESET_D[102]
  PIN SET_VRESET_D[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14698.315 187.44 14698.595 188.44 ;
    END
  END SET_VRESET_D[101]
  PIN SET_VRESET_D[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14558.315 187.44 14558.595 188.44 ;
    END
  END SET_VRESET_D[100]
  PIN SET_VRESET_D[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14418.315 187.44 14418.595 188.44 ;
    END
  END SET_VRESET_D[99]
  PIN SET_VRESET_D[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14278.315 187.44 14278.595 188.44 ;
    END
  END SET_VRESET_D[98]
  PIN SET_VRESET_D[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14138.315 187.44 14138.595 188.44 ;
    END
  END SET_VRESET_D[97]
  PIN SET_VRESET_D[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13998.315 187.44 13998.595 188.44 ;
    END
  END SET_VRESET_D[96]
  PIN SET_VRESET_D[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13858.315 187.44 13858.595 188.44 ;
    END
  END SET_VRESET_D[95]
  PIN SET_VRESET_D[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13718.315 187.44 13718.595 188.44 ;
    END
  END SET_VRESET_D[94]
  PIN SET_VRESET_D[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13578.315 187.44 13578.595 188.44 ;
    END
  END SET_VRESET_D[93]
  PIN SET_VRESET_D[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13438.315 187.44 13438.595 188.44 ;
    END
  END SET_VRESET_D[92]
  PIN SET_VRESET_D[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13298.315 187.44 13298.595 188.44 ;
    END
  END SET_VRESET_D[91]
  PIN SET_VRESET_D[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13158.315 187.44 13158.595 188.44 ;
    END
  END SET_VRESET_D[90]
  PIN SET_VRESET_D[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13018.315 187.44 13018.595 188.44 ;
    END
  END SET_VRESET_D[89]
  PIN SET_VRESET_D[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12878.315 187.44 12878.595 188.44 ;
    END
  END SET_VRESET_D[88]
  PIN SET_VRESET_D[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12738.315 187.44 12738.595 188.44 ;
    END
  END SET_VRESET_D[87]
  PIN SET_VRESET_D[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12598.315 187.44 12598.595 188.44 ;
    END
  END SET_VRESET_D[86]
  PIN SET_VRESET_D[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12458.315 187.44 12458.595 188.44 ;
    END
  END SET_VRESET_D[85]
  PIN SET_VRESET_D[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12318.315 187.44 12318.595 188.44 ;
    END
  END SET_VRESET_D[84]
  PIN SET_VRESET_D[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12178.315 187.44 12178.595 188.44 ;
    END
  END SET_VRESET_D[83]
  PIN SET_VRESET_D[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12038.315 187.44 12038.595 188.44 ;
    END
  END SET_VRESET_D[82]
  PIN SET_VRESET_D[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11898.315 187.44 11898.595 188.44 ;
    END
  END SET_VRESET_D[81]
  PIN SET_VRESET_D[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11758.315 187.44 11758.595 188.44 ;
    END
  END SET_VRESET_D[80]
  PIN SET_VRESET_D[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11618.315 187.44 11618.595 188.44 ;
    END
  END SET_VRESET_D[79]
  PIN SET_VRESET_D[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11478.315 187.44 11478.595 188.44 ;
    END
  END SET_VRESET_D[78]
  PIN SET_VRESET_D[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11338.315 187.44 11338.595 188.44 ;
    END
  END SET_VRESET_D[77]
  PIN SET_VRESET_D[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11198.315 187.44 11198.595 188.44 ;
    END
  END SET_VRESET_D[76]
  PIN SET_VRESET_D[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11058.315 187.44 11058.595 188.44 ;
    END
  END SET_VRESET_D[75]
  PIN SET_VRESET_D[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10918.315 187.44 10918.595 188.44 ;
    END
  END SET_VRESET_D[74]
  PIN SET_VRESET_D[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10778.315 187.44 10778.595 188.44 ;
    END
  END SET_VRESET_D[73]
  PIN SET_VRESET_D[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10638.315 187.44 10638.595 188.44 ;
    END
  END SET_VRESET_D[72]
  PIN SET_VRESET_D[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10498.315 187.44 10498.595 188.44 ;
    END
  END SET_VRESET_D[71]
  PIN SET_VRESET_D[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10358.315 187.44 10358.595 188.44 ;
    END
  END SET_VRESET_D[70]
  PIN SET_VRESET_D[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10218.315 187.44 10218.595 188.44 ;
    END
  END SET_VRESET_D[69]
  PIN SET_VRESET_D[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10078.315 187.44 10078.595 188.44 ;
    END
  END SET_VRESET_D[68]
  PIN SET_VRESET_D[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9938.315 187.44 9938.595 188.44 ;
    END
  END SET_VRESET_D[67]
  PIN SET_VRESET_D[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9798.315 187.44 9798.595 188.44 ;
    END
  END SET_VRESET_D[66]
  PIN SET_VRESET_D[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9658.315 187.44 9658.595 188.44 ;
    END
  END SET_VRESET_D[65]
  PIN SET_VRESET_D[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9518.315 187.44 9518.595 188.44 ;
    END
  END SET_VRESET_D[64]
  PIN SET_VRESET_D[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9378.315 187.44 9378.595 188.44 ;
    END
  END SET_VRESET_D[63]
  PIN SET_VRESET_D[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9238.315 187.44 9238.595 188.44 ;
    END
  END SET_VRESET_D[62]
  PIN SET_VRESET_D[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9098.315 187.44 9098.595 188.44 ;
    END
  END SET_VRESET_D[61]
  PIN SET_VRESET_D[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8958.315 187.44 8958.595 188.44 ;
    END
  END SET_VRESET_D[60]
  PIN SET_VRESET_D[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8818.315 187.44 8818.595 188.44 ;
    END
  END SET_VRESET_D[59]
  PIN SET_VRESET_D[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8678.315 187.44 8678.595 188.44 ;
    END
  END SET_VRESET_D[58]
  PIN SET_VRESET_D[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8538.315 187.44 8538.595 188.44 ;
    END
  END SET_VRESET_D[57]
  PIN SET_VRESET_D[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8398.315 187.44 8398.595 188.44 ;
    END
  END SET_VRESET_D[56]
  PIN SET_VRESET_D[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8258.315 187.44 8258.595 188.44 ;
    END
  END SET_VRESET_D[55]
  PIN SET_VRESET_D[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8118.315 187.44 8118.595 188.44 ;
    END
  END SET_VRESET_D[54]
  PIN SET_VRESET_D[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7978.315 187.44 7978.595 188.44 ;
    END
  END SET_VRESET_D[53]
  PIN SET_VRESET_D[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7838.315 187.44 7838.595 188.44 ;
    END
  END SET_VRESET_D[52]
  PIN SET_VRESET_D[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7698.315 187.44 7698.595 188.44 ;
    END
  END SET_VRESET_D[51]
  PIN SET_VRESET_D[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7558.315 187.44 7558.595 188.44 ;
    END
  END SET_VRESET_D[50]
  PIN SET_VRESET_D[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7418.315 187.44 7418.595 188.44 ;
    END
  END SET_VRESET_D[49]
  PIN SET_VRESET_D[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7278.315 187.44 7278.595 188.44 ;
    END
  END SET_VRESET_D[48]
  PIN SET_VRESET_D[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7138.315 187.44 7138.595 188.44 ;
    END
  END SET_VRESET_D[47]
  PIN SET_VRESET_D[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6998.315 187.44 6998.595 188.44 ;
    END
  END SET_VRESET_D[46]
  PIN SET_VRESET_D[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6858.315 187.44 6858.595 188.44 ;
    END
  END SET_VRESET_D[45]
  PIN SET_VRESET_D[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6718.315 187.44 6718.595 188.44 ;
    END
  END SET_VRESET_D[44]
  PIN SET_VRESET_D[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6578.315 187.44 6578.595 188.44 ;
    END
  END SET_VRESET_D[43]
  PIN SET_VRESET_D[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6438.315 187.44 6438.595 188.44 ;
    END
  END SET_VRESET_D[42]
  PIN SET_VRESET_D[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6298.315 187.44 6298.595 188.44 ;
    END
  END SET_VRESET_D[41]
  PIN SET_VRESET_D[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6158.315 187.44 6158.595 188.44 ;
    END
  END SET_VRESET_D[40]
  PIN SET_VRESET_D[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6018.315 187.44 6018.595 188.44 ;
    END
  END SET_VRESET_D[39]
  PIN SET_VRESET_D[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5878.315 187.44 5878.595 188.44 ;
    END
  END SET_VRESET_D[38]
  PIN SET_VRESET_D[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5738.315 187.44 5738.595 188.44 ;
    END
  END SET_VRESET_D[37]
  PIN SET_VRESET_D[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5598.315 187.44 5598.595 188.44 ;
    END
  END SET_VRESET_D[36]
  PIN SET_VRESET_D[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5458.315 187.44 5458.595 188.44 ;
    END
  END SET_VRESET_D[35]
  PIN SET_VRESET_D[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5318.315 187.44 5318.595 188.44 ;
    END
  END SET_VRESET_D[34]
  PIN SET_VRESET_D[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5178.315 187.44 5178.595 188.44 ;
    END
  END SET_VRESET_D[33]
  PIN SET_VRESET_D[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5038.315 187.44 5038.595 188.44 ;
    END
  END SET_VRESET_D[32]
  PIN SET_VRESET_D[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4898.315 187.44 4898.595 188.44 ;
    END
  END SET_VRESET_D[31]
  PIN SET_VRESET_D[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4758.315 187.44 4758.595 188.44 ;
    END
  END SET_VRESET_D[30]
  PIN SET_VRESET_D[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4618.315 187.44 4618.595 188.44 ;
    END
  END SET_VRESET_D[29]
  PIN SET_VRESET_D[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4478.315 187.44 4478.595 188.44 ;
    END
  END SET_VRESET_D[28]
  PIN SET_VRESET_D[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4338.315 187.44 4338.595 188.44 ;
    END
  END SET_VRESET_D[27]
  PIN SET_VRESET_D[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4198.315 187.44 4198.595 188.44 ;
    END
  END SET_VRESET_D[26]
  PIN SET_VRESET_D[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4058.315 187.44 4058.595 188.44 ;
    END
  END SET_VRESET_D[25]
  PIN SET_VRESET_D[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3918.315 187.44 3918.595 188.44 ;
    END
  END SET_VRESET_D[24]
  PIN SET_VRESET_D[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3778.315 187.44 3778.595 188.44 ;
    END
  END SET_VRESET_D[23]
  PIN SET_VRESET_D[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3638.315 187.44 3638.595 188.44 ;
    END
  END SET_VRESET_D[22]
  PIN SET_VRESET_D[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3498.315 187.44 3498.595 188.44 ;
    END
  END SET_VRESET_D[21]
  PIN SET_VRESET_D[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3358.315 187.44 3358.595 188.44 ;
    END
  END SET_VRESET_D[20]
  PIN SET_VRESET_D[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3218.315 187.44 3218.595 188.44 ;
    END
  END SET_VRESET_D[19]
  PIN SET_VRESET_D[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3078.315 187.44 3078.595 188.44 ;
    END
  END SET_VRESET_D[18]
  PIN SET_VRESET_D[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2938.315 187.44 2938.595 188.44 ;
    END
  END SET_VRESET_D[17]
  PIN SET_VRESET_D[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2798.315 187.44 2798.595 188.44 ;
    END
  END SET_VRESET_D[16]
  PIN SET_VRESET_D[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2658.315 187.44 2658.595 188.44 ;
    END
  END SET_VRESET_D[15]
  PIN SET_VRESET_D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2518.315 187.44 2518.595 188.44 ;
    END
  END SET_VRESET_D[14]
  PIN SET_VRESET_D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2378.315 187.44 2378.595 188.44 ;
    END
  END SET_VRESET_D[13]
  PIN SET_VRESET_D[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2238.315 187.44 2238.595 188.44 ;
    END
  END SET_VRESET_D[12]
  PIN SET_VRESET_D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2098.315 187.44 2098.595 188.44 ;
    END
  END SET_VRESET_D[11]
  PIN SET_VRESET_D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1958.315 187.44 1958.595 188.44 ;
    END
  END SET_VRESET_D[10]
  PIN SET_VRESET_D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1818.315 187.44 1818.595 188.44 ;
    END
  END SET_VRESET_D[9]
  PIN SET_VRESET_D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1678.315 187.44 1678.595 188.44 ;
    END
  END SET_VRESET_D[8]
  PIN SET_VRESET_D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1538.315 187.44 1538.595 188.44 ;
    END
  END SET_VRESET_D[7]
  PIN SET_VRESET_D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1398.315 187.44 1398.595 188.44 ;
    END
  END SET_VRESET_D[6]
  PIN SET_VRESET_D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1258.315 187.44 1258.595 188.44 ;
    END
  END SET_VRESET_D[5]
  PIN SET_VRESET_D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1118.315 187.44 1118.595 188.44 ;
    END
  END SET_VRESET_D[4]
  PIN SET_VRESET_D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 978.315 187.44 978.595 188.44 ;
    END
  END SET_VRESET_D[3]
  PIN SET_VRESET_D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 838.315 187.44 838.595 188.44 ;
    END
  END SET_VRESET_D[2]
  PIN SET_VRESET_D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 698.315 187.44 698.595 188.44 ;
    END
  END SET_VRESET_D[1]
  PIN SET_VRESET_D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 558.315 187.44 558.595 188.44 ;
    END
  END SET_VRESET_D[0]
  PIN SET_ICASN[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18279.235 187.44 18279.515 188.44 ;
    END
  END SET_ICASN[127]
  PIN SET_ICASN[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18139.235 187.44 18139.515 188.44 ;
    END
  END SET_ICASN[126]
  PIN SWCNTL_ITHR
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9409.795 187.44 9410.355 188.44 ;
    END
  END SWCNTL_ITHR
  PIN SET_ICASN[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17999.235 187.44 17999.515 188.44 ;
    END
  END SET_ICASN[125]
  PIN SET_ICASN[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17859.235 187.44 17859.515 188.44 ;
    END
  END SET_ICASN[124]
  PIN SET_ICASN[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17719.235 187.44 17719.515 188.44 ;
    END
  END SET_ICASN[123]
  PIN SET_ICASN[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17579.235 187.44 17579.515 188.44 ;
    END
  END SET_ICASN[122]
  PIN SET_ICASN[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17439.235 187.44 17439.515 188.44 ;
    END
  END SET_ICASN[121]
  PIN SET_ICASN[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17299.235 187.44 17299.515 188.44 ;
    END
  END SET_ICASN[120]
  PIN SET_ICASN[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17159.235 187.44 17159.515 188.44 ;
    END
  END SET_ICASN[119]
  PIN SET_ICASN[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17019.235 187.44 17019.515 188.44 ;
    END
  END SET_ICASN[118]
  PIN SET_ICASN[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16879.235 187.44 16879.515 188.44 ;
    END
  END SET_ICASN[117]
  PIN SET_ICASN[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16739.235 187.44 16739.515 188.44 ;
    END
  END SET_ICASN[116]
  PIN SET_ICASN[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16599.235 187.44 16599.515 188.44 ;
    END
  END SET_ICASN[115]
  PIN SET_ICASN[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16459.235 187.44 16459.515 188.44 ;
    END
  END SET_ICASN[114]
  PIN SET_ICASN[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16319.235 187.44 16319.515 188.44 ;
    END
  END SET_ICASN[113]
  PIN SET_ICASN[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16179.235 187.44 16179.515 188.44 ;
    END
  END SET_ICASN[112]
  PIN SET_ICASN[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16039.235 187.44 16039.515 188.44 ;
    END
  END SET_ICASN[111]
  PIN SET_ICASN[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15899.235 187.44 15899.515 188.44 ;
    END
  END SET_ICASN[110]
  PIN SET_ICASN[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15759.235 187.44 15759.515 188.44 ;
    END
  END SET_ICASN[109]
  PIN SET_ICASN[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15619.235 187.44 15619.515 188.44 ;
    END
  END SET_ICASN[108]
  PIN SET_ICASN[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15479.235 187.44 15479.515 188.44 ;
    END
  END SET_ICASN[107]
  PIN SET_ICASN[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15339.235 187.44 15339.515 188.44 ;
    END
  END SET_ICASN[106]
  PIN SET_ICASN[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15199.235 187.44 15199.515 188.44 ;
    END
  END SET_ICASN[105]
  PIN SET_ICASN[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15059.235 187.44 15059.515 188.44 ;
    END
  END SET_ICASN[104]
  PIN SET_ICASN[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14919.235 187.44 14919.515 188.44 ;
    END
  END SET_ICASN[103]
  PIN SET_ICASN[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14779.235 187.44 14779.515 188.44 ;
    END
  END SET_ICASN[102]
  PIN SET_ICASN[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14639.235 187.44 14639.515 188.44 ;
    END
  END SET_ICASN[101]
  PIN SET_ICASN[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14499.235 187.44 14499.515 188.44 ;
    END
  END SET_ICASN[100]
  PIN SET_ICASN[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14359.235 187.44 14359.515 188.44 ;
    END
  END SET_ICASN[99]
  PIN SET_ICASN[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14219.235 187.44 14219.515 188.44 ;
    END
  END SET_ICASN[98]
  PIN SET_ICASN[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14079.235 187.44 14079.515 188.44 ;
    END
  END SET_ICASN[97]
  PIN SET_ICASN[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13939.235 187.44 13939.515 188.44 ;
    END
  END SET_ICASN[96]
  PIN SET_ICASN[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13799.235 187.44 13799.515 188.44 ;
    END
  END SET_ICASN[95]
  PIN SET_ICASN[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13659.235 187.44 13659.515 188.44 ;
    END
  END SET_ICASN[94]
  PIN SET_ICASN[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13519.235 187.44 13519.515 188.44 ;
    END
  END SET_ICASN[93]
  PIN SET_ICASN[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13379.235 187.44 13379.515 188.44 ;
    END
  END SET_ICASN[92]
  PIN SET_ICASN[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13239.235 187.44 13239.515 188.44 ;
    END
  END SET_ICASN[91]
  PIN SET_ICASN[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13099.235 187.44 13099.515 188.44 ;
    END
  END SET_ICASN[90]
  PIN SET_ICASN[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12959.235 187.44 12959.515 188.44 ;
    END
  END SET_ICASN[89]
  PIN SET_ICASN[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12819.235 187.44 12819.515 188.44 ;
    END
  END SET_ICASN[88]
  PIN SET_ICASN[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12679.235 187.44 12679.515 188.44 ;
    END
  END SET_ICASN[87]
  PIN SET_ICASN[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12539.235 187.44 12539.515 188.44 ;
    END
  END SET_ICASN[86]
  PIN SET_ICASN[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12399.235 187.44 12399.515 188.44 ;
    END
  END SET_ICASN[85]
  PIN SET_ICASN[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12259.235 187.44 12259.515 188.44 ;
    END
  END SET_ICASN[84]
  PIN SET_ICASN[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12119.235 187.44 12119.515 188.44 ;
    END
  END SET_ICASN[83]
  PIN SET_ICASN[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11979.235 187.44 11979.515 188.44 ;
    END
  END SET_ICASN[82]
  PIN SET_ICASN[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11839.235 187.44 11839.515 188.44 ;
    END
  END SET_ICASN[81]
  PIN SET_ICASN[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11699.235 187.44 11699.515 188.44 ;
    END
  END SET_ICASN[80]
  PIN SET_ICASN[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11559.235 187.44 11559.515 188.44 ;
    END
  END SET_ICASN[79]
  PIN SET_ICASN[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11419.235 187.44 11419.515 188.44 ;
    END
  END SET_ICASN[78]
  PIN SET_ICASN[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11279.235 187.44 11279.515 188.44 ;
    END
  END SET_ICASN[77]
  PIN SET_ICASN[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11139.235 187.44 11139.515 188.44 ;
    END
  END SET_ICASN[76]
  PIN SET_ICASN[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10999.235 187.44 10999.515 188.44 ;
    END
  END SET_ICASN[75]
  PIN SET_ICASN[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10859.235 187.44 10859.515 188.44 ;
    END
  END SET_ICASN[74]
  PIN SET_ICASN[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10719.235 187.44 10719.515 188.44 ;
    END
  END SET_ICASN[73]
  PIN SET_ICASN[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10579.235 187.44 10579.515 188.44 ;
    END
  END SET_ICASN[72]
  PIN SET_ICASN[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10439.235 187.44 10439.515 188.44 ;
    END
  END SET_ICASN[71]
  PIN SET_ICASN[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10299.235 187.44 10299.515 188.44 ;
    END
  END SET_ICASN[70]
  PIN SET_ICASN[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10159.235 187.44 10159.515 188.44 ;
    END
  END SET_ICASN[69]
  PIN SET_ICASN[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10019.235 187.44 10019.515 188.44 ;
    END
  END SET_ICASN[68]
  PIN SET_ICASN[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9879.235 187.44 9879.515 188.44 ;
    END
  END SET_ICASN[67]
  PIN SET_ICASN[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9739.235 187.44 9739.515 188.44 ;
    END
  END SET_ICASN[66]
  PIN SET_ICASN[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9599.235 187.44 9599.515 188.44 ;
    END
  END SET_ICASN[65]
  PIN SET_ICASN[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9459.235 187.44 9459.515 188.44 ;
    END
  END SET_ICASN[64]
  PIN SET_ICASN[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9319.235 187.44 9319.515 188.44 ;
    END
  END SET_ICASN[63]
  PIN SET_ICASN[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9179.235 187.44 9179.515 188.44 ;
    END
  END SET_ICASN[62]
  PIN SET_ICASN[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9039.235 187.44 9039.515 188.44 ;
    END
  END SET_ICASN[61]
  PIN SET_ICASN[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8899.235 187.44 8899.515 188.44 ;
    END
  END SET_ICASN[60]
  PIN SET_ICASN[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8759.235 187.44 8759.515 188.44 ;
    END
  END SET_ICASN[59]
  PIN SET_ICASN[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8619.235 187.44 8619.515 188.44 ;
    END
  END SET_ICASN[58]
  PIN SET_ICASN[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8479.235 187.44 8479.515 188.44 ;
    END
  END SET_ICASN[57]
  PIN SET_ICASN[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8339.235 187.44 8339.515 188.44 ;
    END
  END SET_ICASN[56]
  PIN SET_ICASN[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8199.235 187.44 8199.515 188.44 ;
    END
  END SET_ICASN[55]
  PIN SET_ICASN[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8059.235 187.44 8059.515 188.44 ;
    END
  END SET_ICASN[54]
  PIN SET_ICASN[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7919.235 187.44 7919.515 188.44 ;
    END
  END SET_ICASN[53]
  PIN SET_ICASN[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7779.235 187.44 7779.515 188.44 ;
    END
  END SET_ICASN[52]
  PIN SET_ICASN[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7639.235 187.44 7639.515 188.44 ;
    END
  END SET_ICASN[51]
  PIN SET_ICASN[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7499.235 187.44 7499.515 188.44 ;
    END
  END SET_ICASN[50]
  PIN SET_ICASN[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7359.235 187.44 7359.515 188.44 ;
    END
  END SET_ICASN[49]
  PIN SET_ICASN[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7219.235 187.44 7219.515 188.44 ;
    END
  END SET_ICASN[48]
  PIN SET_ICASN[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7079.235 187.44 7079.515 188.44 ;
    END
  END SET_ICASN[47]
  PIN SET_ICASN[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6939.235 187.44 6939.515 188.44 ;
    END
  END SET_ICASN[46]
  PIN SET_ICASN[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6799.235 187.44 6799.515 188.44 ;
    END
  END SET_ICASN[45]
  PIN SET_ICASN[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6659.235 187.44 6659.515 188.44 ;
    END
  END SET_ICASN[44]
  PIN SET_ICASN[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6519.235 187.44 6519.515 188.44 ;
    END
  END SET_ICASN[43]
  PIN SET_ICASN[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6379.235 187.44 6379.515 188.44 ;
    END
  END SET_ICASN[42]
  PIN SET_ICASN[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6239.235 187.44 6239.515 188.44 ;
    END
  END SET_ICASN[41]
  PIN SET_ICASN[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6099.235 187.44 6099.515 188.44 ;
    END
  END SET_ICASN[40]
  PIN SET_ICASN[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5959.235 187.44 5959.515 188.44 ;
    END
  END SET_ICASN[39]
  PIN SET_ICASN[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5819.235 187.44 5819.515 188.44 ;
    END
  END SET_ICASN[38]
  PIN SET_ICASN[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5679.235 187.44 5679.515 188.44 ;
    END
  END SET_ICASN[37]
  PIN SET_ICASN[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5539.235 187.44 5539.515 188.44 ;
    END
  END SET_ICASN[36]
  PIN SET_ICASN[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5399.235 187.44 5399.515 188.44 ;
    END
  END SET_ICASN[35]
  PIN SET_ICASN[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5259.235 187.44 5259.515 188.44 ;
    END
  END SET_ICASN[34]
  PIN SET_ICASN[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5119.235 187.44 5119.515 188.44 ;
    END
  END SET_ICASN[33]
  PIN SET_ICASN[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4979.235 187.44 4979.515 188.44 ;
    END
  END SET_ICASN[32]
  PIN SET_ICASN[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4839.235 187.44 4839.515 188.44 ;
    END
  END SET_ICASN[31]
  PIN SET_ICASN[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4699.235 187.44 4699.515 188.44 ;
    END
  END SET_ICASN[30]
  PIN SET_ICASN[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4559.235 187.44 4559.515 188.44 ;
    END
  END SET_ICASN[29]
  PIN SET_ICASN[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4419.235 187.44 4419.515 188.44 ;
    END
  END SET_ICASN[28]
  PIN SET_ICASN[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4279.235 187.44 4279.515 188.44 ;
    END
  END SET_ICASN[27]
  PIN SET_ICASN[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4139.235 187.44 4139.515 188.44 ;
    END
  END SET_ICASN[26]
  PIN SET_ICASN[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3999.235 187.44 3999.515 188.44 ;
    END
  END SET_ICASN[25]
  PIN SET_ICASN[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3859.235 187.44 3859.515 188.44 ;
    END
  END SET_ICASN[24]
  PIN SET_ICASN[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3719.235 187.44 3719.515 188.44 ;
    END
  END SET_ICASN[23]
  PIN SET_ICASN[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3579.235 187.44 3579.515 188.44 ;
    END
  END SET_ICASN[22]
  PIN SET_ICASN[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3439.235 187.44 3439.515 188.44 ;
    END
  END SET_ICASN[21]
  PIN SET_ICASN[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3299.235 187.44 3299.515 188.44 ;
    END
  END SET_ICASN[20]
  PIN SET_ICASN[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3159.235 187.44 3159.515 188.44 ;
    END
  END SET_ICASN[19]
  PIN SET_ICASN[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3019.235 187.44 3019.515 188.44 ;
    END
  END SET_ICASN[18]
  PIN SET_ICASN[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2879.235 187.44 2879.515 188.44 ;
    END
  END SET_ICASN[17]
  PIN SET_ICASN[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2739.235 187.44 2739.515 188.44 ;
    END
  END SET_ICASN[16]
  PIN SET_ICASN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2599.235 187.44 2599.515 188.44 ;
    END
  END SET_ICASN[15]
  PIN SET_ICASN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2459.235 187.44 2459.515 188.44 ;
    END
  END SET_ICASN[14]
  PIN SET_ICASN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2319.235 187.44 2319.515 188.44 ;
    END
  END SET_ICASN[13]
  PIN SET_ICASN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2179.235 187.44 2179.515 188.44 ;
    END
  END SET_ICASN[12]
  PIN SET_ICASN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2039.235 187.44 2039.515 188.44 ;
    END
  END SET_ICASN[11]
  PIN SET_ICASN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1899.235 187.44 1899.515 188.44 ;
    END
  END SET_ICASN[10]
  PIN SET_ICASN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1759.235 187.44 1759.515 188.44 ;
    END
  END SET_ICASN[9]
  PIN SET_ICASN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1619.235 187.44 1619.515 188.44 ;
    END
  END SET_ICASN[8]
  PIN SET_ICASN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1479.235 187.44 1479.515 188.44 ;
    END
  END SET_ICASN[7]
  PIN SET_ICASN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1339.235 187.44 1339.515 188.44 ;
    END
  END SET_ICASN[6]
  PIN SET_ICASN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1199.235 187.44 1199.515 188.44 ;
    END
  END SET_ICASN[5]
  PIN SET_ICASN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1059.235 187.44 1059.515 188.44 ;
    END
  END SET_ICASN[4]
  PIN SET_ICASN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 919.235 187.44 919.515 188.44 ;
    END
  END SET_ICASN[3]
  PIN SET_ICASN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 779.235 187.44 779.515 188.44 ;
    END
  END SET_ICASN[2]
  PIN SET_ICASN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 639.235 187.44 639.515 188.44 ;
    END
  END SET_ICASN[1]
  PIN SET_ICASN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 499.235 187.44 499.515 188.44 ;
    END
  END SET_ICASN[0]
  PIN SET_IRESET[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18275.315 187.44 18275.595 188.44 ;
    END
  END SET_IRESET[127]
  PIN SET_IRESET[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18135.315 187.44 18135.595 188.44 ;
    END
  END SET_IRESET[126]
  PIN SET_IRESET[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17995.315 187.44 17995.595 188.44 ;
    END
  END SET_IRESET[125]
  PIN SET_IRESET[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17855.315 187.44 17855.595 188.44 ;
    END
  END SET_IRESET[124]
  PIN SET_IRESET[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17715.315 187.44 17715.595 188.44 ;
    END
  END SET_IRESET[123]
  PIN SET_IRESET[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17575.315 187.44 17575.595 188.44 ;
    END
  END SET_IRESET[122]
  PIN SET_IRESET[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17435.315 187.44 17435.595 188.44 ;
    END
  END SET_IRESET[121]
  PIN SET_IRESET[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17295.315 187.44 17295.595 188.44 ;
    END
  END SET_IRESET[120]
  PIN SET_IRESET[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17155.315 187.44 17155.595 188.44 ;
    END
  END SET_IRESET[119]
  PIN SET_IRESET[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17015.315 187.44 17015.595 188.44 ;
    END
  END SET_IRESET[118]
  PIN SET_IRESET[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16875.315 187.44 16875.595 188.44 ;
    END
  END SET_IRESET[117]
  PIN SET_IRESET[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16735.315 187.44 16735.595 188.44 ;
    END
  END SET_IRESET[116]
  PIN SET_IRESET[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16595.315 187.44 16595.595 188.44 ;
    END
  END SET_IRESET[115]
  PIN SET_IRESET[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16455.315 187.44 16455.595 188.44 ;
    END
  END SET_IRESET[114]
  PIN SET_IRESET[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16315.315 187.44 16315.595 188.44 ;
    END
  END SET_IRESET[113]
  PIN SET_IRESET[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16175.315 187.44 16175.595 188.44 ;
    END
  END SET_IRESET[112]
  PIN SET_IRESET[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16035.315 187.44 16035.595 188.44 ;
    END
  END SET_IRESET[111]
  PIN SET_IRESET[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15895.315 187.44 15895.595 188.44 ;
    END
  END SET_IRESET[110]
  PIN SET_IRESET[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15755.315 187.44 15755.595 188.44 ;
    END
  END SET_IRESET[109]
  PIN SET_IRESET[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15615.315 187.44 15615.595 188.44 ;
    END
  END SET_IRESET[108]
  PIN SET_IRESET[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15475.315 187.44 15475.595 188.44 ;
    END
  END SET_IRESET[107]
  PIN SET_IRESET[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15335.315 187.44 15335.595 188.44 ;
    END
  END SET_IRESET[106]
  PIN SET_IRESET[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15195.315 187.44 15195.595 188.44 ;
    END
  END SET_IRESET[105]
  PIN SET_IRESET[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15055.315 187.44 15055.595 188.44 ;
    END
  END SET_IRESET[104]
  PIN SET_IRESET[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14915.315 187.44 14915.595 188.44 ;
    END
  END SET_IRESET[103]
  PIN SET_IRESET[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14775.315 187.44 14775.595 188.44 ;
    END
  END SET_IRESET[102]
  PIN SET_IRESET[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14635.315 187.44 14635.595 188.44 ;
    END
  END SET_IRESET[101]
  PIN SET_IRESET[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14495.315 187.44 14495.595 188.44 ;
    END
  END SET_IRESET[100]
  PIN SET_IRESET[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14355.315 187.44 14355.595 188.44 ;
    END
  END SET_IRESET[99]
  PIN SET_IRESET[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14215.315 187.44 14215.595 188.44 ;
    END
  END SET_IRESET[98]
  PIN SET_IRESET[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14075.315 187.44 14075.595 188.44 ;
    END
  END SET_IRESET[97]
  PIN SET_IRESET[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13935.315 187.44 13935.595 188.44 ;
    END
  END SET_IRESET[96]
  PIN SET_IRESET[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13795.315 187.44 13795.595 188.44 ;
    END
  END SET_IRESET[95]
  PIN SET_IRESET[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13655.315 187.44 13655.595 188.44 ;
    END
  END SET_IRESET[94]
  PIN SET_IRESET[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13515.315 187.44 13515.595 188.44 ;
    END
  END SET_IRESET[93]
  PIN SET_IRESET[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13375.315 187.44 13375.595 188.44 ;
    END
  END SET_IRESET[92]
  PIN SET_IRESET[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13235.315 187.44 13235.595 188.44 ;
    END
  END SET_IRESET[91]
  PIN SET_IRESET[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13095.315 187.44 13095.595 188.44 ;
    END
  END SET_IRESET[90]
  PIN SET_IRESET[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12955.315 187.44 12955.595 188.44 ;
    END
  END SET_IRESET[89]
  PIN SET_IRESET[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12815.315 187.44 12815.595 188.44 ;
    END
  END SET_IRESET[88]
  PIN SET_IRESET[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12675.315 187.44 12675.595 188.44 ;
    END
  END SET_IRESET[87]
  PIN SET_IRESET[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12535.315 187.44 12535.595 188.44 ;
    END
  END SET_IRESET[86]
  PIN SET_IRESET[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12395.315 187.44 12395.595 188.44 ;
    END
  END SET_IRESET[85]
  PIN SET_IRESET[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12255.315 187.44 12255.595 188.44 ;
    END
  END SET_IRESET[84]
  PIN SET_IRESET[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12115.315 187.44 12115.595 188.44 ;
    END
  END SET_IRESET[83]
  PIN SET_IRESET[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11975.315 187.44 11975.595 188.44 ;
    END
  END SET_IRESET[82]
  PIN SET_IRESET[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11835.315 187.44 11835.595 188.44 ;
    END
  END SET_IRESET[81]
  PIN SET_IRESET[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11695.315 187.44 11695.595 188.44 ;
    END
  END SET_IRESET[80]
  PIN SET_IRESET[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11555.315 187.44 11555.595 188.44 ;
    END
  END SET_IRESET[79]
  PIN SET_IRESET[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11415.315 187.44 11415.595 188.44 ;
    END
  END SET_IRESET[78]
  PIN SET_IRESET[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11275.315 187.44 11275.595 188.44 ;
    END
  END SET_IRESET[77]
  PIN SET_IRESET[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11135.315 187.44 11135.595 188.44 ;
    END
  END SET_IRESET[76]
  PIN SET_IRESET[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10995.315 187.44 10995.595 188.44 ;
    END
  END SET_IRESET[75]
  PIN SET_IRESET[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10855.315 187.44 10855.595 188.44 ;
    END
  END SET_IRESET[74]
  PIN SET_IRESET[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10715.315 187.44 10715.595 188.44 ;
    END
  END SET_IRESET[73]
  PIN SET_IRESET[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10575.315 187.44 10575.595 188.44 ;
    END
  END SET_IRESET[72]
  PIN SET_IRESET[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10435.315 187.44 10435.595 188.44 ;
    END
  END SET_IRESET[71]
  PIN SET_IRESET[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10295.315 187.44 10295.595 188.44 ;
    END
  END SET_IRESET[70]
  PIN SET_IRESET[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10155.315 187.44 10155.595 188.44 ;
    END
  END SET_IRESET[69]
  PIN SET_IRESET[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10015.315 187.44 10015.595 188.44 ;
    END
  END SET_IRESET[68]
  PIN SET_IRESET[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9875.315 187.44 9875.595 188.44 ;
    END
  END SET_IRESET[67]
  PIN SET_IRESET[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9735.315 187.44 9735.595 188.44 ;
    END
  END SET_IRESET[66]
  PIN SET_IRESET[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9595.315 187.44 9595.595 188.44 ;
    END
  END SET_IRESET[65]
  PIN SET_IRESET[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9455.315 187.44 9455.595 188.44 ;
    END
  END SET_IRESET[64]
  PIN SET_IRESET[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9315.315 187.44 9315.595 188.44 ;
    END
  END SET_IRESET[63]
  PIN SET_IRESET[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9175.315 187.44 9175.595 188.44 ;
    END
  END SET_IRESET[62]
  PIN SET_IRESET[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9035.315 187.44 9035.595 188.44 ;
    END
  END SET_IRESET[61]
  PIN SET_IRESET[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8895.315 187.44 8895.595 188.44 ;
    END
  END SET_IRESET[60]
  PIN SET_IRESET[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8755.315 187.44 8755.595 188.44 ;
    END
  END SET_IRESET[59]
  PIN SET_IRESET[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8615.315 187.44 8615.595 188.44 ;
    END
  END SET_IRESET[58]
  PIN SET_IRESET[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8475.315 187.44 8475.595 188.44 ;
    END
  END SET_IRESET[57]
  PIN SET_IRESET[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8335.315 187.44 8335.595 188.44 ;
    END
  END SET_IRESET[56]
  PIN SET_IRESET[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8195.315 187.44 8195.595 188.44 ;
    END
  END SET_IRESET[55]
  PIN SET_IRESET[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8055.315 187.44 8055.595 188.44 ;
    END
  END SET_IRESET[54]
  PIN SET_IRESET[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7915.315 187.44 7915.595 188.44 ;
    END
  END SET_IRESET[53]
  PIN SET_IRESET[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7775.315 187.44 7775.595 188.44 ;
    END
  END SET_IRESET[52]
  PIN SET_IRESET[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7635.315 187.44 7635.595 188.44 ;
    END
  END SET_IRESET[51]
  PIN SET_IRESET[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7495.315 187.44 7495.595 188.44 ;
    END
  END SET_IRESET[50]
  PIN SET_IRESET[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7355.315 187.44 7355.595 188.44 ;
    END
  END SET_IRESET[49]
  PIN SET_IRESET[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7215.315 187.44 7215.595 188.44 ;
    END
  END SET_IRESET[48]
  PIN SET_IRESET[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7075.315 187.44 7075.595 188.44 ;
    END
  END SET_IRESET[47]
  PIN SET_IRESET[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6935.315 187.44 6935.595 188.44 ;
    END
  END SET_IRESET[46]
  PIN SET_IRESET[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6795.315 187.44 6795.595 188.44 ;
    END
  END SET_IRESET[45]
  PIN SET_IRESET[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6655.315 187.44 6655.595 188.44 ;
    END
  END SET_IRESET[44]
  PIN SET_IRESET[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6515.315 187.44 6515.595 188.44 ;
    END
  END SET_IRESET[43]
  PIN SET_IRESET[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6375.315 187.44 6375.595 188.44 ;
    END
  END SET_IRESET[42]
  PIN SET_IRESET[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6235.315 187.44 6235.595 188.44 ;
    END
  END SET_IRESET[41]
  PIN SET_IRESET[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6095.315 187.44 6095.595 188.44 ;
    END
  END SET_IRESET[40]
  PIN SET_IRESET[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5955.315 187.44 5955.595 188.44 ;
    END
  END SET_IRESET[39]
  PIN SET_IRESET[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5815.315 187.44 5815.595 188.44 ;
    END
  END SET_IRESET[38]
  PIN SET_IRESET[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5675.315 187.44 5675.595 188.44 ;
    END
  END SET_IRESET[37]
  PIN SET_IRESET[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5535.315 187.44 5535.595 188.44 ;
    END
  END SET_IRESET[36]
  PIN SET_IRESET[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5395.315 187.44 5395.595 188.44 ;
    END
  END SET_IRESET[35]
  PIN SET_IRESET[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5255.315 187.44 5255.595 188.44 ;
    END
  END SET_IRESET[34]
  PIN SET_IRESET[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5115.315 187.44 5115.595 188.44 ;
    END
  END SET_IRESET[33]
  PIN SET_IRESET[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4975.315 187.44 4975.595 188.44 ;
    END
  END SET_IRESET[32]
  PIN SET_IRESET[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4835.315 187.44 4835.595 188.44 ;
    END
  END SET_IRESET[31]
  PIN SET_IRESET[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4695.315 187.44 4695.595 188.44 ;
    END
  END SET_IRESET[30]
  PIN SET_IRESET[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4555.315 187.44 4555.595 188.44 ;
    END
  END SET_IRESET[29]
  PIN SET_IRESET[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4415.315 187.44 4415.595 188.44 ;
    END
  END SET_IRESET[28]
  PIN SET_IRESET[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4275.315 187.44 4275.595 188.44 ;
    END
  END SET_IRESET[27]
  PIN SET_IRESET[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4135.315 187.44 4135.595 188.44 ;
    END
  END SET_IRESET[26]
  PIN SET_IRESET[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3995.315 187.44 3995.595 188.44 ;
    END
  END SET_IRESET[25]
  PIN SET_IRESET[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3855.315 187.44 3855.595 188.44 ;
    END
  END SET_IRESET[24]
  PIN SET_IRESET[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3715.315 187.44 3715.595 188.44 ;
    END
  END SET_IRESET[23]
  PIN SET_IRESET[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3575.315 187.44 3575.595 188.44 ;
    END
  END SET_IRESET[22]
  PIN SET_IRESET[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3435.315 187.44 3435.595 188.44 ;
    END
  END SET_IRESET[21]
  PIN SET_IRESET[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3295.315 187.44 3295.595 188.44 ;
    END
  END SET_IRESET[20]
  PIN SET_IRESET[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3155.315 187.44 3155.595 188.44 ;
    END
  END SET_IRESET[19]
  PIN SET_IRESET[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3015.315 187.44 3015.595 188.44 ;
    END
  END SET_IRESET[18]
  PIN SET_IRESET[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2875.315 187.44 2875.595 188.44 ;
    END
  END SET_IRESET[17]
  PIN SET_IRESET[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2735.315 187.44 2735.595 188.44 ;
    END
  END SET_IRESET[16]
  PIN SET_IRESET[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2595.315 187.44 2595.595 188.44 ;
    END
  END SET_IRESET[15]
  PIN SET_IRESET[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2455.315 187.44 2455.595 188.44 ;
    END
  END SET_IRESET[14]
  PIN SET_IRESET[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2315.315 187.44 2315.595 188.44 ;
    END
  END SET_IRESET[13]
  PIN SET_IRESET[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2175.315 187.44 2175.595 188.44 ;
    END
  END SET_IRESET[12]
  PIN SET_IRESET[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2035.315 187.44 2035.595 188.44 ;
    END
  END SET_IRESET[11]
  PIN SET_IRESET[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1895.315 187.44 1895.595 188.44 ;
    END
  END SET_IRESET[10]
  PIN SET_IRESET[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1755.315 187.44 1755.595 188.44 ;
    END
  END SET_IRESET[9]
  PIN SET_IRESET[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1615.315 187.44 1615.595 188.44 ;
    END
  END SET_IRESET[8]
  PIN SET_IRESET[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1475.315 187.44 1475.595 188.44 ;
    END
  END SET_IRESET[7]
  PIN SET_IRESET[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1335.315 187.44 1335.595 188.44 ;
    END
  END SET_IRESET[6]
  PIN SET_IRESET[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1195.315 187.44 1195.595 188.44 ;
    END
  END SET_IRESET[5]
  PIN SET_IRESET[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1055.315 187.44 1055.595 188.44 ;
    END
  END SET_IRESET[4]
  PIN SET_IRESET[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 915.315 187.44 915.595 188.44 ;
    END
  END SET_IRESET[3]
  PIN SET_IRESET[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 775.315 187.44 775.595 188.44 ;
    END
  END SET_IRESET[2]
  PIN SET_IRESET[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 635.315 187.44 635.595 188.44 ;
    END
  END SET_IRESET[1]
  PIN SET_IRESET[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 495.315 187.44 495.595 188.44 ;
    END
  END SET_IRESET[0]
  PIN SET_IDB[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18271.395 187.44 18271.675 188.44 ;
    END
  END SET_IDB[127]
  PIN SET_IDB[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18131.395 187.44 18131.675 188.44 ;
    END
  END SET_IDB[126]
  PIN SET_IDB[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17991.395 187.44 17991.675 188.44 ;
    END
  END SET_IDB[125]
  PIN SET_IDB[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17851.395 187.44 17851.675 188.44 ;
    END
  END SET_IDB[124]
  PIN SET_IDB[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17711.395 187.44 17711.675 188.44 ;
    END
  END SET_IDB[123]
  PIN SET_IDB[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17571.395 187.44 17571.675 188.44 ;
    END
  END SET_IDB[122]
  PIN SET_IDB[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17431.395 187.44 17431.675 188.44 ;
    END
  END SET_IDB[121]
  PIN SET_IDB[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17291.395 187.44 17291.675 188.44 ;
    END
  END SET_IDB[120]
  PIN SET_IDB[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17151.395 187.44 17151.675 188.44 ;
    END
  END SET_IDB[119]
  PIN SET_IDB[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17011.395 187.44 17011.675 188.44 ;
    END
  END SET_IDB[118]
  PIN SET_IDB[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16871.395 187.44 16871.675 188.44 ;
    END
  END SET_IDB[117]
  PIN SET_IDB[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16731.395 187.44 16731.675 188.44 ;
    END
  END SET_IDB[116]
  PIN SET_IDB[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16591.395 187.44 16591.675 188.44 ;
    END
  END SET_IDB[115]
  PIN SET_IDB[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16451.395 187.44 16451.675 188.44 ;
    END
  END SET_IDB[114]
  PIN SET_IDB[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16311.395 187.44 16311.675 188.44 ;
    END
  END SET_IDB[113]
  PIN SET_IDB[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16171.395 187.44 16171.675 188.44 ;
    END
  END SET_IDB[112]
  PIN SET_IDB[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16031.395 187.44 16031.675 188.44 ;
    END
  END SET_IDB[111]
  PIN SET_IDB[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15891.395 187.44 15891.675 188.44 ;
    END
  END SET_IDB[110]
  PIN SET_IDB[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15751.395 187.44 15751.675 188.44 ;
    END
  END SET_IDB[109]
  PIN SET_IDB[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15611.395 187.44 15611.675 188.44 ;
    END
  END SET_IDB[108]
  PIN SET_IDB[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15471.395 187.44 15471.675 188.44 ;
    END
  END SET_IDB[107]
  PIN SET_IDB[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15331.395 187.44 15331.675 188.44 ;
    END
  END SET_IDB[106]
  PIN SET_IDB[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15191.395 187.44 15191.675 188.44 ;
    END
  END SET_IDB[105]
  PIN SET_IDB[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15051.395 187.44 15051.675 188.44 ;
    END
  END SET_IDB[104]
  PIN SET_IDB[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14911.395 187.44 14911.675 188.44 ;
    END
  END SET_IDB[103]
  PIN SET_IDB[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14771.395 187.44 14771.675 188.44 ;
    END
  END SET_IDB[102]
  PIN SET_IDB[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14631.395 187.44 14631.675 188.44 ;
    END
  END SET_IDB[101]
  PIN SET_IDB[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14491.395 187.44 14491.675 188.44 ;
    END
  END SET_IDB[100]
  PIN SET_IDB[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14351.395 187.44 14351.675 188.44 ;
    END
  END SET_IDB[99]
  PIN SET_IDB[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14211.395 187.44 14211.675 188.44 ;
    END
  END SET_IDB[98]
  PIN SET_IDB[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14071.395 187.44 14071.675 188.44 ;
    END
  END SET_IDB[97]
  PIN SET_IDB[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13931.395 187.44 13931.675 188.44 ;
    END
  END SET_IDB[96]
  PIN SET_IDB[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13791.395 187.44 13791.675 188.44 ;
    END
  END SET_IDB[95]
  PIN SET_IDB[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13651.395 187.44 13651.675 188.44 ;
    END
  END SET_IDB[94]
  PIN SET_IDB[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13511.395 187.44 13511.675 188.44 ;
    END
  END SET_IDB[93]
  PIN SET_IDB[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13371.395 187.44 13371.675 188.44 ;
    END
  END SET_IDB[92]
  PIN SET_IDB[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13231.395 187.44 13231.675 188.44 ;
    END
  END SET_IDB[91]
  PIN SET_IDB[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13091.395 187.44 13091.675 188.44 ;
    END
  END SET_IDB[90]
  PIN SET_IDB[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12951.395 187.44 12951.675 188.44 ;
    END
  END SET_IDB[89]
  PIN SET_IDB[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12811.395 187.44 12811.675 188.44 ;
    END
  END SET_IDB[88]
  PIN SET_IDB[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12671.395 187.44 12671.675 188.44 ;
    END
  END SET_IDB[87]
  PIN SET_IDB[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12531.395 187.44 12531.675 188.44 ;
    END
  END SET_IDB[86]
  PIN SET_IDB[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12391.395 187.44 12391.675 188.44 ;
    END
  END SET_IDB[85]
  PIN SET_IDB[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12251.395 187.44 12251.675 188.44 ;
    END
  END SET_IDB[84]
  PIN SET_IDB[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12111.395 187.44 12111.675 188.44 ;
    END
  END SET_IDB[83]
  PIN SET_IDB[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11971.395 187.44 11971.675 188.44 ;
    END
  END SET_IDB[82]
  PIN SET_IDB[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11831.395 187.44 11831.675 188.44 ;
    END
  END SET_IDB[81]
  PIN SET_IDB[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11691.395 187.44 11691.675 188.44 ;
    END
  END SET_IDB[80]
  PIN SET_IDB[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11551.395 187.44 11551.675 188.44 ;
    END
  END SET_IDB[79]
  PIN SET_IDB[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11411.395 187.44 11411.675 188.44 ;
    END
  END SET_IDB[78]
  PIN SET_IDB[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11271.395 187.44 11271.675 188.44 ;
    END
  END SET_IDB[77]
  PIN SET_IDB[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11131.395 187.44 11131.675 188.44 ;
    END
  END SET_IDB[76]
  PIN SET_IDB[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10991.395 187.44 10991.675 188.44 ;
    END
  END SET_IDB[75]
  PIN SET_IDB[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10851.395 187.44 10851.675 188.44 ;
    END
  END SET_IDB[74]
  PIN SET_IDB[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10711.395 187.44 10711.675 188.44 ;
    END
  END SET_IDB[73]
  PIN SET_IDB[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10571.395 187.44 10571.675 188.44 ;
    END
  END SET_IDB[72]
  PIN SET_IDB[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10431.395 187.44 10431.675 188.44 ;
    END
  END SET_IDB[71]
  PIN SET_IDB[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10291.395 187.44 10291.675 188.44 ;
    END
  END SET_IDB[70]
  PIN SET_IDB[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10151.395 187.44 10151.675 188.44 ;
    END
  END SET_IDB[69]
  PIN SET_IDB[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10011.395 187.44 10011.675 188.44 ;
    END
  END SET_IDB[68]
  PIN SET_IDB[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9871.395 187.44 9871.675 188.44 ;
    END
  END SET_IDB[67]
  PIN SET_IDB[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9731.395 187.44 9731.675 188.44 ;
    END
  END SET_IDB[66]
  PIN SET_IDB[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9591.395 187.44 9591.675 188.44 ;
    END
  END SET_IDB[65]
  PIN SET_IDB[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9451.395 187.44 9451.675 188.44 ;
    END
  END SET_IDB[64]
  PIN SET_IDB[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9311.395 187.44 9311.675 188.44 ;
    END
  END SET_IDB[63]
  PIN SET_IDB[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9171.395 187.44 9171.675 188.44 ;
    END
  END SET_IDB[62]
  PIN SET_IDB[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9031.395 187.44 9031.675 188.44 ;
    END
  END SET_IDB[61]
  PIN SET_IDB[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8891.395 187.44 8891.675 188.44 ;
    END
  END SET_IDB[60]
  PIN SET_IDB[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8751.395 187.44 8751.675 188.44 ;
    END
  END SET_IDB[59]
  PIN SET_IDB[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8611.395 187.44 8611.675 188.44 ;
    END
  END SET_IDB[58]
  PIN SET_IDB[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8471.395 187.44 8471.675 188.44 ;
    END
  END SET_IDB[57]
  PIN SET_IDB[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8331.395 187.44 8331.675 188.44 ;
    END
  END SET_IDB[56]
  PIN SET_IDB[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8191.395 187.44 8191.675 188.44 ;
    END
  END SET_IDB[55]
  PIN SET_IDB[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8051.395 187.44 8051.675 188.44 ;
    END
  END SET_IDB[54]
  PIN SET_IDB[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7911.395 187.44 7911.675 188.44 ;
    END
  END SET_IDB[53]
  PIN SET_IDB[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7771.395 187.44 7771.675 188.44 ;
    END
  END SET_IDB[52]
  PIN SET_IDB[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7631.395 187.44 7631.675 188.44 ;
    END
  END SET_IDB[51]
  PIN SET_IDB[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7491.395 187.44 7491.675 188.44 ;
    END
  END SET_IDB[50]
  PIN SET_IDB[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7351.395 187.44 7351.675 188.44 ;
    END
  END SET_IDB[49]
  PIN SET_IDB[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7211.395 187.44 7211.675 188.44 ;
    END
  END SET_IDB[48]
  PIN SET_IDB[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7071.395 187.44 7071.675 188.44 ;
    END
  END SET_IDB[47]
  PIN SET_IDB[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6931.395 187.44 6931.675 188.44 ;
    END
  END SET_IDB[46]
  PIN SET_IDB[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6791.395 187.44 6791.675 188.44 ;
    END
  END SET_IDB[45]
  PIN SET_IDB[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6651.395 187.44 6651.675 188.44 ;
    END
  END SET_IDB[44]
  PIN SET_IDB[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6511.395 187.44 6511.675 188.44 ;
    END
  END SET_IDB[43]
  PIN SET_IDB[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6371.395 187.44 6371.675 188.44 ;
    END
  END SET_IDB[42]
  PIN SET_IDB[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6231.395 187.44 6231.675 188.44 ;
    END
  END SET_IDB[41]
  PIN SET_IDB[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6091.395 187.44 6091.675 188.44 ;
    END
  END SET_IDB[40]
  PIN SET_IDB[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5951.395 187.44 5951.675 188.44 ;
    END
  END SET_IDB[39]
  PIN SET_IDB[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5811.395 187.44 5811.675 188.44 ;
    END
  END SET_IDB[38]
  PIN SET_IDB[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5671.395 187.44 5671.675 188.44 ;
    END
  END SET_IDB[37]
  PIN SET_IDB[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5531.395 187.44 5531.675 188.44 ;
    END
  END SET_IDB[36]
  PIN SET_IDB[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5391.395 187.44 5391.675 188.44 ;
    END
  END SET_IDB[35]
  PIN SET_IDB[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5251.395 187.44 5251.675 188.44 ;
    END
  END SET_IDB[34]
  PIN SET_IDB[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5111.395 187.44 5111.675 188.44 ;
    END
  END SET_IDB[33]
  PIN SET_IDB[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4971.395 187.44 4971.675 188.44 ;
    END
  END SET_IDB[32]
  PIN SET_IDB[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4831.395 187.44 4831.675 188.44 ;
    END
  END SET_IDB[31]
  PIN SET_IDB[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4691.395 187.44 4691.675 188.44 ;
    END
  END SET_IDB[30]
  PIN SET_IDB[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4551.395 187.44 4551.675 188.44 ;
    END
  END SET_IDB[29]
  PIN SET_IDB[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4411.395 187.44 4411.675 188.44 ;
    END
  END SET_IDB[28]
  PIN SET_IDB[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4271.395 187.44 4271.675 188.44 ;
    END
  END SET_IDB[27]
  PIN SET_IDB[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4131.395 187.44 4131.675 188.44 ;
    END
  END SET_IDB[26]
  PIN SET_IDB[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3991.395 187.44 3991.675 188.44 ;
    END
  END SET_IDB[25]
  PIN SET_IDB[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3851.395 187.44 3851.675 188.44 ;
    END
  END SET_IDB[24]
  PIN SET_IDB[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3711.395 187.44 3711.675 188.44 ;
    END
  END SET_IDB[23]
  PIN SET_IDB[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3571.395 187.44 3571.675 188.44 ;
    END
  END SET_IDB[22]
  PIN SET_IDB[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3431.395 187.44 3431.675 188.44 ;
    END
  END SET_IDB[21]
  PIN SET_IDB[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3291.395 187.44 3291.675 188.44 ;
    END
  END SET_IDB[20]
  PIN SET_IDB[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3151.395 187.44 3151.675 188.44 ;
    END
  END SET_IDB[19]
  PIN SET_IDB[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3011.395 187.44 3011.675 188.44 ;
    END
  END SET_IDB[18]
  PIN SET_IDB[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2871.395 187.44 2871.675 188.44 ;
    END
  END SET_IDB[17]
  PIN SET_IDB[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2731.395 187.44 2731.675 188.44 ;
    END
  END SET_IDB[16]
  PIN SET_IDB[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2591.395 187.44 2591.675 188.44 ;
    END
  END SET_IDB[15]
  PIN SET_IDB[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2451.395 187.44 2451.675 188.44 ;
    END
  END SET_IDB[14]
  PIN SET_IDB[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2311.395 187.44 2311.675 188.44 ;
    END
  END SET_IDB[13]
  PIN SET_IDB[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2171.395 187.44 2171.675 188.44 ;
    END
  END SET_IDB[12]
  PIN SET_IDB[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2031.395 187.44 2031.675 188.44 ;
    END
  END SET_IDB[11]
  PIN SET_IDB[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1891.395 187.44 1891.675 188.44 ;
    END
  END SET_IDB[10]
  PIN SET_IDB[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1751.395 187.44 1751.675 188.44 ;
    END
  END SET_IDB[9]
  PIN SET_IDB[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1611.395 187.44 1611.675 188.44 ;
    END
  END SET_IDB[8]
  PIN SET_IDB[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1471.395 187.44 1471.675 188.44 ;
    END
  END SET_IDB[7]
  PIN SET_IDB[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1331.395 187.44 1331.675 188.44 ;
    END
  END SET_IDB[6]
  PIN SET_IDB[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1191.395 187.44 1191.675 188.44 ;
    END
  END SET_IDB[5]
  PIN SET_IDB[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1051.395 187.44 1051.675 188.44 ;
    END
  END SET_IDB[4]
  PIN SET_IDB[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 911.395 187.44 911.675 188.44 ;
    END
  END SET_IDB[3]
  PIN SET_IDB[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 771.395 187.44 771.675 188.44 ;
    END
  END SET_IDB[2]
  PIN SET_IDB[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 631.395 187.44 631.675 188.44 ;
    END
  END SET_IDB[1]
  PIN SET_IDB[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 491.395 187.44 491.675 188.44 ;
    END
  END SET_IDB[0]
  PIN SET_ITHR[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18267.475 187.44 18267.755 188.44 ;
    END
  END SET_ITHR[127]
  PIN SET_ITHR[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18127.475 187.44 18127.755 188.44 ;
    END
  END SET_ITHR[126]
  PIN SET_ITHR[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17987.475 187.44 17987.755 188.44 ;
    END
  END SET_ITHR[125]
  PIN SET_ITHR[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17847.475 187.44 17847.755 188.44 ;
    END
  END SET_ITHR[124]
  PIN SET_ITHR[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17707.475 187.44 17707.755 188.44 ;
    END
  END SET_ITHR[123]
  PIN SET_ITHR[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17567.475 187.44 17567.755 188.44 ;
    END
  END SET_ITHR[122]
  PIN SET_ITHR[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17427.475 187.44 17427.755 188.44 ;
    END
  END SET_ITHR[121]
  PIN SET_ITHR[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17287.475 187.44 17287.755 188.44 ;
    END
  END SET_ITHR[120]
  PIN SET_ITHR[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17147.475 187.44 17147.755 188.44 ;
    END
  END SET_ITHR[119]
  PIN SET_ITHR[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17007.475 187.44 17007.755 188.44 ;
    END
  END SET_ITHR[118]
  PIN SET_ITHR[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16867.475 187.44 16867.755 188.44 ;
    END
  END SET_ITHR[117]
  PIN SET_ITHR[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16727.475 187.44 16727.755 188.44 ;
    END
  END SET_ITHR[116]
  PIN SET_ITHR[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16587.475 187.44 16587.755 188.44 ;
    END
  END SET_ITHR[115]
  PIN SET_ITHR[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16447.475 187.44 16447.755 188.44 ;
    END
  END SET_ITHR[114]
  PIN SET_ITHR[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16307.475 187.44 16307.755 188.44 ;
    END
  END SET_ITHR[113]
  PIN SET_ITHR[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16167.475 187.44 16167.755 188.44 ;
    END
  END SET_ITHR[112]
  PIN SET_ITHR[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16027.475 187.44 16027.755 188.44 ;
    END
  END SET_ITHR[111]
  PIN SET_ITHR[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15887.475 187.44 15887.755 188.44 ;
    END
  END SET_ITHR[110]
  PIN SET_ITHR[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15747.475 187.44 15747.755 188.44 ;
    END
  END SET_ITHR[109]
  PIN SET_ITHR[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15607.475 187.44 15607.755 188.44 ;
    END
  END SET_ITHR[108]
  PIN SET_ITHR[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15467.475 187.44 15467.755 188.44 ;
    END
  END SET_ITHR[107]
  PIN SET_ITHR[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15327.475 187.44 15327.755 188.44 ;
    END
  END SET_ITHR[106]
  PIN SET_ITHR[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15187.475 187.44 15187.755 188.44 ;
    END
  END SET_ITHR[105]
  PIN SET_ITHR[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15047.475 187.44 15047.755 188.44 ;
    END
  END SET_ITHR[104]
  PIN SET_ITHR[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14907.475 187.44 14907.755 188.44 ;
    END
  END SET_ITHR[103]
  PIN SET_ITHR[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14767.475 187.44 14767.755 188.44 ;
    END
  END SET_ITHR[102]
  PIN SET_ITHR[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14627.475 187.44 14627.755 188.44 ;
    END
  END SET_ITHR[101]
  PIN SET_ITHR[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14487.475 187.44 14487.755 188.44 ;
    END
  END SET_ITHR[100]
  PIN SET_ITHR[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14347.475 187.44 14347.755 188.44 ;
    END
  END SET_ITHR[99]
  PIN SET_ITHR[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14207.475 187.44 14207.755 188.44 ;
    END
  END SET_ITHR[98]
  PIN SET_ITHR[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14067.475 187.44 14067.755 188.44 ;
    END
  END SET_ITHR[97]
  PIN SET_ITHR[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13927.475 187.44 13927.755 188.44 ;
    END
  END SET_ITHR[96]
  PIN SET_ITHR[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13787.475 187.44 13787.755 188.44 ;
    END
  END SET_ITHR[95]
  PIN SET_ITHR[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13647.475 187.44 13647.755 188.44 ;
    END
  END SET_ITHR[94]
  PIN SET_ITHR[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13507.475 187.44 13507.755 188.44 ;
    END
  END SET_ITHR[93]
  PIN SET_ITHR[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13367.475 187.44 13367.755 188.44 ;
    END
  END SET_ITHR[92]
  PIN SET_ITHR[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13227.475 187.44 13227.755 188.44 ;
    END
  END SET_ITHR[91]
  PIN SET_ITHR[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13087.475 187.44 13087.755 188.44 ;
    END
  END SET_ITHR[90]
  PIN SET_ITHR[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12947.475 187.44 12947.755 188.44 ;
    END
  END SET_ITHR[89]
  PIN SET_ITHR[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12807.475 187.44 12807.755 188.44 ;
    END
  END SET_ITHR[88]
  PIN SET_ITHR[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12667.475 187.44 12667.755 188.44 ;
    END
  END SET_ITHR[87]
  PIN SET_ITHR[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12527.475 187.44 12527.755 188.44 ;
    END
  END SET_ITHR[86]
  PIN SET_ITHR[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12387.475 187.44 12387.755 188.44 ;
    END
  END SET_ITHR[85]
  PIN SET_ITHR[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12247.475 187.44 12247.755 188.44 ;
    END
  END SET_ITHR[84]
  PIN SET_ITHR[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12107.475 187.44 12107.755 188.44 ;
    END
  END SET_ITHR[83]
  PIN SET_ITHR[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11967.475 187.44 11967.755 188.44 ;
    END
  END SET_ITHR[82]
  PIN SET_ITHR[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11827.475 187.44 11827.755 188.44 ;
    END
  END SET_ITHR[81]
  PIN SET_ITHR[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11687.475 187.44 11687.755 188.44 ;
    END
  END SET_ITHR[80]
  PIN SET_ITHR[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11547.475 187.44 11547.755 188.44 ;
    END
  END SET_ITHR[79]
  PIN SET_ITHR[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11407.475 187.44 11407.755 188.44 ;
    END
  END SET_ITHR[78]
  PIN SET_ITHR[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11267.475 187.44 11267.755 188.44 ;
    END
  END SET_ITHR[77]
  PIN SET_ITHR[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11127.475 187.44 11127.755 188.44 ;
    END
  END SET_ITHR[76]
  PIN SET_ITHR[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10987.475 187.44 10987.755 188.44 ;
    END
  END SET_ITHR[75]
  PIN SET_ITHR[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10847.475 187.44 10847.755 188.44 ;
    END
  END SET_ITHR[74]
  PIN SET_ITHR[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10707.475 187.44 10707.755 188.44 ;
    END
  END SET_ITHR[73]
  PIN SET_ITHR[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10567.475 187.44 10567.755 188.44 ;
    END
  END SET_ITHR[72]
  PIN SET_ITHR[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10427.475 187.44 10427.755 188.44 ;
    END
  END SET_ITHR[71]
  PIN SET_ITHR[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10287.475 187.44 10287.755 188.44 ;
    END
  END SET_ITHR[70]
  PIN SET_ITHR[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10147.475 187.44 10147.755 188.44 ;
    END
  END SET_ITHR[69]
  PIN SET_ITHR[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10007.475 187.44 10007.755 188.44 ;
    END
  END SET_ITHR[68]
  PIN SET_ITHR[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9867.475 187.44 9867.755 188.44 ;
    END
  END SET_ITHR[67]
  PIN SET_ITHR[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9727.475 187.44 9727.755 188.44 ;
    END
  END SET_ITHR[66]
  PIN SET_ITHR[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9587.475 187.44 9587.755 188.44 ;
    END
  END SET_ITHR[65]
  PIN SET_ITHR[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9447.475 187.44 9447.755 188.44 ;
    END
  END SET_ITHR[64]
  PIN SET_ITHR[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9307.475 187.44 9307.755 188.44 ;
    END
  END SET_ITHR[63]
  PIN SET_ITHR[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9167.475 187.44 9167.755 188.44 ;
    END
  END SET_ITHR[62]
  PIN SET_ITHR[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9027.475 187.44 9027.755 188.44 ;
    END
  END SET_ITHR[61]
  PIN SET_ITHR[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8887.475 187.44 8887.755 188.44 ;
    END
  END SET_ITHR[60]
  PIN SET_ITHR[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8747.475 187.44 8747.755 188.44 ;
    END
  END SET_ITHR[59]
  PIN SET_ITHR[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8607.475 187.44 8607.755 188.44 ;
    END
  END SET_ITHR[58]
  PIN SET_ITHR[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8467.475 187.44 8467.755 188.44 ;
    END
  END SET_ITHR[57]
  PIN SET_ITHR[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8327.475 187.44 8327.755 188.44 ;
    END
  END SET_ITHR[56]
  PIN SET_ITHR[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8187.475 187.44 8187.755 188.44 ;
    END
  END SET_ITHR[55]
  PIN SET_ITHR[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8047.475 187.44 8047.755 188.44 ;
    END
  END SET_ITHR[54]
  PIN SET_ITHR[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7907.475 187.44 7907.755 188.44 ;
    END
  END SET_ITHR[53]
  PIN SET_ITHR[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7767.475 187.44 7767.755 188.44 ;
    END
  END SET_ITHR[52]
  PIN SET_ITHR[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7627.475 187.44 7627.755 188.44 ;
    END
  END SET_ITHR[51]
  PIN SET_ITHR[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7487.475 187.44 7487.755 188.44 ;
    END
  END SET_ITHR[50]
  PIN SET_ITHR[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7347.475 187.44 7347.755 188.44 ;
    END
  END SET_ITHR[49]
  PIN SET_ITHR[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7207.475 187.44 7207.755 188.44 ;
    END
  END SET_ITHR[48]
  PIN SET_ITHR[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7067.475 187.44 7067.755 188.44 ;
    END
  END SET_ITHR[47]
  PIN SET_ITHR[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6927.475 187.44 6927.755 188.44 ;
    END
  END SET_ITHR[46]
  PIN SET_ITHR[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6787.475 187.44 6787.755 188.44 ;
    END
  END SET_ITHR[45]
  PIN SET_ITHR[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6647.475 187.44 6647.755 188.44 ;
    END
  END SET_ITHR[44]
  PIN SET_ITHR[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6507.475 187.44 6507.755 188.44 ;
    END
  END SET_ITHR[43]
  PIN SET_ITHR[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6367.475 187.44 6367.755 188.44 ;
    END
  END SET_ITHR[42]
  PIN SET_ITHR[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6227.475 187.44 6227.755 188.44 ;
    END
  END SET_ITHR[41]
  PIN SET_ITHR[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6087.475 187.44 6087.755 188.44 ;
    END
  END SET_ITHR[40]
  PIN SET_ITHR[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5947.475 187.44 5947.755 188.44 ;
    END
  END SET_ITHR[39]
  PIN SET_ITHR[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5807.475 187.44 5807.755 188.44 ;
    END
  END SET_ITHR[38]
  PIN SET_ITHR[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5667.475 187.44 5667.755 188.44 ;
    END
  END SET_ITHR[37]
  PIN SET_ITHR[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5527.475 187.44 5527.755 188.44 ;
    END
  END SET_ITHR[36]
  PIN SET_ITHR[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5387.475 187.44 5387.755 188.44 ;
    END
  END SET_ITHR[35]
  PIN SET_ITHR[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5247.475 187.44 5247.755 188.44 ;
    END
  END SET_ITHR[34]
  PIN SET_ITHR[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5107.475 187.44 5107.755 188.44 ;
    END
  END SET_ITHR[33]
  PIN SET_ITHR[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4967.475 187.44 4967.755 188.44 ;
    END
  END SET_ITHR[32]
  PIN SET_ITHR[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4827.475 187.44 4827.755 188.44 ;
    END
  END SET_ITHR[31]
  PIN SET_ITHR[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4687.475 187.44 4687.755 188.44 ;
    END
  END SET_ITHR[30]
  PIN SET_ITHR[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4547.475 187.44 4547.755 188.44 ;
    END
  END SET_ITHR[29]
  PIN SET_ITHR[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4407.475 187.44 4407.755 188.44 ;
    END
  END SET_ITHR[28]
  PIN SET_ITHR[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4267.475 187.44 4267.755 188.44 ;
    END
  END SET_ITHR[27]
  PIN SET_ITHR[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4127.475 187.44 4127.755 188.44 ;
    END
  END SET_ITHR[26]
  PIN SET_ITHR[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3987.475 187.44 3987.755 188.44 ;
    END
  END SET_ITHR[25]
  PIN SET_ITHR[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3847.475 187.44 3847.755 188.44 ;
    END
  END SET_ITHR[24]
  PIN SET_ITHR[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3707.475 187.44 3707.755 188.44 ;
    END
  END SET_ITHR[23]
  PIN SET_ITHR[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3567.475 187.44 3567.755 188.44 ;
    END
  END SET_ITHR[22]
  PIN SET_ITHR[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3427.475 187.44 3427.755 188.44 ;
    END
  END SET_ITHR[21]
  PIN SET_ITHR[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3287.475 187.44 3287.755 188.44 ;
    END
  END SET_ITHR[20]
  PIN SET_ITHR[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3147.475 187.44 3147.755 188.44 ;
    END
  END SET_ITHR[19]
  PIN SET_ITHR[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3007.475 187.44 3007.755 188.44 ;
    END
  END SET_ITHR[18]
  PIN SET_ITHR[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2867.475 187.44 2867.755 188.44 ;
    END
  END SET_ITHR[17]
  PIN SET_ITHR[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2727.475 187.44 2727.755 188.44 ;
    END
  END SET_ITHR[16]
  PIN SET_ITHR[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2587.475 187.44 2587.755 188.44 ;
    END
  END SET_ITHR[15]
  PIN SET_ITHR[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2447.475 187.44 2447.755 188.44 ;
    END
  END SET_ITHR[14]
  PIN SET_ITHR[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2307.475 187.44 2307.755 188.44 ;
    END
  END SET_ITHR[13]
  PIN SET_ITHR[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2167.475 187.44 2167.755 188.44 ;
    END
  END SET_ITHR[12]
  PIN SET_ITHR[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2027.475 187.44 2027.755 188.44 ;
    END
  END SET_ITHR[11]
  PIN SET_ITHR[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1887.475 187.44 1887.755 188.44 ;
    END
  END SET_ITHR[10]
  PIN SET_ITHR[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1747.475 187.44 1747.755 188.44 ;
    END
  END SET_ITHR[9]
  PIN SET_ITHR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1607.475 187.44 1607.755 188.44 ;
    END
  END SET_ITHR[8]
  PIN SET_ITHR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1467.475 187.44 1467.755 188.44 ;
    END
  END SET_ITHR[7]
  PIN SET_ITHR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1327.475 187.44 1327.755 188.44 ;
    END
  END SET_ITHR[6]
  PIN SET_ITHR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1187.475 187.44 1187.755 188.44 ;
    END
  END SET_ITHR[5]
  PIN SET_ITHR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1047.475 187.44 1047.755 188.44 ;
    END
  END SET_ITHR[4]
  PIN SET_ITHR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 907.475 187.44 907.755 188.44 ;
    END
  END SET_ITHR[3]
  PIN SET_ITHR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 767.475 187.44 767.755 188.44 ;
    END
  END SET_ITHR[2]
  PIN SET_ITHR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 627.475 187.44 627.755 188.44 ;
    END
  END SET_ITHR[1]
  PIN SET_ITHR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 487.475 187.44 487.755 188.44 ;
    END
  END SET_ITHR[0]
  PIN SWCNTL_IBIAS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9408.115 187.44 9408.675 188.44 ;
    END
  END SWCNTL_IBIAS
  PIN SET_IBIAS[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18263.555 187.44 18263.835 188.44 ;
    END
  END SET_IBIAS[127]
  PIN SET_IBIAS[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18123.555 187.44 18123.835 188.44 ;
    END
  END SET_IBIAS[126]
  PIN SET_IBIAS[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17983.555 187.44 17983.835 188.44 ;
    END
  END SET_IBIAS[125]
  PIN SET_IBIAS[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17843.555 187.44 17843.835 188.44 ;
    END
  END SET_IBIAS[124]
  PIN SET_IBIAS[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17703.555 187.44 17703.835 188.44 ;
    END
  END SET_IBIAS[123]
  PIN SET_IBIAS[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17563.555 187.44 17563.835 188.44 ;
    END
  END SET_IBIAS[122]
  PIN SET_IBIAS[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17423.555 187.44 17423.835 188.44 ;
    END
  END SET_IBIAS[121]
  PIN SET_IBIAS[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17283.555 187.44 17283.835 188.44 ;
    END
  END SET_IBIAS[120]
  PIN SET_IBIAS[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17143.555 187.44 17143.835 188.44 ;
    END
  END SET_IBIAS[119]
  PIN SET_IBIAS[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17003.555 187.44 17003.835 188.44 ;
    END
  END SET_IBIAS[118]
  PIN SET_IBIAS[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16863.555 187.44 16863.835 188.44 ;
    END
  END SET_IBIAS[117]
  PIN SET_IBIAS[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16723.555 187.44 16723.835 188.44 ;
    END
  END SET_IBIAS[116]
  PIN SET_IBIAS[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16583.555 187.44 16583.835 188.44 ;
    END
  END SET_IBIAS[115]
  PIN SET_IBIAS[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16443.555 187.44 16443.835 188.44 ;
    END
  END SET_IBIAS[114]
  PIN SET_IBIAS[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16303.555 187.44 16303.835 188.44 ;
    END
  END SET_IBIAS[113]
  PIN SET_IBIAS[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16163.555 187.44 16163.835 188.44 ;
    END
  END SET_IBIAS[112]
  PIN SET_IBIAS[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16023.555 187.44 16023.835 188.44 ;
    END
  END SET_IBIAS[111]
  PIN SET_IBIAS[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15883.555 187.44 15883.835 188.44 ;
    END
  END SET_IBIAS[110]
  PIN SET_IBIAS[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15743.555 187.44 15743.835 188.44 ;
    END
  END SET_IBIAS[109]
  PIN SET_IBIAS[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15603.555 187.44 15603.835 188.44 ;
    END
  END SET_IBIAS[108]
  PIN SET_IBIAS[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15463.555 187.44 15463.835 188.44 ;
    END
  END SET_IBIAS[107]
  PIN SET_IBIAS[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15323.555 187.44 15323.835 188.44 ;
    END
  END SET_IBIAS[106]
  PIN SET_IBIAS[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15183.555 187.44 15183.835 188.44 ;
    END
  END SET_IBIAS[105]
  PIN SET_IBIAS[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15043.555 187.44 15043.835 188.44 ;
    END
  END SET_IBIAS[104]
  PIN SET_IBIAS[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14903.555 187.44 14903.835 188.44 ;
    END
  END SET_IBIAS[103]
  PIN SET_IBIAS[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14763.555 187.44 14763.835 188.44 ;
    END
  END SET_IBIAS[102]
  PIN SET_IBIAS[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14623.555 187.44 14623.835 188.44 ;
    END
  END SET_IBIAS[101]
  PIN SET_IBIAS[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14483.555 187.44 14483.835 188.44 ;
    END
  END SET_IBIAS[100]
  PIN SET_IBIAS[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14343.555 187.44 14343.835 188.44 ;
    END
  END SET_IBIAS[99]
  PIN SET_IBIAS[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14203.555 187.44 14203.835 188.44 ;
    END
  END SET_IBIAS[98]
  PIN SET_IBIAS[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14063.555 187.44 14063.835 188.44 ;
    END
  END SET_IBIAS[97]
  PIN SET_IBIAS[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13923.555 187.44 13923.835 188.44 ;
    END
  END SET_IBIAS[96]
  PIN SET_IBIAS[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13783.555 187.44 13783.835 188.44 ;
    END
  END SET_IBIAS[95]
  PIN SET_IBIAS[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13643.555 187.44 13643.835 188.44 ;
    END
  END SET_IBIAS[94]
  PIN SET_IBIAS[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13503.555 187.44 13503.835 188.44 ;
    END
  END SET_IBIAS[93]
  PIN SET_IBIAS[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13363.555 187.44 13363.835 188.44 ;
    END
  END SET_IBIAS[92]
  PIN SET_IBIAS[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13223.555 187.44 13223.835 188.44 ;
    END
  END SET_IBIAS[91]
  PIN SET_IBIAS[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13083.555 187.44 13083.835 188.44 ;
    END
  END SET_IBIAS[90]
  PIN SET_IBIAS[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12943.555 187.44 12943.835 188.44 ;
    END
  END SET_IBIAS[89]
  PIN SET_IBIAS[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12803.555 187.44 12803.835 188.44 ;
    END
  END SET_IBIAS[88]
  PIN SET_IBIAS[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12663.555 187.44 12663.835 188.44 ;
    END
  END SET_IBIAS[87]
  PIN SET_IBIAS[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12523.555 187.44 12523.835 188.44 ;
    END
  END SET_IBIAS[86]
  PIN SET_IBIAS[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12383.555 187.44 12383.835 188.44 ;
    END
  END SET_IBIAS[85]
  PIN SET_IBIAS[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12243.555 187.44 12243.835 188.44 ;
    END
  END SET_IBIAS[84]
  PIN SET_IBIAS[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12103.555 187.44 12103.835 188.44 ;
    END
  END SET_IBIAS[83]
  PIN SET_IBIAS[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11963.555 187.44 11963.835 188.44 ;
    END
  END SET_IBIAS[82]
  PIN SET_IBIAS[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11823.555 187.44 11823.835 188.44 ;
    END
  END SET_IBIAS[81]
  PIN SET_IBIAS[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11683.555 187.44 11683.835 188.44 ;
    END
  END SET_IBIAS[80]
  PIN SET_IBIAS[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11543.555 187.44 11543.835 188.44 ;
    END
  END SET_IBIAS[79]
  PIN SET_IBIAS[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11403.555 187.44 11403.835 188.44 ;
    END
  END SET_IBIAS[78]
  PIN SET_IBIAS[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11263.555 187.44 11263.835 188.44 ;
    END
  END SET_IBIAS[77]
  PIN SET_IBIAS[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11123.555 187.44 11123.835 188.44 ;
    END
  END SET_IBIAS[76]
  PIN SET_IBIAS[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10983.555 187.44 10983.835 188.44 ;
    END
  END SET_IBIAS[75]
  PIN SET_IBIAS[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10843.555 187.44 10843.835 188.44 ;
    END
  END SET_IBIAS[74]
  PIN SET_IBIAS[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10703.555 187.44 10703.835 188.44 ;
    END
  END SET_IBIAS[73]
  PIN SET_IBIAS[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10563.555 187.44 10563.835 188.44 ;
    END
  END SET_IBIAS[72]
  PIN SET_IBIAS[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10423.555 187.44 10423.835 188.44 ;
    END
  END SET_IBIAS[71]
  PIN SET_IBIAS[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10283.555 187.44 10283.835 188.44 ;
    END
  END SET_IBIAS[70]
  PIN SET_IBIAS[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10143.555 187.44 10143.835 188.44 ;
    END
  END SET_IBIAS[69]
  PIN SET_IBIAS[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10003.555 187.44 10003.835 188.44 ;
    END
  END SET_IBIAS[68]
  PIN SET_IBIAS[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9863.555 187.44 9863.835 188.44 ;
    END
  END SET_IBIAS[67]
  PIN SET_IBIAS[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9723.555 187.44 9723.835 188.44 ;
    END
  END SET_IBIAS[66]
  PIN SET_IBIAS[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9583.555 187.44 9583.835 188.44 ;
    END
  END SET_IBIAS[65]
  PIN SET_IBIAS[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9443.555 187.44 9443.835 188.44 ;
    END
  END SET_IBIAS[64]
  PIN SET_IBIAS[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9303.555 187.44 9303.835 188.44 ;
    END
  END SET_IBIAS[63]
  PIN SET_IBIAS[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9163.555 187.44 9163.835 188.44 ;
    END
  END SET_IBIAS[62]
  PIN SET_IBIAS[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9023.555 187.44 9023.835 188.44 ;
    END
  END SET_IBIAS[61]
  PIN SET_IBIAS[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8883.555 187.44 8883.835 188.44 ;
    END
  END SET_IBIAS[60]
  PIN SET_IBIAS[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8743.555 187.44 8743.835 188.44 ;
    END
  END SET_IBIAS[59]
  PIN SET_IBIAS[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8603.555 187.44 8603.835 188.44 ;
    END
  END SET_IBIAS[58]
  PIN SET_IBIAS[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8463.555 187.44 8463.835 188.44 ;
    END
  END SET_IBIAS[57]
  PIN SET_IBIAS[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8323.555 187.44 8323.835 188.44 ;
    END
  END SET_IBIAS[56]
  PIN SET_IBIAS[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8183.555 187.44 8183.835 188.44 ;
    END
  END SET_IBIAS[55]
  PIN SET_IBIAS[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8043.555 187.44 8043.835 188.44 ;
    END
  END SET_IBIAS[54]
  PIN SET_IBIAS[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7903.555 187.44 7903.835 188.44 ;
    END
  END SET_IBIAS[53]
  PIN SET_IBIAS[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7763.555 187.44 7763.835 188.44 ;
    END
  END SET_IBIAS[52]
  PIN SET_IBIAS[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7623.555 187.44 7623.835 188.44 ;
    END
  END SET_IBIAS[51]
  PIN SET_IBIAS[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7483.555 187.44 7483.835 188.44 ;
    END
  END SET_IBIAS[50]
  PIN SET_IBIAS[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7343.555 187.44 7343.835 188.44 ;
    END
  END SET_IBIAS[49]
  PIN SET_IBIAS[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7203.555 187.44 7203.835 188.44 ;
    END
  END SET_IBIAS[48]
  PIN SET_IBIAS[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7063.555 187.44 7063.835 188.44 ;
    END
  END SET_IBIAS[47]
  PIN SET_IBIAS[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6923.555 187.44 6923.835 188.44 ;
    END
  END SET_IBIAS[46]
  PIN SET_IBIAS[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6783.555 187.44 6783.835 188.44 ;
    END
  END SET_IBIAS[45]
  PIN SET_IBIAS[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6643.555 187.44 6643.835 188.44 ;
    END
  END SET_IBIAS[44]
  PIN SET_IBIAS[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6503.555 187.44 6503.835 188.44 ;
    END
  END SET_IBIAS[43]
  PIN SET_IBIAS[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6363.555 187.44 6363.835 188.44 ;
    END
  END SET_IBIAS[42]
  PIN SET_IBIAS[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6223.555 187.44 6223.835 188.44 ;
    END
  END SET_IBIAS[41]
  PIN SET_IBIAS[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6083.555 187.44 6083.835 188.44 ;
    END
  END SET_IBIAS[40]
  PIN SET_IBIAS[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5943.555 187.44 5943.835 188.44 ;
    END
  END SET_IBIAS[39]
  PIN SET_IBIAS[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5803.555 187.44 5803.835 188.44 ;
    END
  END SET_IBIAS[38]
  PIN SET_IBIAS[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5663.555 187.44 5663.835 188.44 ;
    END
  END SET_IBIAS[37]
  PIN SET_IBIAS[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5523.555 187.44 5523.835 188.44 ;
    END
  END SET_IBIAS[36]
  PIN SET_IBIAS[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5383.555 187.44 5383.835 188.44 ;
    END
  END SET_IBIAS[35]
  PIN SET_IBIAS[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5243.555 187.44 5243.835 188.44 ;
    END
  END SET_IBIAS[34]
  PIN SET_IBIAS[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5103.555 187.44 5103.835 188.44 ;
    END
  END SET_IBIAS[33]
  PIN SET_IBIAS[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4963.555 187.44 4963.835 188.44 ;
    END
  END SET_IBIAS[32]
  PIN SET_IBIAS[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4823.555 187.44 4823.835 188.44 ;
    END
  END SET_IBIAS[31]
  PIN SET_IBIAS[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4683.555 187.44 4683.835 188.44 ;
    END
  END SET_IBIAS[30]
  PIN SET_IBIAS[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4543.555 187.44 4543.835 188.44 ;
    END
  END SET_IBIAS[29]
  PIN SET_IBIAS[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4403.555 187.44 4403.835 188.44 ;
    END
  END SET_IBIAS[28]
  PIN SET_IBIAS[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4263.555 187.44 4263.835 188.44 ;
    END
  END SET_IBIAS[27]
  PIN SET_IBIAS[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4123.555 187.44 4123.835 188.44 ;
    END
  END SET_IBIAS[26]
  PIN SET_IBIAS[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3983.555 187.44 3983.835 188.44 ;
    END
  END SET_IBIAS[25]
  PIN SET_IBIAS[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3843.555 187.44 3843.835 188.44 ;
    END
  END SET_IBIAS[24]
  PIN SET_IBIAS[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3703.555 187.44 3703.835 188.44 ;
    END
  END SET_IBIAS[23]
  PIN SET_IBIAS[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3563.555 187.44 3563.835 188.44 ;
    END
  END SET_IBIAS[22]
  PIN SET_IBIAS[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3423.555 187.44 3423.835 188.44 ;
    END
  END SET_IBIAS[21]
  PIN SET_IBIAS[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3283.555 187.44 3283.835 188.44 ;
    END
  END SET_IBIAS[20]
  PIN SET_IBIAS[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3143.555 187.44 3143.835 188.44 ;
    END
  END SET_IBIAS[19]
  PIN SET_IBIAS[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3003.555 187.44 3003.835 188.44 ;
    END
  END SET_IBIAS[18]
  PIN SET_IBIAS[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2863.555 187.44 2863.835 188.44 ;
    END
  END SET_IBIAS[17]
  PIN SET_IBIAS[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2723.555 187.44 2723.835 188.44 ;
    END
  END SET_IBIAS[16]
  PIN SET_IBIAS[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2583.555 187.44 2583.835 188.44 ;
    END
  END SET_IBIAS[15]
  PIN SET_IBIAS[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2443.555 187.44 2443.835 188.44 ;
    END
  END SET_IBIAS[14]
  PIN SET_IBIAS[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2303.555 187.44 2303.835 188.44 ;
    END
  END SET_IBIAS[13]
  PIN SET_IBIAS[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2163.555 187.44 2163.835 188.44 ;
    END
  END SET_IBIAS[12]
  PIN SET_IBIAS[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2023.555 187.44 2023.835 188.44 ;
    END
  END SET_IBIAS[11]
  PIN SET_IBIAS[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1883.555 187.44 1883.835 188.44 ;
    END
  END SET_IBIAS[10]
  PIN SET_IBIAS[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1743.555 187.44 1743.835 188.44 ;
    END
  END SET_IBIAS[9]
  PIN SET_IBIAS[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1603.555 187.44 1603.835 188.44 ;
    END
  END SET_IBIAS[8]
  PIN SET_IBIAS[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1463.555 187.44 1463.835 188.44 ;
    END
  END SET_IBIAS[7]
  PIN SET_IBIAS[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1323.555 187.44 1323.835 188.44 ;
    END
  END SET_IBIAS[6]
  PIN SET_IBIAS[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1183.555 187.44 1183.835 188.44 ;
    END
  END SET_IBIAS[5]
  PIN SET_IBIAS[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1043.555 187.44 1043.835 188.44 ;
    END
  END SET_IBIAS[4]
  PIN SET_IBIAS[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 903.555 187.44 903.835 188.44 ;
    END
  END SET_IBIAS[3]
  PIN SET_IBIAS[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 763.555 187.44 763.835 188.44 ;
    END
  END SET_IBIAS[2]
  PIN SET_IBIAS[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 623.555 187.44 623.835 188.44 ;
    END
  END SET_IBIAS[1]
  PIN SET_IBIAS[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 483.555 187.44 483.835 188.44 ;
    END
  END SET_IBIAS[0]
  PIN GNDA_VDAC
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 326.66 309.245 327.66 323.275 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 326.66 196.245 327.66 210.275 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 309.245 18490.46 323.275 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 18489.46 196.245 18490.46 210.275 ;
    END
  END GNDA_VDAC
  PIN SET_IRESET_BIT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9431.635 187.44 9432.195 188.295 ;
    END
  END SET_IRESET_BIT
  PIN VCASN_DAC_MON_L
    DIRECTION OUTPUT ;
    USE ANALOG ;
    PORT
      LAYER M4 ;
        RECT 326.66 8399.58 327.66 8401 ;
    END
  END VCASN_DAC_MON_L
  PIN VCASN_MON_R
    DIRECTION OUTPUT ;
    USE ANALOG ;
    PORT
      LAYER M4 ;
        RECT 18489.46 8438.095 18490.46 8439.515 ;
    END
  END VCASN_MON_R
  PIN VCASN_DAC_MON_R
    DIRECTION OUTPUT ;
    USE ANALOG ;
    PORT
      LAYER M4 ;
        RECT 18489.46 8399.58 18490.46 8401 ;
    END
  END VCASN_DAC_MON_R
  PIN DACMON_VCASN_DAC
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER M5 ;
        RECT 18489.46 259.99 18490.46 261.19 ;
    END
  END DACMON_VCASN_DAC
  PIN GNDP
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 474.56 187.44 502.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 554.56 187.44 582.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 634.56 187.44 662.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 714.56 187.44 742.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 794.56 187.44 822.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 874.56 187.44 902.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 954.56 187.44 982.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1034.56 187.44 1062.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1114.56 187.44 1142.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1194.56 187.44 1222.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1274.56 187.44 1302.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1354.56 187.44 1382.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1434.56 187.44 1462.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1514.56 187.44 1542.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1594.56 187.44 1622.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1674.56 187.44 1702.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1754.56 187.44 1782.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1834.56 187.44 1862.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1914.56 187.44 1942.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1994.56 187.44 2022.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2074.56 187.44 2102.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2154.56 187.44 2182.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2234.56 187.44 2262.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2314.56 187.44 2342.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2394.56 187.44 2422.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2474.56 187.44 2502.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2554.56 187.44 2582.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2634.56 187.44 2662.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2714.56 187.44 2742.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2794.56 187.44 2822.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2874.56 187.44 2902.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2954.56 187.44 2982.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3034.56 187.44 3062.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3114.56 187.44 3142.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3194.56 187.44 3222.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3274.56 187.44 3302.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3354.56 187.44 3382.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3434.56 187.44 3462.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3514.56 187.44 3542.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3594.56 187.44 3622.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3674.56 187.44 3702.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3754.56 187.44 3782.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3834.56 187.44 3862.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3914.56 187.44 3942.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3994.56 187.44 4022.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4074.56 187.44 4102.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4154.56 187.44 4182.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4234.56 187.44 4262.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4314.56 187.44 4342.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4394.56 187.44 4422.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4474.56 187.44 4502.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4554.56 187.44 4582.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4634.56 187.44 4662.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4714.56 187.44 4742.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4794.56 187.44 4822.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4874.56 187.44 4902.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4954.56 187.44 4982.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5034.56 187.44 5062.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5114.56 187.44 5142.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5194.56 187.44 5222.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5274.56 187.44 5302.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5354.56 187.44 5382.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5434.56 187.44 5462.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5514.56 187.44 5542.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5594.56 187.44 5622.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5674.56 187.44 5702.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5754.56 187.44 5782.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5834.56 187.44 5862.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5914.56 187.44 5942.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5994.56 187.44 6022.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6074.56 187.44 6102.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6154.56 187.44 6182.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6234.56 187.44 6262.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6314.56 187.44 6342.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6394.56 187.44 6422.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6474.56 187.44 6502.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6554.56 187.44 6582.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6634.56 187.44 6662.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6714.56 187.44 6742.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6794.56 187.44 6822.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6874.56 187.44 6902.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6954.56 187.44 6982.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7034.56 187.44 7062.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7114.56 187.44 7142.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7194.56 187.44 7222.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7274.56 187.44 7302.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7354.56 187.44 7382.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7434.56 187.44 7462.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7514.56 187.44 7542.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7594.56 187.44 7622.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7674.56 187.44 7702.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7754.56 187.44 7782.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7834.56 187.44 7862.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7914.56 187.44 7942.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7994.56 187.44 8022.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8074.56 187.44 8102.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8154.56 187.44 8182.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8234.56 187.44 8262.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8314.56 187.44 8342.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8394.56 187.44 8422.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8474.56 187.44 8502.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8554.56 187.44 8582.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8634.56 187.44 8662.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8714.56 187.44 8742.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8794.56 187.44 8822.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8874.56 187.44 8902.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8954.56 187.44 8982.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9034.56 187.44 9062.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9114.56 187.44 9142.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9194.56 187.44 9222.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9274.56 187.44 9302.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9354.56 187.44 9382.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9434.56 187.44 9462.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9514.56 187.44 9542.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9594.56 187.44 9622.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9674.56 187.44 9702.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9754.56 187.44 9782.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9834.56 187.44 9862.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9914.56 187.44 9942.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9994.56 187.44 10022.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10074.56 187.44 10102.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10154.56 187.44 10182.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10234.56 187.44 10262.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10314.56 187.44 10342.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10394.56 187.44 10422.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10474.56 187.44 10502.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10554.56 187.44 10582.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10634.56 187.44 10662.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10714.56 187.44 10742.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10794.56 187.44 10822.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10874.56 187.44 10902.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10954.56 187.44 10982.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11034.56 187.44 11062.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11114.56 187.44 11142.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11194.56 187.44 11222.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11274.56 187.44 11302.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11354.56 187.44 11382.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11434.56 187.44 11462.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11514.56 187.44 11542.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11594.56 187.44 11622.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11674.56 187.44 11702.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11754.56 187.44 11782.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11834.56 187.44 11862.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11914.56 187.44 11942.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11994.56 187.44 12022.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12074.56 187.44 12102.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12154.56 187.44 12182.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12234.56 187.44 12262.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12314.56 187.44 12342.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12394.56 187.44 12422.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12474.56 187.44 12502.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12554.56 187.44 12582.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12634.56 187.44 12662.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12714.56 187.44 12742.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12794.56 187.44 12822.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12874.56 187.44 12902.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12954.56 187.44 12982.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13034.56 187.44 13062.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13114.56 187.44 13142.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13194.56 187.44 13222.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13274.56 187.44 13302.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13354.56 187.44 13382.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13434.56 187.44 13462.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13514.56 187.44 13542.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13594.56 187.44 13622.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13674.56 187.44 13702.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13754.56 187.44 13782.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13834.56 187.44 13862.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13914.56 187.44 13942.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13994.56 187.44 14022.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14074.56 187.44 14102.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14154.56 187.44 14182.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14234.56 187.44 14262.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14314.56 187.44 14342.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14394.56 187.44 14422.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14474.56 187.44 14502.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14554.56 187.44 14582.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14634.56 187.44 14662.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14714.56 187.44 14742.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14794.56 187.44 14822.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14874.56 187.44 14902.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14954.56 187.44 14982.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15034.56 187.44 15062.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15114.56 187.44 15142.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15194.56 187.44 15222.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15274.56 187.44 15302.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15354.56 187.44 15382.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15434.56 187.44 15462.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15514.56 187.44 15542.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15594.56 187.44 15622.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15674.56 187.44 15702.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15754.56 187.44 15782.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15834.56 187.44 15862.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15914.56 187.44 15942.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15994.56 187.44 16022.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16074.56 187.44 16102.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16154.56 187.44 16182.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16234.56 187.44 16262.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16314.56 187.44 16342.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16394.56 187.44 16422.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16474.56 187.44 16502.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16554.56 187.44 16582.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16634.56 187.44 16662.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16714.56 187.44 16742.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16794.56 187.44 16822.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16874.56 187.44 16902.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16954.56 187.44 16982.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17034.56 187.44 17062.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17114.56 187.44 17142.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17194.56 187.44 17222.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17274.56 187.44 17302.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17354.56 187.44 17382.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17434.56 187.44 17462.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17514.56 187.44 17542.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17594.56 187.44 17622.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17674.56 187.44 17702.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17754.56 187.44 17782.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17834.56 187.44 17862.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17914.56 187.44 17942.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17994.56 187.44 18022.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 18074.56 187.44 18102.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 18154.56 187.44 18182.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 18234.56 187.44 18262.56 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 18314.56 187.44 18342.56 188.44 ;
    END
  END GNDP
  PIN VPC
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 18489.46 505.445 18490.46 506.445 ;
    END
  END VPC
  PIN VPCNOSF
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 326.66 500.265 327.66 510.265 ;
    END
  END VPCNOSF
  PIN VDDP
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 459.04 187.44 472.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 505.08 187.44 518.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 522.06 187.44 535.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 539.04 187.44 552.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 585.08 187.44 598.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 602.06 187.44 615.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 619.04 187.44 632.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 665.08 187.44 678.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 682.06 187.44 695.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 699.04 187.44 712.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 745.08 187.44 758.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 762.06 187.44 775.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 779.04 187.44 792.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 825.08 187.44 838.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 842.06 187.44 855.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 859.04 187.44 872.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 905.08 187.44 918.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 922.06 187.44 935.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 939.04 187.44 952.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 985.08 187.44 998.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1002.06 187.44 1015.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1019.04 187.44 1032.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1065.08 187.44 1078.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1082.06 187.44 1095.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1099.04 187.44 1112.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1145.08 187.44 1158.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1162.06 187.44 1175.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1179.04 187.44 1192.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1225.08 187.44 1238.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1242.06 187.44 1255.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1259.04 187.44 1272.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1305.08 187.44 1318.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1322.06 187.44 1335.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1339.04 187.44 1352.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1385.08 187.44 1398.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1402.06 187.44 1415.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1419.04 187.44 1432.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1465.08 187.44 1478.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1482.06 187.44 1495.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1499.04 187.44 1512.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1545.08 187.44 1558.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1562.06 187.44 1575.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1579.04 187.44 1592.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1625.08 187.44 1638.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1642.06 187.44 1655.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1659.04 187.44 1672.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1705.08 187.44 1718.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1722.06 187.44 1735.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1739.04 187.44 1752.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1785.08 187.44 1798.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1802.06 187.44 1815.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1819.04 187.44 1832.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1865.08 187.44 1878.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1882.06 187.44 1895.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1899.04 187.44 1912.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1945.08 187.44 1958.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1962.06 187.44 1975.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 1979.04 187.44 1992.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2025.08 187.44 2038.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2042.06 187.44 2055.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2059.04 187.44 2072.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2105.08 187.44 2118.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2122.06 187.44 2135.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2139.04 187.44 2152.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2185.08 187.44 2198.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2202.06 187.44 2215.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2219.04 187.44 2232.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2265.08 187.44 2278.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2282.06 187.44 2295.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2299.04 187.44 2312.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2345.08 187.44 2358.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2362.06 187.44 2375.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2379.04 187.44 2392.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2425.08 187.44 2438.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2442.06 187.44 2455.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2459.04 187.44 2472.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2505.08 187.44 2518.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2522.06 187.44 2535.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2539.04 187.44 2552.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2585.08 187.44 2598.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2602.06 187.44 2615.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2619.04 187.44 2632.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2665.08 187.44 2678.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2682.06 187.44 2695.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2699.04 187.44 2712.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2745.08 187.44 2758.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2762.06 187.44 2775.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2779.04 187.44 2792.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2825.08 187.44 2838.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2842.06 187.44 2855.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2859.04 187.44 2872.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2905.08 187.44 2918.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2922.06 187.44 2935.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2939.04 187.44 2952.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 2985.08 187.44 2998.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3002.06 187.44 3015.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3019.04 187.44 3032.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3065.08 187.44 3078.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3082.06 187.44 3095.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3099.04 187.44 3112.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3145.08 187.44 3158.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3162.06 187.44 3175.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3179.04 187.44 3192.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3225.08 187.44 3238.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3242.06 187.44 3255.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3259.04 187.44 3272.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3305.08 187.44 3318.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3322.06 187.44 3335.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3339.04 187.44 3352.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3385.08 187.44 3398.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3402.06 187.44 3415.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3419.04 187.44 3432.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3465.08 187.44 3478.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3482.06 187.44 3495.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3499.04 187.44 3512.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3545.08 187.44 3558.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3562.06 187.44 3575.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3579.04 187.44 3592.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3625.08 187.44 3638.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3642.06 187.44 3655.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3659.04 187.44 3672.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3705.08 187.44 3718.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3722.06 187.44 3735.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3739.04 187.44 3752.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3785.08 187.44 3798.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3802.06 187.44 3815.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3819.04 187.44 3832.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3865.08 187.44 3878.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3882.06 187.44 3895.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3899.04 187.44 3912.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3945.08 187.44 3958.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3962.06 187.44 3975.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 3979.04 187.44 3992.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4025.08 187.44 4038.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4042.06 187.44 4055.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4059.04 187.44 4072.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4105.08 187.44 4118.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4122.06 187.44 4135.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4139.04 187.44 4152.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4185.08 187.44 4198.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4202.06 187.44 4215.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4219.04 187.44 4232.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4265.08 187.44 4278.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4282.06 187.44 4295.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4299.04 187.44 4312.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4345.08 187.44 4358.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4362.06 187.44 4375.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4379.04 187.44 4392.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4425.08 187.44 4438.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4442.06 187.44 4455.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4459.04 187.44 4472.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4505.08 187.44 4518.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4522.06 187.44 4535.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4539.04 187.44 4552.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4585.08 187.44 4598.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4602.06 187.44 4615.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4619.04 187.44 4632.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4665.08 187.44 4678.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4682.06 187.44 4695.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4699.04 187.44 4712.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4745.08 187.44 4758.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4762.06 187.44 4775.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4779.04 187.44 4792.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4825.08 187.44 4838.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4842.06 187.44 4855.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4859.04 187.44 4872.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4905.08 187.44 4918.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4922.06 187.44 4935.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4939.04 187.44 4952.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 4985.08 187.44 4998.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5002.06 187.44 5015.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5019.04 187.44 5032.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5065.08 187.44 5078.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5082.06 187.44 5095.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5099.04 187.44 5112.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5145.08 187.44 5158.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5162.06 187.44 5175.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5179.04 187.44 5192.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5225.08 187.44 5238.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5242.06 187.44 5255.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5259.04 187.44 5272.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5305.08 187.44 5318.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5322.06 187.44 5335.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5339.04 187.44 5352.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5385.08 187.44 5398.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5402.06 187.44 5415.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5419.04 187.44 5432.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5465.08 187.44 5478.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5482.06 187.44 5495.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5499.04 187.44 5512.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5545.08 187.44 5558.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5562.06 187.44 5575.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5579.04 187.44 5592.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5625.08 187.44 5638.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5642.06 187.44 5655.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5659.04 187.44 5672.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5705.08 187.44 5718.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5722.06 187.44 5735.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5739.04 187.44 5752.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5785.08 187.44 5798.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5802.06 187.44 5815.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5819.04 187.44 5832.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5865.08 187.44 5878.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5882.06 187.44 5895.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5899.04 187.44 5912.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5945.08 187.44 5958.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5962.06 187.44 5975.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 5979.04 187.44 5992.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6025.08 187.44 6038.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6042.06 187.44 6055.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6059.04 187.44 6072.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6105.08 187.44 6118.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6122.06 187.44 6135.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6139.04 187.44 6152.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6185.08 187.44 6198.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6202.06 187.44 6215.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6219.04 187.44 6232.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6265.08 187.44 6278.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6282.06 187.44 6295.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6299.04 187.44 6312.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6345.08 187.44 6358.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6362.06 187.44 6375.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6379.04 187.44 6392.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6425.08 187.44 6438.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6442.06 187.44 6455.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6459.04 187.44 6472.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6505.08 187.44 6518.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6522.06 187.44 6535.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6539.04 187.44 6552.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6585.08 187.44 6598.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6602.06 187.44 6615.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6619.04 187.44 6632.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6665.08 187.44 6678.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6682.06 187.44 6695.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6699.04 187.44 6712.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6745.08 187.44 6758.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6762.06 187.44 6775.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6779.04 187.44 6792.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6825.08 187.44 6838.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6842.06 187.44 6855.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6859.04 187.44 6872.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6905.08 187.44 6918.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6922.06 187.44 6935.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6939.04 187.44 6952.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 6985.08 187.44 6998.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7002.06 187.44 7015.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7019.04 187.44 7032.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7065.08 187.44 7078.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7082.06 187.44 7095.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7099.04 187.44 7112.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7145.08 187.44 7158.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7162.06 187.44 7175.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7179.04 187.44 7192.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7225.08 187.44 7238.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7242.06 187.44 7255.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7259.04 187.44 7272.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7305.08 187.44 7318.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7322.06 187.44 7335.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7339.04 187.44 7352.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7385.08 187.44 7398.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7402.06 187.44 7415.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7419.04 187.44 7432.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7465.08 187.44 7478.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7482.06 187.44 7495.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7499.04 187.44 7512.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7545.08 187.44 7558.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7562.06 187.44 7575.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7579.04 187.44 7592.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7625.08 187.44 7638.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7642.06 187.44 7655.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7659.04 187.44 7672.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7705.08 187.44 7718.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7722.06 187.44 7735.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7739.04 187.44 7752.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7785.08 187.44 7798.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7802.06 187.44 7815.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7819.04 187.44 7832.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7865.08 187.44 7878.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7882.06 187.44 7895.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7899.04 187.44 7912.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7945.08 187.44 7958.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7962.06 187.44 7975.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 7979.04 187.44 7992.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8025.08 187.44 8038.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8042.06 187.44 8055.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8059.04 187.44 8072.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8105.08 187.44 8118.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8122.06 187.44 8135.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8139.04 187.44 8152.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8185.08 187.44 8198.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8202.06 187.44 8215.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8219.04 187.44 8232.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8265.08 187.44 8278.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8282.06 187.44 8295.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8299.04 187.44 8312.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8345.08 187.44 8358.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8362.06 187.44 8375.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8379.04 187.44 8392.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8425.08 187.44 8438.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8442.06 187.44 8455.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8459.04 187.44 8472.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8505.08 187.44 8518.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8522.06 187.44 8535.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8539.04 187.44 8552.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8585.08 187.44 8598.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8602.06 187.44 8615.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8619.04 187.44 8632.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8665.08 187.44 8678.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8682.06 187.44 8695.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8699.04 187.44 8712.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8745.08 187.44 8758.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8762.06 187.44 8775.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8779.04 187.44 8792.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8825.08 187.44 8838.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8842.06 187.44 8855.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8859.04 187.44 8872.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8905.08 187.44 8918.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8922.06 187.44 8935.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8939.04 187.44 8952.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 8985.08 187.44 8998.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9002.06 187.44 9015.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9019.04 187.44 9032.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9065.08 187.44 9078.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9082.06 187.44 9095.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9099.04 187.44 9112.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9145.08 187.44 9158.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9162.06 187.44 9175.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9179.04 187.44 9192.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9225.08 187.44 9238.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9242.06 187.44 9255.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9259.04 187.44 9272.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9305.08 187.44 9318.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9322.06 187.44 9335.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9339.04 187.44 9352.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9385.08 187.44 9398.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9402.06 187.44 9415.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9419.04 187.44 9432.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9465.08 187.44 9478.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9482.06 187.44 9495.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9499.04 187.44 9512.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9545.08 187.44 9558.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9562.06 187.44 9575.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9579.04 187.44 9592.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9625.08 187.44 9638.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9642.06 187.44 9655.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9659.04 187.44 9672.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9705.08 187.44 9718.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9722.06 187.44 9735.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9739.04 187.44 9752.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9785.08 187.44 9798.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9802.06 187.44 9815.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9819.04 187.44 9832.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9865.08 187.44 9878.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9882.06 187.44 9895.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9899.04 187.44 9912.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9945.08 187.44 9958.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9962.06 187.44 9975.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 9979.04 187.44 9992.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10025.08 187.44 10038.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10042.06 187.44 10055.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10059.04 187.44 10072.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10105.08 187.44 10118.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10122.06 187.44 10135.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10139.04 187.44 10152.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10185.08 187.44 10198.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10202.06 187.44 10215.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10219.04 187.44 10232.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10265.08 187.44 10278.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10282.06 187.44 10295.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10299.04 187.44 10312.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10345.08 187.44 10358.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10362.06 187.44 10375.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10379.04 187.44 10392.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10425.08 187.44 10438.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10442.06 187.44 10455.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10459.04 187.44 10472.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10505.08 187.44 10518.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10522.06 187.44 10535.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10539.04 187.44 10552.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10585.08 187.44 10598.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10602.06 187.44 10615.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10619.04 187.44 10632.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10665.08 187.44 10678.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10682.06 187.44 10695.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10699.04 187.44 10712.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10745.08 187.44 10758.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10762.06 187.44 10775.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10779.04 187.44 10792.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10825.08 187.44 10838.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10842.06 187.44 10855.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10859.04 187.44 10872.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10905.08 187.44 10918.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10922.06 187.44 10935.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10939.04 187.44 10952.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 10985.08 187.44 10998.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11002.06 187.44 11015.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11019.04 187.44 11032.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11065.08 187.44 11078.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11082.06 187.44 11095.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11099.04 187.44 11112.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11145.08 187.44 11158.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11162.06 187.44 11175.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11179.04 187.44 11192.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11225.08 187.44 11238.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11242.06 187.44 11255.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11259.04 187.44 11272.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11305.08 187.44 11318.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11322.06 187.44 11335.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11339.04 187.44 11352.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11385.08 187.44 11398.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11402.06 187.44 11415.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11419.04 187.44 11432.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11465.08 187.44 11478.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11482.06 187.44 11495.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11499.04 187.44 11512.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11545.08 187.44 11558.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11562.06 187.44 11575.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11579.04 187.44 11592.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11625.08 187.44 11638.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11642.06 187.44 11655.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11659.04 187.44 11672.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11705.08 187.44 11718.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11722.06 187.44 11735.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11739.04 187.44 11752.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11785.08 187.44 11798.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11802.06 187.44 11815.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11819.04 187.44 11832.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11865.08 187.44 11878.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11882.06 187.44 11895.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11899.04 187.44 11912.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11945.08 187.44 11958.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11962.06 187.44 11975.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 11979.04 187.44 11992.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12025.08 187.44 12038.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12042.06 187.44 12055.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12059.04 187.44 12072.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12105.08 187.44 12118.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12122.06 187.44 12135.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12139.04 187.44 12152.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12185.08 187.44 12198.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12202.06 187.44 12215.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12219.04 187.44 12232.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12265.08 187.44 12278.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12282.06 187.44 12295.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12299.04 187.44 12312.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12345.08 187.44 12358.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12362.06 187.44 12375.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12379.04 187.44 12392.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12425.08 187.44 12438.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12442.06 187.44 12455.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12459.04 187.44 12472.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12505.08 187.44 12518.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12522.06 187.44 12535.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12539.04 187.44 12552.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12585.08 187.44 12598.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12602.06 187.44 12615.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12619.04 187.44 12632.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12665.08 187.44 12678.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12682.06 187.44 12695.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12699.04 187.44 12712.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12745.08 187.44 12758.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12762.06 187.44 12775.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12779.04 187.44 12792.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12825.08 187.44 12838.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12842.06 187.44 12855.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12859.04 187.44 12872.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12905.08 187.44 12918.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12922.06 187.44 12935.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12939.04 187.44 12952.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 12985.08 187.44 12998.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13002.06 187.44 13015.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13019.04 187.44 13032.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13065.08 187.44 13078.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13082.06 187.44 13095.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13099.04 187.44 13112.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13145.08 187.44 13158.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13162.06 187.44 13175.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13179.04 187.44 13192.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13225.08 187.44 13238.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13242.06 187.44 13255.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13259.04 187.44 13272.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13305.08 187.44 13318.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13322.06 187.44 13335.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13339.04 187.44 13352.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13385.08 187.44 13398.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13402.06 187.44 13415.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13419.04 187.44 13432.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13465.08 187.44 13478.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13482.06 187.44 13495.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13499.04 187.44 13512.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13545.08 187.44 13558.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13562.06 187.44 13575.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13579.04 187.44 13592.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13625.08 187.44 13638.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13642.06 187.44 13655.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13659.04 187.44 13672.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13705.08 187.44 13718.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13722.06 187.44 13735.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13739.04 187.44 13752.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13785.08 187.44 13798.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13802.06 187.44 13815.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13819.04 187.44 13832.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13865.08 187.44 13878.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13882.06 187.44 13895.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13899.04 187.44 13912.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13945.08 187.44 13958.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13962.06 187.44 13975.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 13979.04 187.44 13992.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14025.08 187.44 14038.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14042.06 187.44 14055.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14059.04 187.44 14072.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14105.08 187.44 14118.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14122.06 187.44 14135.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14139.04 187.44 14152.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14185.08 187.44 14198.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14202.06 187.44 14215.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14219.04 187.44 14232.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14265.08 187.44 14278.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14282.06 187.44 14295.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14299.04 187.44 14312.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14345.08 187.44 14358.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14362.06 187.44 14375.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14379.04 187.44 14392.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14425.08 187.44 14438.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14442.06 187.44 14455.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14459.04 187.44 14472.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14505.08 187.44 14518.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14522.06 187.44 14535.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14539.04 187.44 14552.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14585.08 187.44 14598.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14602.06 187.44 14615.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14619.04 187.44 14632.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14665.08 187.44 14678.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14682.06 187.44 14695.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14699.04 187.44 14712.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14745.08 187.44 14758.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14762.06 187.44 14775.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14779.04 187.44 14792.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14825.08 187.44 14838.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14842.06 187.44 14855.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14859.04 187.44 14872.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14905.08 187.44 14918.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14922.06 187.44 14935.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14939.04 187.44 14952.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 14985.08 187.44 14998.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15002.06 187.44 15015.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15019.04 187.44 15032.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15065.08 187.44 15078.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15082.06 187.44 15095.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15099.04 187.44 15112.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15145.08 187.44 15158.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15162.06 187.44 15175.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15179.04 187.44 15192.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15225.08 187.44 15238.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15242.06 187.44 15255.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15259.04 187.44 15272.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15305.08 187.44 15318.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15322.06 187.44 15335.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15339.04 187.44 15352.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15385.08 187.44 15398.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15402.06 187.44 15415.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15419.04 187.44 15432.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15465.08 187.44 15478.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15482.06 187.44 15495.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15499.04 187.44 15512.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15545.08 187.44 15558.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15562.06 187.44 15575.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15579.04 187.44 15592.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15625.08 187.44 15638.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15642.06 187.44 15655.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15659.04 187.44 15672.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15705.08 187.44 15718.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15722.06 187.44 15735.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15739.04 187.44 15752.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15785.08 187.44 15798.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15802.06 187.44 15815.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15819.04 187.44 15832.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15865.08 187.44 15878.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15882.06 187.44 15895.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15899.04 187.44 15912.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15945.08 187.44 15958.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15962.06 187.44 15975.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 15979.04 187.44 15992.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16025.08 187.44 16038.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16042.06 187.44 16055.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16059.04 187.44 16072.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16105.08 187.44 16118.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16122.06 187.44 16135.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16139.04 187.44 16152.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16185.08 187.44 16198.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16202.06 187.44 16215.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16219.04 187.44 16232.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16265.08 187.44 16278.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16282.06 187.44 16295.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16299.04 187.44 16312.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16345.08 187.44 16358.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16362.06 187.44 16375.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16379.04 187.44 16392.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16425.08 187.44 16438.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16442.06 187.44 16455.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16459.04 187.44 16472.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16505.08 187.44 16518.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16522.06 187.44 16535.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16539.04 187.44 16552.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16585.08 187.44 16598.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16602.06 187.44 16615.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16619.04 187.44 16632.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16665.08 187.44 16678.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16682.06 187.44 16695.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16699.04 187.44 16712.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16745.08 187.44 16758.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16762.06 187.44 16775.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16779.04 187.44 16792.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16825.08 187.44 16838.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16842.06 187.44 16855.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16859.04 187.44 16872.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16905.08 187.44 16918.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16922.06 187.44 16935.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16939.04 187.44 16952.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 16985.08 187.44 16998.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17002.06 187.44 17015.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17019.04 187.44 17032.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17065.08 187.44 17078.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17082.06 187.44 17095.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17099.04 187.44 17112.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17145.08 187.44 17158.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17162.06 187.44 17175.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17179.04 187.44 17192.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17225.08 187.44 17238.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17242.06 187.44 17255.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17259.04 187.44 17272.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17305.08 187.44 17318.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17322.06 187.44 17335.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17339.04 187.44 17352.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17385.08 187.44 17398.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17402.06 187.44 17415.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17419.04 187.44 17432.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17465.08 187.44 17478.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17482.06 187.44 17495.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17499.04 187.44 17512.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17545.08 187.44 17558.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17562.06 187.44 17575.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17579.04 187.44 17592.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17625.08 187.44 17638.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17642.06 187.44 17655.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17659.04 187.44 17672.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17705.08 187.44 17718.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17722.06 187.44 17735.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17739.04 187.44 17752.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17785.08 187.44 17798.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17802.06 187.44 17815.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17819.04 187.44 17832.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17865.08 187.44 17878.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17882.06 187.44 17895.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17899.04 187.44 17912.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17945.08 187.44 17958.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17962.06 187.44 17975.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 17979.04 187.44 17992.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 18025.08 187.44 18038.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 18042.06 187.44 18055.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 18059.04 187.44 18072.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 18105.08 187.44 18118.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 18122.06 187.44 18135.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 18139.04 187.44 18152.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 18185.08 187.44 18198.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 18202.06 187.44 18215.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 18219.04 187.44 18232.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 18265.08 187.44 18278.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 18282.06 187.44 18295.06 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 18299.04 187.44 18312.04 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 18345.08 187.44 18358.08 188.44 ;
    END
    PORT
      LAYER M5 ;
        RECT 18362.06 187.44 18375.06 188.44 ;
    END
  END VDDP
  PIN SET_IBUFN_L[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 332.405 187.44 332.685 188.44 ;
    END
  END SET_IBUFN_L[3]
  PIN SET_IBUFN_L[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 332.965 187.44 333.245 188.44 ;
    END
  END SET_IBUFN_L[2]
  PIN SET_IBUFN_L[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 333.525 187.44 333.805 188.44 ;
    END
  END SET_IBUFN_L[1]
  PIN SET_IBUFN_L[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 334.085 187.44 334.365 188.44 ;
    END
  END SET_IBUFN_L[0]
  PIN SET_IBUFP_L[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 334.645 187.44 334.925 188.44 ;
    END
  END SET_IBUFP_L[3]
  PIN SET_IBUFP_L[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 335.205 187.44 335.485 188.44 ;
    END
  END SET_IBUFP_L[2]
  PIN SET_IBUFP_L[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 335.765 187.44 336.045 188.44 ;
    END
  END SET_IBUFP_L[1]
  PIN SET_IBUFP_L[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 336.325 187.44 336.605 188.44 ;
    END
  END SET_IBUFP_L[0]
  PIN SET_IBUFP_R[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18480.515 187.44 18480.795 188.44 ;
    END
  END SET_IBUFP_R[0]
  PIN SET_IBUFP_R[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18481.075 187.44 18481.355 188.44 ;
    END
  END SET_IBUFP_R[1]
  PIN SET_IBUFP_R[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18481.635 187.44 18481.915 188.44 ;
    END
  END SET_IBUFP_R[2]
  PIN SET_IBUFP_R[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18482.195 187.44 18482.475 188.44 ;
    END
  END SET_IBUFP_R[3]
  PIN SET_IBUFN_R[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18482.755 187.44 18483.035 188.44 ;
    END
  END SET_IBUFN_R[0]
  PIN SET_IBUFN_R[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18483.315 187.44 18483.595 188.44 ;
    END
  END SET_IBUFN_R[1]
  PIN SET_IBUFN_R[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18483.875 187.44 18484.155 188.44 ;
    END
  END SET_IBUFN_R[2]
  PIN SET_IBUFN_R[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18484.435 187.44 18484.715 188.44 ;
    END
  END SET_IBUFN_R[3]
  PIN BcidMtx[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 973.065 187.44 973.345 188.44 ;
    END
  END BcidMtx[39]
  PIN BcidMtx[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 970.265 187.44 970.545 188.44 ;
    END
  END BcidMtx[36]
  PIN BcidMtx[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 894.665 187.44 894.945 188.44 ;
    END
  END BcidMtx[32]
  PIN BcidMtx[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 827.465 187.44 827.745 188.44 ;
    END
  END BcidMtx[29]
  PIN BcidMtx[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 824.105 187.44 824.385 188.44 ;
    END
  END BcidMtx[25]
  PIN BcidMtx[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 748.785 187.44 749.065 188.44 ;
    END
  END BcidMtx[23]
  PIN BcidMtx[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 720.505 187.44 720.785 188.44 ;
    END
  END BcidMtx[20]
  PIN BcidMtx[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 719.385 187.44 719.665 188.44 ;
    END
  END BcidMtx[18]
  PIN BcidMtx[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 640.425 187.44 640.705 188.44 ;
    END
  END BcidMtx[15]
  PIN BcidMtx[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 575.465 187.44 575.745 188.44 ;
    END
  END BcidMtx[10]
  PIN BcidMtx[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 572.665 187.44 572.945 188.44 ;
    END
  END BcidMtx[7]
  PIN BcidMtx[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1533.625 187.44 1533.905 188.44 ;
    END
  END BcidMtx[82]
  PIN BcidMtx[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1531.385 187.44 1531.665 188.44 ;
    END
  END BcidMtx[80]
  PIN BcidMtx[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1530.265 187.44 1530.545 188.44 ;
    END
  END BcidMtx[78]
  PIN BcidMtx[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1456.905 187.44 1457.185 188.44 ;
    END
  END BcidMtx[76]
  PIN BcidMtx[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1454.105 187.44 1454.385 188.44 ;
    END
  END BcidMtx[73]
  PIN BcidMtx[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1453.545 187.44 1453.825 188.44 ;
    END
  END BcidMtx[72]
  PIN BcidMtx[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1386.345 187.44 1386.625 188.44 ;
    END
  END BcidMtx[69]
  PIN BcidMtx[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1383.545 187.44 1383.825 188.44 ;
    END
  END BcidMtx[66]
  PIN BcidMtx[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1308.225 187.44 1308.505 188.44 ;
    END
  END BcidMtx[64]
  PIN BcidMtx[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1280.505 187.44 1280.785 188.44 ;
    END
  END BcidMtx[62]
  PIN BcidMtx[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1201.545 187.44 1201.825 188.44 ;
    END
  END BcidMtx[59]
  PIN BcidMtx[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1136.025 187.44 1136.305 188.44 ;
    END
  END BcidMtx[53]
  PIN BcidMtx[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1133.225 187.44 1133.505 188.44 ;
    END
  END BcidMtx[50]
  PIN BcidMtx[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1132.105 187.44 1132.385 188.44 ;
    END
  END BcidMtx[48]
  PIN BcidMtx[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1052.585 187.44 1052.865 188.44 ;
    END
  END BcidMtx[45]
  PIN BcidMtx[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1050.905 187.44 1051.185 188.44 ;
    END
  END BcidMtx[44]
  PIN BcidMtx[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2093.065 187.44 2093.345 188.44 ;
    END
  END BcidMtx[123]
  PIN BcidMtx[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2091.385 187.44 2091.665 188.44 ;
    END
  END BcidMtx[122]
  PIN BcidMtx[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2017.465 187.44 2017.745 188.44 ;
    END
  END BcidMtx[119]
  PIN BcidMtx[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2014.105 187.44 2014.385 188.44 ;
    END
  END BcidMtx[115]
  PIN BcidMtx[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1947.465 187.44 1947.745 188.44 ;
    END
  END BcidMtx[113]
  PIN BcidMtx[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1946.345 187.44 1946.625 188.44 ;
    END
  END BcidMtx[111]
  PIN BcidMtx[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1943.545 187.44 1943.825 188.44 ;
    END
  END BcidMtx[108]
  PIN BcidMtx[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1868.225 187.44 1868.505 188.44 ;
    END
  END BcidMtx[106]
  PIN BcidMtx[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1760.425 187.44 1760.705 188.44 ;
    END
  END BcidMtx[99]
  PIN BcidMtx[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1758.745 187.44 1759.025 188.44 ;
    END
  END BcidMtx[98]
  PIN BcidMtx[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1696.025 187.44 1696.305 188.44 ;
    END
  END BcidMtx[95]
  PIN BcidMtx[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1692.105 187.44 1692.385 188.44 ;
    END
  END BcidMtx[90]
  PIN BcidMtx[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1613.705 187.44 1613.985 188.44 ;
    END
  END BcidMtx[89]
  PIN BcidMtx[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1610.345 187.44 1610.625 188.44 ;
    END
  END BcidMtx[85]
  PIN BcidMtx[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2653.625 187.44 2653.905 188.44 ;
    END
  END BcidMtx[166]
  PIN BcidMtx[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2650.265 187.44 2650.545 188.44 ;
    END
  END BcidMtx[162]
  PIN BcidMtx[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2576.905 187.44 2577.185 188.44 ;
    END
  END BcidMtx[160]
  PIN BcidMtx[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2574.105 187.44 2574.385 188.44 ;
    END
  END BcidMtx[157]
  PIN BcidMtx[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2507.465 187.44 2507.745 188.44 ;
    END
  END BcidMtx[155]
  PIN BcidMtx[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2504.105 187.44 2504.385 188.44 ;
    END
  END BcidMtx[151]
  PIN BcidMtx[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2428.225 187.44 2428.505 188.44 ;
    END
  END BcidMtx[148]
  PIN BcidMtx[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2400.505 187.44 2400.785 188.44 ;
    END
  END BcidMtx[146]
  PIN BcidMtx[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2320.985 187.44 2321.265 188.44 ;
    END
  END BcidMtx[142]
  PIN BcidMtx[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2317.625 187.44 2317.905 188.44 ;
    END
  END BcidMtx[138]
  PIN BcidMtx[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2256.025 187.44 2256.305 188.44 ;
    END
  END BcidMtx[137]
  PIN BcidMtx[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2253.225 187.44 2253.505 188.44 ;
    END
  END BcidMtx[134]
  PIN BcidMtx[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2252.105 187.44 2252.385 188.44 ;
    END
  END BcidMtx[132]
  PIN BcidMtx[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2173.705 187.44 2173.985 188.44 ;
    END
  END BcidMtx[131]
  PIN BcidMtx[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3214.185 187.44 3214.465 188.44 ;
    END
  END BcidMtx[209]
  PIN BcidMtx[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3210.825 187.44 3211.105 188.44 ;
    END
  END BcidMtx[205]
  PIN BcidMtx[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3136.905 187.44 3137.185 188.44 ;
    END
  END BcidMtx[202]
  PIN BcidMtx[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3133.545 187.44 3133.825 188.44 ;
    END
  END BcidMtx[198]
  PIN BcidMtx[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3066.905 187.44 3067.185 188.44 ;
    END
  END BcidMtx[196]
  PIN BcidMtx[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3063.545 187.44 3063.825 188.44 ;
    END
  END BcidMtx[192]
  PIN BcidMtx[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2987.665 187.44 2987.945 188.44 ;
    END
  END BcidMtx[189]
  PIN BcidMtx[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2959.945 187.44 2960.225 188.44 ;
    END
  END BcidMtx[187]
  PIN BcidMtx[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2881.545 187.44 2881.825 188.44 ;
    END
  END BcidMtx[185]
  PIN BcidMtx[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2880.425 187.44 2880.705 188.44 ;
    END
  END BcidMtx[183]
  PIN BcidMtx[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2877.625 187.44 2877.905 188.44 ;
    END
  END BcidMtx[180]
  PIN BcidMtx[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2815.465 187.44 2815.745 188.44 ;
    END
  END BcidMtx[178]
  PIN BcidMtx[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2812.665 187.44 2812.945 188.44 ;
    END
  END BcidMtx[175]
  PIN BcidMtx[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2733.145 187.44 2733.425 188.44 ;
    END
  END BcidMtx[172]
  PIN BcidMtx[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3773.625 187.44 3773.905 188.44 ;
    END
  END BcidMtx[250]
  PIN BcidMtx[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3696.345 187.44 3696.625 188.44 ;
    END
  END BcidMtx[243]
  PIN BcidMtx[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3694.105 187.44 3694.385 188.44 ;
    END
  END BcidMtx[241]
  PIN BcidMtx[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3627.465 187.44 3627.745 188.44 ;
    END
  END BcidMtx[239]
  PIN BcidMtx[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3624.105 187.44 3624.385 188.44 ;
    END
  END BcidMtx[235]
  PIN BcidMtx[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3548.225 187.44 3548.505 188.44 ;
    END
  END BcidMtx[232]
  PIN BcidMtx[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3519.945 187.44 3520.225 188.44 ;
    END
  END BcidMtx[229]
  PIN BcidMtx[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3441.545 187.44 3441.825 188.44 ;
    END
  END BcidMtx[227]
  PIN BcidMtx[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3375.465 187.44 3375.745 188.44 ;
    END
  END BcidMtx[220]
  PIN BcidMtx[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3372.665 187.44 3372.945 188.44 ;
    END
  END BcidMtx[217]
  PIN BcidMtx[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3293.705 187.44 3293.985 188.44 ;
    END
  END BcidMtx[215]
  PIN BcidMtx[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3292.585 187.44 3292.865 188.44 ;
    END
  END BcidMtx[213]
  PIN BcidMtx[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3290.905 187.44 3291.185 188.44 ;
    END
  END BcidMtx[212]
  PIN BcidMtx[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4334.185 187.44 4334.465 188.44 ;
    END
  END BcidMtx[293]
  PIN BcidMtx[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4330.265 187.44 4330.545 188.44 ;
    END
  END BcidMtx[288]
  PIN BcidMtx[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4257.465 187.44 4257.745 188.44 ;
    END
  END BcidMtx[287]
  PIN BcidMtx[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4186.905 187.44 4187.185 188.44 ;
    END
  END BcidMtx[280]
  PIN BcidMtx[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4186.345 187.44 4186.625 188.44 ;
    END
  END BcidMtx[279]
  PIN BcidMtx[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4184.665 187.44 4184.945 188.44 ;
    END
  END BcidMtx[278]
  PIN BcidMtx[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4107.665 187.44 4107.945 188.44 ;
    END
  END BcidMtx[273]
  PIN BcidMtx[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4079.385 187.44 4079.665 188.44 ;
    END
  END BcidMtx[270]
  PIN BcidMtx[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4001.545 187.44 4001.825 188.44 ;
    END
  END BcidMtx[269]
  PIN BcidMtx[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3998.745 187.44 3999.025 188.44 ;
    END
  END BcidMtx[266]
  PIN BcidMtx[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3998.185 187.44 3998.465 188.44 ;
    END
  END BcidMtx[265]
  PIN BcidMtx[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3934.905 187.44 3935.185 188.44 ;
    END
  END BcidMtx[261]
  PIN BcidMtx[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3932.105 187.44 3932.385 188.44 ;
    END
  END BcidMtx[258]
  PIN BcidMtx[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3850.345 187.44 3850.625 188.44 ;
    END
  END BcidMtx[253]
  PIN BcidMtx[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3849.785 187.44 3850.065 188.44 ;
    END
  END BcidMtx[252]
  PIN BcidMtx[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4893.625 187.44 4893.905 188.44 ;
    END
  END BcidMtx[334]
  PIN BcidMtx[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4890.825 187.44 4891.105 188.44 ;
    END
  END BcidMtx[331]
  PIN BcidMtx[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4890.265 187.44 4890.545 188.44 ;
    END
  END BcidMtx[330]
  PIN BcidMtx[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4817.465 187.44 4817.745 188.44 ;
    END
  END BcidMtx[329]
  PIN BcidMtx[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4747.465 187.44 4747.745 188.44 ;
    END
  END BcidMtx[323]
  PIN BcidMtx[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4668.225 187.44 4668.505 188.44 ;
    END
  END BcidMtx[316]
  PIN BcidMtx[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4667.665 187.44 4667.945 188.44 ;
    END
  END BcidMtx[315]
  PIN BcidMtx[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4639.945 187.44 4640.225 188.44 ;
    END
  END BcidMtx[313]
  PIN BcidMtx[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4560.425 187.44 4560.705 188.44 ;
    END
  END BcidMtx[309]
  PIN BcidMtx[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4558.185 187.44 4558.465 188.44 ;
    END
  END BcidMtx[307]
  PIN BcidMtx[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4494.905 187.44 4495.185 188.44 ;
    END
  END BcidMtx[303]
  PIN BcidMtx[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4493.225 187.44 4493.505 188.44 ;
    END
  END BcidMtx[302]
  PIN BcidMtx[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4412.585 187.44 4412.865 188.44 ;
    END
  END BcidMtx[297]
  PIN BcidMtx[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4410.345 187.44 4410.625 188.44 ;
    END
  END BcidMtx[295]
  PIN BcidMtx[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5453.625 187.44 5453.905 188.44 ;
    END
  END BcidMtx[376]
  PIN BcidMtx[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5450.825 187.44 5451.105 188.44 ;
    END
  END BcidMtx[373]
  PIN BcidMtx[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5377.465 187.44 5377.745 188.44 ;
    END
  END BcidMtx[371]
  PIN BcidMtx[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5373.545 187.44 5373.825 188.44 ;
    END
  END BcidMtx[366]
  PIN BcidMtx[1331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18187.465 187.44 18187.745 188.44 ;
    END
  END BcidMtx[1331]
  PIN BcidMtx[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5306.905 187.44 5307.185 188.44 ;
    END
  END BcidMtx[364]
  PIN BcidMtx[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5228.225 187.44 5228.505 188.44 ;
    END
  END BcidMtx[358]
  PIN BcidMtx[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5199.385 187.44 5199.665 188.44 ;
    END
  END BcidMtx[354]
  PIN BcidMtx[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5120.985 187.44 5121.265 188.44 ;
    END
  END BcidMtx[352]
  PIN BcidMtx[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5117.625 187.44 5117.905 188.44 ;
    END
  END BcidMtx[348]
  PIN BcidMtx[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5054.905 187.44 5055.185 188.44 ;
    END
  END BcidMtx[345]
  PIN BcidMtx[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5052.105 187.44 5052.385 188.44 ;
    END
  END BcidMtx[342]
  PIN BcidMtx[1330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18186.905 187.44 18187.185 188.44 ;
    END
  END BcidMtx[1330]
  PIN BcidMtx[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4973.145 187.44 4973.425 188.44 ;
    END
  END BcidMtx[340]
  PIN BcidMtx[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4970.345 187.44 4970.625 188.44 ;
    END
  END BcidMtx[337]
  PIN BcidMtx[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6013.065 187.44 6013.345 188.44 ;
    END
  END BcidMtx[417]
  PIN BcidMtx[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6011.385 187.44 6011.665 188.44 ;
    END
  END BcidMtx[416]
  PIN BcidMtx[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5937.465 187.44 5937.745 188.44 ;
    END
  END BcidMtx[413]
  PIN BcidMtx[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5934.105 187.44 5934.385 188.44 ;
    END
  END BcidMtx[409]
  PIN BcidMtx[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5866.345 187.44 5866.625 188.44 ;
    END
  END BcidMtx[405]
  PIN BcidMtx[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5863.545 187.44 5863.825 188.44 ;
    END
  END BcidMtx[402]
  PIN BcidMtx[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5788.785 187.44 5789.065 188.44 ;
    END
  END BcidMtx[401]
  PIN BcidMtx[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5760.505 187.44 5760.785 188.44 ;
    END
  END BcidMtx[398]
  PIN BcidMtx[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5759.385 187.44 5759.665 188.44 ;
    END
  END BcidMtx[396]
  PIN BcidMtx[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5681.545 187.44 5681.825 188.44 ;
    END
  END BcidMtx[395]
  PIN BcidMtx[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5678.185 187.44 5678.465 188.44 ;
    END
  END BcidMtx[391]
  PIN BcidMtx[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5614.905 187.44 5615.185 188.44 ;
    END
  END BcidMtx[387]
  PIN BcidMtx[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5613.225 187.44 5613.505 188.44 ;
    END
  END BcidMtx[386]
  PIN BcidMtx[1327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18184.105 187.44 18184.385 188.44 ;
    END
  END BcidMtx[1327]
  PIN BcidMtx[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5533.145 187.44 5533.425 188.44 ;
    END
  END BcidMtx[382]
  PIN BcidMtx[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5530.345 187.44 5530.625 188.44 ;
    END
  END BcidMtx[379]
  PIN BcidMtx[459]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6573.065 187.44 6573.345 188.44 ;
    END
  END BcidMtx[459]
  PIN BcidMtx[458]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6571.385 187.44 6571.665 188.44 ;
    END
  END BcidMtx[458]
  PIN BcidMtx[453]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6496.345 187.44 6496.625 188.44 ;
    END
  END BcidMtx[453]
  PIN BcidMtx[450]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6493.545 187.44 6493.825 188.44 ;
    END
  END BcidMtx[450]
  PIN BcidMtx[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6424.665 187.44 6424.945 188.44 ;
    END
  END BcidMtx[446]
  PIN BcidMtx[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6348.225 187.44 6348.505 188.44 ;
    END
  END BcidMtx[442]
  PIN BcidMtx[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6319.945 187.44 6320.225 188.44 ;
    END
  END BcidMtx[439]
  PIN BcidMtx[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6240.985 187.44 6241.265 188.44 ;
    END
  END BcidMtx[436]
  PIN BcidMtx[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6237.625 187.44 6237.905 188.44 ;
    END
  END BcidMtx[432]
  PIN BcidMtx[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6175.465 187.44 6175.745 188.44 ;
    END
  END BcidMtx[430]
  PIN BcidMtx[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6093.145 187.44 6093.425 188.44 ;
    END
  END BcidMtx[424]
  PIN BcidMtx[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6090.345 187.44 6090.625 188.44 ;
    END
  END BcidMtx[421]
  PIN BcidMtx[503]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7134.185 187.44 7134.465 188.44 ;
    END
  END BcidMtx[503]
  PIN BcidMtx[501]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7133.065 187.44 7133.345 188.44 ;
    END
  END BcidMtx[501]
  PIN BcidMtx[500]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7131.385 187.44 7131.665 188.44 ;
    END
  END BcidMtx[500]
  PIN BcidMtx[496]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7056.905 187.44 7057.185 188.44 ;
    END
  END BcidMtx[496]
  PIN BcidMtx[493]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7054.105 187.44 7054.385 188.44 ;
    END
  END BcidMtx[493]
  PIN BcidMtx[489]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6986.345 187.44 6986.625 188.44 ;
    END
  END BcidMtx[489]
  PIN BcidMtx[486]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6983.545 187.44 6983.825 188.44 ;
    END
  END BcidMtx[486]
  PIN BcidMtx[485]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6908.785 187.44 6909.065 188.44 ;
    END
  END BcidMtx[485]
  PIN BcidMtx[482]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6880.505 187.44 6880.785 188.44 ;
    END
  END BcidMtx[482]
  PIN BcidMtx[480]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6879.385 187.44 6879.665 188.44 ;
    END
  END BcidMtx[480]
  PIN BcidMtx[479]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6801.545 187.44 6801.825 188.44 ;
    END
  END BcidMtx[479]
  PIN BcidMtx[475]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6798.185 187.44 6798.465 188.44 ;
    END
  END BcidMtx[475]
  PIN BcidMtx[472]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6735.465 187.44 6735.745 188.44 ;
    END
  END BcidMtx[472]
  PIN BcidMtx[470]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6733.225 187.44 6733.505 188.44 ;
    END
  END BcidMtx[470]
  PIN BcidMtx[467]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6653.705 187.44 6653.985 188.44 ;
    END
  END BcidMtx[467]
  PIN BcidMtx[465]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6652.585 187.44 6652.865 188.44 ;
    END
  END BcidMtx[465]
  PIN BcidMtx[464]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6650.905 187.44 6651.185 188.44 ;
    END
  END BcidMtx[464]
  PIN BcidMtx[542]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7691.385 187.44 7691.665 188.44 ;
    END
  END BcidMtx[542]
  PIN BcidMtx[538]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7616.905 187.44 7617.185 188.44 ;
    END
  END BcidMtx[538]
  PIN BcidMtx[536]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7614.665 187.44 7614.945 188.44 ;
    END
  END BcidMtx[536]
  PIN BcidMtx[531]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7546.345 187.44 7546.625 188.44 ;
    END
  END BcidMtx[531]
  PIN BcidMtx[528]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7543.545 187.44 7543.825 188.44 ;
    END
  END BcidMtx[528]
  PIN BcidMtx[527]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7468.785 187.44 7469.065 188.44 ;
    END
  END BcidMtx[527]
  PIN BcidMtx[525]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7467.665 187.44 7467.945 188.44 ;
    END
  END BcidMtx[525]
  PIN BcidMtx[523]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7439.945 187.44 7440.225 188.44 ;
    END
  END BcidMtx[523]
  PIN BcidMtx[518]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7358.745 187.44 7359.025 188.44 ;
    END
  END BcidMtx[518]
  PIN BcidMtx[514]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7295.465 187.44 7295.745 188.44 ;
    END
  END BcidMtx[514]
  PIN BcidMtx[512]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7293.225 187.44 7293.505 188.44 ;
    END
  END BcidMtx[512]
  PIN BcidMtx[508]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7213.145 187.44 7213.425 188.44 ;
    END
  END BcidMtx[508]
  PIN BcidMtx[505]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7210.345 187.44 7210.625 188.44 ;
    END
  END BcidMtx[505]
  PIN BcidMtx[504]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7209.785 187.44 7210.065 188.44 ;
    END
  END BcidMtx[504]
  PIN BcidMtx[587]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8254.185 187.44 8254.465 188.44 ;
    END
  END BcidMtx[587]
  PIN BcidMtx[584]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8251.385 187.44 8251.665 188.44 ;
    END
  END BcidMtx[584]
  PIN BcidMtx[581]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8177.465 187.44 8177.745 188.44 ;
    END
  END BcidMtx[581]
  PIN BcidMtx[577]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8174.105 187.44 8174.385 188.44 ;
    END
  END BcidMtx[577]
  PIN BcidMtx[573]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8106.345 187.44 8106.625 188.44 ;
    END
  END BcidMtx[573]
  PIN BcidMtx[572]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8104.665 187.44 8104.945 188.44 ;
    END
  END BcidMtx[572]
  PIN BcidMtx[568]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8028.225 187.44 8028.505 188.44 ;
    END
  END BcidMtx[568]
  PIN BcidMtx[566]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8000.505 187.44 8000.785 188.44 ;
    END
  END BcidMtx[566]
  PIN BcidMtx[565]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7999.945 187.44 8000.225 188.44 ;
    END
  END BcidMtx[565]
  PIN BcidMtx[563]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7921.545 187.44 7921.825 188.44 ;
    END
  END BcidMtx[563]
  PIN BcidMtx[559]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7918.185 187.44 7918.465 188.44 ;
    END
  END BcidMtx[559]
  PIN BcidMtx[556]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7855.465 187.44 7855.745 188.44 ;
    END
  END BcidMtx[556]
  PIN BcidMtx[553]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7852.665 187.44 7852.945 188.44 ;
    END
  END BcidMtx[553]
  PIN BcidMtx[551]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7773.705 187.44 7773.985 188.44 ;
    END
  END BcidMtx[551]
  PIN BcidMtx[549]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7772.585 187.44 7772.865 188.44 ;
    END
  END BcidMtx[549]
  PIN BcidMtx[547]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7770.345 187.44 7770.625 188.44 ;
    END
  END BcidMtx[547]
  PIN BcidMtx[628]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8813.625 187.44 8813.905 188.44 ;
    END
  END BcidMtx[628]
  PIN BcidMtx[624]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8810.265 187.44 8810.545 188.44 ;
    END
  END BcidMtx[624]
  PIN BcidMtx[621]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8736.345 187.44 8736.625 188.44 ;
    END
  END BcidMtx[621]
  PIN BcidMtx[620]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8734.665 187.44 8734.945 188.44 ;
    END
  END BcidMtx[620]
  PIN BcidMtx[617]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8667.465 187.44 8667.745 188.44 ;
    END
  END BcidMtx[617]
  PIN BcidMtx[613]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8664.105 187.44 8664.385 188.44 ;
    END
  END BcidMtx[613]
  PIN BcidMtx[609]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8587.665 187.44 8587.945 188.44 ;
    END
  END BcidMtx[609]
  PIN BcidMtx[607]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8559.945 187.44 8560.225 188.44 ;
    END
  END BcidMtx[607]
  PIN BcidMtx[604]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8480.985 187.44 8481.265 188.44 ;
    END
  END BcidMtx[604]
  PIN BcidMtx[600]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8477.625 187.44 8477.905 188.44 ;
    END
  END BcidMtx[600]
  PIN BcidMtx[598]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8415.465 187.44 8415.745 188.44 ;
    END
  END BcidMtx[598]
  PIN BcidMtx[594]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8412.105 187.44 8412.385 188.44 ;
    END
  END BcidMtx[594]
  PIN BcidMtx[593]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8333.705 187.44 8333.985 188.44 ;
    END
  END BcidMtx[593]
  PIN BcidMtx[588]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8329.785 187.44 8330.065 188.44 ;
    END
  END BcidMtx[588]
  PIN BcidMtx[671]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9374.185 187.44 9374.465 188.44 ;
    END
  END BcidMtx[671]
  PIN BcidMtx[666]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9370.265 187.44 9370.545 188.44 ;
    END
  END BcidMtx[666]
  PIN BcidMtx[664]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9296.905 187.44 9297.185 188.44 ;
    END
  END BcidMtx[664]
  PIN BcidMtx[658]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9226.905 187.44 9227.185 188.44 ;
    END
  END BcidMtx[658]
  PIN BcidMtx[655]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9224.105 187.44 9224.385 188.44 ;
    END
  END BcidMtx[655]
  PIN BcidMtx[651]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9147.665 187.44 9147.945 188.44 ;
    END
  END BcidMtx[651]
  PIN BcidMtx[649]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9119.945 187.44 9120.225 188.44 ;
    END
  END BcidMtx[649]
  PIN BcidMtx[647]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9041.545 187.44 9041.825 188.44 ;
    END
  END BcidMtx[647]
  PIN BcidMtx[643]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9038.185 187.44 9038.465 188.44 ;
    END
  END BcidMtx[643]
  PIN BcidMtx[640]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8975.465 187.44 8975.745 188.44 ;
    END
  END BcidMtx[640]
  PIN BcidMtx[638]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8973.225 187.44 8973.505 188.44 ;
    END
  END BcidMtx[638]
  PIN BcidMtx[633]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8892.585 187.44 8892.865 188.44 ;
    END
  END BcidMtx[633]
  PIN BcidMtx[630]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8889.785 187.44 8890.065 188.44 ;
    END
  END BcidMtx[630]
  PIN BcidMtx[712]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9933.625 187.44 9933.905 188.44 ;
    END
  END BcidMtx[712]
  PIN BcidMtx[710]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9931.385 187.44 9931.665 188.44 ;
    END
  END BcidMtx[710]
  PIN BcidMtx[705]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9856.345 187.44 9856.625 188.44 ;
    END
  END BcidMtx[705]
  PIN BcidMtx[703]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9854.105 187.44 9854.385 188.44 ;
    END
  END BcidMtx[703]
  PIN BcidMtx[701]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9787.465 187.44 9787.745 188.44 ;
    END
  END BcidMtx[701]
  PIN BcidMtx[698]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9784.665 187.44 9784.945 188.44 ;
    END
  END BcidMtx[698]
  PIN BcidMtx[696]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9783.545 187.44 9783.825 188.44 ;
    END
  END BcidMtx[696]
  PIN BcidMtx[695]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9708.785 187.44 9709.065 188.44 ;
    END
  END BcidMtx[695]
  PIN BcidMtx[693]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9707.665 187.44 9707.945 188.44 ;
    END
  END BcidMtx[693]
  PIN BcidMtx[689]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9601.545 187.44 9601.825 188.44 ;
    END
  END BcidMtx[689]
  PIN BcidMtx[687]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9600.425 187.44 9600.705 188.44 ;
    END
  END BcidMtx[687]
  PIN BcidMtx[683]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9536.025 187.44 9536.305 188.44 ;
    END
  END BcidMtx[683]
  PIN BcidMtx[676]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9453.145 187.44 9453.425 188.44 ;
    END
  END BcidMtx[676]
  PIN BcidMtx[755]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10494.185 187.44 10494.465 188.44 ;
    END
  END BcidMtx[755]
  PIN BcidMtx[753]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10493.065 187.44 10493.345 188.44 ;
    END
  END BcidMtx[753]
  PIN BcidMtx[752]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10491.385 187.44 10491.665 188.44 ;
    END
  END BcidMtx[752]
  PIN BcidMtx[748]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10416.905 187.44 10417.185 188.44 ;
    END
  END BcidMtx[748]
  PIN BcidMtx[747]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10416.345 187.44 10416.625 188.44 ;
    END
  END BcidMtx[747]
  PIN BcidMtx[746]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10414.665 187.44 10414.945 188.44 ;
    END
  END BcidMtx[746]
  PIN BcidMtx[738]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10343.545 187.44 10343.825 188.44 ;
    END
  END BcidMtx[738]
  PIN BcidMtx[737]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10268.785 187.44 10269.065 188.44 ;
    END
  END BcidMtx[737]
  PIN BcidMtx[733]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10239.945 187.44 10240.225 188.44 ;
    END
  END BcidMtx[733]
  PIN BcidMtx[732]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10239.385 187.44 10239.665 188.44 ;
    END
  END BcidMtx[732]
  PIN BcidMtx[730]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10160.985 187.44 10161.265 188.44 ;
    END
  END BcidMtx[730]
  PIN BcidMtx[727]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10158.185 187.44 10158.465 188.44 ;
    END
  END BcidMtx[727]
  PIN BcidMtx[726]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10157.625 187.44 10157.905 188.44 ;
    END
  END BcidMtx[726]
  PIN BcidMtx[724]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10095.465 187.44 10095.745 188.44 ;
    END
  END BcidMtx[724]
  PIN BcidMtx[721]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10092.665 187.44 10092.945 188.44 ;
    END
  END BcidMtx[721]
  PIN BcidMtx[720]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10092.105 187.44 10092.385 188.44 ;
    END
  END BcidMtx[720]
  PIN BcidMtx[719]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10013.705 187.44 10013.985 188.44 ;
    END
  END BcidMtx[719]
  PIN BcidMtx[716]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10010.905 187.44 10011.185 188.44 ;
    END
  END BcidMtx[716]
  PIN BcidMtx[715]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10010.345 187.44 10010.625 188.44 ;
    END
  END BcidMtx[715]
  PIN BcidMtx[796]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11053.625 187.44 11053.905 188.44 ;
    END
  END BcidMtx[796]
  PIN BcidMtx[793]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11050.825 187.44 11051.105 188.44 ;
    END
  END BcidMtx[793]
  PIN BcidMtx[792]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11050.265 187.44 11050.545 188.44 ;
    END
  END BcidMtx[792]
  PIN BcidMtx[791]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10977.465 187.44 10977.745 188.44 ;
    END
  END BcidMtx[791]
  PIN BcidMtx[784]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10906.905 187.44 10907.185 188.44 ;
    END
  END BcidMtx[784]
  PIN BcidMtx[783]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10906.345 187.44 10906.625 188.44 ;
    END
  END BcidMtx[783]
  PIN BcidMtx[782]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10904.665 187.44 10904.945 188.44 ;
    END
  END BcidMtx[782]
  PIN BcidMtx[776]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10800.505 187.44 10800.785 188.44 ;
    END
  END BcidMtx[776]
  PIN BcidMtx[772]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10720.985 187.44 10721.265 188.44 ;
    END
  END BcidMtx[772]
  PIN BcidMtx[769]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10718.185 187.44 10718.465 188.44 ;
    END
  END BcidMtx[769]
  PIN BcidMtx[766]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10655.465 187.44 10655.745 188.44 ;
    END
  END BcidMtx[766]
  PIN BcidMtx[763]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10652.665 187.44 10652.945 188.44 ;
    END
  END BcidMtx[763]
  PIN BcidMtx[762]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10652.105 187.44 10652.385 188.44 ;
    END
  END BcidMtx[762]
  PIN BcidMtx[759]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10572.585 187.44 10572.865 188.44 ;
    END
  END BcidMtx[759]
  PIN BcidMtx[758]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10570.905 187.44 10571.185 188.44 ;
    END
  END BcidMtx[758]
  PIN BcidMtx[756]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10569.785 187.44 10570.065 188.44 ;
    END
  END BcidMtx[756]
  PIN BcidMtx[837]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11613.065 187.44 11613.345 188.44 ;
    END
  END BcidMtx[837]
  PIN BcidMtx[836]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11611.385 187.44 11611.665 188.44 ;
    END
  END BcidMtx[836]
  PIN BcidMtx[829]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11534.105 187.44 11534.385 188.44 ;
    END
  END BcidMtx[829]
  PIN BcidMtx[825]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11466.345 187.44 11466.625 188.44 ;
    END
  END BcidMtx[825]
  PIN BcidMtx[824]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11464.665 187.44 11464.945 188.44 ;
    END
  END BcidMtx[824]
  PIN BcidMtx[820]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11388.225 187.44 11388.505 188.44 ;
    END
  END BcidMtx[820]
  PIN BcidMtx[816]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11359.385 187.44 11359.665 188.44 ;
    END
  END BcidMtx[816]
  PIN BcidMtx[815]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11281.545 187.44 11281.825 188.44 ;
    END
  END BcidMtx[815]
  PIN BcidMtx[811]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11278.185 187.44 11278.465 188.44 ;
    END
  END BcidMtx[811]
  PIN BcidMtx[801]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11132.585 187.44 11132.865 188.44 ;
    END
  END BcidMtx[801]
  PIN BcidMtx[798]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11129.785 187.44 11130.065 188.44 ;
    END
  END BcidMtx[798]
  PIN BcidMtx[877]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12170.825 187.44 12171.105 188.44 ;
    END
  END BcidMtx[877]
  PIN BcidMtx[876]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12170.265 187.44 12170.545 188.44 ;
    END
  END BcidMtx[876]
  PIN BcidMtx[874]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12096.905 187.44 12097.185 188.44 ;
    END
  END BcidMtx[874]
  PIN BcidMtx[871]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12094.105 187.44 12094.385 188.44 ;
    END
  END BcidMtx[871]
  PIN BcidMtx[869]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12027.465 187.44 12027.745 188.44 ;
    END
  END BcidMtx[869]
  PIN BcidMtx[864]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12023.545 187.44 12023.825 188.44 ;
    END
  END BcidMtx[864]
  PIN BcidMtx[862]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11948.225 187.44 11948.505 188.44 ;
    END
  END BcidMtx[862]
  PIN BcidMtx[860]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11920.505 187.44 11920.785 188.44 ;
    END
  END BcidMtx[860]
  PIN BcidMtx[857]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11841.545 187.44 11841.825 188.44 ;
    END
  END BcidMtx[857]
  PIN BcidMtx[853]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11838.185 187.44 11838.465 188.44 ;
    END
  END BcidMtx[853]
  PIN BcidMtx[850]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11775.465 187.44 11775.745 188.44 ;
    END
  END BcidMtx[850]
  PIN BcidMtx[846]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11772.105 187.44 11772.385 188.44 ;
    END
  END BcidMtx[846]
  PIN BcidMtx[842]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11690.905 187.44 11691.185 188.44 ;
    END
  END BcidMtx[842]
  PIN BcidMtx[920]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12731.385 187.44 12731.665 188.44 ;
    END
  END BcidMtx[920]
  PIN BcidMtx[916]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12656.905 187.44 12657.185 188.44 ;
    END
  END BcidMtx[916]
  PIN BcidMtx[914]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12654.665 187.44 12654.945 188.44 ;
    END
  END BcidMtx[914]
  PIN BcidMtx[912]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12653.545 187.44 12653.825 188.44 ;
    END
  END BcidMtx[912]
  PIN BcidMtx[911]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12587.465 187.44 12587.745 188.44 ;
    END
  END BcidMtx[911]
  PIN BcidMtx[907]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12584.105 187.44 12584.385 188.44 ;
    END
  END BcidMtx[907]
  PIN BcidMtx[905]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12508.785 187.44 12509.065 188.44 ;
    END
  END BcidMtx[905]
  PIN BcidMtx[899]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12401.545 187.44 12401.825 188.44 ;
    END
  END BcidMtx[899]
  PIN BcidMtx[894]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12397.625 187.44 12397.905 188.44 ;
    END
  END BcidMtx[894]
  PIN BcidMtx[891]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12334.905 187.44 12335.185 188.44 ;
    END
  END BcidMtx[891]
  PIN BcidMtx[889]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12332.665 187.44 12332.945 188.44 ;
    END
  END BcidMtx[889]
  PIN BcidMtx[886]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12253.145 187.44 12253.425 188.44 ;
    END
  END BcidMtx[886]
  PIN BcidMtx[964]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13293.625 187.44 13293.905 188.44 ;
    END
  END BcidMtx[964]
  PIN BcidMtx[958]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13216.905 187.44 13217.185 188.44 ;
    END
  END BcidMtx[958]
  PIN BcidMtx[955]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13214.105 187.44 13214.385 188.44 ;
    END
  END BcidMtx[955]
  PIN BcidMtx[950]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13144.665 187.44 13144.945 188.44 ;
    END
  END BcidMtx[950]
  PIN BcidMtx[946]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13068.225 187.44 13068.505 188.44 ;
    END
  END BcidMtx[946]
  PIN BcidMtx[943]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13039.945 187.44 13040.225 188.44 ;
    END
  END BcidMtx[943]
  PIN BcidMtx[939]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12960.425 187.44 12960.705 188.44 ;
    END
  END BcidMtx[939]
  PIN BcidMtx[937]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12958.185 187.44 12958.465 188.44 ;
    END
  END BcidMtx[937]
  PIN BcidMtx[933]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12894.905 187.44 12895.185 188.44 ;
    END
  END BcidMtx[933]
  PIN BcidMtx[931]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12892.665 187.44 12892.945 188.44 ;
    END
  END BcidMtx[931]
  PIN BcidMtx[929]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12813.705 187.44 12813.985 188.44 ;
    END
  END BcidMtx[929]
  PIN BcidMtx[925]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12810.345 187.44 12810.625 188.44 ;
    END
  END BcidMtx[925]
  PIN BcidMtx[1313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17936.025 187.44 17936.305 188.44 ;
    END
  END BcidMtx[1313]
  PIN BcidMtx[1006]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13853.625 187.44 13853.905 188.44 ;
    END
  END BcidMtx[1006]
  PIN BcidMtx[1002]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13850.265 187.44 13850.545 188.44 ;
    END
  END BcidMtx[1002]
  PIN BcidMtx[999]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13776.345 187.44 13776.625 188.44 ;
    END
  END BcidMtx[999]
  PIN BcidMtx[997]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13774.105 187.44 13774.385 188.44 ;
    END
  END BcidMtx[997]
  PIN BcidMtx[994]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13706.905 187.44 13707.185 188.44 ;
    END
  END BcidMtx[994]
  PIN BcidMtx[988]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13628.225 187.44 13628.505 188.44 ;
    END
  END BcidMtx[988]
  PIN BcidMtx[984]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13599.385 187.44 13599.665 188.44 ;
    END
  END BcidMtx[984]
  PIN BcidMtx[1312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17935.465 187.44 17935.745 188.44 ;
    END
  END BcidMtx[1312]
  PIN BcidMtx[980]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13518.745 187.44 13519.025 188.44 ;
    END
  END BcidMtx[980]
  PIN BcidMtx[977]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13456.025 187.44 13456.305 188.44 ;
    END
  END BcidMtx[977]
  PIN BcidMtx[973]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13452.665 187.44 13452.945 188.44 ;
    END
  END BcidMtx[973]
  PIN BcidMtx[970]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13373.145 187.44 13373.425 188.44 ;
    END
  END BcidMtx[970]
  PIN BcidMtx[967]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13370.345 187.44 13370.625 188.44 ;
    END
  END BcidMtx[967]
  PIN BcidMtx[1045]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14410.825 187.44 14411.105 188.44 ;
    END
  END BcidMtx[1045]
  PIN BcidMtx[1044]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14410.265 187.44 14410.545 188.44 ;
    END
  END BcidMtx[1044]
  PIN BcidMtx[1043]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14337.465 187.44 14337.745 188.44 ;
    END
  END BcidMtx[1043]
  PIN BcidMtx[1042]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14336.905 187.44 14337.185 188.44 ;
    END
  END BcidMtx[1042]
  PIN BcidMtx[1039]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14334.105 187.44 14334.385 188.44 ;
    END
  END BcidMtx[1039]
  PIN BcidMtx[1035]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14266.345 187.44 14266.625 188.44 ;
    END
  END BcidMtx[1035]
  PIN BcidMtx[1034]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14264.665 187.44 14264.945 188.44 ;
    END
  END BcidMtx[1034]
  PIN BcidMtx[1031]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14188.785 187.44 14189.065 188.44 ;
    END
  END BcidMtx[1031]
  PIN BcidMtx[1028]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14160.505 187.44 14160.785 188.44 ;
    END
  END BcidMtx[1028]
  PIN BcidMtx[1025]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14081.545 187.44 14081.825 188.44 ;
    END
  END BcidMtx[1025]
  PIN BcidMtx[1021]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14078.185 187.44 14078.465 188.44 ;
    END
  END BcidMtx[1021]
  PIN BcidMtx[1019]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14016.025 187.44 14016.305 188.44 ;
    END
  END BcidMtx[1019]
  PIN BcidMtx[1016]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14013.225 187.44 14013.505 188.44 ;
    END
  END BcidMtx[1016]
  PIN BcidMtx[1014]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14012.105 187.44 14012.385 188.44 ;
    END
  END BcidMtx[1014]
  PIN BcidMtx[1013]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13933.705 187.44 13933.985 188.44 ;
    END
  END BcidMtx[1013]
  PIN BcidMtx[1008]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13929.785 187.44 13930.065 188.44 ;
    END
  END BcidMtx[1008]
  PIN BcidMtx[1090]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14973.625 187.44 14973.905 188.44 ;
    END
  END BcidMtx[1090]
  PIN BcidMtx[1086]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14970.265 187.44 14970.545 188.44 ;
    END
  END BcidMtx[1086]
  PIN BcidMtx[1085]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14897.465 187.44 14897.745 188.44 ;
    END
  END BcidMtx[1085]
  PIN BcidMtx[1079]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14827.465 187.44 14827.745 188.44 ;
    END
  END BcidMtx[1079]
  PIN BcidMtx[1077]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14826.345 187.44 14826.625 188.44 ;
    END
  END BcidMtx[1077]
  PIN BcidMtx[1076]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14824.665 187.44 14824.945 188.44 ;
    END
  END BcidMtx[1076]
  PIN BcidMtx[1075]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14824.105 187.44 14824.385 188.44 ;
    END
  END BcidMtx[1075]
  PIN BcidMtx[1071]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14747.665 187.44 14747.945 188.44 ;
    END
  END BcidMtx[1071]
  PIN BcidMtx[1065]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14640.425 187.44 14640.705 188.44 ;
    END
  END BcidMtx[1065]
  PIN BcidMtx[1062]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14637.625 187.44 14637.905 188.44 ;
    END
  END BcidMtx[1062]
  PIN BcidMtx[1060]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14575.465 187.44 14575.745 188.44 ;
    END
  END BcidMtx[1060]
  PIN BcidMtx[1056]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14572.105 187.44 14572.385 188.44 ;
    END
  END BcidMtx[1056]
  PIN BcidMtx[1055]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14493.705 187.44 14493.985 188.44 ;
    END
  END BcidMtx[1055]
  PIN BcidMtx[1051]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14490.345 187.44 14490.625 188.44 ;
    END
  END BcidMtx[1051]
  PIN BcidMtx[1133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15534.185 187.44 15534.465 188.44 ;
    END
  END BcidMtx[1133]
  PIN BcidMtx[1129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15530.825 187.44 15531.105 188.44 ;
    END
  END BcidMtx[1129]
  PIN BcidMtx[1125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15456.345 187.44 15456.625 188.44 ;
    END
  END BcidMtx[1125]
  PIN BcidMtx[1123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15454.105 187.44 15454.385 188.44 ;
    END
  END BcidMtx[1123]
  PIN BcidMtx[1120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15386.905 187.44 15387.185 188.44 ;
    END
  END BcidMtx[1120]
  PIN BcidMtx[1116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15383.545 187.44 15383.825 188.44 ;
    END
  END BcidMtx[1116]
  PIN BcidMtx[1107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15200.425 187.44 15200.705 188.44 ;
    END
  END BcidMtx[1107]
  PIN BcidMtx[1104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15197.625 187.44 15197.905 188.44 ;
    END
  END BcidMtx[1104]
  PIN BcidMtx[1103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15136.025 187.44 15136.305 188.44 ;
    END
  END BcidMtx[1103]
  PIN BcidMtx[1101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15134.905 187.44 15135.185 188.44 ;
    END
  END BcidMtx[1101]
  PIN BcidMtx[1100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15133.225 187.44 15133.505 188.44 ;
    END
  END BcidMtx[1100]
  PIN BcidMtx[1096]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15053.145 187.44 15053.425 188.44 ;
    END
  END BcidMtx[1096]
  PIN BcidMtx[1093]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15050.345 187.44 15050.625 188.44 ;
    END
  END BcidMtx[1093]
  PIN BcidMtx[1174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16093.625 187.44 16093.905 188.44 ;
    END
  END BcidMtx[1174]
  PIN BcidMtx[1170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16090.265 187.44 16090.545 188.44 ;
    END
  END BcidMtx[1170]
  PIN BcidMtx[1169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16017.465 187.44 16017.745 188.44 ;
    END
  END BcidMtx[1169]
  PIN BcidMtx[1167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16016.345 187.44 16016.625 188.44 ;
    END
  END BcidMtx[1167]
  PIN BcidMtx[1166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16014.665 187.44 16014.945 188.44 ;
    END
  END BcidMtx[1166]
  PIN BcidMtx[1163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15947.465 187.44 15947.745 188.44 ;
    END
  END BcidMtx[1163]
  PIN BcidMtx[1161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15946.345 187.44 15946.625 188.44 ;
    END
  END BcidMtx[1161]
  PIN BcidMtx[1158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15943.545 187.44 15943.825 188.44 ;
    END
  END BcidMtx[1158]
  PIN BcidMtx[1157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15868.785 187.44 15869.065 188.44 ;
    END
  END BcidMtx[1157]
  PIN BcidMtx[1155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15867.665 187.44 15867.945 188.44 ;
    END
  END BcidMtx[1155]
  PIN BcidMtx[1151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15761.545 187.44 15761.825 188.44 ;
    END
  END BcidMtx[1151]
  PIN BcidMtx[1149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15760.425 187.44 15760.705 188.44 ;
    END
  END BcidMtx[1149]
  PIN BcidMtx[1143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15694.905 187.44 15695.185 188.44 ;
    END
  END BcidMtx[1143]
  PIN BcidMtx[1141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15692.665 187.44 15692.945 188.44 ;
    END
  END BcidMtx[1141]
  PIN BcidMtx[1136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15610.905 187.44 15611.185 188.44 ;
    END
  END BcidMtx[1136]
  PIN BcidMtx[1214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16651.385 187.44 16651.665 188.44 ;
    END
  END BcidMtx[1214]
  PIN BcidMtx[1209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16576.345 187.44 16576.625 188.44 ;
    END
  END BcidMtx[1209]
  PIN BcidMtx[1206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16573.545 187.44 16573.825 188.44 ;
    END
  END BcidMtx[1206]
  PIN BcidMtx[1205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16507.465 187.44 16507.745 188.44 ;
    END
  END BcidMtx[1205]
  PIN BcidMtx[1198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16428.225 187.44 16428.505 188.44 ;
    END
  END BcidMtx[1198]
  PIN BcidMtx[1197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16427.665 187.44 16427.945 188.44 ;
    END
  END BcidMtx[1197]
  PIN BcidMtx[1195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16399.945 187.44 16400.225 188.44 ;
    END
  END BcidMtx[1195]
  PIN BcidMtx[1319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18001.545 187.44 18001.825 188.44 ;
    END
  END BcidMtx[1319]
  PIN BcidMtx[1318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18000.985 187.44 18001.265 188.44 ;
    END
  END BcidMtx[1318]
  PIN BcidMtx[1191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16320.425 187.44 16320.705 188.44 ;
    END
  END BcidMtx[1191]
  PIN BcidMtx[1189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16318.185 187.44 16318.465 188.44 ;
    END
  END BcidMtx[1189]
  PIN BcidMtx[1317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18000.425 187.44 18000.705 188.44 ;
    END
  END BcidMtx[1317]
  PIN BcidMtx[1182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16252.105 187.44 16252.385 188.44 ;
    END
  END BcidMtx[1182]
  PIN BcidMtx[1178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16170.905 187.44 16171.185 188.44 ;
    END
  END BcidMtx[1178]
  PIN BcidMtx[1256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17211.385 187.44 17211.665 188.44 ;
    END
  END BcidMtx[1256]
  PIN BcidMtx[1252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17136.905 187.44 17137.185 188.44 ;
    END
  END BcidMtx[1252]
  PIN BcidMtx[1249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17134.105 187.44 17134.385 188.44 ;
    END
  END BcidMtx[1249]
  PIN BcidMtx[1248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17133.545 187.44 17133.825 188.44 ;
    END
  END BcidMtx[1248]
  PIN BcidMtx[1245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17066.345 187.44 17066.625 188.44 ;
    END
  END BcidMtx[1245]
  PIN BcidMtx[1242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17063.545 187.44 17063.825 188.44 ;
    END
  END BcidMtx[1242]
  PIN BcidMtx[1239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16987.665 187.44 16987.945 188.44 ;
    END
  END BcidMtx[1239]
  PIN BcidMtx[1316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17998.745 187.44 17999.025 188.44 ;
    END
  END BcidMtx[1316]
  PIN BcidMtx[1314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17997.625 187.44 17997.905 188.44 ;
    END
  END BcidMtx[1314]
  PIN BcidMtx[1233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16880.425 187.44 16880.705 188.44 ;
    END
  END BcidMtx[1233]
  PIN BcidMtx[1230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16877.625 187.44 16877.905 188.44 ;
    END
  END BcidMtx[1230]
  PIN BcidMtx[1229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16816.025 187.44 16816.305 188.44 ;
    END
  END BcidMtx[1229]
  PIN BcidMtx[1228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16815.465 187.44 16815.745 188.44 ;
    END
  END BcidMtx[1228]
  PIN BcidMtx[1221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16732.585 187.44 16732.865 188.44 ;
    END
  END BcidMtx[1221]
  PIN BcidMtx[1219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16730.345 187.44 16730.625 188.44 ;
    END
  END BcidMtx[1219]
  PIN BcidMtx[1300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17773.625 187.44 17773.905 188.44 ;
    END
  END BcidMtx[1300]
  PIN BcidMtx[1296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17770.265 187.44 17770.545 188.44 ;
    END
  END BcidMtx[1296]
  PIN BcidMtx[1295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17697.465 187.44 17697.745 188.44 ;
    END
  END BcidMtx[1295]
  PIN BcidMtx[1291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17694.105 187.44 17694.385 188.44 ;
    END
  END BcidMtx[1291]
  PIN BcidMtx[1289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17627.465 187.44 17627.745 188.44 ;
    END
  END BcidMtx[1289]
  PIN BcidMtx[1285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17624.105 187.44 17624.385 188.44 ;
    END
  END BcidMtx[1285]
  PIN BcidMtx[1278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17519.385 187.44 17519.665 188.44 ;
    END
  END BcidMtx[1278]
  PIN BcidMtx[1276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17440.985 187.44 17441.265 188.44 ;
    END
  END BcidMtx[1276]
  PIN BcidMtx[1273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17438.185 187.44 17438.465 188.44 ;
    END
  END BcidMtx[1273]
  PIN BcidMtx[1271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17376.025 187.44 17376.305 188.44 ;
    END
  END BcidMtx[1271]
  PIN BcidMtx[1269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17374.905 187.44 17375.185 188.44 ;
    END
  END BcidMtx[1269]
  PIN BcidMtx[1266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17372.105 187.44 17372.385 188.44 ;
    END
  END BcidMtx[1266]
  PIN BcidMtx[1263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17292.585 187.44 17292.865 188.44 ;
    END
  END BcidMtx[1263]
  PIN BcidMtx[1261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17290.345 187.44 17290.625 188.44 ;
    END
  END BcidMtx[1261]
  PIN BcidMtx[1342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18333.625 187.44 18333.905 188.44 ;
    END
  END BcidMtx[1342]
  PIN BcidMtx[1335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18256.345 187.44 18256.625 188.44 ;
    END
  END BcidMtx[1335]
  PIN BcidMtx[1333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18254.105 187.44 18254.385 188.44 ;
    END
  END BcidMtx[1333]
  PIN BcidMtx[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 973.625 187.44 973.905 188.44 ;
    END
  END BcidMtx[40]
  PIN BcidMtx[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 971.385 187.44 971.665 188.44 ;
    END
  END BcidMtx[38]
  PIN BcidMtx[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 897.465 187.44 897.745 188.44 ;
    END
  END BcidMtx[35]
  PIN BcidMtx[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 896.345 187.44 896.625 188.44 ;
    END
  END BcidMtx[33]
  PIN BcidMtx[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 894.105 187.44 894.385 188.44 ;
    END
  END BcidMtx[31]
  PIN BcidMtx[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 826.905 187.44 827.185 188.44 ;
    END
  END BcidMtx[28]
  PIN BcidMtx[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 823.545 187.44 823.825 188.44 ;
    END
  END BcidMtx[24]
  PIN BcidMtx[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 638.745 187.44 639.025 188.44 ;
    END
  END BcidMtx[14]
  PIN BcidMtx[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 748.225 187.44 748.505 188.44 ;
    END
  END BcidMtx[22]
  PIN BcidMtx[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 641.545 187.44 641.825 188.44 ;
    END
  END BcidMtx[17]
  PIN BcidMtx[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 638.185 187.44 638.465 188.44 ;
    END
  END BcidMtx[13]
  PIN BcidMtx[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 574.905 187.44 575.185 188.44 ;
    END
  END BcidMtx[9]
  PIN BcidMtx[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 572.105 187.44 572.385 188.44 ;
    END
  END BcidMtx[6]
  PIN BcidMtx[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1533.065 187.44 1533.345 188.44 ;
    END
  END BcidMtx[81]
  PIN BcidMtx[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1530.825 187.44 1531.105 188.44 ;
    END
  END BcidMtx[79]
  PIN BcidMtx[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1456.345 187.44 1456.625 188.44 ;
    END
  END BcidMtx[75]
  PIN BcidMtx[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1454.665 187.44 1454.945 188.44 ;
    END
  END BcidMtx[74]
  PIN BcidMtx[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1387.465 187.44 1387.745 188.44 ;
    END
  END BcidMtx[71]
  PIN BcidMtx[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1384.665 187.44 1384.945 188.44 ;
    END
  END BcidMtx[68]
  PIN BcidMtx[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1308.785 187.44 1309.065 188.44 ;
    END
  END BcidMtx[65]
  PIN BcidMtx[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1307.665 187.44 1307.945 188.44 ;
    END
  END BcidMtx[63]
  PIN BcidMtx[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1279.945 187.44 1280.225 188.44 ;
    END
  END BcidMtx[61]
  PIN BcidMtx[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1200.985 187.44 1201.265 188.44 ;
    END
  END BcidMtx[58]
  PIN BcidMtx[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1198.745 187.44 1199.025 188.44 ;
    END
  END BcidMtx[56]
  PIN BcidMtx[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1197.625 187.44 1197.905 188.44 ;
    END
  END BcidMtx[54]
  PIN BcidMtx[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1135.465 187.44 1135.745 188.44 ;
    END
  END BcidMtx[52]
  PIN BcidMtx[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1053.705 187.44 1053.985 188.44 ;
    END
  END BcidMtx[47]
  PIN BcidMtx[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1050.345 187.44 1050.625 188.44 ;
    END
  END BcidMtx[43]
  PIN BcidMtx[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2094.185 187.44 2094.465 188.44 ;
    END
  END BcidMtx[125]
  PIN BcidMtx[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2090.825 187.44 2091.105 188.44 ;
    END
  END BcidMtx[121]
  PIN BcidMtx[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2016.905 187.44 2017.185 188.44 ;
    END
  END BcidMtx[118]
  PIN BcidMtx[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2013.545 187.44 2013.825 188.44 ;
    END
  END BcidMtx[114]
  PIN BcidMtx[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1944.665 187.44 1944.945 188.44 ;
    END
  END BcidMtx[110]
  PIN BcidMtx[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1867.665 187.44 1867.945 188.44 ;
    END
  END BcidMtx[105]
  PIN BcidMtx[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1839.945 187.44 1840.225 188.44 ;
    END
  END BcidMtx[103]
  PIN BcidMtx[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1760.985 187.44 1761.265 188.44 ;
    END
  END BcidMtx[100]
  PIN BcidMtx[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1758.185 187.44 1758.465 188.44 ;
    END
  END BcidMtx[97]
  PIN BcidMtx[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1695.465 187.44 1695.745 188.44 ;
    END
  END BcidMtx[94]
  PIN BcidMtx[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1694.905 187.44 1695.185 188.44 ;
    END
  END BcidMtx[93]
  PIN BcidMtx[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1693.225 187.44 1693.505 188.44 ;
    END
  END BcidMtx[92]
  PIN BcidMtx[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1612.585 187.44 1612.865 188.44 ;
    END
  END BcidMtx[87]
  PIN BcidMtx[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1610.905 187.44 1611.185 188.44 ;
    END
  END BcidMtx[86]
  PIN BcidMtx[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1609.785 187.44 1610.065 188.44 ;
    END
  END BcidMtx[84]
  PIN BcidMtx[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2651.385 187.44 2651.665 188.44 ;
    END
  END BcidMtx[164]
  PIN BcidMtx[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2573.545 187.44 2573.825 188.44 ;
    END
  END BcidMtx[156]
  PIN BcidMtx[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2506.905 187.44 2507.185 188.44 ;
    END
  END BcidMtx[154]
  PIN BcidMtx[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2428.785 187.44 2429.065 188.44 ;
    END
  END BcidMtx[149]
  PIN BcidMtx[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2427.665 187.44 2427.945 188.44 ;
    END
  END BcidMtx[147]
  PIN BcidMtx[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2399.945 187.44 2400.225 188.44 ;
    END
  END BcidMtx[145]
  PIN BcidMtx[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2320.425 187.44 2320.705 188.44 ;
    END
  END BcidMtx[141]
  PIN BcidMtx[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2318.745 187.44 2319.025 188.44 ;
    END
  END BcidMtx[140]
  PIN BcidMtx[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2255.465 187.44 2255.745 188.44 ;
    END
  END BcidMtx[136]
  PIN BcidMtx[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2173.145 187.44 2173.425 188.44 ;
    END
  END BcidMtx[130]
  PIN BcidMtx[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2170.345 187.44 2170.625 188.44 ;
    END
  END BcidMtx[127]
  PIN BcidMtx[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3213.625 187.44 3213.905 188.44 ;
    END
  END BcidMtx[208]
  PIN BcidMtx[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3136.345 187.44 3136.625 188.44 ;
    END
  END BcidMtx[201]
  PIN BcidMtx[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3134.105 187.44 3134.385 188.44 ;
    END
  END BcidMtx[199]
  PIN BcidMtx[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3066.345 187.44 3066.625 188.44 ;
    END
  END BcidMtx[195]
  PIN BcidMtx[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3064.105 187.44 3064.385 188.44 ;
    END
  END BcidMtx[193]
  PIN BcidMtx[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2988.785 187.44 2989.065 188.44 ;
    END
  END BcidMtx[191]
  PIN BcidMtx[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2880.985 187.44 2881.265 188.44 ;
    END
  END BcidMtx[184]
  PIN BcidMtx[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2878.745 187.44 2879.025 188.44 ;
    END
  END BcidMtx[182]
  PIN BcidMtx[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2814.905 187.44 2815.185 188.44 ;
    END
  END BcidMtx[177]
  PIN BcidMtx[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2812.105 187.44 2812.385 188.44 ;
    END
  END BcidMtx[174]
  PIN BcidMtx[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2730.905 187.44 2731.185 188.44 ;
    END
  END BcidMtx[170]
  PIN BcidMtx[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2729.785 187.44 2730.065 188.44 ;
    END
  END BcidMtx[168]
  PIN BcidMtx[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3771.385 187.44 3771.665 188.44 ;
    END
  END BcidMtx[248]
  PIN BcidMtx[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3770.265 187.44 3770.545 188.44 ;
    END
  END BcidMtx[246]
  PIN BcidMtx[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3697.465 187.44 3697.745 188.44 ;
    END
  END BcidMtx[245]
  PIN BcidMtx[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3694.665 187.44 3694.945 188.44 ;
    END
  END BcidMtx[242]
  PIN BcidMtx[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3693.545 187.44 3693.825 188.44 ;
    END
  END BcidMtx[240]
  PIN BcidMtx[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3626.905 187.44 3627.185 188.44 ;
    END
  END BcidMtx[238]
  PIN BcidMtx[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3623.545 187.44 3623.825 188.44 ;
    END
  END BcidMtx[234]
  PIN BcidMtx[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3547.665 187.44 3547.945 188.44 ;
    END
  END BcidMtx[231]
  PIN BcidMtx[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3520.505 187.44 3520.785 188.44 ;
    END
  END BcidMtx[230]
  PIN BcidMtx[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3440.985 187.44 3441.265 188.44 ;
    END
  END BcidMtx[226]
  PIN BcidMtx[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3438.185 187.44 3438.465 188.44 ;
    END
  END BcidMtx[223]
  PIN BcidMtx[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3376.025 187.44 3376.305 188.44 ;
    END
  END BcidMtx[221]
  PIN BcidMtx[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3372.105 187.44 3372.385 188.44 ;
    END
  END BcidMtx[216]
  PIN BcidMtx[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3290.345 187.44 3290.625 188.44 ;
    END
  END BcidMtx[211]
  PIN BcidMtx[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3289.785 187.44 3290.065 188.44 ;
    END
  END BcidMtx[210]
  PIN BcidMtx[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4333.625 187.44 4333.905 188.44 ;
    END
  END BcidMtx[292]
  PIN BcidMtx[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4330.825 187.44 4331.105 188.44 ;
    END
  END BcidMtx[289]
  PIN BcidMtx[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4256.905 187.44 4257.185 188.44 ;
    END
  END BcidMtx[286]
  PIN BcidMtx[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4254.105 187.44 4254.385 188.44 ;
    END
  END BcidMtx[283]
  PIN BcidMtx[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4184.105 187.44 4184.385 188.44 ;
    END
  END BcidMtx[277]
  PIN BcidMtx[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4108.785 187.44 4109.065 188.44 ;
    END
  END BcidMtx[275]
  PIN BcidMtx[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4080.505 187.44 4080.785 188.44 ;
    END
  END BcidMtx[272]
  PIN BcidMtx[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4000.985 187.44 4001.265 188.44 ;
    END
  END BcidMtx[268]
  PIN BcidMtx[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3997.625 187.44 3997.905 188.44 ;
    END
  END BcidMtx[264]
  PIN BcidMtx[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3936.025 187.44 3936.305 188.44 ;
    END
  END BcidMtx[263]
  PIN BcidMtx[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3933.225 187.44 3933.505 188.44 ;
    END
  END BcidMtx[260]
  PIN BcidMtx[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3853.705 187.44 3853.985 188.44 ;
    END
  END BcidMtx[257]
  PIN BcidMtx[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3852.585 187.44 3852.865 188.44 ;
    END
  END BcidMtx[255]
  PIN BcidMtx[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4893.065 187.44 4893.345 188.44 ;
    END
  END BcidMtx[333]
  PIN BcidMtx[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4816.905 187.44 4817.185 188.44 ;
    END
  END BcidMtx[328]
  PIN BcidMtx[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4814.105 187.44 4814.385 188.44 ;
    END
  END BcidMtx[325]
  PIN BcidMtx[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4746.905 187.44 4747.185 188.44 ;
    END
  END BcidMtx[322]
  PIN BcidMtx[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4744.105 187.44 4744.385 188.44 ;
    END
  END BcidMtx[319]
  PIN BcidMtx[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4639.385 187.44 4639.665 188.44 ;
    END
  END BcidMtx[312]
  PIN BcidMtx[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4561.545 187.44 4561.825 188.44 ;
    END
  END BcidMtx[311]
  PIN BcidMtx[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4557.625 187.44 4557.905 188.44 ;
    END
  END BcidMtx[306]
  PIN BcidMtx[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4496.025 187.44 4496.305 188.44 ;
    END
  END BcidMtx[305]
  PIN BcidMtx[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4492.665 187.44 4492.945 188.44 ;
    END
  END BcidMtx[301]
  PIN BcidMtx[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4413.705 187.44 4413.985 188.44 ;
    END
  END BcidMtx[299]
  PIN BcidMtx[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4410.905 187.44 4411.185 188.44 ;
    END
  END BcidMtx[296]
  PIN BcidMtx[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4409.785 187.44 4410.065 188.44 ;
    END
  END BcidMtx[294]
  PIN BcidMtx[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5453.065 187.44 5453.345 188.44 ;
    END
  END BcidMtx[375]
  PIN BcidMtx[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5450.265 187.44 5450.545 188.44 ;
    END
  END BcidMtx[372]
  PIN BcidMtx[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5376.905 187.44 5377.185 188.44 ;
    END
  END BcidMtx[370]
  PIN BcidMtx[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5307.465 187.44 5307.745 188.44 ;
    END
  END BcidMtx[365]
  PIN BcidMtx[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5306.345 187.44 5306.625 188.44 ;
    END
  END BcidMtx[363]
  PIN BcidMtx[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5304.665 187.44 5304.945 188.44 ;
    END
  END BcidMtx[362]
  PIN BcidMtx[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5227.665 187.44 5227.945 188.44 ;
    END
  END BcidMtx[357]
  PIN BcidMtx[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5200.505 187.44 5200.785 188.44 ;
    END
  END BcidMtx[356]
  PIN BcidMtx[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5120.425 187.44 5120.705 188.44 ;
    END
  END BcidMtx[351]
  PIN BcidMtx[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5118.745 187.44 5119.025 188.44 ;
    END
  END BcidMtx[350]
  PIN BcidMtx[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5055.465 187.44 5055.745 188.44 ;
    END
  END BcidMtx[346]
  PIN BcidMtx[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5053.225 187.44 5053.505 188.44 ;
    END
  END BcidMtx[344]
  PIN BcidMtx[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4972.585 187.44 4972.865 188.44 ;
    END
  END BcidMtx[339]
  PIN BcidMtx[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4970.905 187.44 4971.185 188.44 ;
    END
  END BcidMtx[338]
  PIN BcidMtx[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4969.785 187.44 4970.065 188.44 ;
    END
  END BcidMtx[336]
  PIN BcidMtx[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6014.185 187.44 6014.465 188.44 ;
    END
  END BcidMtx[419]
  PIN BcidMtx[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6010.825 187.44 6011.105 188.44 ;
    END
  END BcidMtx[415]
  PIN BcidMtx[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5936.905 187.44 5937.185 188.44 ;
    END
  END BcidMtx[412]
  PIN BcidMtx[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5933.545 187.44 5933.825 188.44 ;
    END
  END BcidMtx[408]
  PIN BcidMtx[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5864.665 187.44 5864.945 188.44 ;
    END
  END BcidMtx[404]
  PIN BcidMtx[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5788.225 187.44 5788.505 188.44 ;
    END
  END BcidMtx[400]
  PIN BcidMtx[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5680.985 187.44 5681.265 188.44 ;
    END
  END BcidMtx[394]
  PIN BcidMtx[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5677.625 187.44 5677.905 188.44 ;
    END
  END BcidMtx[390]
  PIN BcidMtx[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5616.025 187.44 5616.305 188.44 ;
    END
  END BcidMtx[389]
  PIN BcidMtx[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5612.665 187.44 5612.945 188.44 ;
    END
  END BcidMtx[385]
  PIN BcidMtx[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5533.705 187.44 5533.985 188.44 ;
    END
  END BcidMtx[383]
  PIN BcidMtx[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5529.785 187.44 5530.065 188.44 ;
    END
  END BcidMtx[378]
  PIN BcidMtx[461]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6574.185 187.44 6574.465 188.44 ;
    END
  END BcidMtx[461]
  PIN BcidMtx[457]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6570.825 187.44 6571.105 188.44 ;
    END
  END BcidMtx[457]
  PIN BcidMtx[454]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6496.905 187.44 6497.185 188.44 ;
    END
  END BcidMtx[454]
  PIN BcidMtx[452]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6494.665 187.44 6494.945 188.44 ;
    END
  END BcidMtx[452]
  PIN BcidMtx[449]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6427.465 187.44 6427.745 188.44 ;
    END
  END BcidMtx[449]
  PIN BcidMtx[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6426.345 187.44 6426.625 188.44 ;
    END
  END BcidMtx[447]
  PIN BcidMtx[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6424.105 187.44 6424.385 188.44 ;
    END
  END BcidMtx[445]
  PIN BcidMtx[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6347.665 187.44 6347.945 188.44 ;
    END
  END BcidMtx[441]
  PIN BcidMtx[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6320.505 187.44 6320.785 188.44 ;
    END
  END BcidMtx[440]
  PIN BcidMtx[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6240.425 187.44 6240.705 188.44 ;
    END
  END BcidMtx[435]
  PIN BcidMtx[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6238.745 187.44 6239.025 188.44 ;
    END
  END BcidMtx[434]
  PIN BcidMtx[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6238.185 187.44 6238.465 188.44 ;
    END
  END BcidMtx[433]
  PIN BcidMtx[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6174.905 187.44 6175.185 188.44 ;
    END
  END BcidMtx[429]
  PIN BcidMtx[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6173.225 187.44 6173.505 188.44 ;
    END
  END BcidMtx[428]
  PIN BcidMtx[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6172.105 187.44 6172.385 188.44 ;
    END
  END BcidMtx[426]
  PIN BcidMtx[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6093.705 187.44 6093.985 188.44 ;
    END
  END BcidMtx[425]
  PIN BcidMtx[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6089.785 187.44 6090.065 188.44 ;
    END
  END BcidMtx[420]
  PIN BcidMtx[499]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7130.825 187.44 7131.105 188.44 ;
    END
  END BcidMtx[499]
  PIN BcidMtx[497]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7057.465 187.44 7057.745 188.44 ;
    END
  END BcidMtx[497]
  PIN BcidMtx[492]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7053.545 187.44 7053.825 188.44 ;
    END
  END BcidMtx[492]
  PIN BcidMtx[490]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6986.905 187.44 6987.185 188.44 ;
    END
  END BcidMtx[490]
  PIN BcidMtx[488]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6984.665 187.44 6984.945 188.44 ;
    END
  END BcidMtx[488]
  PIN BcidMtx[484]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6908.225 187.44 6908.505 188.44 ;
    END
  END BcidMtx[484]
  PIN BcidMtx[478]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6800.985 187.44 6801.265 188.44 ;
    END
  END BcidMtx[478]
  PIN BcidMtx[474]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6797.625 187.44 6797.905 188.44 ;
    END
  END BcidMtx[474]
  PIN BcidMtx[473]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6736.025 187.44 6736.305 188.44 ;
    END
  END BcidMtx[473]
  PIN BcidMtx[469]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6732.665 187.44 6732.945 188.44 ;
    END
  END BcidMtx[469]
  PIN BcidMtx[463]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6650.345 187.44 6650.625 188.44 ;
    END
  END BcidMtx[463]
  PIN BcidMtx[545]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7694.185 187.44 7694.465 188.44 ;
    END
  END BcidMtx[545]
  PIN BcidMtx[541]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7690.825 187.44 7691.105 188.44 ;
    END
  END BcidMtx[541]
  PIN BcidMtx[537]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7616.345 187.44 7616.625 188.44 ;
    END
  END BcidMtx[537]
  PIN BcidMtx[535]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7614.105 187.44 7614.385 188.44 ;
    END
  END BcidMtx[535]
  PIN BcidMtx[534]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7613.545 187.44 7613.825 188.44 ;
    END
  END BcidMtx[534]
  PIN BcidMtx[533]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7547.465 187.44 7547.745 188.44 ;
    END
  END BcidMtx[533]
  PIN BcidMtx[530]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7544.665 187.44 7544.945 188.44 ;
    END
  END BcidMtx[530]
  PIN BcidMtx[526]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7468.225 187.44 7468.505 188.44 ;
    END
  END BcidMtx[526]
  PIN BcidMtx[521]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7361.545 187.44 7361.825 188.44 ;
    END
  END BcidMtx[521]
  PIN BcidMtx[517]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7358.185 187.44 7358.465 188.44 ;
    END
  END BcidMtx[517]
  PIN BcidMtx[515]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7296.025 187.44 7296.305 188.44 ;
    END
  END BcidMtx[515]
  PIN BcidMtx[513]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7294.905 187.44 7295.185 188.44 ;
    END
  END BcidMtx[513]
  PIN BcidMtx[511]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7292.665 187.44 7292.945 188.44 ;
    END
  END BcidMtx[511]
  PIN BcidMtx[509]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7213.705 187.44 7213.985 188.44 ;
    END
  END BcidMtx[509]
  PIN BcidMtx[507]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7212.585 187.44 7212.865 188.44 ;
    END
  END BcidMtx[507]
  PIN BcidMtx[586]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8253.625 187.44 8253.905 188.44 ;
    END
  END BcidMtx[586]
  PIN BcidMtx[583]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8250.825 187.44 8251.105 188.44 ;
    END
  END BcidMtx[583]
  PIN BcidMtx[580]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8176.905 187.44 8177.185 188.44 ;
    END
  END BcidMtx[580]
  PIN BcidMtx[576]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8173.545 187.44 8173.825 188.44 ;
    END
  END BcidMtx[576]
  PIN BcidMtx[575]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8107.465 187.44 8107.745 188.44 ;
    END
  END BcidMtx[575]
  PIN BcidMtx[571]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8104.105 187.44 8104.385 188.44 ;
    END
  END BcidMtx[571]
  PIN BcidMtx[567]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8027.665 187.44 8027.945 188.44 ;
    END
  END BcidMtx[567]
  PIN BcidMtx[564]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7999.385 187.44 7999.665 188.44 ;
    END
  END BcidMtx[564]
  PIN BcidMtx[562]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7920.985 187.44 7921.265 188.44 ;
    END
  END BcidMtx[562]
  PIN BcidMtx[555]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7854.905 187.44 7855.185 188.44 ;
    END
  END BcidMtx[555]
  PIN BcidMtx[552]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7852.105 187.44 7852.385 188.44 ;
    END
  END BcidMtx[552]
  PIN BcidMtx[548]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7770.905 187.44 7771.185 188.44 ;
    END
  END BcidMtx[548]
  PIN BcidMtx[546]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7769.785 187.44 7770.065 188.44 ;
    END
  END BcidMtx[546]
  PIN BcidMtx[626]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8811.385 187.44 8811.665 188.44 ;
    END
  END BcidMtx[626]
  PIN BcidMtx[623]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8737.465 187.44 8737.745 188.44 ;
    END
  END BcidMtx[623]
  PIN BcidMtx[619]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8734.105 187.44 8734.385 188.44 ;
    END
  END BcidMtx[619]
  PIN BcidMtx[616]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8666.905 187.44 8667.185 188.44 ;
    END
  END BcidMtx[616]
  PIN BcidMtx[610]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8588.225 187.44 8588.505 188.44 ;
    END
  END BcidMtx[610]
  PIN BcidMtx[606]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8559.385 187.44 8559.665 188.44 ;
    END
  END BcidMtx[606]
  PIN BcidMtx[603]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8480.425 187.44 8480.705 188.44 ;
    END
  END BcidMtx[603]
  PIN BcidMtx[602]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8478.745 187.44 8479.025 188.44 ;
    END
  END BcidMtx[602]
  PIN BcidMtx[596]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8413.225 187.44 8413.505 188.44 ;
    END
  END BcidMtx[596]
  PIN BcidMtx[592]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8333.145 187.44 8333.425 188.44 ;
    END
  END BcidMtx[592]
  PIN BcidMtx[589]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8330.345 187.44 8330.625 188.44 ;
    END
  END BcidMtx[589]
  PIN BcidMtx[670]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9373.625 187.44 9373.905 188.44 ;
    END
  END BcidMtx[670]
  PIN BcidMtx[667]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9370.825 187.44 9371.105 188.44 ;
    END
  END BcidMtx[667]
  PIN BcidMtx[663]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9296.345 187.44 9296.625 188.44 ;
    END
  END BcidMtx[663]
  PIN BcidMtx[662]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9294.665 187.44 9294.945 188.44 ;
    END
  END BcidMtx[662]
  PIN BcidMtx[660]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9293.545 187.44 9293.825 188.44 ;
    END
  END BcidMtx[660]
  PIN BcidMtx[659]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9227.465 187.44 9227.745 188.44 ;
    END
  END BcidMtx[659]
  PIN BcidMtx[657]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9226.345 187.44 9226.625 188.44 ;
    END
  END BcidMtx[657]
  PIN BcidMtx[654]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9223.545 187.44 9223.825 188.44 ;
    END
  END BcidMtx[654]
  PIN BcidMtx[652]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9148.225 187.44 9148.505 188.44 ;
    END
  END BcidMtx[652]
  PIN BcidMtx[648]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9119.385 187.44 9119.665 188.44 ;
    END
  END BcidMtx[648]
  PIN BcidMtx[645]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9040.425 187.44 9040.705 188.44 ;
    END
  END BcidMtx[645]
  PIN BcidMtx[642]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9037.625 187.44 9037.905 188.44 ;
    END
  END BcidMtx[642]
  PIN BcidMtx[637]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8972.665 187.44 8972.945 188.44 ;
    END
  END BcidMtx[637]
  PIN BcidMtx[632]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8890.905 187.44 8891.185 188.44 ;
    END
  END BcidMtx[632]
  PIN BcidMtx[709]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9930.825 187.44 9931.105 188.44 ;
    END
  END BcidMtx[709]
  PIN BcidMtx[707]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9857.465 187.44 9857.745 188.44 ;
    END
  END BcidMtx[707]
  PIN BcidMtx[704]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9854.665 187.44 9854.945 188.44 ;
    END
  END BcidMtx[704]
  PIN BcidMtx[702]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9853.545 187.44 9853.825 188.44 ;
    END
  END BcidMtx[702]
  PIN BcidMtx[700]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9786.905 187.44 9787.185 188.44 ;
    END
  END BcidMtx[700]
  PIN BcidMtx[694]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9708.225 187.44 9708.505 188.44 ;
    END
  END BcidMtx[694]
  PIN BcidMtx[691]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9679.945 187.44 9680.225 188.44 ;
    END
  END BcidMtx[691]
  PIN BcidMtx[686]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9598.745 187.44 9599.025 188.44 ;
    END
  END BcidMtx[686]
  PIN BcidMtx[684]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9597.625 187.44 9597.905 188.44 ;
    END
  END BcidMtx[684]
  PIN BcidMtx[682]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9535.465 187.44 9535.745 188.44 ;
    END
  END BcidMtx[682]
  PIN BcidMtx[679]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9532.665 187.44 9532.945 188.44 ;
    END
  END BcidMtx[679]
  PIN BcidMtx[675]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9452.585 187.44 9452.865 188.44 ;
    END
  END BcidMtx[675]
  PIN BcidMtx[674]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9450.905 187.44 9451.185 188.44 ;
    END
  END BcidMtx[674]
  PIN BcidMtx[672]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9449.785 187.44 9450.065 188.44 ;
    END
  END BcidMtx[672]
  PIN BcidMtx[751]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10490.825 187.44 10491.105 188.44 ;
    END
  END BcidMtx[751]
  PIN BcidMtx[745]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10414.105 187.44 10414.385 188.44 ;
    END
  END BcidMtx[745]
  PIN BcidMtx[742]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10346.905 187.44 10347.185 188.44 ;
    END
  END BcidMtx[742]
  PIN BcidMtx[740]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10344.665 187.44 10344.945 188.44 ;
    END
  END BcidMtx[740]
  PIN BcidMtx[736]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10268.225 187.44 10268.505 188.44 ;
    END
  END BcidMtx[736]
  PIN BcidMtx[729]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10160.425 187.44 10160.705 188.44 ;
    END
  END BcidMtx[729]
  PIN BcidMtx[723]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10094.905 187.44 10095.185 188.44 ;
    END
  END BcidMtx[723]
  PIN BcidMtx[718]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10013.145 187.44 10013.425 188.44 ;
    END
  END BcidMtx[718]
  PIN BcidMtx[714]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10009.785 187.44 10010.065 188.44 ;
    END
  END BcidMtx[714]
  PIN BcidMtx[795]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11053.065 187.44 11053.345 188.44 ;
    END
  END BcidMtx[795]
  PIN BcidMtx[790]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10976.905 187.44 10977.185 188.44 ;
    END
  END BcidMtx[790]
  PIN BcidMtx[787]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10974.105 187.44 10974.385 188.44 ;
    END
  END BcidMtx[787]
  PIN BcidMtx[781]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10904.105 187.44 10904.385 188.44 ;
    END
  END BcidMtx[781]
  PIN BcidMtx[778]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10828.225 187.44 10828.505 188.44 ;
    END
  END BcidMtx[778]
  PIN BcidMtx[775]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10799.945 187.44 10800.225 188.44 ;
    END
  END BcidMtx[775]
  PIN BcidMtx[771]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10720.425 187.44 10720.705 188.44 ;
    END
  END BcidMtx[771]
  PIN BcidMtx[1325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18108.785 187.44 18109.065 188.44 ;
    END
  END BcidMtx[1325]
  PIN BcidMtx[765]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10654.905 187.44 10655.185 188.44 ;
    END
  END BcidMtx[765]
  PIN BcidMtx[761]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10573.705 187.44 10573.985 188.44 ;
    END
  END BcidMtx[761]
  PIN BcidMtx[757]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10570.345 187.44 10570.625 188.44 ;
    END
  END BcidMtx[757]
  PIN BcidMtx[839]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11614.185 187.44 11614.465 188.44 ;
    END
  END BcidMtx[839]
  PIN BcidMtx[835]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11610.825 187.44 11611.105 188.44 ;
    END
  END BcidMtx[835]
  PIN BcidMtx[833]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11537.465 187.44 11537.745 188.44 ;
    END
  END BcidMtx[833]
  PIN BcidMtx[832]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11536.905 187.44 11537.185 188.44 ;
    END
  END BcidMtx[832]
  PIN BcidMtx[826]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11466.905 187.44 11467.185 188.44 ;
    END
  END BcidMtx[826]
  PIN BcidMtx[823]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11464.105 187.44 11464.385 188.44 ;
    END
  END BcidMtx[823]
  PIN BcidMtx[819]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11387.665 187.44 11387.945 188.44 ;
    END
  END BcidMtx[819]
  PIN BcidMtx[818]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11360.505 187.44 11360.785 188.44 ;
    END
  END BcidMtx[818]
  PIN BcidMtx[814]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11280.985 187.44 11281.265 188.44 ;
    END
  END BcidMtx[814]
  PIN BcidMtx[812]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11278.745 187.44 11279.025 188.44 ;
    END
  END BcidMtx[812]
  PIN BcidMtx[810]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11277.625 187.44 11277.905 188.44 ;
    END
  END BcidMtx[810]
  PIN BcidMtx[808]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11215.465 187.44 11215.745 188.44 ;
    END
  END BcidMtx[808]
  PIN BcidMtx[1320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18079.385 187.44 18079.665 188.44 ;
    END
  END BcidMtx[1320]
  PIN BcidMtx[805]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11212.665 187.44 11212.945 188.44 ;
    END
  END BcidMtx[805]
  PIN BcidMtx[803]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11133.705 187.44 11133.985 188.44 ;
    END
  END BcidMtx[803]
  PIN BcidMtx[800]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11130.905 187.44 11131.185 188.44 ;
    END
  END BcidMtx[800]
  PIN BcidMtx[881]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12174.185 187.44 12174.465 188.44 ;
    END
  END BcidMtx[881]
  PIN BcidMtx[875]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12097.465 187.44 12097.745 188.44 ;
    END
  END BcidMtx[875]
  PIN BcidMtx[873]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12096.345 187.44 12096.625 188.44 ;
    END
  END BcidMtx[873]
  PIN BcidMtx[868]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12026.905 187.44 12027.185 188.44 ;
    END
  END BcidMtx[868]
  PIN BcidMtx[861]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11947.665 187.44 11947.945 188.44 ;
    END
  END BcidMtx[861]
  PIN BcidMtx[859]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11919.945 187.44 11920.225 188.44 ;
    END
  END BcidMtx[859]
  PIN BcidMtx[856]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11840.985 187.44 11841.265 188.44 ;
    END
  END BcidMtx[856]
  PIN BcidMtx[852]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11837.625 187.44 11837.905 188.44 ;
    END
  END BcidMtx[852]
  PIN BcidMtx[849]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11774.905 187.44 11775.185 188.44 ;
    END
  END BcidMtx[849]
  PIN BcidMtx[848]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11773.225 187.44 11773.505 188.44 ;
    END
  END BcidMtx[848]
  PIN BcidMtx[845]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11693.705 187.44 11693.985 188.44 ;
    END
  END BcidMtx[845]
  PIN BcidMtx[843]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11692.585 187.44 11692.865 188.44 ;
    END
  END BcidMtx[843]
  PIN BcidMtx[841]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11690.345 187.44 11690.625 188.44 ;
    END
  END BcidMtx[841]
  PIN BcidMtx[923]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12734.185 187.44 12734.465 188.44 ;
    END
  END BcidMtx[923]
  PIN BcidMtx[921]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12733.065 187.44 12733.345 188.44 ;
    END
  END BcidMtx[921]
  PIN BcidMtx[919]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12730.825 187.44 12731.105 188.44 ;
    END
  END BcidMtx[919]
  PIN BcidMtx[915]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12656.345 187.44 12656.625 188.44 ;
    END
  END BcidMtx[915]
  PIN BcidMtx[910]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12586.905 187.44 12587.185 188.44 ;
    END
  END BcidMtx[910]
  PIN BcidMtx[906]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12583.545 187.44 12583.825 188.44 ;
    END
  END BcidMtx[906]
  PIN BcidMtx[904]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12508.225 187.44 12508.505 188.44 ;
    END
  END BcidMtx[904]
  PIN BcidMtx[902]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12480.505 187.44 12480.785 188.44 ;
    END
  END BcidMtx[902]
  PIN BcidMtx[900]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12479.385 187.44 12479.665 188.44 ;
    END
  END BcidMtx[900]
  PIN BcidMtx[898]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12400.985 187.44 12401.265 188.44 ;
    END
  END BcidMtx[898]
  PIN BcidMtx[895]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12398.185 187.44 12398.465 188.44 ;
    END
  END BcidMtx[895]
  PIN BcidMtx[893]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12336.025 187.44 12336.305 188.44 ;
    END
  END BcidMtx[893]
  PIN BcidMtx[890]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12333.225 187.44 12333.505 188.44 ;
    END
  END BcidMtx[890]
  PIN BcidMtx[885]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12252.585 187.44 12252.865 188.44 ;
    END
  END BcidMtx[885]
  PIN BcidMtx[884]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12250.905 187.44 12251.185 188.44 ;
    END
  END BcidMtx[884]
  PIN BcidMtx[882]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12249.785 187.44 12250.065 188.44 ;
    END
  END BcidMtx[882]
  PIN BcidMtx[963]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13293.065 187.44 13293.345 188.44 ;
    END
  END BcidMtx[963]
  PIN BcidMtx[962]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13291.385 187.44 13291.665 188.44 ;
    END
  END BcidMtx[962]
  PIN BcidMtx[960]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13290.265 187.44 13290.545 188.44 ;
    END
  END BcidMtx[960]
  PIN BcidMtx[959]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13217.465 187.44 13217.745 188.44 ;
    END
  END BcidMtx[959]
  PIN BcidMtx[954]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13213.545 187.44 13213.825 188.44 ;
    END
  END BcidMtx[954]
  PIN BcidMtx[953]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13147.465 187.44 13147.745 188.44 ;
    END
  END BcidMtx[953]
  PIN BcidMtx[951]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13146.345 187.44 13146.625 188.44 ;
    END
  END BcidMtx[951]
  PIN BcidMtx[949]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13144.105 187.44 13144.385 188.44 ;
    END
  END BcidMtx[949]
  PIN BcidMtx[945]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13067.665 187.44 13067.945 188.44 ;
    END
  END BcidMtx[945]
  PIN BcidMtx[944]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13040.505 187.44 13040.785 188.44 ;
    END
  END BcidMtx[944]
  PIN BcidMtx[941]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12961.545 187.44 12961.825 188.44 ;
    END
  END BcidMtx[941]
  PIN BcidMtx[938]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12958.745 187.44 12959.025 188.44 ;
    END
  END BcidMtx[938]
  PIN BcidMtx[935]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12896.025 187.44 12896.305 188.44 ;
    END
  END BcidMtx[935]
  PIN BcidMtx[932]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12893.225 187.44 12893.505 188.44 ;
    END
  END BcidMtx[932]
  PIN BcidMtx[928]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12813.145 187.44 12813.425 188.44 ;
    END
  END BcidMtx[928]
  PIN BcidMtx[926]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12810.905 187.44 12811.185 188.44 ;
    END
  END BcidMtx[926]
  PIN BcidMtx[924]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12809.785 187.44 12810.065 188.44 ;
    END
  END BcidMtx[924]
  PIN BcidMtx[1005]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13853.065 187.44 13853.345 188.44 ;
    END
  END BcidMtx[1005]
  PIN BcidMtx[1004]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13851.385 187.44 13851.665 188.44 ;
    END
  END BcidMtx[1004]
  PIN BcidMtx[1001]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13777.465 187.44 13777.745 188.44 ;
    END
  END BcidMtx[1001]
  PIN BcidMtx[996]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13773.545 187.44 13773.825 188.44 ;
    END
  END BcidMtx[996]
  PIN BcidMtx[995]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13707.465 187.44 13707.745 188.44 ;
    END
  END BcidMtx[995]
  PIN BcidMtx[993]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13706.345 187.44 13706.625 188.44 ;
    END
  END BcidMtx[993]
  PIN BcidMtx[992]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13704.665 187.44 13704.945 188.44 ;
    END
  END BcidMtx[992]
  PIN BcidMtx[987]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13627.665 187.44 13627.945 188.44 ;
    END
  END BcidMtx[987]
  PIN BcidMtx[986]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13600.505 187.44 13600.785 188.44 ;
    END
  END BcidMtx[986]
  PIN BcidMtx[983]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13521.545 187.44 13521.825 188.44 ;
    END
  END BcidMtx[983]
  PIN BcidMtx[979]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13518.185 187.44 13518.465 188.44 ;
    END
  END BcidMtx[979]
  PIN BcidMtx[976]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13455.465 187.44 13455.745 188.44 ;
    END
  END BcidMtx[976]
  PIN BcidMtx[974]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13453.225 187.44 13453.505 188.44 ;
    END
  END BcidMtx[974]
  PIN BcidMtx[972]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13452.105 187.44 13452.385 188.44 ;
    END
  END BcidMtx[972]
  PIN BcidMtx[969]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13372.585 187.44 13372.865 188.44 ;
    END
  END BcidMtx[969]
  PIN BcidMtx[966]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13369.785 187.44 13370.065 188.44 ;
    END
  END BcidMtx[966]
  PIN BcidMtx[1048]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14413.625 187.44 14413.905 188.44 ;
    END
  END BcidMtx[1048]
  PIN BcidMtx[1041]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14336.345 187.44 14336.625 188.44 ;
    END
  END BcidMtx[1041]
  PIN BcidMtx[1038]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14333.545 187.44 14333.825 188.44 ;
    END
  END BcidMtx[1038]
  PIN BcidMtx[1037]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14267.465 187.44 14267.745 188.44 ;
    END
  END BcidMtx[1037]
  PIN BcidMtx[1033]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14264.105 187.44 14264.385 188.44 ;
    END
  END BcidMtx[1033]
  PIN BcidMtx[1030]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14188.225 187.44 14188.505 188.44 ;
    END
  END BcidMtx[1030]
  PIN BcidMtx[1027]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14159.945 187.44 14160.225 188.44 ;
    END
  END BcidMtx[1027]
  PIN BcidMtx[1024]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14080.985 187.44 14081.265 188.44 ;
    END
  END BcidMtx[1024]
  PIN BcidMtx[1020]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14077.625 187.44 14077.905 188.44 ;
    END
  END BcidMtx[1020]
  PIN BcidMtx[1018]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14015.465 187.44 14015.745 188.44 ;
    END
  END BcidMtx[1018]
  PIN BcidMtx[1015]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14012.665 187.44 14012.945 188.44 ;
    END
  END BcidMtx[1015]
  PIN BcidMtx[1011]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13932.585 187.44 13932.865 188.44 ;
    END
  END BcidMtx[1011]
  PIN BcidMtx[1010]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13930.905 187.44 13931.185 188.44 ;
    END
  END BcidMtx[1010]
  PIN BcidMtx[1088]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14971.385 187.44 14971.665 188.44 ;
    END
  END BcidMtx[1088]
  PIN BcidMtx[1084]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14896.905 187.44 14897.185 188.44 ;
    END
  END BcidMtx[1084]
  PIN BcidMtx[1081]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14894.105 187.44 14894.385 188.44 ;
    END
  END BcidMtx[1081]
  PIN BcidMtx[1078]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14826.905 187.44 14827.185 188.44 ;
    END
  END BcidMtx[1078]
  PIN BcidMtx[1073]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14748.785 187.44 14749.065 188.44 ;
    END
  END BcidMtx[1073]
  PIN BcidMtx[1069]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14719.945 187.44 14720.225 188.44 ;
    END
  END BcidMtx[1069]
  PIN BcidMtx[1067]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14641.545 187.44 14641.825 188.44 ;
    END
  END BcidMtx[1067]
  PIN BcidMtx[1064]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14638.745 187.44 14639.025 188.44 ;
    END
  END BcidMtx[1064]
  PIN BcidMtx[1061]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14576.025 187.44 14576.305 188.44 ;
    END
  END BcidMtx[1061]
  PIN BcidMtx[1059]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14574.905 187.44 14575.185 188.44 ;
    END
  END BcidMtx[1059]
  PIN BcidMtx[1058]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14573.225 187.44 14573.505 188.44 ;
    END
  END BcidMtx[1058]
  PIN BcidMtx[1053]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14492.585 187.44 14492.865 188.44 ;
    END
  END BcidMtx[1053]
  PIN BcidMtx[1050]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14489.785 187.44 14490.065 188.44 ;
    END
  END BcidMtx[1050]
  PIN BcidMtx[1132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15533.625 187.44 15533.905 188.44 ;
    END
  END BcidMtx[1132]
  PIN BcidMtx[1128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15530.265 187.44 15530.545 188.44 ;
    END
  END BcidMtx[1128]
  PIN BcidMtx[1127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15457.465 187.44 15457.745 188.44 ;
    END
  END BcidMtx[1127]
  PIN BcidMtx[1124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15454.665 187.44 15454.945 188.44 ;
    END
  END BcidMtx[1124]
  PIN BcidMtx[1119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15386.345 187.44 15386.625 188.44 ;
    END
  END BcidMtx[1119]
  PIN BcidMtx[1118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15384.665 187.44 15384.945 188.44 ;
    END
  END BcidMtx[1118]
  PIN BcidMtx[1114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15308.225 187.44 15308.505 188.44 ;
    END
  END BcidMtx[1114]
  PIN BcidMtx[1112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15280.505 187.44 15280.785 188.44 ;
    END
  END BcidMtx[1112]
  PIN BcidMtx[1110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15279.385 187.44 15279.665 188.44 ;
    END
  END BcidMtx[1110]
  PIN BcidMtx[1109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15201.545 187.44 15201.825 188.44 ;
    END
  END BcidMtx[1109]
  PIN BcidMtx[1105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15198.185 187.44 15198.465 188.44 ;
    END
  END BcidMtx[1105]
  PIN BcidMtx[1102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15135.465 187.44 15135.745 188.44 ;
    END
  END BcidMtx[1102]
  PIN BcidMtx[1098]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15132.105 187.44 15132.385 188.44 ;
    END
  END BcidMtx[1098]
  PIN BcidMtx[1097]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15053.705 187.44 15053.985 188.44 ;
    END
  END BcidMtx[1097]
  PIN BcidMtx[1095]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15052.585 187.44 15052.865 188.44 ;
    END
  END BcidMtx[1095]
  PIN BcidMtx[1094]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15050.905 187.44 15051.185 188.44 ;
    END
  END BcidMtx[1094]
  PIN BcidMtx[1175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16094.185 187.44 16094.465 188.44 ;
    END
  END BcidMtx[1175]
  PIN BcidMtx[1173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16093.065 187.44 16093.345 188.44 ;
    END
  END BcidMtx[1173]
  PIN BcidMtx[1168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16016.905 187.44 16017.185 188.44 ;
    END
  END BcidMtx[1168]
  PIN BcidMtx[1165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16014.105 187.44 16014.385 188.44 ;
    END
  END BcidMtx[1165]
  PIN BcidMtx[1310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17933.225 187.44 17933.505 188.44 ;
    END
  END BcidMtx[1310]
  PIN BcidMtx[1162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15946.905 187.44 15947.185 188.44 ;
    END
  END BcidMtx[1162]
  PIN BcidMtx[1160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15944.665 187.44 15944.945 188.44 ;
    END
  END BcidMtx[1160]
  PIN BcidMtx[1308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17932.105 187.44 17932.385 188.44 ;
    END
  END BcidMtx[1308]
  PIN BcidMtx[1156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15868.225 187.44 15868.505 188.44 ;
    END
  END BcidMtx[1156]
  PIN BcidMtx[1153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15839.945 187.44 15840.225 188.44 ;
    END
  END BcidMtx[1153]
  PIN BcidMtx[1148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15758.745 187.44 15759.025 188.44 ;
    END
  END BcidMtx[1148]
  PIN BcidMtx[1146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15757.625 187.44 15757.905 188.44 ;
    END
  END BcidMtx[1146]
  PIN BcidMtx[1145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15696.025 187.44 15696.305 188.44 ;
    END
  END BcidMtx[1145]
  PIN BcidMtx[1142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15693.225 187.44 15693.505 188.44 ;
    END
  END BcidMtx[1142]
  PIN BcidMtx[1140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15692.105 187.44 15692.385 188.44 ;
    END
  END BcidMtx[1140]
  PIN BcidMtx[1138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15613.145 187.44 15613.425 188.44 ;
    END
  END BcidMtx[1138]
  PIN BcidMtx[1135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15610.345 187.44 15610.625 188.44 ;
    END
  END BcidMtx[1135]
  PIN BcidMtx[1217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16654.185 187.44 16654.465 188.44 ;
    END
  END BcidMtx[1217]
  PIN BcidMtx[1215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16653.065 187.44 16653.345 188.44 ;
    END
  END BcidMtx[1215]
  PIN BcidMtx[1213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16650.825 187.44 16651.105 188.44 ;
    END
  END BcidMtx[1213]
  PIN BcidMtx[1211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16577.465 187.44 16577.745 188.44 ;
    END
  END BcidMtx[1211]
  PIN BcidMtx[1208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16574.665 187.44 16574.945 188.44 ;
    END
  END BcidMtx[1208]
  PIN BcidMtx[1204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16506.905 187.44 16507.185 188.44 ;
    END
  END BcidMtx[1204]
  PIN BcidMtx[1201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16504.105 187.44 16504.385 188.44 ;
    END
  END BcidMtx[1201]
  PIN BcidMtx[1194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16399.385 187.44 16399.665 188.44 ;
    END
  END BcidMtx[1194]
  PIN BcidMtx[1193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16321.545 187.44 16321.825 188.44 ;
    END
  END BcidMtx[1193]
  PIN BcidMtx[1188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16317.625 187.44 16317.905 188.44 ;
    END
  END BcidMtx[1188]
  PIN BcidMtx[1186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16255.465 187.44 16255.745 188.44 ;
    END
  END BcidMtx[1186]
  PIN BcidMtx[1184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16253.225 187.44 16253.505 188.44 ;
    END
  END BcidMtx[1184]
  PIN BcidMtx[1181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16173.705 187.44 16173.985 188.44 ;
    END
  END BcidMtx[1181]
  PIN BcidMtx[1179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16172.585 187.44 16172.865 188.44 ;
    END
  END BcidMtx[1179]
  PIN BcidMtx[1177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16170.345 187.44 16170.625 188.44 ;
    END
  END BcidMtx[1177]
  PIN BcidMtx[1259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17214.185 187.44 17214.465 188.44 ;
    END
  END BcidMtx[1259]
  PIN BcidMtx[1257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17213.065 187.44 17213.345 188.44 ;
    END
  END BcidMtx[1257]
  PIN BcidMtx[1255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17210.825 187.44 17211.105 188.44 ;
    END
  END BcidMtx[1255]
  PIN BcidMtx[1251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17136.345 187.44 17136.625 188.44 ;
    END
  END BcidMtx[1251]
  PIN BcidMtx[1247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17067.465 187.44 17067.745 188.44 ;
    END
  END BcidMtx[1247]
  PIN BcidMtx[1244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17064.665 187.44 17064.945 188.44 ;
    END
  END BcidMtx[1244]
  PIN BcidMtx[1241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16988.785 187.44 16989.065 188.44 ;
    END
  END BcidMtx[1241]
  PIN BcidMtx[1237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16959.945 187.44 16960.225 188.44 ;
    END
  END BcidMtx[1237]
  PIN BcidMtx[1235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16881.545 187.44 16881.825 188.44 ;
    END
  END BcidMtx[1235]
  PIN BcidMtx[1232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16878.745 187.44 16879.025 188.44 ;
    END
  END BcidMtx[1232]
  PIN BcidMtx[1227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16814.905 187.44 16815.185 188.44 ;
    END
  END BcidMtx[1227]
  PIN BcidMtx[1226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16813.225 187.44 16813.505 188.44 ;
    END
  END BcidMtx[1226]
  PIN BcidMtx[1224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16812.105 187.44 16812.385 188.44 ;
    END
  END BcidMtx[1224]
  PIN BcidMtx[1223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16733.705 187.44 16733.985 188.44 ;
    END
  END BcidMtx[1223]
  PIN BcidMtx[1218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16729.785 187.44 16730.065 188.44 ;
    END
  END BcidMtx[1218]
  PIN BcidMtx[1299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17773.065 187.44 17773.345 188.44 ;
    END
  END BcidMtx[1299]
  PIN BcidMtx[1298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17771.385 187.44 17771.665 188.44 ;
    END
  END BcidMtx[1298]
  PIN BcidMtx[1294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17696.905 187.44 17697.185 188.44 ;
    END
  END BcidMtx[1294]
  PIN BcidMtx[1290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17693.545 187.44 17693.825 188.44 ;
    END
  END BcidMtx[1290]
  PIN BcidMtx[1288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17626.905 187.44 17627.185 188.44 ;
    END
  END BcidMtx[1288]
  PIN BcidMtx[1283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17548.785 187.44 17549.065 188.44 ;
    END
  END BcidMtx[1283]
  PIN BcidMtx[1282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17548.225 187.44 17548.505 188.44 ;
    END
  END BcidMtx[1282]
  PIN BcidMtx[1280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17520.505 187.44 17520.785 188.44 ;
    END
  END BcidMtx[1280]
  PIN BcidMtx[1275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17440.425 187.44 17440.705 188.44 ;
    END
  END BcidMtx[1275]
  PIN BcidMtx[1272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17437.625 187.44 17437.905 188.44 ;
    END
  END BcidMtx[1272]
  PIN BcidMtx[1268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17373.225 187.44 17373.505 188.44 ;
    END
  END BcidMtx[1268]
  PIN BcidMtx[1265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17293.705 187.44 17293.985 188.44 ;
    END
  END BcidMtx[1265]
  PIN BcidMtx[1260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17289.785 187.44 17290.065 188.44 ;
    END
  END BcidMtx[1260]
  PIN BcidMtx[1341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18333.065 187.44 18333.345 188.44 ;
    END
  END BcidMtx[1341]
  PIN BcidMtx[1339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18330.825 187.44 18331.105 188.44 ;
    END
  END BcidMtx[1339]
  PIN BcidMtx[1337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18257.465 187.44 18257.745 188.44 ;
    END
  END BcidMtx[1337]
  PIN BcidMtx[1332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18253.545 187.44 18253.825 188.44 ;
    END
  END BcidMtx[1332]
  PIN BcidMtx[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 974.185 187.44 974.465 188.44 ;
    END
  END BcidMtx[41]
  PIN BcidMtx[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 970.825 187.44 971.105 188.44 ;
    END
  END BcidMtx[37]
  PIN BcidMtx[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 896.905 187.44 897.185 188.44 ;
    END
  END BcidMtx[34]
  PIN BcidMtx[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 893.545 187.44 893.825 188.44 ;
    END
  END BcidMtx[30]
  PIN BcidMtx[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 826.345 187.44 826.625 188.44 ;
    END
  END BcidMtx[27]
  PIN BcidMtx[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 824.665 187.44 824.945 188.44 ;
    END
  END BcidMtx[26]
  PIN BcidMtx[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 747.665 187.44 747.945 188.44 ;
    END
  END BcidMtx[21]
  PIN BcidMtx[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 719.945 187.44 720.225 188.44 ;
    END
  END BcidMtx[19]
  PIN BcidMtx[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 640.985 187.44 641.265 188.44 ;
    END
  END BcidMtx[16]
  PIN BcidMtx[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 637.625 187.44 637.905 188.44 ;
    END
  END BcidMtx[12]
  PIN BcidMtx[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 576.025 187.44 576.305 188.44 ;
    END
  END BcidMtx[11]
  PIN BcidMtx[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 573.225 187.44 573.505 188.44 ;
    END
  END BcidMtx[8]
  PIN BcidMtx[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1534.185 187.44 1534.465 188.44 ;
    END
  END BcidMtx[83]
  PIN BcidMtx[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1457.465 187.44 1457.745 188.44 ;
    END
  END BcidMtx[77]
  PIN BcidMtx[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1386.905 187.44 1387.185 188.44 ;
    END
  END BcidMtx[70]
  PIN BcidMtx[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1384.105 187.44 1384.385 188.44 ;
    END
  END BcidMtx[67]
  PIN BcidMtx[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1279.385 187.44 1279.665 188.44 ;
    END
  END BcidMtx[60]
  PIN BcidMtx[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1200.425 187.44 1200.705 188.44 ;
    END
  END BcidMtx[57]
  PIN BcidMtx[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1198.185 187.44 1198.465 188.44 ;
    END
  END BcidMtx[55]
  PIN BcidMtx[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1134.905 187.44 1135.185 188.44 ;
    END
  END BcidMtx[51]
  PIN BcidMtx[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1132.665 187.44 1132.945 188.44 ;
    END
  END BcidMtx[49]
  PIN BcidMtx[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1053.145 187.44 1053.425 188.44 ;
    END
  END BcidMtx[46]
  PIN BcidMtx[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1049.785 187.44 1050.065 188.44 ;
    END
  END BcidMtx[42]
  PIN BcidMtx[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2093.625 187.44 2093.905 188.44 ;
    END
  END BcidMtx[124]
  PIN BcidMtx[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2090.265 187.44 2090.545 188.44 ;
    END
  END BcidMtx[120]
  PIN BcidMtx[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2016.345 187.44 2016.625 188.44 ;
    END
  END BcidMtx[117]
  PIN BcidMtx[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2014.665 187.44 2014.945 188.44 ;
    END
  END BcidMtx[116]
  PIN BcidMtx[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1946.905 187.44 1947.185 188.44 ;
    END
  END BcidMtx[112]
  PIN BcidMtx[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1944.105 187.44 1944.385 188.44 ;
    END
  END BcidMtx[109]
  PIN BcidMtx[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1868.785 187.44 1869.065 188.44 ;
    END
  END BcidMtx[107]
  PIN BcidMtx[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1840.505 187.44 1840.785 188.44 ;
    END
  END BcidMtx[104]
  PIN BcidMtx[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1839.385 187.44 1839.665 188.44 ;
    END
  END BcidMtx[102]
  PIN BcidMtx[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1761.545 187.44 1761.825 188.44 ;
    END
  END BcidMtx[101]
  PIN BcidMtx[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1757.625 187.44 1757.905 188.44 ;
    END
  END BcidMtx[96]
  PIN BcidMtx[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1692.665 187.44 1692.945 188.44 ;
    END
  END BcidMtx[91]
  PIN BcidMtx[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1613.145 187.44 1613.425 188.44 ;
    END
  END BcidMtx[88]
  PIN BcidMtx[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2654.185 187.44 2654.465 188.44 ;
    END
  END BcidMtx[167]
  PIN BcidMtx[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2653.065 187.44 2653.345 188.44 ;
    END
  END BcidMtx[165]
  PIN BcidMtx[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2650.825 187.44 2651.105 188.44 ;
    END
  END BcidMtx[163]
  PIN BcidMtx[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2577.465 187.44 2577.745 188.44 ;
    END
  END BcidMtx[161]
  PIN BcidMtx[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2576.345 187.44 2576.625 188.44 ;
    END
  END BcidMtx[159]
  PIN BcidMtx[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2574.665 187.44 2574.945 188.44 ;
    END
  END BcidMtx[158]
  PIN BcidMtx[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2506.345 187.44 2506.625 188.44 ;
    END
  END BcidMtx[153]
  PIN BcidMtx[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2504.665 187.44 2504.945 188.44 ;
    END
  END BcidMtx[152]
  PIN BcidMtx[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2503.545 187.44 2503.825 188.44 ;
    END
  END BcidMtx[150]
  PIN BcidMtx[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2399.385 187.44 2399.665 188.44 ;
    END
  END BcidMtx[144]
  PIN BcidMtx[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2321.545 187.44 2321.825 188.44 ;
    END
  END BcidMtx[143]
  PIN BcidMtx[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2318.185 187.44 2318.465 188.44 ;
    END
  END BcidMtx[139]
  PIN BcidMtx[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2254.905 187.44 2255.185 188.44 ;
    END
  END BcidMtx[135]
  PIN BcidMtx[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2252.665 187.44 2252.945 188.44 ;
    END
  END BcidMtx[133]
  PIN BcidMtx[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2172.585 187.44 2172.865 188.44 ;
    END
  END BcidMtx[129]
  PIN BcidMtx[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2170.905 187.44 2171.185 188.44 ;
    END
  END BcidMtx[128]
  PIN BcidMtx[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2169.785 187.44 2170.065 188.44 ;
    END
  END BcidMtx[126]
  PIN BcidMtx[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3213.065 187.44 3213.345 188.44 ;
    END
  END BcidMtx[207]
  PIN BcidMtx[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3211.385 187.44 3211.665 188.44 ;
    END
  END BcidMtx[206]
  PIN BcidMtx[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3210.265 187.44 3210.545 188.44 ;
    END
  END BcidMtx[204]
  PIN BcidMtx[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3137.465 187.44 3137.745 188.44 ;
    END
  END BcidMtx[203]
  PIN BcidMtx[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3134.665 187.44 3134.945 188.44 ;
    END
  END BcidMtx[200]
  PIN BcidMtx[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3067.465 187.44 3067.745 188.44 ;
    END
  END BcidMtx[197]
  PIN BcidMtx[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3064.665 187.44 3064.945 188.44 ;
    END
  END BcidMtx[194]
  PIN BcidMtx[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2988.225 187.44 2988.505 188.44 ;
    END
  END BcidMtx[190]
  PIN BcidMtx[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2960.505 187.44 2960.785 188.44 ;
    END
  END BcidMtx[188]
  PIN BcidMtx[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2959.385 187.44 2959.665 188.44 ;
    END
  END BcidMtx[186]
  PIN BcidMtx[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2878.185 187.44 2878.465 188.44 ;
    END
  END BcidMtx[181]
  PIN BcidMtx[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2816.025 187.44 2816.305 188.44 ;
    END
  END BcidMtx[179]
  PIN BcidMtx[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2813.225 187.44 2813.505 188.44 ;
    END
  END BcidMtx[176]
  PIN BcidMtx[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2733.705 187.44 2733.985 188.44 ;
    END
  END BcidMtx[173]
  PIN BcidMtx[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2732.585 187.44 2732.865 188.44 ;
    END
  END BcidMtx[171]
  PIN BcidMtx[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2730.345 187.44 2730.625 188.44 ;
    END
  END BcidMtx[169]
  PIN BcidMtx[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3774.185 187.44 3774.465 188.44 ;
    END
  END BcidMtx[251]
  PIN BcidMtx[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3773.065 187.44 3773.345 188.44 ;
    END
  END BcidMtx[249]
  PIN BcidMtx[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3770.825 187.44 3771.105 188.44 ;
    END
  END BcidMtx[247]
  PIN BcidMtx[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3696.905 187.44 3697.185 188.44 ;
    END
  END BcidMtx[244]
  PIN BcidMtx[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3626.345 187.44 3626.625 188.44 ;
    END
  END BcidMtx[237]
  PIN BcidMtx[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3624.665 187.44 3624.945 188.44 ;
    END
  END BcidMtx[236]
  PIN BcidMtx[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3548.785 187.44 3549.065 188.44 ;
    END
  END BcidMtx[233]
  PIN BcidMtx[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3519.385 187.44 3519.665 188.44 ;
    END
  END BcidMtx[228]
  PIN BcidMtx[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3440.425 187.44 3440.705 188.44 ;
    END
  END BcidMtx[225]
  PIN BcidMtx[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3438.745 187.44 3439.025 188.44 ;
    END
  END BcidMtx[224]
  PIN BcidMtx[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3437.625 187.44 3437.905 188.44 ;
    END
  END BcidMtx[222]
  PIN BcidMtx[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3374.905 187.44 3375.185 188.44 ;
    END
  END BcidMtx[219]
  PIN BcidMtx[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3373.225 187.44 3373.505 188.44 ;
    END
  END BcidMtx[218]
  PIN BcidMtx[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3293.145 187.44 3293.425 188.44 ;
    END
  END BcidMtx[214]
  PIN BcidMtx[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4333.065 187.44 4333.345 188.44 ;
    END
  END BcidMtx[291]
  PIN BcidMtx[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4331.385 187.44 4331.665 188.44 ;
    END
  END BcidMtx[290]
  PIN BcidMtx[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4256.345 187.44 4256.625 188.44 ;
    END
  END BcidMtx[285]
  PIN BcidMtx[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4254.665 187.44 4254.945 188.44 ;
    END
  END BcidMtx[284]
  PIN BcidMtx[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4253.545 187.44 4253.825 188.44 ;
    END
  END BcidMtx[282]
  PIN BcidMtx[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4187.465 187.44 4187.745 188.44 ;
    END
  END BcidMtx[281]
  PIN BcidMtx[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4183.545 187.44 4183.825 188.44 ;
    END
  END BcidMtx[276]
  PIN BcidMtx[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4108.225 187.44 4108.505 188.44 ;
    END
  END BcidMtx[274]
  PIN BcidMtx[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4079.945 187.44 4080.225 188.44 ;
    END
  END BcidMtx[271]
  PIN BcidMtx[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4000.425 187.44 4000.705 188.44 ;
    END
  END BcidMtx[267]
  PIN BcidMtx[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3935.465 187.44 3935.745 188.44 ;
    END
  END BcidMtx[262]
  PIN BcidMtx[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3932.665 187.44 3932.945 188.44 ;
    END
  END BcidMtx[259]
  PIN BcidMtx[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3853.145 187.44 3853.425 188.44 ;
    END
  END BcidMtx[256]
  PIN BcidMtx[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3850.905 187.44 3851.185 188.44 ;
    END
  END BcidMtx[254]
  PIN BcidMtx[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4894.185 187.44 4894.465 188.44 ;
    END
  END BcidMtx[335]
  PIN BcidMtx[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4891.385 187.44 4891.665 188.44 ;
    END
  END BcidMtx[332]
  PIN BcidMtx[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4816.345 187.44 4816.625 188.44 ;
    END
  END BcidMtx[327]
  PIN BcidMtx[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4814.665 187.44 4814.945 188.44 ;
    END
  END BcidMtx[326]
  PIN BcidMtx[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4813.545 187.44 4813.825 188.44 ;
    END
  END BcidMtx[324]
  PIN BcidMtx[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4746.345 187.44 4746.625 188.44 ;
    END
  END BcidMtx[321]
  PIN BcidMtx[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4744.665 187.44 4744.945 188.44 ;
    END
  END BcidMtx[320]
  PIN BcidMtx[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4743.545 187.44 4743.825 188.44 ;
    END
  END BcidMtx[318]
  PIN BcidMtx[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4668.785 187.44 4669.065 188.44 ;
    END
  END BcidMtx[317]
  PIN BcidMtx[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4640.505 187.44 4640.785 188.44 ;
    END
  END BcidMtx[314]
  PIN BcidMtx[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4560.985 187.44 4561.265 188.44 ;
    END
  END BcidMtx[310]
  PIN BcidMtx[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4558.745 187.44 4559.025 188.44 ;
    END
  END BcidMtx[308]
  PIN BcidMtx[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4495.465 187.44 4495.745 188.44 ;
    END
  END BcidMtx[304]
  PIN BcidMtx[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4492.105 187.44 4492.385 188.44 ;
    END
  END BcidMtx[300]
  PIN BcidMtx[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4413.145 187.44 4413.425 188.44 ;
    END
  END BcidMtx[298]
  PIN BcidMtx[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5454.185 187.44 5454.465 188.44 ;
    END
  END BcidMtx[377]
  PIN BcidMtx[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5451.385 187.44 5451.665 188.44 ;
    END
  END BcidMtx[374]
  PIN BcidMtx[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5376.345 187.44 5376.625 188.44 ;
    END
  END BcidMtx[369]
  PIN BcidMtx[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5374.665 187.44 5374.945 188.44 ;
    END
  END BcidMtx[368]
  PIN BcidMtx[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5374.105 187.44 5374.385 188.44 ;
    END
  END BcidMtx[367]
  PIN BcidMtx[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5304.105 187.44 5304.385 188.44 ;
    END
  END BcidMtx[361]
  PIN BcidMtx[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5303.545 187.44 5303.825 188.44 ;
    END
  END BcidMtx[360]
  PIN BcidMtx[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5228.785 187.44 5229.065 188.44 ;
    END
  END BcidMtx[359]
  PIN BcidMtx[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5199.945 187.44 5200.225 188.44 ;
    END
  END BcidMtx[355]
  PIN BcidMtx[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5121.545 187.44 5121.825 188.44 ;
    END
  END BcidMtx[353]
  PIN BcidMtx[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5118.185 187.44 5118.465 188.44 ;
    END
  END BcidMtx[349]
  PIN BcidMtx[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5056.025 187.44 5056.305 188.44 ;
    END
  END BcidMtx[347]
  PIN BcidMtx[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5052.665 187.44 5052.945 188.44 ;
    END
  END BcidMtx[343]
  PIN BcidMtx[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4973.705 187.44 4973.985 188.44 ;
    END
  END BcidMtx[341]
  PIN BcidMtx[1329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18186.345 187.44 18186.625 188.44 ;
    END
  END BcidMtx[1329]
  PIN BcidMtx[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6013.625 187.44 6013.905 188.44 ;
    END
  END BcidMtx[418]
  PIN BcidMtx[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6010.265 187.44 6010.545 188.44 ;
    END
  END BcidMtx[414]
  PIN BcidMtx[1328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18184.665 187.44 18184.945 188.44 ;
    END
  END BcidMtx[1328]
  PIN BcidMtx[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5936.345 187.44 5936.625 188.44 ;
    END
  END BcidMtx[411]
  PIN BcidMtx[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5934.665 187.44 5934.945 188.44 ;
    END
  END BcidMtx[410]
  PIN BcidMtx[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5867.465 187.44 5867.745 188.44 ;
    END
  END BcidMtx[407]
  PIN BcidMtx[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5866.905 187.44 5867.185 188.44 ;
    END
  END BcidMtx[406]
  PIN BcidMtx[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5864.105 187.44 5864.385 188.44 ;
    END
  END BcidMtx[403]
  PIN BcidMtx[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5787.665 187.44 5787.945 188.44 ;
    END
  END BcidMtx[399]
  PIN BcidMtx[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5759.945 187.44 5760.225 188.44 ;
    END
  END BcidMtx[397]
  PIN BcidMtx[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5680.425 187.44 5680.705 188.44 ;
    END
  END BcidMtx[393]
  PIN BcidMtx[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5678.745 187.44 5679.025 188.44 ;
    END
  END BcidMtx[392]
  PIN BcidMtx[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5615.465 187.44 5615.745 188.44 ;
    END
  END BcidMtx[388]
  PIN BcidMtx[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5612.105 187.44 5612.385 188.44 ;
    END
  END BcidMtx[384]
  PIN BcidMtx[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5532.585 187.44 5532.865 188.44 ;
    END
  END BcidMtx[381]
  PIN BcidMtx[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5530.905 187.44 5531.185 188.44 ;
    END
  END BcidMtx[380]
  PIN BcidMtx[460]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6573.625 187.44 6573.905 188.44 ;
    END
  END BcidMtx[460]
  PIN BcidMtx[456]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6570.265 187.44 6570.545 188.44 ;
    END
  END BcidMtx[456]
  PIN BcidMtx[455]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6497.465 187.44 6497.745 188.44 ;
    END
  END BcidMtx[455]
  PIN BcidMtx[451]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6494.105 187.44 6494.385 188.44 ;
    END
  END BcidMtx[451]
  PIN BcidMtx[448]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6426.905 187.44 6427.185 188.44 ;
    END
  END BcidMtx[448]
  PIN BcidMtx[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6423.545 187.44 6423.825 188.44 ;
    END
  END BcidMtx[444]
  PIN BcidMtx[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6348.785 187.44 6349.065 188.44 ;
    END
  END BcidMtx[443]
  PIN BcidMtx[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6319.385 187.44 6319.665 188.44 ;
    END
  END BcidMtx[438]
  PIN BcidMtx[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6241.545 187.44 6241.825 188.44 ;
    END
  END BcidMtx[437]
  PIN BcidMtx[1326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18183.545 187.44 18183.825 188.44 ;
    END
  END BcidMtx[1326]
  PIN BcidMtx[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6176.025 187.44 6176.305 188.44 ;
    END
  END BcidMtx[431]
  PIN BcidMtx[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6172.665 187.44 6172.945 188.44 ;
    END
  END BcidMtx[427]
  PIN BcidMtx[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6092.585 187.44 6092.865 188.44 ;
    END
  END BcidMtx[423]
  PIN BcidMtx[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6090.905 187.44 6091.185 188.44 ;
    END
  END BcidMtx[422]
  PIN BcidMtx[502]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7133.625 187.44 7133.905 188.44 ;
    END
  END BcidMtx[502]
  PIN BcidMtx[498]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7130.265 187.44 7130.545 188.44 ;
    END
  END BcidMtx[498]
  PIN BcidMtx[495]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7056.345 187.44 7056.625 188.44 ;
    END
  END BcidMtx[495]
  PIN BcidMtx[494]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7054.665 187.44 7054.945 188.44 ;
    END
  END BcidMtx[494]
  PIN BcidMtx[491]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6987.465 187.44 6987.745 188.44 ;
    END
  END BcidMtx[491]
  PIN BcidMtx[487]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6984.105 187.44 6984.385 188.44 ;
    END
  END BcidMtx[487]
  PIN BcidMtx[483]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6907.665 187.44 6907.945 188.44 ;
    END
  END BcidMtx[483]
  PIN BcidMtx[481]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6879.945 187.44 6880.225 188.44 ;
    END
  END BcidMtx[481]
  PIN BcidMtx[477]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6800.425 187.44 6800.705 188.44 ;
    END
  END BcidMtx[477]
  PIN BcidMtx[476]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6798.745 187.44 6799.025 188.44 ;
    END
  END BcidMtx[476]
  PIN BcidMtx[471]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6734.905 187.44 6735.185 188.44 ;
    END
  END BcidMtx[471]
  PIN BcidMtx[468]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6732.105 187.44 6732.385 188.44 ;
    END
  END BcidMtx[468]
  PIN BcidMtx[466]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6653.145 187.44 6653.425 188.44 ;
    END
  END BcidMtx[466]
  PIN BcidMtx[462]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6649.785 187.44 6650.065 188.44 ;
    END
  END BcidMtx[462]
  PIN BcidMtx[544]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7693.625 187.44 7693.905 188.44 ;
    END
  END BcidMtx[544]
  PIN BcidMtx[543]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7693.065 187.44 7693.345 188.44 ;
    END
  END BcidMtx[543]
  PIN BcidMtx[540]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7690.265 187.44 7690.545 188.44 ;
    END
  END BcidMtx[540]
  PIN BcidMtx[539]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7617.465 187.44 7617.745 188.44 ;
    END
  END BcidMtx[539]
  PIN BcidMtx[532]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7546.905 187.44 7547.185 188.44 ;
    END
  END BcidMtx[532]
  PIN BcidMtx[529]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7544.105 187.44 7544.385 188.44 ;
    END
  END BcidMtx[529]
  PIN BcidMtx[524]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7440.505 187.44 7440.785 188.44 ;
    END
  END BcidMtx[524]
  PIN BcidMtx[522]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7439.385 187.44 7439.665 188.44 ;
    END
  END BcidMtx[522]
  PIN BcidMtx[520]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7360.985 187.44 7361.265 188.44 ;
    END
  END BcidMtx[520]
  PIN BcidMtx[519]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7360.425 187.44 7360.705 188.44 ;
    END
  END BcidMtx[519]
  PIN BcidMtx[516]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7357.625 187.44 7357.905 188.44 ;
    END
  END BcidMtx[516]
  PIN BcidMtx[510]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7292.105 187.44 7292.385 188.44 ;
    END
  END BcidMtx[510]
  PIN BcidMtx[506]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7210.905 187.44 7211.185 188.44 ;
    END
  END BcidMtx[506]
  PIN BcidMtx[585]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8253.065 187.44 8253.345 188.44 ;
    END
  END BcidMtx[585]
  PIN BcidMtx[582]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8250.265 187.44 8250.545 188.44 ;
    END
  END BcidMtx[582]
  PIN BcidMtx[579]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8176.345 187.44 8176.625 188.44 ;
    END
  END BcidMtx[579]
  PIN BcidMtx[578]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8174.665 187.44 8174.945 188.44 ;
    END
  END BcidMtx[578]
  PIN BcidMtx[574]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8106.905 187.44 8107.185 188.44 ;
    END
  END BcidMtx[574]
  PIN BcidMtx[570]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8103.545 187.44 8103.825 188.44 ;
    END
  END BcidMtx[570]
  PIN BcidMtx[569]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8028.785 187.44 8029.065 188.44 ;
    END
  END BcidMtx[569]
  PIN BcidMtx[561]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7920.425 187.44 7920.705 188.44 ;
    END
  END BcidMtx[561]
  PIN BcidMtx[560]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7918.745 187.44 7919.025 188.44 ;
    END
  END BcidMtx[560]
  PIN BcidMtx[558]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7917.625 187.44 7917.905 188.44 ;
    END
  END BcidMtx[558]
  PIN BcidMtx[557]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7856.025 187.44 7856.305 188.44 ;
    END
  END BcidMtx[557]
  PIN BcidMtx[554]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7853.225 187.44 7853.505 188.44 ;
    END
  END BcidMtx[554]
  PIN BcidMtx[550]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7773.145 187.44 7773.425 188.44 ;
    END
  END BcidMtx[550]
  PIN BcidMtx[629]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8814.185 187.44 8814.465 188.44 ;
    END
  END BcidMtx[629]
  PIN BcidMtx[627]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8813.065 187.44 8813.345 188.44 ;
    END
  END BcidMtx[627]
  PIN BcidMtx[625]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8810.825 187.44 8811.105 188.44 ;
    END
  END BcidMtx[625]
  PIN BcidMtx[622]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8736.905 187.44 8737.185 188.44 ;
    END
  END BcidMtx[622]
  PIN BcidMtx[618]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8733.545 187.44 8733.825 188.44 ;
    END
  END BcidMtx[618]
  PIN BcidMtx[615]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8666.345 187.44 8666.625 188.44 ;
    END
  END BcidMtx[615]
  PIN BcidMtx[614]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8664.665 187.44 8664.945 188.44 ;
    END
  END BcidMtx[614]
  PIN BcidMtx[612]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8663.545 187.44 8663.825 188.44 ;
    END
  END BcidMtx[612]
  PIN BcidMtx[611]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8588.785 187.44 8589.065 188.44 ;
    END
  END BcidMtx[611]
  PIN BcidMtx[608]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8560.505 187.44 8560.785 188.44 ;
    END
  END BcidMtx[608]
  PIN BcidMtx[605]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8481.545 187.44 8481.825 188.44 ;
    END
  END BcidMtx[605]
  PIN BcidMtx[601]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8478.185 187.44 8478.465 188.44 ;
    END
  END BcidMtx[601]
  PIN BcidMtx[599]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8416.025 187.44 8416.305 188.44 ;
    END
  END BcidMtx[599]
  PIN BcidMtx[597]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8414.905 187.44 8415.185 188.44 ;
    END
  END BcidMtx[597]
  PIN BcidMtx[595]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8412.665 187.44 8412.945 188.44 ;
    END
  END BcidMtx[595]
  PIN BcidMtx[591]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8332.585 187.44 8332.865 188.44 ;
    END
  END BcidMtx[591]
  PIN BcidMtx[590]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8330.905 187.44 8331.185 188.44 ;
    END
  END BcidMtx[590]
  PIN BcidMtx[669]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9373.065 187.44 9373.345 188.44 ;
    END
  END BcidMtx[669]
  PIN BcidMtx[668]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9371.385 187.44 9371.665 188.44 ;
    END
  END BcidMtx[668]
  PIN BcidMtx[665]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9297.465 187.44 9297.745 188.44 ;
    END
  END BcidMtx[665]
  PIN BcidMtx[661]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9294.105 187.44 9294.385 188.44 ;
    END
  END BcidMtx[661]
  PIN BcidMtx[656]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9224.665 187.44 9224.945 188.44 ;
    END
  END BcidMtx[656]
  PIN BcidMtx[653]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9148.785 187.44 9149.065 188.44 ;
    END
  END BcidMtx[653]
  PIN BcidMtx[650]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9120.505 187.44 9120.785 188.44 ;
    END
  END BcidMtx[650]
  PIN BcidMtx[646]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9040.985 187.44 9041.265 188.44 ;
    END
  END BcidMtx[646]
  PIN BcidMtx[644]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9038.745 187.44 9039.025 188.44 ;
    END
  END BcidMtx[644]
  PIN BcidMtx[641]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8976.025 187.44 8976.305 188.44 ;
    END
  END BcidMtx[641]
  PIN BcidMtx[639]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8974.905 187.44 8975.185 188.44 ;
    END
  END BcidMtx[639]
  PIN BcidMtx[636]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8972.105 187.44 8972.385 188.44 ;
    END
  END BcidMtx[636]
  PIN BcidMtx[635]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8893.705 187.44 8893.985 188.44 ;
    END
  END BcidMtx[635]
  PIN BcidMtx[634]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8893.145 187.44 8893.425 188.44 ;
    END
  END BcidMtx[634]
  PIN BcidMtx[631]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8890.345 187.44 8890.625 188.44 ;
    END
  END BcidMtx[631]
  PIN BcidMtx[713]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9934.185 187.44 9934.465 188.44 ;
    END
  END BcidMtx[713]
  PIN BcidMtx[711]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9933.065 187.44 9933.345 188.44 ;
    END
  END BcidMtx[711]
  PIN BcidMtx[708]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9930.265 187.44 9930.545 188.44 ;
    END
  END BcidMtx[708]
  PIN BcidMtx[706]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9856.905 187.44 9857.185 188.44 ;
    END
  END BcidMtx[706]
  PIN BcidMtx[699]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9786.345 187.44 9786.625 188.44 ;
    END
  END BcidMtx[699]
  PIN BcidMtx[697]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9784.105 187.44 9784.385 188.44 ;
    END
  END BcidMtx[697]
  PIN BcidMtx[692]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9680.505 187.44 9680.785 188.44 ;
    END
  END BcidMtx[692]
  PIN BcidMtx[690]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9679.385 187.44 9679.665 188.44 ;
    END
  END BcidMtx[690]
  PIN BcidMtx[688]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9600.985 187.44 9601.265 188.44 ;
    END
  END BcidMtx[688]
  PIN BcidMtx[685]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9598.185 187.44 9598.465 188.44 ;
    END
  END BcidMtx[685]
  PIN BcidMtx[681]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9534.905 187.44 9535.185 188.44 ;
    END
  END BcidMtx[681]
  PIN BcidMtx[680]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9533.225 187.44 9533.505 188.44 ;
    END
  END BcidMtx[680]
  PIN BcidMtx[678]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9532.105 187.44 9532.385 188.44 ;
    END
  END BcidMtx[678]
  PIN BcidMtx[677]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9453.705 187.44 9453.985 188.44 ;
    END
  END BcidMtx[677]
  PIN BcidMtx[673]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9450.345 187.44 9450.625 188.44 ;
    END
  END BcidMtx[673]
  PIN BcidMtx[754]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10493.625 187.44 10493.905 188.44 ;
    END
  END BcidMtx[754]
  PIN BcidMtx[750]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10490.265 187.44 10490.545 188.44 ;
    END
  END BcidMtx[750]
  PIN BcidMtx[749]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10417.465 187.44 10417.745 188.44 ;
    END
  END BcidMtx[749]
  PIN BcidMtx[744]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10413.545 187.44 10413.825 188.44 ;
    END
  END BcidMtx[744]
  PIN BcidMtx[743]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10347.465 187.44 10347.745 188.44 ;
    END
  END BcidMtx[743]
  PIN BcidMtx[741]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10346.345 187.44 10346.625 188.44 ;
    END
  END BcidMtx[741]
  PIN BcidMtx[739]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10344.105 187.44 10344.385 188.44 ;
    END
  END BcidMtx[739]
  PIN BcidMtx[735]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10267.665 187.44 10267.945 188.44 ;
    END
  END BcidMtx[735]
  PIN BcidMtx[734]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10240.505 187.44 10240.785 188.44 ;
    END
  END BcidMtx[734]
  PIN BcidMtx[731]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10161.545 187.44 10161.825 188.44 ;
    END
  END BcidMtx[731]
  PIN BcidMtx[728]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10158.745 187.44 10159.025 188.44 ;
    END
  END BcidMtx[728]
  PIN BcidMtx[725]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10096.025 187.44 10096.305 188.44 ;
    END
  END BcidMtx[725]
  PIN BcidMtx[722]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10093.225 187.44 10093.505 188.44 ;
    END
  END BcidMtx[722]
  PIN BcidMtx[717]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10012.585 187.44 10012.865 188.44 ;
    END
  END BcidMtx[717]
  PIN BcidMtx[797]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11054.185 187.44 11054.465 188.44 ;
    END
  END BcidMtx[797]
  PIN BcidMtx[794]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11051.385 187.44 11051.665 188.44 ;
    END
  END BcidMtx[794]
  PIN BcidMtx[789]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10976.345 187.44 10976.625 188.44 ;
    END
  END BcidMtx[789]
  PIN BcidMtx[788]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10974.665 187.44 10974.945 188.44 ;
    END
  END BcidMtx[788]
  PIN BcidMtx[786]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10973.545 187.44 10973.825 188.44 ;
    END
  END BcidMtx[786]
  PIN BcidMtx[785]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10907.465 187.44 10907.745 188.44 ;
    END
  END BcidMtx[785]
  PIN BcidMtx[780]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10903.545 187.44 10903.825 188.44 ;
    END
  END BcidMtx[780]
  PIN BcidMtx[779]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10828.785 187.44 10829.065 188.44 ;
    END
  END BcidMtx[779]
  PIN BcidMtx[777]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10827.665 187.44 10827.945 188.44 ;
    END
  END BcidMtx[777]
  PIN BcidMtx[774]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10799.385 187.44 10799.665 188.44 ;
    END
  END BcidMtx[774]
  PIN BcidMtx[773]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10721.545 187.44 10721.825 188.44 ;
    END
  END BcidMtx[773]
  PIN BcidMtx[770]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10718.745 187.44 10719.025 188.44 ;
    END
  END BcidMtx[770]
  PIN BcidMtx[768]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10717.625 187.44 10717.905 188.44 ;
    END
  END BcidMtx[768]
  PIN BcidMtx[767]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10656.025 187.44 10656.305 188.44 ;
    END
  END BcidMtx[767]
  PIN BcidMtx[764]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10653.225 187.44 10653.505 188.44 ;
    END
  END BcidMtx[764]
  PIN BcidMtx[1324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18108.225 187.44 18108.505 188.44 ;
    END
  END BcidMtx[1324]
  PIN BcidMtx[760]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10573.145 187.44 10573.425 188.44 ;
    END
  END BcidMtx[760]
  PIN BcidMtx[1323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18107.665 187.44 18107.945 188.44 ;
    END
  END BcidMtx[1323]
  PIN BcidMtx[838]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11613.625 187.44 11613.905 188.44 ;
    END
  END BcidMtx[838]
  PIN BcidMtx[834]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11610.265 187.44 11610.545 188.44 ;
    END
  END BcidMtx[834]
  PIN BcidMtx[831]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11536.345 187.44 11536.625 188.44 ;
    END
  END BcidMtx[831]
  PIN BcidMtx[830]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11534.665 187.44 11534.945 188.44 ;
    END
  END BcidMtx[830]
  PIN BcidMtx[828]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11533.545 187.44 11533.825 188.44 ;
    END
  END BcidMtx[828]
  PIN BcidMtx[827]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11467.465 187.44 11467.745 188.44 ;
    END
  END BcidMtx[827]
  PIN BcidMtx[822]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11463.545 187.44 11463.825 188.44 ;
    END
  END BcidMtx[822]
  PIN BcidMtx[821]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11388.785 187.44 11389.065 188.44 ;
    END
  END BcidMtx[821]
  PIN BcidMtx[817]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11359.945 187.44 11360.225 188.44 ;
    END
  END BcidMtx[817]
  PIN BcidMtx[1321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18079.945 187.44 18080.225 188.44 ;
    END
  END BcidMtx[1321]
  PIN BcidMtx[813]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11280.425 187.44 11280.705 188.44 ;
    END
  END BcidMtx[813]
  PIN BcidMtx[809]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11216.025 187.44 11216.305 188.44 ;
    END
  END BcidMtx[809]
  PIN BcidMtx[807]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11214.905 187.44 11215.185 188.44 ;
    END
  END BcidMtx[807]
  PIN BcidMtx[806]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11213.225 187.44 11213.505 188.44 ;
    END
  END BcidMtx[806]
  PIN BcidMtx[804]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11212.105 187.44 11212.385 188.44 ;
    END
  END BcidMtx[804]
  PIN BcidMtx[802]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11133.145 187.44 11133.425 188.44 ;
    END
  END BcidMtx[802]
  PIN BcidMtx[799]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11130.345 187.44 11130.625 188.44 ;
    END
  END BcidMtx[799]
  PIN BcidMtx[880]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12173.625 187.44 12173.905 188.44 ;
    END
  END BcidMtx[880]
  PIN BcidMtx[879]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12173.065 187.44 12173.345 188.44 ;
    END
  END BcidMtx[879]
  PIN BcidMtx[878]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12171.385 187.44 12171.665 188.44 ;
    END
  END BcidMtx[878]
  PIN BcidMtx[872]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12094.665 187.44 12094.945 188.44 ;
    END
  END BcidMtx[872]
  PIN BcidMtx[870]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12093.545 187.44 12093.825 188.44 ;
    END
  END BcidMtx[870]
  PIN BcidMtx[867]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12026.345 187.44 12026.625 188.44 ;
    END
  END BcidMtx[867]
  PIN BcidMtx[866]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12024.665 187.44 12024.945 188.44 ;
    END
  END BcidMtx[866]
  PIN BcidMtx[865]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12024.105 187.44 12024.385 188.44 ;
    END
  END BcidMtx[865]
  PIN BcidMtx[1322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18080.505 187.44 18080.785 188.44 ;
    END
  END BcidMtx[1322]
  PIN BcidMtx[863]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11948.785 187.44 11949.065 188.44 ;
    END
  END BcidMtx[863]
  PIN BcidMtx[858]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11919.385 187.44 11919.665 188.44 ;
    END
  END BcidMtx[858]
  PIN BcidMtx[855]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11840.425 187.44 11840.705 188.44 ;
    END
  END BcidMtx[855]
  PIN BcidMtx[854]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11838.745 187.44 11839.025 188.44 ;
    END
  END BcidMtx[854]
  PIN BcidMtx[851]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11776.025 187.44 11776.305 188.44 ;
    END
  END BcidMtx[851]
  PIN BcidMtx[847]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11772.665 187.44 11772.945 188.44 ;
    END
  END BcidMtx[847]
  PIN BcidMtx[844]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11693.145 187.44 11693.425 188.44 ;
    END
  END BcidMtx[844]
  PIN BcidMtx[840]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11689.785 187.44 11690.065 188.44 ;
    END
  END BcidMtx[840]
  PIN BcidMtx[922]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12733.625 187.44 12733.905 188.44 ;
    END
  END BcidMtx[922]
  PIN BcidMtx[918]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12730.265 187.44 12730.545 188.44 ;
    END
  END BcidMtx[918]
  PIN BcidMtx[917]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12657.465 187.44 12657.745 188.44 ;
    END
  END BcidMtx[917]
  PIN BcidMtx[913]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12654.105 187.44 12654.385 188.44 ;
    END
  END BcidMtx[913]
  PIN BcidMtx[909]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12586.345 187.44 12586.625 188.44 ;
    END
  END BcidMtx[909]
  PIN BcidMtx[908]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12584.665 187.44 12584.945 188.44 ;
    END
  END BcidMtx[908]
  PIN BcidMtx[903]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12507.665 187.44 12507.945 188.44 ;
    END
  END BcidMtx[903]
  PIN BcidMtx[901]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12479.945 187.44 12480.225 188.44 ;
    END
  END BcidMtx[901]
  PIN BcidMtx[897]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12400.425 187.44 12400.705 188.44 ;
    END
  END BcidMtx[897]
  PIN BcidMtx[896]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12398.745 187.44 12399.025 188.44 ;
    END
  END BcidMtx[896]
  PIN BcidMtx[892]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12335.465 187.44 12335.745 188.44 ;
    END
  END BcidMtx[892]
  PIN BcidMtx[888]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12332.105 187.44 12332.385 188.44 ;
    END
  END BcidMtx[888]
  PIN BcidMtx[887]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12253.705 187.44 12253.985 188.44 ;
    END
  END BcidMtx[887]
  PIN BcidMtx[883]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12250.345 187.44 12250.625 188.44 ;
    END
  END BcidMtx[883]
  PIN BcidMtx[965]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13294.185 187.44 13294.465 188.44 ;
    END
  END BcidMtx[965]
  PIN BcidMtx[961]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13290.825 187.44 13291.105 188.44 ;
    END
  END BcidMtx[961]
  PIN BcidMtx[957]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13216.345 187.44 13216.625 188.44 ;
    END
  END BcidMtx[957]
  PIN BcidMtx[956]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13214.665 187.44 13214.945 188.44 ;
    END
  END BcidMtx[956]
  PIN BcidMtx[952]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13146.905 187.44 13147.185 188.44 ;
    END
  END BcidMtx[952]
  PIN BcidMtx[948]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13143.545 187.44 13143.825 188.44 ;
    END
  END BcidMtx[948]
  PIN BcidMtx[947]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13068.785 187.44 13069.065 188.44 ;
    END
  END BcidMtx[947]
  PIN BcidMtx[942]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13039.385 187.44 13039.665 188.44 ;
    END
  END BcidMtx[942]
  PIN BcidMtx[940]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12960.985 187.44 12961.265 188.44 ;
    END
  END BcidMtx[940]
  PIN BcidMtx[936]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12957.625 187.44 12957.905 188.44 ;
    END
  END BcidMtx[936]
  PIN BcidMtx[934]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12895.465 187.44 12895.745 188.44 ;
    END
  END BcidMtx[934]
  PIN BcidMtx[930]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12892.105 187.44 12892.385 188.44 ;
    END
  END BcidMtx[930]
  PIN BcidMtx[927]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12812.585 187.44 12812.865 188.44 ;
    END
  END BcidMtx[927]
  PIN BcidMtx[1007]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13854.185 187.44 13854.465 188.44 ;
    END
  END BcidMtx[1007]
  PIN BcidMtx[1003]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13850.825 187.44 13851.105 188.44 ;
    END
  END BcidMtx[1003]
  PIN BcidMtx[1000]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13776.905 187.44 13777.185 188.44 ;
    END
  END BcidMtx[1000]
  PIN BcidMtx[998]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13774.665 187.44 13774.945 188.44 ;
    END
  END BcidMtx[998]
  PIN BcidMtx[991]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13704.105 187.44 13704.385 188.44 ;
    END
  END BcidMtx[991]
  PIN BcidMtx[990]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13703.545 187.44 13703.825 188.44 ;
    END
  END BcidMtx[990]
  PIN BcidMtx[989]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13628.785 187.44 13629.065 188.44 ;
    END
  END BcidMtx[989]
  PIN BcidMtx[985]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13599.945 187.44 13600.225 188.44 ;
    END
  END BcidMtx[985]
  PIN BcidMtx[982]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13520.985 187.44 13521.265 188.44 ;
    END
  END BcidMtx[982]
  PIN BcidMtx[981]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13520.425 187.44 13520.705 188.44 ;
    END
  END BcidMtx[981]
  PIN BcidMtx[978]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13517.625 187.44 13517.905 188.44 ;
    END
  END BcidMtx[978]
  PIN BcidMtx[975]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13454.905 187.44 13455.185 188.44 ;
    END
  END BcidMtx[975]
  PIN BcidMtx[971]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13373.705 187.44 13373.985 188.44 ;
    END
  END BcidMtx[971]
  PIN BcidMtx[968]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13370.905 187.44 13371.185 188.44 ;
    END
  END BcidMtx[968]
  PIN BcidMtx[1049]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14414.185 187.44 14414.465 188.44 ;
    END
  END BcidMtx[1049]
  PIN BcidMtx[1047]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14413.065 187.44 14413.345 188.44 ;
    END
  END BcidMtx[1047]
  PIN BcidMtx[1046]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14411.385 187.44 14411.665 188.44 ;
    END
  END BcidMtx[1046]
  PIN BcidMtx[1040]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14334.665 187.44 14334.945 188.44 ;
    END
  END BcidMtx[1040]
  PIN BcidMtx[1036]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14266.905 187.44 14267.185 188.44 ;
    END
  END BcidMtx[1036]
  PIN BcidMtx[1032]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14263.545 187.44 14263.825 188.44 ;
    END
  END BcidMtx[1032]
  PIN BcidMtx[1029]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14187.665 187.44 14187.945 188.44 ;
    END
  END BcidMtx[1029]
  PIN BcidMtx[1026]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14159.385 187.44 14159.665 188.44 ;
    END
  END BcidMtx[1026]
  PIN BcidMtx[1023]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14080.425 187.44 14080.705 188.44 ;
    END
  END BcidMtx[1023]
  PIN BcidMtx[1022]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14078.745 187.44 14079.025 188.44 ;
    END
  END BcidMtx[1022]
  PIN BcidMtx[1017]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14014.905 187.44 14015.185 188.44 ;
    END
  END BcidMtx[1017]
  PIN BcidMtx[1012]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13933.145 187.44 13933.425 188.44 ;
    END
  END BcidMtx[1012]
  PIN BcidMtx[1009]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13930.345 187.44 13930.625 188.44 ;
    END
  END BcidMtx[1009]
  PIN BcidMtx[1091]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14974.185 187.44 14974.465 188.44 ;
    END
  END BcidMtx[1091]
  PIN BcidMtx[1089]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14973.065 187.44 14973.345 188.44 ;
    END
  END BcidMtx[1089]
  PIN BcidMtx[1087]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14970.825 187.44 14971.105 188.44 ;
    END
  END BcidMtx[1087]
  PIN BcidMtx[1083]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14896.345 187.44 14896.625 188.44 ;
    END
  END BcidMtx[1083]
  PIN BcidMtx[1082]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14894.665 187.44 14894.945 188.44 ;
    END
  END BcidMtx[1082]
  PIN BcidMtx[1080]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14893.545 187.44 14893.825 188.44 ;
    END
  END BcidMtx[1080]
  PIN BcidMtx[1311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17934.905 187.44 17935.185 188.44 ;
    END
  END BcidMtx[1311]
  PIN BcidMtx[1074]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14823.545 187.44 14823.825 188.44 ;
    END
  END BcidMtx[1074]
  PIN BcidMtx[1072]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14748.225 187.44 14748.505 188.44 ;
    END
  END BcidMtx[1072]
  PIN BcidMtx[1070]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14720.505 187.44 14720.785 188.44 ;
    END
  END BcidMtx[1070]
  PIN BcidMtx[1068]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14719.385 187.44 14719.665 188.44 ;
    END
  END BcidMtx[1068]
  PIN BcidMtx[1066]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14640.985 187.44 14641.265 188.44 ;
    END
  END BcidMtx[1066]
  PIN BcidMtx[1063]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14638.185 187.44 14638.465 188.44 ;
    END
  END BcidMtx[1063]
  PIN BcidMtx[1057]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14572.665 187.44 14572.945 188.44 ;
    END
  END BcidMtx[1057]
  PIN BcidMtx[1054]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14493.145 187.44 14493.425 188.44 ;
    END
  END BcidMtx[1054]
  PIN BcidMtx[1052]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14490.905 187.44 14491.185 188.44 ;
    END
  END BcidMtx[1052]
  PIN BcidMtx[1131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15533.065 187.44 15533.345 188.44 ;
    END
  END BcidMtx[1131]
  PIN BcidMtx[1130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15531.385 187.44 15531.665 188.44 ;
    END
  END BcidMtx[1130]
  PIN BcidMtx[1126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15456.905 187.44 15457.185 188.44 ;
    END
  END BcidMtx[1126]
  PIN BcidMtx[1122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15453.545 187.44 15453.825 188.44 ;
    END
  END BcidMtx[1122]
  PIN BcidMtx[1121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15387.465 187.44 15387.745 188.44 ;
    END
  END BcidMtx[1121]
  PIN BcidMtx[1117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15384.105 187.44 15384.385 188.44 ;
    END
  END BcidMtx[1117]
  PIN BcidMtx[1115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15308.785 187.44 15309.065 188.44 ;
    END
  END BcidMtx[1115]
  PIN BcidMtx[1113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15307.665 187.44 15307.945 188.44 ;
    END
  END BcidMtx[1113]
  PIN BcidMtx[1111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15279.945 187.44 15280.225 188.44 ;
    END
  END BcidMtx[1111]
  PIN BcidMtx[1108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15200.985 187.44 15201.265 188.44 ;
    END
  END BcidMtx[1108]
  PIN BcidMtx[1106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15198.745 187.44 15199.025 188.44 ;
    END
  END BcidMtx[1106]
  PIN BcidMtx[1099]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15132.665 187.44 15132.945 188.44 ;
    END
  END BcidMtx[1099]
  PIN BcidMtx[1309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17932.665 187.44 17932.945 188.44 ;
    END
  END BcidMtx[1309]
  PIN BcidMtx[1092]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15049.785 187.44 15050.065 188.44 ;
    END
  END BcidMtx[1092]
  PIN BcidMtx[1172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16091.385 187.44 16091.665 188.44 ;
    END
  END BcidMtx[1172]
  PIN BcidMtx[1171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16090.825 187.44 16091.105 188.44 ;
    END
  END BcidMtx[1171]
  PIN BcidMtx[1164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16013.545 187.44 16013.825 188.44 ;
    END
  END BcidMtx[1164]
  PIN BcidMtx[1159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15944.105 187.44 15944.385 188.44 ;
    END
  END BcidMtx[1159]
  PIN BcidMtx[1154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15840.505 187.44 15840.785 188.44 ;
    END
  END BcidMtx[1154]
  PIN BcidMtx[1152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15839.385 187.44 15839.665 188.44 ;
    END
  END BcidMtx[1152]
  PIN BcidMtx[1150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15760.985 187.44 15761.265 188.44 ;
    END
  END BcidMtx[1150]
  PIN BcidMtx[1147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15758.185 187.44 15758.465 188.44 ;
    END
  END BcidMtx[1147]
  PIN BcidMtx[1144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15695.465 187.44 15695.745 188.44 ;
    END
  END BcidMtx[1144]
  PIN BcidMtx[1139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15613.705 187.44 15613.985 188.44 ;
    END
  END BcidMtx[1139]
  PIN BcidMtx[1137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15612.585 187.44 15612.865 188.44 ;
    END
  END BcidMtx[1137]
  PIN BcidMtx[1134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15609.785 187.44 15610.065 188.44 ;
    END
  END BcidMtx[1134]
  PIN BcidMtx[1216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16653.625 187.44 16653.905 188.44 ;
    END
  END BcidMtx[1216]
  PIN BcidMtx[1212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16650.265 187.44 16650.545 188.44 ;
    END
  END BcidMtx[1212]
  PIN BcidMtx[1210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16576.905 187.44 16577.185 188.44 ;
    END
  END BcidMtx[1210]
  PIN BcidMtx[1207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16574.105 187.44 16574.385 188.44 ;
    END
  END BcidMtx[1207]
  PIN BcidMtx[1203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16506.345 187.44 16506.625 188.44 ;
    END
  END BcidMtx[1203]
  PIN BcidMtx[1202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16504.665 187.44 16504.945 188.44 ;
    END
  END BcidMtx[1202]
  PIN BcidMtx[1200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16503.545 187.44 16503.825 188.44 ;
    END
  END BcidMtx[1200]
  PIN BcidMtx[1199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16428.785 187.44 16429.065 188.44 ;
    END
  END BcidMtx[1199]
  PIN BcidMtx[1196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16400.505 187.44 16400.785 188.44 ;
    END
  END BcidMtx[1196]
  PIN BcidMtx[1192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16320.985 187.44 16321.265 188.44 ;
    END
  END BcidMtx[1192]
  PIN BcidMtx[1190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16318.745 187.44 16319.025 188.44 ;
    END
  END BcidMtx[1190]
  PIN BcidMtx[1187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16256.025 187.44 16256.305 188.44 ;
    END
  END BcidMtx[1187]
  PIN BcidMtx[1185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16254.905 187.44 16255.185 188.44 ;
    END
  END BcidMtx[1185]
  PIN BcidMtx[1183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16252.665 187.44 16252.945 188.44 ;
    END
  END BcidMtx[1183]
  PIN BcidMtx[1180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16173.145 187.44 16173.425 188.44 ;
    END
  END BcidMtx[1180]
  PIN BcidMtx[1176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16169.785 187.44 16170.065 188.44 ;
    END
  END BcidMtx[1176]
  PIN BcidMtx[1258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17213.625 187.44 17213.905 188.44 ;
    END
  END BcidMtx[1258]
  PIN BcidMtx[1254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17210.265 187.44 17210.545 188.44 ;
    END
  END BcidMtx[1254]
  PIN BcidMtx[1253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17137.465 187.44 17137.745 188.44 ;
    END
  END BcidMtx[1253]
  PIN BcidMtx[1250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17134.665 187.44 17134.945 188.44 ;
    END
  END BcidMtx[1250]
  PIN BcidMtx[1246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17066.905 187.44 17067.185 188.44 ;
    END
  END BcidMtx[1246]
  PIN BcidMtx[1243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17064.105 187.44 17064.385 188.44 ;
    END
  END BcidMtx[1243]
  PIN BcidMtx[1315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17998.185 187.44 17998.465 188.44 ;
    END
  END BcidMtx[1315]
  PIN BcidMtx[1240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16988.225 187.44 16988.505 188.44 ;
    END
  END BcidMtx[1240]
  PIN BcidMtx[1238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16960.505 187.44 16960.785 188.44 ;
    END
  END BcidMtx[1238]
  PIN BcidMtx[1236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16959.385 187.44 16959.665 188.44 ;
    END
  END BcidMtx[1236]
  PIN BcidMtx[1234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16880.985 187.44 16881.265 188.44 ;
    END
  END BcidMtx[1234]
  PIN BcidMtx[1231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16878.185 187.44 16878.465 188.44 ;
    END
  END BcidMtx[1231]
  PIN BcidMtx[1225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16812.665 187.44 16812.945 188.44 ;
    END
  END BcidMtx[1225]
  PIN BcidMtx[1222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16733.145 187.44 16733.425 188.44 ;
    END
  END BcidMtx[1222]
  PIN BcidMtx[1220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16730.905 187.44 16731.185 188.44 ;
    END
  END BcidMtx[1220]
  PIN BcidMtx[1301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17774.185 187.44 17774.465 188.44 ;
    END
  END BcidMtx[1301]
  PIN BcidMtx[1297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17770.825 187.44 17771.105 188.44 ;
    END
  END BcidMtx[1297]
  PIN BcidMtx[1293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17696.345 187.44 17696.625 188.44 ;
    END
  END BcidMtx[1293]
  PIN BcidMtx[1292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17694.665 187.44 17694.945 188.44 ;
    END
  END BcidMtx[1292]
  PIN BcidMtx[1287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17626.345 187.44 17626.625 188.44 ;
    END
  END BcidMtx[1287]
  PIN BcidMtx[1286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17624.665 187.44 17624.945 188.44 ;
    END
  END BcidMtx[1286]
  PIN BcidMtx[1284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17623.545 187.44 17623.825 188.44 ;
    END
  END BcidMtx[1284]
  PIN BcidMtx[1281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17547.665 187.44 17547.945 188.44 ;
    END
  END BcidMtx[1281]
  PIN BcidMtx[1279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17519.945 187.44 17520.225 188.44 ;
    END
  END BcidMtx[1279]
  PIN BcidMtx[1277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17441.545 187.44 17441.825 188.44 ;
    END
  END BcidMtx[1277]
  PIN BcidMtx[1274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17438.745 187.44 17439.025 188.44 ;
    END
  END BcidMtx[1274]
  PIN BcidMtx[1270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17375.465 187.44 17375.745 188.44 ;
    END
  END BcidMtx[1270]
  PIN BcidMtx[1267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17372.665 187.44 17372.945 188.44 ;
    END
  END BcidMtx[1267]
  PIN BcidMtx[1264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17293.145 187.44 17293.425 188.44 ;
    END
  END BcidMtx[1264]
  PIN BcidMtx[1262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17290.905 187.44 17291.185 188.44 ;
    END
  END BcidMtx[1262]
  PIN BcidMtx[1343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18334.185 187.44 18334.465 188.44 ;
    END
  END BcidMtx[1343]
  PIN BcidMtx[1340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18331.385 187.44 18331.665 188.44 ;
    END
  END BcidMtx[1340]
  PIN BcidMtx[1338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18330.265 187.44 18330.545 188.44 ;
    END
  END BcidMtx[1338]
  PIN BcidMtx[1336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18256.905 187.44 18257.185 188.44 ;
    END
  END BcidMtx[1336]
  PIN BcidMtx[1334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18254.665 187.44 18254.945 188.44 ;
    END
  END BcidMtx[1334]
  PIN BcidMtx[1304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17850.905 187.44 17851.185 188.44 ;
    END
  END BcidMtx[1304]
  PIN BcidMtx[1303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17850.345 187.44 17850.625 188.44 ;
    END
  END BcidMtx[1303]
  PIN BcidMtx[1302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17849.785 187.44 17850.065 188.44 ;
    END
  END BcidMtx[1302]
  PIN BcidMtx[1307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17853.705 187.44 17853.985 188.44 ;
    END
  END BcidMtx[1307]
  PIN BcidMtx[1306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17853.145 187.44 17853.425 188.44 ;
    END
  END BcidMtx[1306]
  PIN BcidMtx[1305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17852.585 187.44 17852.865 188.44 ;
    END
  END BcidMtx[1305]
  PIN SET_VCASN[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18356.515 187.44 18356.795 188.44 ;
    END
  END SET_VCASN[127]
  PIN DIG_MON_PMOS_NOSF[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 998.265 187.44 998.545 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[13]
  PIN Data_PMOS_NOSF[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 996.025 187.44 996.305 188.44 ;
    END
  END Data_PMOS_NOSF[144]
  PIN Data_PMOS_NOSF[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 995.465 187.44 995.745 188.44 ;
    END
  END Data_PMOS_NOSF[134]
  PIN Data_PMOS_NOSF[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 994.905 187.44 995.185 188.44 ;
    END
  END Data_PMOS_NOSF[138]
  PIN Data_PMOS_NOSF[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 994.345 187.44 994.625 188.44 ;
    END
  END Data_PMOS_NOSF[145]
  PIN Data_PMOS_NOSF[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 993.785 187.44 994.065 188.44 ;
    END
  END Data_PMOS_NOSF[131]
  PIN Data_PMOS_NOSF[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 993.225 187.44 993.505 188.44 ;
    END
  END Data_PMOS_NOSF[139]
  PIN Data_PMOS_NOSF[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 992.665 187.44 992.945 188.44 ;
    END
  END Data_PMOS_NOSF[146]
  PIN Data_PMOS_NOSF[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 992.105 187.44 992.385 188.44 ;
    END
  END Data_PMOS_NOSF[140]
  PIN Data_PMOS_NOSF[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 991.545 187.44 991.825 188.44 ;
    END
  END Data_PMOS_NOSF[133]
  PIN Data_PMOS_NOSF[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 990.985 187.44 991.265 188.44 ;
    END
  END Data_PMOS_NOSF[132]
  PIN nTOK_PMOS_NOSF[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 988.745 187.44 989.025 188.44 ;
    END
  END nTOK_PMOS_NOSF[6]
  PIN FREEZE_PMOS_NOSF[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 972.505 187.44 972.785 188.44 ;
    END
  END FREEZE_PMOS_NOSF[6]
  PIN Read_PMOS_NOSF[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 971.945 187.44 972.225 188.44 ;
    END
  END Read_PMOS_NOSF[6]
  PIN Data_PMOS_NOSF[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 968.025 187.44 968.305 188.44 ;
    END
  END Data_PMOS_NOSF[129]
  PIN Data_PMOS_NOSF[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 967.465 187.44 967.745 188.44 ;
    END
  END Data_PMOS_NOSF[128]
  PIN Data_PMOS_NOSF[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 966.905 187.44 967.185 188.44 ;
    END
  END Data_PMOS_NOSF[135]
  PIN Data_PMOS_NOSF[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 966.345 187.44 966.625 188.44 ;
    END
  END Data_PMOS_NOSF[141]
  PIN Data_PMOS_NOSF[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 965.785 187.44 966.065 188.44 ;
    END
  END Data_PMOS_NOSF[136]
  PIN Data_PMOS_NOSF[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 965.225 187.44 965.505 188.44 ;
    END
  END Data_PMOS_NOSF[130]
  PIN Data_PMOS_NOSF[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 964.665 187.44 964.945 188.44 ;
    END
  END Data_PMOS_NOSF[142]
  PIN Data_PMOS_NOSF[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 964.105 187.44 964.385 188.44 ;
    END
  END Data_PMOS_NOSF[137]
  PIN Data_PMOS_NOSF[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 963.545 187.44 963.825 188.44 ;
    END
  END Data_PMOS_NOSF[127]
  PIN Data_PMOS_NOSF[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 962.985 187.44 963.265 188.44 ;
    END
  END Data_PMOS_NOSF[126]
  PIN Data_PMOS_NOSF[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 962.425 187.44 962.705 188.44 ;
    END
  END Data_PMOS_NOSF[143]
  PIN DIG_MON_PMOS_NOSF[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 920.985 187.44 921.265 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[12]
  PIN DIG_MON_PMOS_NOSF[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 916.505 187.44 916.785 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[11]
  PIN Data_PMOS_NOSF[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 914.265 187.44 914.545 188.44 ;
    END
  END Data_PMOS_NOSF[123]
  PIN Data_PMOS_NOSF[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 913.705 187.44 913.985 188.44 ;
    END
  END Data_PMOS_NOSF[113]
  PIN Data_PMOS_NOSF[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 913.145 187.44 913.425 188.44 ;
    END
  END Data_PMOS_NOSF[117]
  PIN Data_PMOS_NOSF[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 912.585 187.44 912.865 188.44 ;
    END
  END Data_PMOS_NOSF[124]
  PIN Data_PMOS_NOSF[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 912.025 187.44 912.305 188.44 ;
    END
  END Data_PMOS_NOSF[110]
  PIN Data_PMOS_NOSF[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 911.465 187.44 911.745 188.44 ;
    END
  END Data_PMOS_NOSF[118]
  PIN Data_PMOS_NOSF[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 910.905 187.44 911.185 188.44 ;
    END
  END Data_PMOS_NOSF[125]
  PIN Data_PMOS_NOSF[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 910.345 187.44 910.625 188.44 ;
    END
  END Data_PMOS_NOSF[119]
  PIN Data_PMOS_NOSF[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 909.785 187.44 910.065 188.44 ;
    END
  END Data_PMOS_NOSF[112]
  PIN Data_PMOS_NOSF[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 900.825 187.44 901.105 188.44 ;
    END
  END Data_PMOS_NOSF[111]
  PIN nTOK_PMOS_NOSF[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 898.585 187.44 898.865 188.44 ;
    END
  END nTOK_PMOS_NOSF[5]
  PIN FREEZE_PMOS_NOSF[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 895.785 187.44 896.065 188.44 ;
    END
  END FREEZE_PMOS_NOSF[5]
  PIN Read_PMOS_NOSF[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 895.225 187.44 895.505 188.44 ;
    END
  END Read_PMOS_NOSF[5]
  PIN Data_PMOS_NOSF[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 889.345 187.44 889.625 188.44 ;
    END
  END Data_PMOS_NOSF[108]
  PIN Data_PMOS_NOSF[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 888.785 187.44 889.065 188.44 ;
    END
  END Data_PMOS_NOSF[107]
  PIN Data_PMOS_NOSF[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 888.225 187.44 888.505 188.44 ;
    END
  END Data_PMOS_NOSF[114]
  PIN Data_PMOS_NOSF[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 887.665 187.44 887.945 188.44 ;
    END
  END Data_PMOS_NOSF[120]
  PIN Data_PMOS_NOSF[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 887.105 187.44 887.385 188.44 ;
    END
  END Data_PMOS_NOSF[115]
  PIN Data_PMOS_NOSF[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 861.065 187.44 861.345 188.44 ;
    END
  END Data_PMOS_NOSF[109]
  PIN Data_PMOS_NOSF[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 860.505 187.44 860.785 188.44 ;
    END
  END Data_PMOS_NOSF[121]
  PIN Data_PMOS_NOSF[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 859.945 187.44 860.225 188.44 ;
    END
  END Data_PMOS_NOSF[116]
  PIN Data_PMOS_NOSF[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 859.385 187.44 859.665 188.44 ;
    END
  END Data_PMOS_NOSF[106]
  PIN Data_PMOS_NOSF[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 858.825 187.44 859.105 188.44 ;
    END
  END Data_PMOS_NOSF[105]
  PIN Data_PMOS_NOSF[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 858.265 187.44 858.545 188.44 ;
    END
  END Data_PMOS_NOSF[122]
  PIN DIG_MON_PMOS_NOSF[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 855.465 187.44 855.745 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[10]
  PIN DIG_MON_PMOS_NOSF[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 850.985 187.44 851.265 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[9]
  PIN Data_PMOS_NOSF[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 848.745 187.44 849.025 188.44 ;
    END
  END Data_PMOS_NOSF[102]
  PIN Data_PMOS_NOSF[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 848.185 187.44 848.465 188.44 ;
    END
  END Data_PMOS_NOSF[92]
  PIN Data_PMOS_NOSF[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 834.745 187.44 835.025 188.44 ;
    END
  END Data_PMOS_NOSF[96]
  PIN Data_PMOS_NOSF[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 834.185 187.44 834.465 188.44 ;
    END
  END Data_PMOS_NOSF[103]
  PIN Data_PMOS_NOSF[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 833.625 187.44 833.905 188.44 ;
    END
  END Data_PMOS_NOSF[89]
  PIN Data_PMOS_NOSF[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 833.065 187.44 833.345 188.44 ;
    END
  END Data_PMOS_NOSF[97]
  PIN Data_PMOS_NOSF[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 832.505 187.44 832.785 188.44 ;
    END
  END Data_PMOS_NOSF[104]
  PIN Data_PMOS_NOSF[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 831.945 187.44 832.225 188.44 ;
    END
  END Data_PMOS_NOSF[98]
  PIN Data_PMOS_NOSF[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 831.385 187.44 831.665 188.44 ;
    END
  END Data_PMOS_NOSF[91]
  PIN Data_PMOS_NOSF[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 830.825 187.44 831.105 188.44 ;
    END
  END Data_PMOS_NOSF[90]
  PIN nTOK_PMOS_NOSF[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 828.585 187.44 828.865 188.44 ;
    END
  END nTOK_PMOS_NOSF[4]
  PIN FREEZE_PMOS_NOSF[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 825.785 187.44 826.065 188.44 ;
    END
  END FREEZE_PMOS_NOSF[4]
  PIN Read_PMOS_NOSF[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 825.225 187.44 825.505 188.44 ;
    END
  END Read_PMOS_NOSF[4]
  PIN Data_PMOS_NOSF[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 782.665 187.44 782.945 188.44 ;
    END
  END Data_PMOS_NOSF[87]
  PIN Data_PMOS_NOSF[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 782.105 187.44 782.385 188.44 ;
    END
  END Data_PMOS_NOSF[86]
  PIN Data_PMOS_NOSF[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 781.545 187.44 781.825 188.44 ;
    END
  END Data_PMOS_NOSF[93]
  PIN Data_PMOS_NOSF[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 780.985 187.44 781.265 188.44 ;
    END
  END Data_PMOS_NOSF[99]
  PIN Data_PMOS_NOSF[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 780.425 187.44 780.705 188.44 ;
    END
  END Data_PMOS_NOSF[94]
  PIN Data_PMOS_NOSF[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 779.865 187.44 780.145 188.44 ;
    END
  END Data_PMOS_NOSF[88]
  PIN Data_PMOS_NOSF[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 779.305 187.44 779.585 188.44 ;
    END
  END Data_PMOS_NOSF[100]
  PIN Data_PMOS_NOSF[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 778.745 187.44 779.025 188.44 ;
    END
  END Data_PMOS_NOSF[95]
  PIN Data_PMOS_NOSF[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 778.185 187.44 778.465 188.44 ;
    END
  END Data_PMOS_NOSF[85]
  PIN Data_PMOS_NOSF[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 777.625 187.44 777.905 188.44 ;
    END
  END Data_PMOS_NOSF[84]
  PIN Data_PMOS_NOSF[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 777.065 187.44 777.345 188.44 ;
    END
  END Data_PMOS_NOSF[101]
  PIN DIG_MON_PMOS_NOSF[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 774.265 187.44 774.545 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[8]
  PIN DIG_MON_PMOS_NOSF[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 769.785 187.44 770.065 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[7]
  PIN Data_PMOS_NOSF[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 759.145 187.44 759.425 188.44 ;
    END
  END Data_PMOS_NOSF[81]
  PIN Data_PMOS_NOSF[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 758.585 187.44 758.865 188.44 ;
    END
  END Data_PMOS_NOSF[71]
  PIN Data_PMOS_NOSF[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 758.025 187.44 758.305 188.44 ;
    END
  END Data_PMOS_NOSF[75]
  PIN Data_PMOS_NOSF[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 757.465 187.44 757.745 188.44 ;
    END
  END Data_PMOS_NOSF[82]
  PIN Data_PMOS_NOSF[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 756.345 187.44 756.625 188.44 ;
    END
  END Data_PMOS_NOSF[76]
  PIN Data_PMOS_NOSF[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 756.905 187.44 757.185 188.44 ;
    END
  END Data_PMOS_NOSF[68]
  PIN Data_PMOS_NOSF[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 755.785 187.44 756.065 188.44 ;
    END
  END Data_PMOS_NOSF[83]
  PIN Data_PMOS_NOSF[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 755.225 187.44 755.505 188.44 ;
    END
  END Data_PMOS_NOSF[77]
  PIN Data_PMOS_NOSF[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 754.665 187.44 754.945 188.44 ;
    END
  END Data_PMOS_NOSF[70]
  PIN Data_PMOS_NOSF[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 754.105 187.44 754.385 188.44 ;
    END
  END Data_PMOS_NOSF[69]
  PIN nTOK_PMOS_NOSF[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 749.905 187.44 750.185 188.44 ;
    END
  END nTOK_PMOS_NOSF[3]
  PIN Read_PMOS_NOSF[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 721.065 187.44 721.345 188.44 ;
    END
  END Read_PMOS_NOSF[3]
  PIN Data_PMOS_NOSF[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 717.145 187.44 717.425 188.44 ;
    END
  END Data_PMOS_NOSF[66]
  PIN Data_PMOS_NOSF[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 716.585 187.44 716.865 188.44 ;
    END
  END Data_PMOS_NOSF[65]
  PIN Data_PMOS_NOSF[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 716.025 187.44 716.305 188.44 ;
    END
  END Data_PMOS_NOSF[72]
  PIN Data_PMOS_NOSF[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 715.465 187.44 715.745 188.44 ;
    END
  END Data_PMOS_NOSF[78]
  PIN Data_PMOS_NOSF[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 714.905 187.44 715.185 188.44 ;
    END
  END Data_PMOS_NOSF[73]
  PIN Data_PMOS_NOSF[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 714.345 187.44 714.625 188.44 ;
    END
  END Data_PMOS_NOSF[67]
  PIN Data_PMOS_NOSF[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 713.225 187.44 713.505 188.44 ;
    END
  END Data_PMOS_NOSF[74]
  PIN Data_PMOS_NOSF[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 713.785 187.44 714.065 188.44 ;
    END
  END Data_PMOS_NOSF[79]
  PIN Data_PMOS_NOSF[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 712.665 187.44 712.945 188.44 ;
    END
  END Data_PMOS_NOSF[64]
  PIN Data_PMOS_NOSF[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 712.105 187.44 712.385 188.44 ;
    END
  END Data_PMOS_NOSF[63]
  PIN Data_PMOS_NOSF[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 711.545 187.44 711.825 188.44 ;
    END
  END Data_PMOS_NOSF[80]
  PIN DIG_MON_PMOS_NOSF[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 708.745 187.44 709.025 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[6]
  PIN DIG_MON_PMOS_NOSF[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 691.385 187.44 691.665 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[5]
  PIN Data_PMOS_NOSF[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 689.145 187.44 689.425 188.44 ;
    END
  END Data_PMOS_NOSF[60]
  PIN Data_PMOS_NOSF[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 688.585 187.44 688.865 188.44 ;
    END
  END Data_PMOS_NOSF[50]
  PIN Data_PMOS_NOSF[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 688.025 187.44 688.305 188.44 ;
    END
  END Data_PMOS_NOSF[54]
  PIN Data_PMOS_NOSF[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 687.465 187.44 687.745 188.44 ;
    END
  END Data_PMOS_NOSF[61]
  PIN Data_PMOS_NOSF[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 686.905 187.44 687.185 188.44 ;
    END
  END Data_PMOS_NOSF[47]
  PIN Data_PMOS_NOSF[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 686.345 187.44 686.625 188.44 ;
    END
  END Data_PMOS_NOSF[55]
  PIN Data_PMOS_NOSF[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 685.785 187.44 686.065 188.44 ;
    END
  END Data_PMOS_NOSF[62]
  PIN Data_PMOS_NOSF[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 684.665 187.44 684.945 188.44 ;
    END
  END Data_PMOS_NOSF[49]
  PIN Data_PMOS_NOSF[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 684.105 187.44 684.385 188.44 ;
    END
  END Data_PMOS_NOSF[48]
  PIN nTOK_PMOS_NOSF[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 642.665 187.44 642.945 188.44 ;
    END
  END nTOK_PMOS_NOSF[2]
  PIN Data_PMOS_NOSF[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 685.225 187.44 685.505 188.44 ;
    END
  END Data_PMOS_NOSF[56]
  PIN FREEZE_PMOS_NOSF[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 639.865 187.44 640.145 188.44 ;
    END
  END FREEZE_PMOS_NOSF[2]
  PIN Read_PMOS_NOSF[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 639.305 187.44 639.585 188.44 ;
    END
  END Read_PMOS_NOSF[2]
  PIN Data_PMOS_NOSF[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 635.385 187.44 635.665 188.44 ;
    END
  END Data_PMOS_NOSF[45]
  PIN Data_PMOS_NOSF[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 634.825 187.44 635.105 188.44 ;
    END
  END Data_PMOS_NOSF[44]
  PIN Data_PMOS_NOSF[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 634.265 187.44 634.545 188.44 ;
    END
  END Data_PMOS_NOSF[51]
  PIN Data_PMOS_NOSF[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 633.705 187.44 633.985 188.44 ;
    END
  END Data_PMOS_NOSF[57]
  PIN Data_PMOS_NOSF[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 633.145 187.44 633.425 188.44 ;
    END
  END Data_PMOS_NOSF[52]
  PIN Data_PMOS_NOSF[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 632.585 187.44 632.865 188.44 ;
    END
  END Data_PMOS_NOSF[46]
  PIN Data_PMOS_NOSF[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 632.025 187.44 632.305 188.44 ;
    END
  END Data_PMOS_NOSF[58]
  PIN Data_PMOS_NOSF[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 631.465 187.44 631.745 188.44 ;
    END
  END Data_PMOS_NOSF[53]
  PIN Data_PMOS_NOSF[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 630.905 187.44 631.185 188.44 ;
    END
  END Data_PMOS_NOSF[43]
  PIN Data_PMOS_NOSF[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 630.345 187.44 630.625 188.44 ;
    END
  END Data_PMOS_NOSF[42]
  PIN Data_PMOS_NOSF[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 629.785 187.44 630.065 188.44 ;
    END
  END Data_PMOS_NOSF[59]
  PIN DIG_MON_PMOS_NOSF[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 618.585 187.44 618.865 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[4]
  PIN DIG_MON_PMOS_NOSF[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 614.105 187.44 614.385 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[3]
  PIN Data_PMOS_NOSF[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 609.905 187.44 610.185 188.44 ;
    END
  END Data_PMOS_NOSF[39]
  PIN Data_PMOS_NOSF[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 609.345 187.44 609.625 188.44 ;
    END
  END Data_PMOS_NOSF[29]
  PIN Data_PMOS_NOSF[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 608.785 187.44 609.065 188.44 ;
    END
  END Data_PMOS_NOSF[33]
  PIN Data_PMOS_NOSF[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 608.225 187.44 608.505 188.44 ;
    END
  END Data_PMOS_NOSF[40]
  PIN Data_PMOS_NOSF[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 607.665 187.44 607.945 188.44 ;
    END
  END Data_PMOS_NOSF[26]
  PIN Data_PMOS_NOSF[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 581.625 187.44 581.905 188.44 ;
    END
  END Data_PMOS_NOSF[34]
  PIN Data_PMOS_NOSF[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 581.065 187.44 581.345 188.44 ;
    END
  END Data_PMOS_NOSF[41]
  PIN Data_PMOS_NOSF[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 580.505 187.44 580.785 188.44 ;
    END
  END Data_PMOS_NOSF[35]
  PIN Data_PMOS_NOSF[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 579.945 187.44 580.225 188.44 ;
    END
  END Data_PMOS_NOSF[28]
  PIN Data_PMOS_NOSF[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 579.385 187.44 579.665 188.44 ;
    END
  END Data_PMOS_NOSF[27]
  PIN nTOK_PMOS_NOSF[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 577.145 187.44 577.425 188.44 ;
    END
  END nTOK_PMOS_NOSF[1]
  PIN FREEZE_PMOS_NOSF[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 574.345 187.44 574.625 188.44 ;
    END
  END FREEZE_PMOS_NOSF[1]
  PIN Read_PMOS_NOSF[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 573.785 187.44 574.065 188.44 ;
    END
  END Read_PMOS_NOSF[1]
  PIN Data_PMOS_NOSF[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 569.865 187.44 570.145 188.44 ;
    END
  END Data_PMOS_NOSF[24]
  PIN Data_PMOS_NOSF[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 569.305 187.44 569.585 188.44 ;
    END
  END Data_PMOS_NOSF[23]
  PIN Data_PMOS_NOSF[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 568.745 187.44 569.025 188.44 ;
    END
  END Data_PMOS_NOSF[30]
  PIN Data_PMOS_NOSF[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 554.745 187.44 555.025 188.44 ;
    END
  END Data_PMOS_NOSF[31]
  PIN Data_PMOS_NOSF[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 555.305 187.44 555.585 188.44 ;
    END
  END Data_PMOS_NOSF[36]
  PIN Data_PMOS_NOSF[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 554.185 187.44 554.465 188.44 ;
    END
  END Data_PMOS_NOSF[25]
  PIN Data_PMOS_NOSF[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 553.625 187.44 553.905 188.44 ;
    END
  END Data_PMOS_NOSF[37]
  PIN Data_PMOS_NOSF[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 552.505 187.44 552.785 188.44 ;
    END
  END Data_PMOS_NOSF[22]
  PIN Data_PMOS_NOSF[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 553.065 187.44 553.345 188.44 ;
    END
  END Data_PMOS_NOSF[32]
  PIN Data_PMOS_NOSF[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 551.945 187.44 552.225 188.44 ;
    END
  END Data_PMOS_NOSF[21]
  PIN Data_PMOS_NOSF[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 551.385 187.44 551.665 188.44 ;
    END
  END Data_PMOS_NOSF[38]
  PIN DIG_MON_PMOS_NOSF[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 548.585 187.44 548.865 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[2]
  PIN DIG_MON_PMOS_NOSF[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 544.105 187.44 544.385 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[1]
  PIN Data_PMOS_NOSF[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 502.105 187.44 502.385 188.44 ;
    END
  END Data_PMOS_NOSF[18]
  PIN Data_PMOS_NOSF[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 501.545 187.44 501.825 188.44 ;
    END
  END Data_PMOS_NOSF[8]
  PIN Data_PMOS_NOSF[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 500.985 187.44 501.265 188.44 ;
    END
  END Data_PMOS_NOSF[12]
  PIN Data_PMOS_NOSF[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 500.425 187.44 500.705 188.44 ;
    END
  END Data_PMOS_NOSF[19]
  PIN Data_PMOS_NOSF[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 499.865 187.44 500.145 188.44 ;
    END
  END Data_PMOS_NOSF[5]
  PIN Data_PMOS_NOSF[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 499.305 187.44 499.585 188.44 ;
    END
  END Data_PMOS_NOSF[13]
  PIN Data_PMOS_NOSF[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 498.745 187.44 499.025 188.44 ;
    END
  END Data_PMOS_NOSF[20]
  PIN Data_PMOS_NOSF[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 498.185 187.44 498.465 188.44 ;
    END
  END Data_PMOS_NOSF[14]
  PIN Data_PMOS_NOSF[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 497.625 187.44 497.905 188.44 ;
    END
  END Data_PMOS_NOSF[7]
  PIN Data_PMOS_NOSF[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 497.065 187.44 497.345 188.44 ;
    END
  END Data_PMOS_NOSF[6]
  PIN nTOK_PMOS_NOSF[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 494.825 187.44 495.105 188.44 ;
    END
  END nTOK_PMOS_NOSF[0]
  PIN FREEZE_PMOS_NOSF[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 492.025 187.44 492.305 188.44 ;
    END
  END FREEZE_PMOS_NOSF[0]
  PIN Read_PMOS_NOSF[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 491.465 187.44 491.745 188.44 ;
    END
  END Read_PMOS_NOSF[0]
  PIN Data_PMOS_NOSF[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 479.145 187.44 479.425 188.44 ;
    END
  END Data_PMOS_NOSF[3]
  PIN Data_PMOS_NOSF[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 478.585 187.44 478.865 188.44 ;
    END
  END Data_PMOS_NOSF[2]
  PIN Data_PMOS_NOSF[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 478.025 187.44 478.305 188.44 ;
    END
  END Data_PMOS_NOSF[9]
  PIN Data_PMOS_NOSF[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 477.465 187.44 477.745 188.44 ;
    END
  END Data_PMOS_NOSF[15]
  PIN Data_PMOS_NOSF[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 476.905 187.44 477.185 188.44 ;
    END
  END Data_PMOS_NOSF[10]
  PIN Data_PMOS_NOSF[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 476.345 187.44 476.625 188.44 ;
    END
  END Data_PMOS_NOSF[4]
  PIN Data_PMOS_NOSF[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 475.785 187.44 476.065 188.44 ;
    END
  END Data_PMOS_NOSF[16]
  PIN Data_PMOS_NOSF[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 475.225 187.44 475.505 188.44 ;
    END
  END Data_PMOS_NOSF[11]
  PIN Data_PMOS_NOSF[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 474.665 187.44 474.945 188.44 ;
    END
  END Data_PMOS_NOSF[1]
  PIN Data_PMOS_NOSF[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 474.105 187.44 474.385 188.44 ;
    END
  END Data_PMOS_NOSF[0]
  PIN Data_PMOS_NOSF[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 473.545 187.44 473.825 188.44 ;
    END
  END Data_PMOS_NOSF[17]
  PIN DIG_MON_PMOS_NOSF[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 468.785 187.44 469.065 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[0]
  PIN Data_PMOS_NOSF[206]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1189.785 187.44 1190.065 188.44 ;
    END
  END Data_PMOS_NOSF[206]
  PIN FREEZE_PMOS_NOSF[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 721.625 187.44 721.905 188.44 ;
    END
  END FREEZE_PMOS_NOSF[3]
  PIN DIG_MON_PMOS_NOSF[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1558.265 187.44 1558.545 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[27]
  PIN Data_PMOS_NOSF[291]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1556.025 187.44 1556.305 188.44 ;
    END
  END Data_PMOS_NOSF[291]
  PIN Data_PMOS_NOSF[281]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1555.465 187.44 1555.745 188.44 ;
    END
  END Data_PMOS_NOSF[281]
  PIN Data_PMOS_NOSF[292]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1554.345 187.44 1554.625 188.44 ;
    END
  END Data_PMOS_NOSF[292]
  PIN Data_PMOS_NOSF[285]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1554.905 187.44 1555.185 188.44 ;
    END
  END Data_PMOS_NOSF[285]
  PIN Data_PMOS_NOSF[278]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1553.785 187.44 1554.065 188.44 ;
    END
  END Data_PMOS_NOSF[278]
  PIN Data_PMOS_NOSF[293]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1552.665 187.44 1552.945 188.44 ;
    END
  END Data_PMOS_NOSF[293]
  PIN Data_PMOS_NOSF[286]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1553.225 187.44 1553.505 188.44 ;
    END
  END Data_PMOS_NOSF[286]
  PIN Data_PMOS_NOSF[287]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1552.105 187.44 1552.385 188.44 ;
    END
  END Data_PMOS_NOSF[287]
  PIN Data_PMOS_NOSF[280]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1551.545 187.44 1551.825 188.44 ;
    END
  END Data_PMOS_NOSF[280]
  PIN Data_PMOS_NOSF[279]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1550.985 187.44 1551.265 188.44 ;
    END
  END Data_PMOS_NOSF[279]
  PIN nTOK_PMOS_NOSF[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1548.745 187.44 1549.025 188.44 ;
    END
  END nTOK_PMOS_NOSF[13]
  PIN FREEZE_PMOS_NOSF[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1532.505 187.44 1532.785 188.44 ;
    END
  END FREEZE_PMOS_NOSF[13]
  PIN Read_PMOS_NOSF[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1531.945 187.44 1532.225 188.44 ;
    END
  END Read_PMOS_NOSF[13]
  PIN Data_PMOS_NOSF[276]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1528.025 187.44 1528.305 188.44 ;
    END
  END Data_PMOS_NOSF[276]
  PIN Data_PMOS_NOSF[275]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1527.465 187.44 1527.745 188.44 ;
    END
  END Data_PMOS_NOSF[275]
  PIN Data_PMOS_NOSF[282]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1526.905 187.44 1527.185 188.44 ;
    END
  END Data_PMOS_NOSF[282]
  PIN Data_PMOS_NOSF[283]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1525.785 187.44 1526.065 188.44 ;
    END
  END Data_PMOS_NOSF[283]
  PIN Data_PMOS_NOSF[288]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1526.345 187.44 1526.625 188.44 ;
    END
  END Data_PMOS_NOSF[288]
  PIN Data_PMOS_NOSF[277]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1525.225 187.44 1525.505 188.44 ;
    END
  END Data_PMOS_NOSF[277]
  PIN Data_PMOS_NOSF[289]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1524.665 187.44 1524.945 188.44 ;
    END
  END Data_PMOS_NOSF[289]
  PIN Data_PMOS_NOSF[284]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1524.105 187.44 1524.385 188.44 ;
    END
  END Data_PMOS_NOSF[284]
  PIN Data_PMOS_NOSF[274]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1523.545 187.44 1523.825 188.44 ;
    END
  END Data_PMOS_NOSF[274]
  PIN Data_PMOS_NOSF[273]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1522.985 187.44 1523.265 188.44 ;
    END
  END Data_PMOS_NOSF[273]
  PIN Data_PMOS_NOSF[290]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1522.425 187.44 1522.705 188.44 ;
    END
  END Data_PMOS_NOSF[290]
  PIN DIG_MON_PMOS_NOSF[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1480.985 187.44 1481.265 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[26]
  PIN DIG_MON_PMOS_NOSF[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1476.505 187.44 1476.785 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[25]
  PIN Data_PMOS_NOSF[270]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1474.265 187.44 1474.545 188.44 ;
    END
  END Data_PMOS_NOSF[270]
  PIN Data_PMOS_NOSF[260]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1473.705 187.44 1473.985 188.44 ;
    END
  END Data_PMOS_NOSF[260]
  PIN Data_PMOS_NOSF[271]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1472.585 187.44 1472.865 188.44 ;
    END
  END Data_PMOS_NOSF[271]
  PIN Data_PMOS_NOSF[264]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1473.145 187.44 1473.425 188.44 ;
    END
  END Data_PMOS_NOSF[264]
  PIN Data_PMOS_NOSF[265]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1471.465 187.44 1471.745 188.44 ;
    END
  END Data_PMOS_NOSF[265]
  PIN Data_PMOS_NOSF[272]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1470.905 187.44 1471.185 188.44 ;
    END
  END Data_PMOS_NOSF[272]
  PIN Data_PMOS_NOSF[257]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1472.025 187.44 1472.305 188.44 ;
    END
  END Data_PMOS_NOSF[257]
  PIN Data_PMOS_NOSF[259]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1469.785 187.44 1470.065 188.44 ;
    END
  END Data_PMOS_NOSF[259]
  PIN Data_PMOS_NOSF[266]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1470.345 187.44 1470.625 188.44 ;
    END
  END Data_PMOS_NOSF[266]
  PIN Data_PMOS_NOSF[258]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1460.825 187.44 1461.105 188.44 ;
    END
  END Data_PMOS_NOSF[258]
  PIN nTOK_PMOS_NOSF[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1458.585 187.44 1458.865 188.44 ;
    END
  END nTOK_PMOS_NOSF[12]
  PIN FREEZE_PMOS_NOSF[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1455.785 187.44 1456.065 188.44 ;
    END
  END FREEZE_PMOS_NOSF[12]
  PIN Read_PMOS_NOSF[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1455.225 187.44 1455.505 188.44 ;
    END
  END Read_PMOS_NOSF[12]
  PIN Data_PMOS_NOSF[255]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1449.345 187.44 1449.625 188.44 ;
    END
  END Data_PMOS_NOSF[255]
  PIN Data_PMOS_NOSF[261]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1448.225 187.44 1448.505 188.44 ;
    END
  END Data_PMOS_NOSF[261]
  PIN Data_PMOS_NOSF[254]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1448.785 187.44 1449.065 188.44 ;
    END
  END Data_PMOS_NOSF[254]
  PIN Data_PMOS_NOSF[262]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1447.105 187.44 1447.385 188.44 ;
    END
  END Data_PMOS_NOSF[262]
  PIN Data_PMOS_NOSF[267]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1447.665 187.44 1447.945 188.44 ;
    END
  END Data_PMOS_NOSF[267]
  PIN Data_PMOS_NOSF[268]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1420.505 187.44 1420.785 188.44 ;
    END
  END Data_PMOS_NOSF[268]
  PIN Data_PMOS_NOSF[256]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1421.065 187.44 1421.345 188.44 ;
    END
  END Data_PMOS_NOSF[256]
  PIN Data_PMOS_NOSF[263]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1419.945 187.44 1420.225 188.44 ;
    END
  END Data_PMOS_NOSF[263]
  PIN Data_PMOS_NOSF[253]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1419.385 187.44 1419.665 188.44 ;
    END
  END Data_PMOS_NOSF[253]
  PIN Data_PMOS_NOSF[252]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1418.825 187.44 1419.105 188.44 ;
    END
  END Data_PMOS_NOSF[252]
  PIN Data_PMOS_NOSF[269]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1418.265 187.44 1418.545 188.44 ;
    END
  END Data_PMOS_NOSF[269]
  PIN DIG_MON_PMOS_NOSF[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1415.465 187.44 1415.745 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[24]
  PIN DIG_MON_PMOS_NOSF[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1410.985 187.44 1411.265 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[23]
  PIN Data_PMOS_NOSF[249]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1408.745 187.44 1409.025 188.44 ;
    END
  END Data_PMOS_NOSF[249]
  PIN Data_PMOS_NOSF[239]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1408.185 187.44 1408.465 188.44 ;
    END
  END Data_PMOS_NOSF[239]
  PIN Data_PMOS_NOSF[243]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1394.745 187.44 1395.025 188.44 ;
    END
  END Data_PMOS_NOSF[243]
  PIN Data_PMOS_NOSF[250]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1394.185 187.44 1394.465 188.44 ;
    END
  END Data_PMOS_NOSF[250]
  PIN Data_PMOS_NOSF[236]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1393.625 187.44 1393.905 188.44 ;
    END
  END Data_PMOS_NOSF[236]
  PIN Data_PMOS_NOSF[244]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1393.065 187.44 1393.345 188.44 ;
    END
  END Data_PMOS_NOSF[244]
  PIN Data_PMOS_NOSF[251]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1392.505 187.44 1392.785 188.44 ;
    END
  END Data_PMOS_NOSF[251]
  PIN Data_PMOS_NOSF[238]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1391.385 187.44 1391.665 188.44 ;
    END
  END Data_PMOS_NOSF[238]
  PIN Data_PMOS_NOSF[245]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1391.945 187.44 1392.225 188.44 ;
    END
  END Data_PMOS_NOSF[245]
  PIN Data_PMOS_NOSF[237]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1390.825 187.44 1391.105 188.44 ;
    END
  END Data_PMOS_NOSF[237]
  PIN nTOK_PMOS_NOSF[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1388.585 187.44 1388.865 188.44 ;
    END
  END nTOK_PMOS_NOSF[11]
  PIN Read_PMOS_NOSF[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1385.225 187.44 1385.505 188.44 ;
    END
  END Read_PMOS_NOSF[11]
  PIN FREEZE_PMOS_NOSF[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1385.785 187.44 1386.065 188.44 ;
    END
  END FREEZE_PMOS_NOSF[11]
  PIN Data_PMOS_NOSF[234]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1342.665 187.44 1342.945 188.44 ;
    END
  END Data_PMOS_NOSF[234]
  PIN Data_PMOS_NOSF[233]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1342.105 187.44 1342.385 188.44 ;
    END
  END Data_PMOS_NOSF[233]
  PIN Data_PMOS_NOSF[240]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1341.545 187.44 1341.825 188.44 ;
    END
  END Data_PMOS_NOSF[240]
  PIN Data_PMOS_NOSF[246]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1340.985 187.44 1341.265 188.44 ;
    END
  END Data_PMOS_NOSF[246]
  PIN Data_PMOS_NOSF[241]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1340.425 187.44 1340.705 188.44 ;
    END
  END Data_PMOS_NOSF[241]
  PIN Data_PMOS_NOSF[247]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1339.305 187.44 1339.585 188.44 ;
    END
  END Data_PMOS_NOSF[247]
  PIN Data_PMOS_NOSF[235]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1339.865 187.44 1340.145 188.44 ;
    END
  END Data_PMOS_NOSF[235]
  PIN Data_PMOS_NOSF[242]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1338.745 187.44 1339.025 188.44 ;
    END
  END Data_PMOS_NOSF[242]
  PIN Data_PMOS_NOSF[232]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1338.185 187.44 1338.465 188.44 ;
    END
  END Data_PMOS_NOSF[232]
  PIN Data_PMOS_NOSF[231]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1337.625 187.44 1337.905 188.44 ;
    END
  END Data_PMOS_NOSF[231]
  PIN Data_PMOS_NOSF[248]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1337.065 187.44 1337.345 188.44 ;
    END
  END Data_PMOS_NOSF[248]
  PIN DIG_MON_PMOS_NOSF[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1334.265 187.44 1334.545 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[22]
  PIN DIG_MON_PMOS_NOSF[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1329.785 187.44 1330.065 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[21]
  PIN Data_PMOS_NOSF[228]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1319.145 187.44 1319.425 188.44 ;
    END
  END Data_PMOS_NOSF[228]
  PIN Data_PMOS_NOSF[218]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1318.585 187.44 1318.865 188.44 ;
    END
  END Data_PMOS_NOSF[218]
  PIN Data_PMOS_NOSF[222]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1318.025 187.44 1318.305 188.44 ;
    END
  END Data_PMOS_NOSF[222]
  PIN Data_PMOS_NOSF[229]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1317.465 187.44 1317.745 188.44 ;
    END
  END Data_PMOS_NOSF[229]
  PIN Data_PMOS_NOSF[215]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1316.905 187.44 1317.185 188.44 ;
    END
  END Data_PMOS_NOSF[215]
  PIN Data_PMOS_NOSF[223]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1316.345 187.44 1316.625 188.44 ;
    END
  END Data_PMOS_NOSF[223]
  PIN Data_PMOS_NOSF[230]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1315.785 187.44 1316.065 188.44 ;
    END
  END Data_PMOS_NOSF[230]
  PIN Data_PMOS_NOSF[224]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1315.225 187.44 1315.505 188.44 ;
    END
  END Data_PMOS_NOSF[224]
  PIN Data_PMOS_NOSF[217]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1314.665 187.44 1314.945 188.44 ;
    END
  END Data_PMOS_NOSF[217]
  PIN Data_PMOS_NOSF[216]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1314.105 187.44 1314.385 188.44 ;
    END
  END Data_PMOS_NOSF[216]
  PIN nTOK_PMOS_NOSF[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1309.905 187.44 1310.185 188.44 ;
    END
  END nTOK_PMOS_NOSF[10]
  PIN Read_PMOS_NOSF[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1281.065 187.44 1281.345 188.44 ;
    END
  END Read_PMOS_NOSF[10]
  PIN Data_PMOS_NOSF[213]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1277.145 187.44 1277.425 188.44 ;
    END
  END Data_PMOS_NOSF[213]
  PIN Data_PMOS_NOSF[212]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1276.585 187.44 1276.865 188.44 ;
    END
  END Data_PMOS_NOSF[212]
  PIN Data_PMOS_NOSF[219]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1276.025 187.44 1276.305 188.44 ;
    END
  END Data_PMOS_NOSF[219]
  PIN Data_PMOS_NOSF[225]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1275.465 187.44 1275.745 188.44 ;
    END
  END Data_PMOS_NOSF[225]
  PIN Data_PMOS_NOSF[220]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1274.905 187.44 1275.185 188.44 ;
    END
  END Data_PMOS_NOSF[220]
  PIN Data_PMOS_NOSF[214]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1274.345 187.44 1274.625 188.44 ;
    END
  END Data_PMOS_NOSF[214]
  PIN Data_PMOS_NOSF[226]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1273.785 187.44 1274.065 188.44 ;
    END
  END Data_PMOS_NOSF[226]
  PIN Data_PMOS_NOSF[221]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1273.225 187.44 1273.505 188.44 ;
    END
  END Data_PMOS_NOSF[221]
  PIN Data_PMOS_NOSF[211]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1272.665 187.44 1272.945 188.44 ;
    END
  END Data_PMOS_NOSF[211]
  PIN Data_PMOS_NOSF[210]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1272.105 187.44 1272.385 188.44 ;
    END
  END Data_PMOS_NOSF[210]
  PIN Data_PMOS_NOSF[227]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1271.545 187.44 1271.825 188.44 ;
    END
  END Data_PMOS_NOSF[227]
  PIN DIG_MON_PMOS_NOSF[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1268.745 187.44 1269.025 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[20]
  PIN DIG_MON_PMOS_NOSF[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1251.385 187.44 1251.665 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[19]
  PIN Data_PMOS_NOSF[207]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1249.145 187.44 1249.425 188.44 ;
    END
  END Data_PMOS_NOSF[207]
  PIN Data_PMOS_NOSF[197]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1248.585 187.44 1248.865 188.44 ;
    END
  END Data_PMOS_NOSF[197]
  PIN Data_PMOS_NOSF[201]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1248.025 187.44 1248.305 188.44 ;
    END
  END Data_PMOS_NOSF[201]
  PIN Data_PMOS_NOSF[208]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1247.465 187.44 1247.745 188.44 ;
    END
  END Data_PMOS_NOSF[208]
  PIN Data_PMOS_NOSF[194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1246.905 187.44 1247.185 188.44 ;
    END
  END Data_PMOS_NOSF[194]
  PIN Data_PMOS_NOSF[202]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1246.345 187.44 1246.625 188.44 ;
    END
  END Data_PMOS_NOSF[202]
  PIN Data_PMOS_NOSF[209]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1245.785 187.44 1246.065 188.44 ;
    END
  END Data_PMOS_NOSF[209]
  PIN Data_PMOS_NOSF[203]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1245.225 187.44 1245.505 188.44 ;
    END
  END Data_PMOS_NOSF[203]
  PIN Data_PMOS_NOSF[196]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1244.665 187.44 1244.945 188.44 ;
    END
  END Data_PMOS_NOSF[196]
  PIN Data_PMOS_NOSF[195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1244.105 187.44 1244.385 188.44 ;
    END
  END Data_PMOS_NOSF[195]
  PIN nTOK_PMOS_NOSF[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1202.665 187.44 1202.945 188.44 ;
    END
  END nTOK_PMOS_NOSF[9]
  PIN FREEZE_PMOS_NOSF[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1199.865 187.44 1200.145 188.44 ;
    END
  END FREEZE_PMOS_NOSF[9]
  PIN Read_PMOS_NOSF[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1199.305 187.44 1199.585 188.44 ;
    END
  END Read_PMOS_NOSF[9]
  PIN Data_PMOS_NOSF[192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1195.385 187.44 1195.665 188.44 ;
    END
  END Data_PMOS_NOSF[192]
  PIN Data_PMOS_NOSF[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1194.825 187.44 1195.105 188.44 ;
    END
  END Data_PMOS_NOSF[191]
  PIN Data_PMOS_NOSF[198]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1194.265 187.44 1194.545 188.44 ;
    END
  END Data_PMOS_NOSF[198]
  PIN Data_PMOS_NOSF[204]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1193.705 187.44 1193.985 188.44 ;
    END
  END Data_PMOS_NOSF[204]
  PIN Data_PMOS_NOSF[199]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1193.145 187.44 1193.425 188.44 ;
    END
  END Data_PMOS_NOSF[199]
  PIN Data_PMOS_NOSF[193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1192.585 187.44 1192.865 188.44 ;
    END
  END Data_PMOS_NOSF[193]
  PIN Data_PMOS_NOSF[205]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1192.025 187.44 1192.305 188.44 ;
    END
  END Data_PMOS_NOSF[205]
  PIN Data_PMOS_NOSF[200]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1191.465 187.44 1191.745 188.44 ;
    END
  END Data_PMOS_NOSF[200]
  PIN Data_PMOS_NOSF[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1190.905 187.44 1191.185 188.44 ;
    END
  END Data_PMOS_NOSF[190]
  PIN Data_PMOS_NOSF[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1190.345 187.44 1190.625 188.44 ;
    END
  END Data_PMOS_NOSF[189]
  PIN Data_PMOS_NOSF[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1036.345 187.44 1036.625 188.44 ;
    END
  END Data_PMOS_NOSF[151]
  PIN DIG_MON_PMOS_NOSF[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1178.585 187.44 1178.865 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[18]
  PIN DIG_MON_PMOS_NOSF[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1174.105 187.44 1174.385 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[17]
  PIN Data_PMOS_NOSF[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1169.905 187.44 1170.185 188.44 ;
    END
  END Data_PMOS_NOSF[186]
  PIN Data_PMOS_NOSF[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1169.345 187.44 1169.625 188.44 ;
    END
  END Data_PMOS_NOSF[176]
  PIN Data_PMOS_NOSF[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1168.785 187.44 1169.065 188.44 ;
    END
  END Data_PMOS_NOSF[180]
  PIN Data_PMOS_NOSF[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1168.225 187.44 1168.505 188.44 ;
    END
  END Data_PMOS_NOSF[187]
  PIN Data_PMOS_NOSF[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1167.665 187.44 1167.945 188.44 ;
    END
  END Data_PMOS_NOSF[173]
  PIN Data_PMOS_NOSF[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1141.625 187.44 1141.905 188.44 ;
    END
  END Data_PMOS_NOSF[181]
  PIN Data_PMOS_NOSF[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1140.505 187.44 1140.785 188.44 ;
    END
  END Data_PMOS_NOSF[182]
  PIN Data_PMOS_NOSF[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1141.065 187.44 1141.345 188.44 ;
    END
  END Data_PMOS_NOSF[188]
  PIN Data_PMOS_NOSF[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1139.945 187.44 1140.225 188.44 ;
    END
  END Data_PMOS_NOSF[175]
  PIN Data_PMOS_NOSF[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1139.385 187.44 1139.665 188.44 ;
    END
  END Data_PMOS_NOSF[174]
  PIN nTOK_PMOS_NOSF[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1137.145 187.44 1137.425 188.44 ;
    END
  END nTOK_PMOS_NOSF[8]
  PIN FREEZE_PMOS_NOSF[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1134.345 187.44 1134.625 188.44 ;
    END
  END FREEZE_PMOS_NOSF[8]
  PIN Read_PMOS_NOSF[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1133.785 187.44 1134.065 188.44 ;
    END
  END Read_PMOS_NOSF[8]
  PIN Data_PMOS_NOSF[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1129.865 187.44 1130.145 188.44 ;
    END
  END Data_PMOS_NOSF[171]
  PIN Data_PMOS_NOSF[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1128.745 187.44 1129.025 188.44 ;
    END
  END Data_PMOS_NOSF[177]
  PIN Data_PMOS_NOSF[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1129.305 187.44 1129.585 188.44 ;
    END
  END Data_PMOS_NOSF[170]
  PIN Data_PMOS_NOSF[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1115.305 187.44 1115.585 188.44 ;
    END
  END Data_PMOS_NOSF[183]
  PIN Data_PMOS_NOSF[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1114.745 187.44 1115.025 188.44 ;
    END
  END Data_PMOS_NOSF[178]
  PIN Data_PMOS_NOSF[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1114.185 187.44 1114.465 188.44 ;
    END
  END Data_PMOS_NOSF[172]
  PIN Data_PMOS_NOSF[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1113.625 187.44 1113.905 188.44 ;
    END
  END Data_PMOS_NOSF[184]
  PIN Data_PMOS_NOSF[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1113.065 187.44 1113.345 188.44 ;
    END
  END Data_PMOS_NOSF[179]
  PIN Data_PMOS_NOSF[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1112.505 187.44 1112.785 188.44 ;
    END
  END Data_PMOS_NOSF[169]
  PIN Data_PMOS_NOSF[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1111.945 187.44 1112.225 188.44 ;
    END
  END Data_PMOS_NOSF[168]
  PIN Data_PMOS_NOSF[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1111.385 187.44 1111.665 188.44 ;
    END
  END Data_PMOS_NOSF[185]
  PIN DIG_MON_PMOS_NOSF[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1108.585 187.44 1108.865 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[16]
  PIN DIG_MON_PMOS_NOSF[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1104.105 187.44 1104.385 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[15]
  PIN Data_PMOS_NOSF[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1062.105 187.44 1062.385 188.44 ;
    END
  END Data_PMOS_NOSF[165]
  PIN Data_PMOS_NOSF[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1061.545 187.44 1061.825 188.44 ;
    END
  END Data_PMOS_NOSF[155]
  PIN Data_PMOS_NOSF[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1060.985 187.44 1061.265 188.44 ;
    END
  END Data_PMOS_NOSF[159]
  PIN Data_PMOS_NOSF[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1060.425 187.44 1060.705 188.44 ;
    END
  END Data_PMOS_NOSF[166]
  PIN Data_PMOS_NOSF[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1059.865 187.44 1060.145 188.44 ;
    END
  END Data_PMOS_NOSF[152]
  PIN Data_PMOS_NOSF[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1059.305 187.44 1059.585 188.44 ;
    END
  END Data_PMOS_NOSF[160]
  PIN Data_PMOS_NOSF[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1058.745 187.44 1059.025 188.44 ;
    END
  END Data_PMOS_NOSF[167]
  PIN Data_PMOS_NOSF[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1058.185 187.44 1058.465 188.44 ;
    END
  END Data_PMOS_NOSF[161]
  PIN Data_PMOS_NOSF[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1057.625 187.44 1057.905 188.44 ;
    END
  END Data_PMOS_NOSF[154]
  PIN Data_PMOS_NOSF[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1057.065 187.44 1057.345 188.44 ;
    END
  END Data_PMOS_NOSF[153]
  PIN nTOK_PMOS_NOSF[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1054.825 187.44 1055.105 188.44 ;
    END
  END nTOK_PMOS_NOSF[7]
  PIN FREEZE_PMOS_NOSF[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1052.025 187.44 1052.305 188.44 ;
    END
  END FREEZE_PMOS_NOSF[7]
  PIN Read_PMOS_NOSF[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1051.465 187.44 1051.745 188.44 ;
    END
  END Read_PMOS_NOSF[7]
  PIN Data_PMOS_NOSF[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1039.145 187.44 1039.425 188.44 ;
    END
  END Data_PMOS_NOSF[150]
  PIN Data_PMOS_NOSF[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1038.585 187.44 1038.865 188.44 ;
    END
  END Data_PMOS_NOSF[149]
  PIN Data_PMOS_NOSF[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1038.025 187.44 1038.305 188.44 ;
    END
  END Data_PMOS_NOSF[156]
  PIN Data_PMOS_NOSF[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1037.465 187.44 1037.745 188.44 ;
    END
  END Data_PMOS_NOSF[162]
  PIN Data_PMOS_NOSF[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1036.905 187.44 1037.185 188.44 ;
    END
  END Data_PMOS_NOSF[157]
  PIN Data_PMOS_NOSF[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1035.785 187.44 1036.065 188.44 ;
    END
  END Data_PMOS_NOSF[163]
  PIN Data_PMOS_NOSF[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1035.225 187.44 1035.505 188.44 ;
    END
  END Data_PMOS_NOSF[158]
  PIN Data_PMOS_NOSF[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1034.665 187.44 1034.945 188.44 ;
    END
  END Data_PMOS_NOSF[148]
  PIN Data_PMOS_NOSF[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1034.105 187.44 1034.385 188.44 ;
    END
  END Data_PMOS_NOSF[147]
  PIN Data_PMOS_NOSF[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1033.545 187.44 1033.825 188.44 ;
    END
  END Data_PMOS_NOSF[164]
  PIN Data_PMOS_NOSF[351]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1753.705 187.44 1753.985 188.44 ;
    END
  END Data_PMOS_NOSF[351]
  PIN DIG_MON_PMOS_NOSF[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1028.785 187.44 1029.065 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[14]
  PIN FREEZE_PMOS_NOSF[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1281.625 187.44 1281.905 188.44 ;
    END
  END FREEZE_PMOS_NOSF[10]
  PIN DIG_MON_PMOS_NOSF[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2118.265 187.44 2118.545 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[41]
  PIN Data_PMOS_NOSF[438]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2116.025 187.44 2116.305 188.44 ;
    END
  END Data_PMOS_NOSF[438]
  PIN Data_PMOS_NOSF[428]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2115.465 187.44 2115.745 188.44 ;
    END
  END Data_PMOS_NOSF[428]
  PIN Data_PMOS_NOSF[432]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2114.905 187.44 2115.185 188.44 ;
    END
  END Data_PMOS_NOSF[432]
  PIN Data_PMOS_NOSF[439]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2114.345 187.44 2114.625 188.44 ;
    END
  END Data_PMOS_NOSF[439]
  PIN Data_PMOS_NOSF[425]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2113.785 187.44 2114.065 188.44 ;
    END
  END Data_PMOS_NOSF[425]
  PIN Data_PMOS_NOSF[433]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2113.225 187.44 2113.505 188.44 ;
    END
  END Data_PMOS_NOSF[433]
  PIN Data_PMOS_NOSF[440]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2112.665 187.44 2112.945 188.44 ;
    END
  END Data_PMOS_NOSF[440]
  PIN Data_PMOS_NOSF[434]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2112.105 187.44 2112.385 188.44 ;
    END
  END Data_PMOS_NOSF[434]
  PIN Data_PMOS_NOSF[427]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2111.545 187.44 2111.825 188.44 ;
    END
  END Data_PMOS_NOSF[427]
  PIN Data_PMOS_NOSF[426]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2110.985 187.44 2111.265 188.44 ;
    END
  END Data_PMOS_NOSF[426]
  PIN nTOK_PMOS_NOSF[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2108.745 187.44 2109.025 188.44 ;
    END
  END nTOK_PMOS_NOSF[20]
  PIN Read_PMOS_NOSF[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2091.945 187.44 2092.225 188.44 ;
    END
  END Read_PMOS_NOSF[20]
  PIN FREEZE_PMOS_NOSF[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2092.505 187.44 2092.785 188.44 ;
    END
  END FREEZE_PMOS_NOSF[20]
  PIN Data_PMOS_NOSF[423]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2088.025 187.44 2088.305 188.44 ;
    END
  END Data_PMOS_NOSF[423]
  PIN Data_PMOS_NOSF[422]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2087.465 187.44 2087.745 188.44 ;
    END
  END Data_PMOS_NOSF[422]
  PIN Data_PMOS_NOSF[429]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2086.905 187.44 2087.185 188.44 ;
    END
  END Data_PMOS_NOSF[429]
  PIN Data_PMOS_NOSF[430]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2085.785 187.44 2086.065 188.44 ;
    END
  END Data_PMOS_NOSF[430]
  PIN Data_PMOS_NOSF[435]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2086.345 187.44 2086.625 188.44 ;
    END
  END Data_PMOS_NOSF[435]
  PIN Data_PMOS_NOSF[436]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2084.665 187.44 2084.945 188.44 ;
    END
  END Data_PMOS_NOSF[436]
  PIN Data_PMOS_NOSF[431]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2084.105 187.44 2084.385 188.44 ;
    END
  END Data_PMOS_NOSF[431]
  PIN Data_PMOS_NOSF[421]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2083.545 187.44 2083.825 188.44 ;
    END
  END Data_PMOS_NOSF[421]
  PIN Data_PMOS_NOSF[420]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2082.985 187.44 2083.265 188.44 ;
    END
  END Data_PMOS_NOSF[420]
  PIN Data_PMOS_NOSF[437]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2082.425 187.44 2082.705 188.44 ;
    END
  END Data_PMOS_NOSF[437]
  PIN Data_PMOS_NOSF[424]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2085.225 187.44 2085.505 188.44 ;
    END
  END Data_PMOS_NOSF[424]
  PIN DIG_MON_PMOS_NOSF[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2040.985 187.44 2041.265 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[40]
  PIN DIG_MON_PMOS_NOSF[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2036.505 187.44 2036.785 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[39]
  PIN Data_PMOS_NOSF[417]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2034.265 187.44 2034.545 188.44 ;
    END
  END Data_PMOS_NOSF[417]
  PIN Data_PMOS_NOSF[407]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2033.705 187.44 2033.985 188.44 ;
    END
  END Data_PMOS_NOSF[407]
  PIN Data_PMOS_NOSF[418]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2032.585 187.44 2032.865 188.44 ;
    END
  END Data_PMOS_NOSF[418]
  PIN Data_PMOS_NOSF[404]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2032.025 187.44 2032.305 188.44 ;
    END
  END Data_PMOS_NOSF[404]
  PIN Data_PMOS_NOSF[419]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2030.905 187.44 2031.185 188.44 ;
    END
  END Data_PMOS_NOSF[419]
  PIN Data_PMOS_NOSF[412]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2031.465 187.44 2031.745 188.44 ;
    END
  END Data_PMOS_NOSF[412]
  PIN Data_PMOS_NOSF[406]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2029.785 187.44 2030.065 188.44 ;
    END
  END Data_PMOS_NOSF[406]
  PIN Data_PMOS_NOSF[411]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2033.145 187.44 2033.425 188.44 ;
    END
  END Data_PMOS_NOSF[411]
  PIN Data_PMOS_NOSF[413]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2030.345 187.44 2030.625 188.44 ;
    END
  END Data_PMOS_NOSF[413]
  PIN Data_PMOS_NOSF[405]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2020.825 187.44 2021.105 188.44 ;
    END
  END Data_PMOS_NOSF[405]
  PIN nTOK_PMOS_NOSF[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2018.585 187.44 2018.865 188.44 ;
    END
  END nTOK_PMOS_NOSF[19]
  PIN FREEZE_PMOS_NOSF[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2015.785 187.44 2016.065 188.44 ;
    END
  END FREEZE_PMOS_NOSF[19]
  PIN Read_PMOS_NOSF[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2015.225 187.44 2015.505 188.44 ;
    END
  END Read_PMOS_NOSF[19]
  PIN Data_PMOS_NOSF[402]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2009.345 187.44 2009.625 188.44 ;
    END
  END Data_PMOS_NOSF[402]
  PIN Data_PMOS_NOSF[355]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1807.465 187.44 1807.745 188.44 ;
    END
  END Data_PMOS_NOSF[355]
  PIN Data_PMOS_NOSF[401]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2008.785 187.44 2009.065 188.44 ;
    END
  END Data_PMOS_NOSF[401]
  PIN Data_PMOS_NOSF[408]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2008.225 187.44 2008.505 188.44 ;
    END
  END Data_PMOS_NOSF[408]
  PIN Data_PMOS_NOSF[409]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2007.105 187.44 2007.385 188.44 ;
    END
  END Data_PMOS_NOSF[409]
  PIN Data_PMOS_NOSF[414]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2007.665 187.44 2007.945 188.44 ;
    END
  END Data_PMOS_NOSF[414]
  PIN Data_PMOS_NOSF[415]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1980.505 187.44 1980.785 188.44 ;
    END
  END Data_PMOS_NOSF[415]
  PIN Data_PMOS_NOSF[403]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1981.065 187.44 1981.345 188.44 ;
    END
  END Data_PMOS_NOSF[403]
  PIN Data_PMOS_NOSF[410]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1979.945 187.44 1980.225 188.44 ;
    END
  END Data_PMOS_NOSF[410]
  PIN Data_PMOS_NOSF[400]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1979.385 187.44 1979.665 188.44 ;
    END
  END Data_PMOS_NOSF[400]
  PIN Data_PMOS_NOSF[399]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1978.825 187.44 1979.105 188.44 ;
    END
  END Data_PMOS_NOSF[399]
  PIN Data_PMOS_NOSF[416]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1978.265 187.44 1978.545 188.44 ;
    END
  END Data_PMOS_NOSF[416]
  PIN DIG_MON_PMOS_NOSF[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1975.465 187.44 1975.745 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[38]
  PIN DIG_MON_PMOS_NOSF[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1970.985 187.44 1971.265 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[37]
  PIN Data_PMOS_NOSF[386]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1968.185 187.44 1968.465 188.44 ;
    END
  END Data_PMOS_NOSF[386]
  PIN Data_PMOS_NOSF[396]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1968.745 187.44 1969.025 188.44 ;
    END
  END Data_PMOS_NOSF[396]
  PIN Data_PMOS_NOSF[390]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1954.745 187.44 1955.025 188.44 ;
    END
  END Data_PMOS_NOSF[390]
  PIN Data_PMOS_NOSF[397]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1954.185 187.44 1954.465 188.44 ;
    END
  END Data_PMOS_NOSF[397]
  PIN Data_PMOS_NOSF[383]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1953.625 187.44 1953.905 188.44 ;
    END
  END Data_PMOS_NOSF[383]
  PIN Data_PMOS_NOSF[391]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1953.065 187.44 1953.345 188.44 ;
    END
  END Data_PMOS_NOSF[391]
  PIN Data_PMOS_NOSF[398]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1952.505 187.44 1952.785 188.44 ;
    END
  END Data_PMOS_NOSF[398]
  PIN Data_PMOS_NOSF[392]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1951.945 187.44 1952.225 188.44 ;
    END
  END Data_PMOS_NOSF[392]
  PIN Data_PMOS_NOSF[385]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1951.385 187.44 1951.665 188.44 ;
    END
  END Data_PMOS_NOSF[385]
  PIN Data_PMOS_NOSF[384]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1950.825 187.44 1951.105 188.44 ;
    END
  END Data_PMOS_NOSF[384]
  PIN nTOK_PMOS_NOSF[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1948.585 187.44 1948.865 188.44 ;
    END
  END nTOK_PMOS_NOSF[18]
  PIN FREEZE_PMOS_NOSF[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1945.785 187.44 1946.065 188.44 ;
    END
  END FREEZE_PMOS_NOSF[18]
  PIN Read_PMOS_NOSF[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1945.225 187.44 1945.505 188.44 ;
    END
  END Read_PMOS_NOSF[18]
  PIN Data_PMOS_NOSF[381]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1902.665 187.44 1902.945 188.44 ;
    END
  END Data_PMOS_NOSF[381]
  PIN Data_PMOS_NOSF[380]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1902.105 187.44 1902.385 188.44 ;
    END
  END Data_PMOS_NOSF[380]
  PIN Data_PMOS_NOSF[387]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1901.545 187.44 1901.825 188.44 ;
    END
  END Data_PMOS_NOSF[387]
  PIN Data_PMOS_NOSF[393]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1900.985 187.44 1901.265 188.44 ;
    END
  END Data_PMOS_NOSF[393]
  PIN Data_PMOS_NOSF[388]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1900.425 187.44 1900.705 188.44 ;
    END
  END Data_PMOS_NOSF[388]
  PIN Data_PMOS_NOSF[382]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1899.865 187.44 1900.145 188.44 ;
    END
  END Data_PMOS_NOSF[382]
  PIN Data_PMOS_NOSF[394]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1899.305 187.44 1899.585 188.44 ;
    END
  END Data_PMOS_NOSF[394]
  PIN Data_PMOS_NOSF[389]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1898.745 187.44 1899.025 188.44 ;
    END
  END Data_PMOS_NOSF[389]
  PIN Data_PMOS_NOSF[379]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1898.185 187.44 1898.465 188.44 ;
    END
  END Data_PMOS_NOSF[379]
  PIN Data_PMOS_NOSF[378]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1897.625 187.44 1897.905 188.44 ;
    END
  END Data_PMOS_NOSF[378]
  PIN Data_PMOS_NOSF[395]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1897.065 187.44 1897.345 188.44 ;
    END
  END Data_PMOS_NOSF[395]
  PIN DIG_MON_PMOS_NOSF[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1894.265 187.44 1894.545 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[36]
  PIN DIG_MON_PMOS_NOSF[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1889.785 187.44 1890.065 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[35]
  PIN Data_PMOS_NOSF[375]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1879.145 187.44 1879.425 188.44 ;
    END
  END Data_PMOS_NOSF[375]
  PIN Data_PMOS_NOSF[365]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1878.585 187.44 1878.865 188.44 ;
    END
  END Data_PMOS_NOSF[365]
  PIN Data_PMOS_NOSF[369]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1878.025 187.44 1878.305 188.44 ;
    END
  END Data_PMOS_NOSF[369]
  PIN Data_PMOS_NOSF[376]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1877.465 187.44 1877.745 188.44 ;
    END
  END Data_PMOS_NOSF[376]
  PIN Data_PMOS_NOSF[362]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1876.905 187.44 1877.185 188.44 ;
    END
  END Data_PMOS_NOSF[362]
  PIN Data_PMOS_NOSF[370]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1876.345 187.44 1876.625 188.44 ;
    END
  END Data_PMOS_NOSF[370]
  PIN Data_PMOS_NOSF[377]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1875.785 187.44 1876.065 188.44 ;
    END
  END Data_PMOS_NOSF[377]
  PIN Data_PMOS_NOSF[371]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1875.225 187.44 1875.505 188.44 ;
    END
  END Data_PMOS_NOSF[371]
  PIN Data_PMOS_NOSF[364]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1874.665 187.44 1874.945 188.44 ;
    END
  END Data_PMOS_NOSF[364]
  PIN Data_PMOS_NOSF[363]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1874.105 187.44 1874.385 188.44 ;
    END
  END Data_PMOS_NOSF[363]
  PIN nTOK_PMOS_NOSF[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1869.905 187.44 1870.185 188.44 ;
    END
  END nTOK_PMOS_NOSF[17]
  PIN Read_PMOS_NOSF[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1841.065 187.44 1841.345 188.44 ;
    END
  END Read_PMOS_NOSF[17]
  PIN Data_PMOS_NOSF[360]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1837.145 187.44 1837.425 188.44 ;
    END
  END Data_PMOS_NOSF[360]
  PIN Data_PMOS_NOSF[359]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1836.585 187.44 1836.865 188.44 ;
    END
  END Data_PMOS_NOSF[359]
  PIN Data_PMOS_NOSF[366]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1836.025 187.44 1836.305 188.44 ;
    END
  END Data_PMOS_NOSF[366]
  PIN Data_PMOS_NOSF[372]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1835.465 187.44 1835.745 188.44 ;
    END
  END Data_PMOS_NOSF[372]
  PIN Data_PMOS_NOSF[367]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1834.905 187.44 1835.185 188.44 ;
    END
  END Data_PMOS_NOSF[367]
  PIN Data_PMOS_NOSF[361]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1834.345 187.44 1834.625 188.44 ;
    END
  END Data_PMOS_NOSF[361]
  PIN Data_PMOS_NOSF[368]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1833.225 187.44 1833.505 188.44 ;
    END
  END Data_PMOS_NOSF[368]
  PIN Data_PMOS_NOSF[358]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1832.665 187.44 1832.945 188.44 ;
    END
  END Data_PMOS_NOSF[358]
  PIN Data_PMOS_NOSF[357]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1832.105 187.44 1832.385 188.44 ;
    END
  END Data_PMOS_NOSF[357]
  PIN Data_PMOS_NOSF[374]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1831.545 187.44 1831.825 188.44 ;
    END
  END Data_PMOS_NOSF[374]
  PIN Data_PMOS_NOSF[373]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1833.785 187.44 1834.065 188.44 ;
    END
  END Data_PMOS_NOSF[373]
  PIN DIG_MON_PMOS_NOSF[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1828.745 187.44 1829.025 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[34]
  PIN DIG_MON_PMOS_NOSF[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1811.385 187.44 1811.665 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[33]
  PIN Data_PMOS_NOSF[344]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1808.585 187.44 1808.865 188.44 ;
    END
  END Data_PMOS_NOSF[344]
  PIN Data_PMOS_NOSF[354]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1809.145 187.44 1809.425 188.44 ;
    END
  END Data_PMOS_NOSF[354]
  PIN Data_PMOS_NOSF[341]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1806.905 187.44 1807.185 188.44 ;
    END
  END Data_PMOS_NOSF[341]
  PIN Data_PMOS_NOSF[349]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1806.345 187.44 1806.625 188.44 ;
    END
  END Data_PMOS_NOSF[349]
  PIN Data_PMOS_NOSF[350]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1805.225 187.44 1805.505 188.44 ;
    END
  END Data_PMOS_NOSF[350]
  PIN Data_PMOS_NOSF[356]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1805.785 187.44 1806.065 188.44 ;
    END
  END Data_PMOS_NOSF[356]
  PIN Data_PMOS_NOSF[343]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1804.665 187.44 1804.945 188.44 ;
    END
  END Data_PMOS_NOSF[343]
  PIN Data_PMOS_NOSF[342]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1804.105 187.44 1804.385 188.44 ;
    END
  END Data_PMOS_NOSF[342]
  PIN Data_PMOS_NOSF[348]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1808.025 187.44 1808.305 188.44 ;
    END
  END Data_PMOS_NOSF[348]
  PIN nTOK_PMOS_NOSF[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1762.665 187.44 1762.945 188.44 ;
    END
  END nTOK_PMOS_NOSF[16]
  PIN FREEZE_PMOS_NOSF[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1759.865 187.44 1760.145 188.44 ;
    END
  END FREEZE_PMOS_NOSF[16]
  PIN Read_PMOS_NOSF[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1759.305 187.44 1759.585 188.44 ;
    END
  END Read_PMOS_NOSF[16]
  PIN Data_PMOS_NOSF[339]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1755.385 187.44 1755.665 188.44 ;
    END
  END Data_PMOS_NOSF[339]
  PIN Data_PMOS_NOSF[338]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1754.825 187.44 1755.105 188.44 ;
    END
  END Data_PMOS_NOSF[338]
  PIN Data_PMOS_NOSF[345]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1754.265 187.44 1754.545 188.44 ;
    END
  END Data_PMOS_NOSF[345]
  PIN Data_PMOS_NOSF[346]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1753.145 187.44 1753.425 188.44 ;
    END
  END Data_PMOS_NOSF[346]
  PIN Data_PMOS_NOSF[340]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1752.585 187.44 1752.865 188.44 ;
    END
  END Data_PMOS_NOSF[340]
  PIN Data_PMOS_NOSF[347]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1751.465 187.44 1751.745 188.44 ;
    END
  END Data_PMOS_NOSF[347]
  PIN Data_PMOS_NOSF[352]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1752.025 187.44 1752.305 188.44 ;
    END
  END Data_PMOS_NOSF[352]
  PIN Data_PMOS_NOSF[337]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1750.905 187.44 1751.185 188.44 ;
    END
  END Data_PMOS_NOSF[337]
  PIN Data_PMOS_NOSF[336]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1750.345 187.44 1750.625 188.44 ;
    END
  END Data_PMOS_NOSF[336]
  PIN Data_PMOS_NOSF[353]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1749.785 187.44 1750.065 188.44 ;
    END
  END Data_PMOS_NOSF[353]
  PIN DIG_MON_PMOS_NOSF[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1738.585 187.44 1738.865 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[32]
  PIN DIG_MON_PMOS_NOSF[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1734.105 187.44 1734.385 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[31]
  PIN Data_PMOS_NOSF[333]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1729.905 187.44 1730.185 188.44 ;
    END
  END Data_PMOS_NOSF[333]
  PIN Data_PMOS_NOSF[323]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1729.345 187.44 1729.625 188.44 ;
    END
  END Data_PMOS_NOSF[323]
  PIN Data_PMOS_NOSF[334]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1728.225 187.44 1728.505 188.44 ;
    END
  END Data_PMOS_NOSF[334]
  PIN Data_PMOS_NOSF[327]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1728.785 187.44 1729.065 188.44 ;
    END
  END Data_PMOS_NOSF[327]
  PIN Data_PMOS_NOSF[328]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1701.625 187.44 1701.905 188.44 ;
    END
  END Data_PMOS_NOSF[328]
  PIN Data_PMOS_NOSF[335]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1701.065 187.44 1701.345 188.44 ;
    END
  END Data_PMOS_NOSF[335]
  PIN Data_PMOS_NOSF[320]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1727.665 187.44 1727.945 188.44 ;
    END
  END Data_PMOS_NOSF[320]
  PIN Data_PMOS_NOSF[322]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1699.945 187.44 1700.225 188.44 ;
    END
  END Data_PMOS_NOSF[322]
  PIN Data_PMOS_NOSF[321]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1699.385 187.44 1699.665 188.44 ;
    END
  END Data_PMOS_NOSF[321]
  PIN nTOK_PMOS_NOSF[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1697.145 187.44 1697.425 188.44 ;
    END
  END nTOK_PMOS_NOSF[15]
  PIN Data_PMOS_NOSF[329]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1700.505 187.44 1700.785 188.44 ;
    END
  END Data_PMOS_NOSF[329]
  PIN FREEZE_PMOS_NOSF[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1694.345 187.44 1694.625 188.44 ;
    END
  END FREEZE_PMOS_NOSF[15]
  PIN Read_PMOS_NOSF[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1693.785 187.44 1694.065 188.44 ;
    END
  END Read_PMOS_NOSF[15]
  PIN Data_PMOS_NOSF[318]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1689.865 187.44 1690.145 188.44 ;
    END
  END Data_PMOS_NOSF[318]
  PIN Data_PMOS_NOSF[317]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1689.305 187.44 1689.585 188.44 ;
    END
  END Data_PMOS_NOSF[317]
  PIN Data_PMOS_NOSF[324]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1688.745 187.44 1689.025 188.44 ;
    END
  END Data_PMOS_NOSF[324]
  PIN Data_PMOS_NOSF[325]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1674.745 187.44 1675.025 188.44 ;
    END
  END Data_PMOS_NOSF[325]
  PIN Data_PMOS_NOSF[330]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1675.305 187.44 1675.585 188.44 ;
    END
  END Data_PMOS_NOSF[330]
  PIN Data_PMOS_NOSF[319]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1674.185 187.44 1674.465 188.44 ;
    END
  END Data_PMOS_NOSF[319]
  PIN Data_PMOS_NOSF[331]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1673.625 187.44 1673.905 188.44 ;
    END
  END Data_PMOS_NOSF[331]
  PIN Data_PMOS_NOSF[326]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1673.065 187.44 1673.345 188.44 ;
    END
  END Data_PMOS_NOSF[326]
  PIN Data_PMOS_NOSF[316]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1672.505 187.44 1672.785 188.44 ;
    END
  END Data_PMOS_NOSF[316]
  PIN Data_PMOS_NOSF[332]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1671.385 187.44 1671.665 188.44 ;
    END
  END Data_PMOS_NOSF[332]
  PIN Data_PMOS_NOSF[315]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1671.945 187.44 1672.225 188.44 ;
    END
  END Data_PMOS_NOSF[315]
  PIN DIG_MON_PMOS_NOSF[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1668.585 187.44 1668.865 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[30]
  PIN DIG_MON_PMOS_NOSF[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1664.105 187.44 1664.385 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[29]
  PIN Data_PMOS_NOSF[312]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1622.105 187.44 1622.385 188.44 ;
    END
  END Data_PMOS_NOSF[312]
  PIN Data_PMOS_NOSF[302]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1621.545 187.44 1621.825 188.44 ;
    END
  END Data_PMOS_NOSF[302]
  PIN Data_PMOS_NOSF[306]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1620.985 187.44 1621.265 188.44 ;
    END
  END Data_PMOS_NOSF[306]
  PIN Data_PMOS_NOSF[313]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1620.425 187.44 1620.705 188.44 ;
    END
  END Data_PMOS_NOSF[313]
  PIN Data_PMOS_NOSF[299]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1619.865 187.44 1620.145 188.44 ;
    END
  END Data_PMOS_NOSF[299]
  PIN Data_PMOS_NOSF[307]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1619.305 187.44 1619.585 188.44 ;
    END
  END Data_PMOS_NOSF[307]
  PIN Data_PMOS_NOSF[314]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1618.745 187.44 1619.025 188.44 ;
    END
  END Data_PMOS_NOSF[314]
  PIN Data_PMOS_NOSF[308]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1618.185 187.44 1618.465 188.44 ;
    END
  END Data_PMOS_NOSF[308]
  PIN Data_PMOS_NOSF[301]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1617.625 187.44 1617.905 188.44 ;
    END
  END Data_PMOS_NOSF[301]
  PIN Data_PMOS_NOSF[300]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1617.065 187.44 1617.345 188.44 ;
    END
  END Data_PMOS_NOSF[300]
  PIN nTOK_PMOS_NOSF[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1614.825 187.44 1615.105 188.44 ;
    END
  END nTOK_PMOS_NOSF[14]
  PIN FREEZE_PMOS_NOSF[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1612.025 187.44 1612.305 188.44 ;
    END
  END FREEZE_PMOS_NOSF[14]
  PIN Read_PMOS_NOSF[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1611.465 187.44 1611.745 188.44 ;
    END
  END Read_PMOS_NOSF[14]
  PIN Data_PMOS_NOSF[297]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1599.145 187.44 1599.425 188.44 ;
    END
  END Data_PMOS_NOSF[297]
  PIN Data_PMOS_NOSF[296]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1598.585 187.44 1598.865 188.44 ;
    END
  END Data_PMOS_NOSF[296]
  PIN Data_PMOS_NOSF[309]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1597.465 187.44 1597.745 188.44 ;
    END
  END Data_PMOS_NOSF[309]
  PIN Data_PMOS_NOSF[303]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1598.025 187.44 1598.305 188.44 ;
    END
  END Data_PMOS_NOSF[303]
  PIN Data_PMOS_NOSF[304]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1596.905 187.44 1597.185 188.44 ;
    END
  END Data_PMOS_NOSF[304]
  PIN Data_PMOS_NOSF[298]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1596.345 187.44 1596.625 188.44 ;
    END
  END Data_PMOS_NOSF[298]
  PIN Data_PMOS_NOSF[310]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1595.785 187.44 1596.065 188.44 ;
    END
  END Data_PMOS_NOSF[310]
  PIN Data_PMOS_NOSF[305]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1595.225 187.44 1595.505 188.44 ;
    END
  END Data_PMOS_NOSF[305]
  PIN Data_PMOS_NOSF[295]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1594.665 187.44 1594.945 188.44 ;
    END
  END Data_PMOS_NOSF[295]
  PIN Data_PMOS_NOSF[294]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1594.105 187.44 1594.385 188.44 ;
    END
  END Data_PMOS_NOSF[294]
  PIN Data_PMOS_NOSF[311]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1593.545 187.44 1593.825 188.44 ;
    END
  END Data_PMOS_NOSF[311]
  PIN DIG_MON_PMOS_NOSF[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1588.785 187.44 1589.065 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[28]
  PIN FREEZE_PMOS_NOSF[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1841.625 187.44 1841.905 188.44 ;
    END
  END FREEZE_PMOS_NOSF[17]
  PIN DIG_MON_PMOS_NOSF[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2678.265 187.44 2678.545 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[55]
  PIN Data_PMOS_NOSF[585]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2676.025 187.44 2676.305 188.44 ;
    END
  END Data_PMOS_NOSF[585]
  PIN Data_PMOS_NOSF[575]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2675.465 187.44 2675.745 188.44 ;
    END
  END Data_PMOS_NOSF[575]
  PIN Data_PMOS_NOSF[579]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2674.905 187.44 2675.185 188.44 ;
    END
  END Data_PMOS_NOSF[579]
  PIN Data_PMOS_NOSF[586]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2674.345 187.44 2674.625 188.44 ;
    END
  END Data_PMOS_NOSF[586]
  PIN Data_PMOS_NOSF[572]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2673.785 187.44 2674.065 188.44 ;
    END
  END Data_PMOS_NOSF[572]
  PIN Data_PMOS_NOSF[580]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2673.225 187.44 2673.505 188.44 ;
    END
  END Data_PMOS_NOSF[580]
  PIN Data_PMOS_NOSF[587]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2672.665 187.44 2672.945 188.44 ;
    END
  END Data_PMOS_NOSF[587]
  PIN Data_PMOS_NOSF[581]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2672.105 187.44 2672.385 188.44 ;
    END
  END Data_PMOS_NOSF[581]
  PIN Data_PMOS_NOSF[574]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2671.545 187.44 2671.825 188.44 ;
    END
  END Data_PMOS_NOSF[574]
  PIN Data_PMOS_NOSF[573]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2670.985 187.44 2671.265 188.44 ;
    END
  END Data_PMOS_NOSF[573]
  PIN nTOK_PMOS_NOSF[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2668.745 187.44 2669.025 188.44 ;
    END
  END nTOK_PMOS_NOSF[27]
  PIN FREEZE_PMOS_NOSF[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2652.505 187.44 2652.785 188.44 ;
    END
  END FREEZE_PMOS_NOSF[27]
  PIN Read_PMOS_NOSF[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2651.945 187.44 2652.225 188.44 ;
    END
  END Read_PMOS_NOSF[27]
  PIN Data_PMOS_NOSF[569]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2647.465 187.44 2647.745 188.44 ;
    END
  END Data_PMOS_NOSF[569]
  PIN Data_PMOS_NOSF[576]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2646.905 187.44 2647.185 188.44 ;
    END
  END Data_PMOS_NOSF[576]
  PIN Data_PMOS_NOSF[582]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2646.345 187.44 2646.625 188.44 ;
    END
  END Data_PMOS_NOSF[582]
  PIN Data_PMOS_NOSF[577]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2645.785 187.44 2646.065 188.44 ;
    END
  END Data_PMOS_NOSF[577]
  PIN Data_PMOS_NOSF[571]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2645.225 187.44 2645.505 188.44 ;
    END
  END Data_PMOS_NOSF[571]
  PIN Data_PMOS_NOSF[583]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2644.665 187.44 2644.945 188.44 ;
    END
  END Data_PMOS_NOSF[583]
  PIN Data_PMOS_NOSF[570]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2648.025 187.44 2648.305 188.44 ;
    END
  END Data_PMOS_NOSF[570]
  PIN Data_PMOS_NOSF[568]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2643.545 187.44 2643.825 188.44 ;
    END
  END Data_PMOS_NOSF[568]
  PIN Data_PMOS_NOSF[567]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2642.985 187.44 2643.265 188.44 ;
    END
  END Data_PMOS_NOSF[567]
  PIN Data_PMOS_NOSF[584]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2642.425 187.44 2642.705 188.44 ;
    END
  END Data_PMOS_NOSF[584]
  PIN DIG_MON_PMOS_NOSF[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2600.985 187.44 2601.265 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[54]
  PIN Data_PMOS_NOSF[578]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2644.105 187.44 2644.385 188.44 ;
    END
  END Data_PMOS_NOSF[578]
  PIN DIG_MON_PMOS_NOSF[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2596.505 187.44 2596.785 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[53]
  PIN Data_PMOS_NOSF[564]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2594.265 187.44 2594.545 188.44 ;
    END
  END Data_PMOS_NOSF[564]
  PIN Data_PMOS_NOSF[554]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2593.705 187.44 2593.985 188.44 ;
    END
  END Data_PMOS_NOSF[554]
  PIN Data_PMOS_NOSF[558]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2593.145 187.44 2593.425 188.44 ;
    END
  END Data_PMOS_NOSF[558]
  PIN Data_PMOS_NOSF[565]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2592.585 187.44 2592.865 188.44 ;
    END
  END Data_PMOS_NOSF[565]
  PIN Data_PMOS_NOSF[551]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2592.025 187.44 2592.305 188.44 ;
    END
  END Data_PMOS_NOSF[551]
  PIN Data_PMOS_NOSF[559]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2591.465 187.44 2591.745 188.44 ;
    END
  END Data_PMOS_NOSF[559]
  PIN Data_PMOS_NOSF[566]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2590.905 187.44 2591.185 188.44 ;
    END
  END Data_PMOS_NOSF[566]
  PIN Data_PMOS_NOSF[560]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2590.345 187.44 2590.625 188.44 ;
    END
  END Data_PMOS_NOSF[560]
  PIN Data_PMOS_NOSF[553]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2589.785 187.44 2590.065 188.44 ;
    END
  END Data_PMOS_NOSF[553]
  PIN Data_PMOS_NOSF[552]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2580.825 187.44 2581.105 188.44 ;
    END
  END Data_PMOS_NOSF[552]
  PIN nTOK_PMOS_NOSF[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2578.585 187.44 2578.865 188.44 ;
    END
  END nTOK_PMOS_NOSF[26]
  PIN FREEZE_PMOS_NOSF[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2575.785 187.44 2576.065 188.44 ;
    END
  END FREEZE_PMOS_NOSF[26]
  PIN Read_PMOS_NOSF[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2575.225 187.44 2575.505 188.44 ;
    END
  END Read_PMOS_NOSF[26]
  PIN Data_PMOS_NOSF[549]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2569.345 187.44 2569.625 188.44 ;
    END
  END Data_PMOS_NOSF[549]
  PIN Data_PMOS_NOSF[548]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2568.785 187.44 2569.065 188.44 ;
    END
  END Data_PMOS_NOSF[548]
  PIN Data_PMOS_NOSF[555]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2568.225 187.44 2568.505 188.44 ;
    END
  END Data_PMOS_NOSF[555]
  PIN Data_PMOS_NOSF[561]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2567.665 187.44 2567.945 188.44 ;
    END
  END Data_PMOS_NOSF[561]
  PIN Data_PMOS_NOSF[556]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2567.105 187.44 2567.385 188.44 ;
    END
  END Data_PMOS_NOSF[556]
  PIN Data_PMOS_NOSF[550]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2541.065 187.44 2541.345 188.44 ;
    END
  END Data_PMOS_NOSF[550]
  PIN Data_PMOS_NOSF[562]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2540.505 187.44 2540.785 188.44 ;
    END
  END Data_PMOS_NOSF[562]
  PIN Data_PMOS_NOSF[557]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2539.945 187.44 2540.225 188.44 ;
    END
  END Data_PMOS_NOSF[557]
  PIN Data_PMOS_NOSF[547]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2539.385 187.44 2539.665 188.44 ;
    END
  END Data_PMOS_NOSF[547]
  PIN Data_PMOS_NOSF[546]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2538.825 187.44 2539.105 188.44 ;
    END
  END Data_PMOS_NOSF[546]
  PIN Data_PMOS_NOSF[563]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2538.265 187.44 2538.545 188.44 ;
    END
  END Data_PMOS_NOSF[563]
  PIN DIG_MON_PMOS_NOSF[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2535.465 187.44 2535.745 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[52]
  PIN DIG_MON_PMOS_NOSF[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2530.985 187.44 2531.265 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[51]
  PIN Data_PMOS_NOSF[543]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2528.745 187.44 2529.025 188.44 ;
    END
  END Data_PMOS_NOSF[543]
  PIN Data_PMOS_NOSF[533]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2528.185 187.44 2528.465 188.44 ;
    END
  END Data_PMOS_NOSF[533]
  PIN Data_PMOS_NOSF[537]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2514.745 187.44 2515.025 188.44 ;
    END
  END Data_PMOS_NOSF[537]
  PIN Data_PMOS_NOSF[544]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2514.185 187.44 2514.465 188.44 ;
    END
  END Data_PMOS_NOSF[544]
  PIN Data_PMOS_NOSF[530]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2513.625 187.44 2513.905 188.44 ;
    END
  END Data_PMOS_NOSF[530]
  PIN Data_PMOS_NOSF[538]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2513.065 187.44 2513.345 188.44 ;
    END
  END Data_PMOS_NOSF[538]
  PIN Data_PMOS_NOSF[545]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2512.505 187.44 2512.785 188.44 ;
    END
  END Data_PMOS_NOSF[545]
  PIN Data_PMOS_NOSF[539]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2511.945 187.44 2512.225 188.44 ;
    END
  END Data_PMOS_NOSF[539]
  PIN Data_PMOS_NOSF[532]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2511.385 187.44 2511.665 188.44 ;
    END
  END Data_PMOS_NOSF[532]
  PIN Data_PMOS_NOSF[531]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2510.825 187.44 2511.105 188.44 ;
    END
  END Data_PMOS_NOSF[531]
  PIN nTOK_PMOS_NOSF[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2508.585 187.44 2508.865 188.44 ;
    END
  END nTOK_PMOS_NOSF[25]
  PIN FREEZE_PMOS_NOSF[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2505.785 187.44 2506.065 188.44 ;
    END
  END FREEZE_PMOS_NOSF[25]
  PIN Read_PMOS_NOSF[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2505.225 187.44 2505.505 188.44 ;
    END
  END Read_PMOS_NOSF[25]
  PIN Data_PMOS_NOSF[528]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2462.665 187.44 2462.945 188.44 ;
    END
  END Data_PMOS_NOSF[528]
  PIN Data_PMOS_NOSF[527]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2462.105 187.44 2462.385 188.44 ;
    END
  END Data_PMOS_NOSF[527]
  PIN Data_PMOS_NOSF[534]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2461.545 187.44 2461.825 188.44 ;
    END
  END Data_PMOS_NOSF[534]
  PIN Data_PMOS_NOSF[540]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2460.985 187.44 2461.265 188.44 ;
    END
  END Data_PMOS_NOSF[540]
  PIN Data_PMOS_NOSF[535]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2460.425 187.44 2460.705 188.44 ;
    END
  END Data_PMOS_NOSF[535]
  PIN Data_PMOS_NOSF[529]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2459.865 187.44 2460.145 188.44 ;
    END
  END Data_PMOS_NOSF[529]
  PIN Data_PMOS_NOSF[541]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2459.305 187.44 2459.585 188.44 ;
    END
  END Data_PMOS_NOSF[541]
  PIN Data_PMOS_NOSF[536]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2458.745 187.44 2459.025 188.44 ;
    END
  END Data_PMOS_NOSF[536]
  PIN Data_PMOS_NOSF[526]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2458.185 187.44 2458.465 188.44 ;
    END
  END Data_PMOS_NOSF[526]
  PIN Data_PMOS_NOSF[525]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2457.625 187.44 2457.905 188.44 ;
    END
  END Data_PMOS_NOSF[525]
  PIN Data_PMOS_NOSF[542]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2457.065 187.44 2457.345 188.44 ;
    END
  END Data_PMOS_NOSF[542]
  PIN DIG_MON_PMOS_NOSF[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2454.265 187.44 2454.545 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[50]
  PIN DIG_MON_PMOS_NOSF[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2449.785 187.44 2450.065 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[49]
  PIN Data_PMOS_NOSF[522]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2439.145 187.44 2439.425 188.44 ;
    END
  END Data_PMOS_NOSF[522]
  PIN Data_PMOS_NOSF[512]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2438.585 187.44 2438.865 188.44 ;
    END
  END Data_PMOS_NOSF[512]
  PIN Data_PMOS_NOSF[516]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2438.025 187.44 2438.305 188.44 ;
    END
  END Data_PMOS_NOSF[516]
  PIN Data_PMOS_NOSF[523]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2437.465 187.44 2437.745 188.44 ;
    END
  END Data_PMOS_NOSF[523]
  PIN Data_PMOS_NOSF[509]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2436.905 187.44 2437.185 188.44 ;
    END
  END Data_PMOS_NOSF[509]
  PIN Data_PMOS_NOSF[517]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2436.345 187.44 2436.625 188.44 ;
    END
  END Data_PMOS_NOSF[517]
  PIN Data_PMOS_NOSF[524]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2435.785 187.44 2436.065 188.44 ;
    END
  END Data_PMOS_NOSF[524]
  PIN Data_PMOS_NOSF[518]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2435.225 187.44 2435.505 188.44 ;
    END
  END Data_PMOS_NOSF[518]
  PIN Data_PMOS_NOSF[511]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2434.665 187.44 2434.945 188.44 ;
    END
  END Data_PMOS_NOSF[511]
  PIN Data_PMOS_NOSF[510]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2434.105 187.44 2434.385 188.44 ;
    END
  END Data_PMOS_NOSF[510]
  PIN nTOK_PMOS_NOSF[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2429.905 187.44 2430.185 188.44 ;
    END
  END nTOK_PMOS_NOSF[24]
  PIN Read_PMOS_NOSF[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2401.065 187.44 2401.345 188.44 ;
    END
  END Read_PMOS_NOSF[24]
  PIN Data_PMOS_NOSF[507]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2397.145 187.44 2397.425 188.44 ;
    END
  END Data_PMOS_NOSF[507]
  PIN Data_PMOS_NOSF[506]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2396.585 187.44 2396.865 188.44 ;
    END
  END Data_PMOS_NOSF[506]
  PIN Data_PMOS_NOSF[513]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2396.025 187.44 2396.305 188.44 ;
    END
  END Data_PMOS_NOSF[513]
  PIN Data_PMOS_NOSF[519]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2395.465 187.44 2395.745 188.44 ;
    END
  END Data_PMOS_NOSF[519]
  PIN Data_PMOS_NOSF[514]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2394.905 187.44 2395.185 188.44 ;
    END
  END Data_PMOS_NOSF[514]
  PIN Data_PMOS_NOSF[508]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2394.345 187.44 2394.625 188.44 ;
    END
  END Data_PMOS_NOSF[508]
  PIN Data_PMOS_NOSF[520]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2393.785 187.44 2394.065 188.44 ;
    END
  END Data_PMOS_NOSF[520]
  PIN Data_PMOS_NOSF[515]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2393.225 187.44 2393.505 188.44 ;
    END
  END Data_PMOS_NOSF[515]
  PIN Data_PMOS_NOSF[505]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2392.665 187.44 2392.945 188.44 ;
    END
  END Data_PMOS_NOSF[505]
  PIN Data_PMOS_NOSF[504]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2392.105 187.44 2392.385 188.44 ;
    END
  END Data_PMOS_NOSF[504]
  PIN Data_PMOS_NOSF[521]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2391.545 187.44 2391.825 188.44 ;
    END
  END Data_PMOS_NOSF[521]
  PIN DIG_MON_PMOS_NOSF[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2388.745 187.44 2389.025 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[48]
  PIN DIG_MON_PMOS_NOSF[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2371.385 187.44 2371.665 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[47]
  PIN Data_PMOS_NOSF[501]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2369.145 187.44 2369.425 188.44 ;
    END
  END Data_PMOS_NOSF[501]
  PIN Data_PMOS_NOSF[491]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2368.585 187.44 2368.865 188.44 ;
    END
  END Data_PMOS_NOSF[491]
  PIN Data_PMOS_NOSF[495]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2368.025 187.44 2368.305 188.44 ;
    END
  END Data_PMOS_NOSF[495]
  PIN Data_PMOS_NOSF[502]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2367.465 187.44 2367.745 188.44 ;
    END
  END Data_PMOS_NOSF[502]
  PIN Data_PMOS_NOSF[488]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2366.905 187.44 2367.185 188.44 ;
    END
  END Data_PMOS_NOSF[488]
  PIN Data_PMOS_NOSF[496]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2366.345 187.44 2366.625 188.44 ;
    END
  END Data_PMOS_NOSF[496]
  PIN Data_PMOS_NOSF[503]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2365.785 187.44 2366.065 188.44 ;
    END
  END Data_PMOS_NOSF[503]
  PIN Data_PMOS_NOSF[497]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2365.225 187.44 2365.505 188.44 ;
    END
  END Data_PMOS_NOSF[497]
  PIN Data_PMOS_NOSF[490]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2364.665 187.44 2364.945 188.44 ;
    END
  END Data_PMOS_NOSF[490]
  PIN Data_PMOS_NOSF[489]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2364.105 187.44 2364.385 188.44 ;
    END
  END Data_PMOS_NOSF[489]
  PIN nTOK_PMOS_NOSF[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2322.665 187.44 2322.945 188.44 ;
    END
  END nTOK_PMOS_NOSF[23]
  PIN FREEZE_PMOS_NOSF[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2319.865 187.44 2320.145 188.44 ;
    END
  END FREEZE_PMOS_NOSF[23]
  PIN Read_PMOS_NOSF[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2319.305 187.44 2319.585 188.44 ;
    END
  END Read_PMOS_NOSF[23]
  PIN Data_PMOS_NOSF[486]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2315.385 187.44 2315.665 188.44 ;
    END
  END Data_PMOS_NOSF[486]
  PIN Data_PMOS_NOSF[485]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2314.825 187.44 2315.105 188.44 ;
    END
  END Data_PMOS_NOSF[485]
  PIN Data_PMOS_NOSF[492]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2314.265 187.44 2314.545 188.44 ;
    END
  END Data_PMOS_NOSF[492]
  PIN Data_PMOS_NOSF[498]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2313.705 187.44 2313.985 188.44 ;
    END
  END Data_PMOS_NOSF[498]
  PIN Data_PMOS_NOSF[493]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2313.145 187.44 2313.425 188.44 ;
    END
  END Data_PMOS_NOSF[493]
  PIN Data_PMOS_NOSF[487]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2312.585 187.44 2312.865 188.44 ;
    END
  END Data_PMOS_NOSF[487]
  PIN Data_PMOS_NOSF[499]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2312.025 187.44 2312.305 188.44 ;
    END
  END Data_PMOS_NOSF[499]
  PIN Data_PMOS_NOSF[494]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2311.465 187.44 2311.745 188.44 ;
    END
  END Data_PMOS_NOSF[494]
  PIN Data_PMOS_NOSF[484]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2310.905 187.44 2311.185 188.44 ;
    END
  END Data_PMOS_NOSF[484]
  PIN Data_PMOS_NOSF[483]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2310.345 187.44 2310.625 188.44 ;
    END
  END Data_PMOS_NOSF[483]
  PIN Data_PMOS_NOSF[500]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2309.785 187.44 2310.065 188.44 ;
    END
  END Data_PMOS_NOSF[500]
  PIN DIG_MON_PMOS_NOSF[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2298.585 187.44 2298.865 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[46]
  PIN DIG_MON_PMOS_NOSF[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2294.105 187.44 2294.385 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[45]
  PIN Data_PMOS_NOSF[480]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2289.905 187.44 2290.185 188.44 ;
    END
  END Data_PMOS_NOSF[480]
  PIN Data_PMOS_NOSF[470]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2289.345 187.44 2289.625 188.44 ;
    END
  END Data_PMOS_NOSF[470]
  PIN Data_PMOS_NOSF[474]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2288.785 187.44 2289.065 188.44 ;
    END
  END Data_PMOS_NOSF[474]
  PIN Data_PMOS_NOSF[481]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2288.225 187.44 2288.505 188.44 ;
    END
  END Data_PMOS_NOSF[481]
  PIN Data_PMOS_NOSF[467]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2287.665 187.44 2287.945 188.44 ;
    END
  END Data_PMOS_NOSF[467]
  PIN Data_PMOS_NOSF[475]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2261.625 187.44 2261.905 188.44 ;
    END
  END Data_PMOS_NOSF[475]
  PIN Data_PMOS_NOSF[482]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2261.065 187.44 2261.345 188.44 ;
    END
  END Data_PMOS_NOSF[482]
  PIN Data_PMOS_NOSF[476]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2260.505 187.44 2260.785 188.44 ;
    END
  END Data_PMOS_NOSF[476]
  PIN Data_PMOS_NOSF[469]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2259.945 187.44 2260.225 188.44 ;
    END
  END Data_PMOS_NOSF[469]
  PIN Data_PMOS_NOSF[468]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2259.385 187.44 2259.665 188.44 ;
    END
  END Data_PMOS_NOSF[468]
  PIN nTOK_PMOS_NOSF[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2257.145 187.44 2257.425 188.44 ;
    END
  END nTOK_PMOS_NOSF[22]
  PIN FREEZE_PMOS_NOSF[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2254.345 187.44 2254.625 188.44 ;
    END
  END FREEZE_PMOS_NOSF[22]
  PIN Read_PMOS_NOSF[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2253.785 187.44 2254.065 188.44 ;
    END
  END Read_PMOS_NOSF[22]
  PIN Data_PMOS_NOSF[465]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2249.865 187.44 2250.145 188.44 ;
    END
  END Data_PMOS_NOSF[465]
  PIN Data_PMOS_NOSF[464]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2249.305 187.44 2249.585 188.44 ;
    END
  END Data_PMOS_NOSF[464]
  PIN Data_PMOS_NOSF[471]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2248.745 187.44 2249.025 188.44 ;
    END
  END Data_PMOS_NOSF[471]
  PIN Data_PMOS_NOSF[477]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2235.305 187.44 2235.585 188.44 ;
    END
  END Data_PMOS_NOSF[477]
  PIN Data_PMOS_NOSF[472]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2234.745 187.44 2235.025 188.44 ;
    END
  END Data_PMOS_NOSF[472]
  PIN Data_PMOS_NOSF[466]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2234.185 187.44 2234.465 188.44 ;
    END
  END Data_PMOS_NOSF[466]
  PIN Data_PMOS_NOSF[478]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2233.625 187.44 2233.905 188.44 ;
    END
  END Data_PMOS_NOSF[478]
  PIN Data_PMOS_NOSF[473]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2233.065 187.44 2233.345 188.44 ;
    END
  END Data_PMOS_NOSF[473]
  PIN Data_PMOS_NOSF[463]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2232.505 187.44 2232.785 188.44 ;
    END
  END Data_PMOS_NOSF[463]
  PIN Data_PMOS_NOSF[462]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2231.945 187.44 2232.225 188.44 ;
    END
  END Data_PMOS_NOSF[462]
  PIN Data_PMOS_NOSF[479]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2231.385 187.44 2231.665 188.44 ;
    END
  END Data_PMOS_NOSF[479]
  PIN DIG_MON_PMOS_NOSF[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2228.585 187.44 2228.865 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[44]
  PIN DIG_MON_PMOS_NOSF[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2224.105 187.44 2224.385 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[43]
  PIN Data_PMOS_NOSF[459]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2182.105 187.44 2182.385 188.44 ;
    END
  END Data_PMOS_NOSF[459]
  PIN Data_PMOS_NOSF[449]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2181.545 187.44 2181.825 188.44 ;
    END
  END Data_PMOS_NOSF[449]
  PIN Data_PMOS_NOSF[453]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2180.985 187.44 2181.265 188.44 ;
    END
  END Data_PMOS_NOSF[453]
  PIN Data_PMOS_NOSF[460]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2180.425 187.44 2180.705 188.44 ;
    END
  END Data_PMOS_NOSF[460]
  PIN Data_PMOS_NOSF[446]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2179.865 187.44 2180.145 188.44 ;
    END
  END Data_PMOS_NOSF[446]
  PIN Data_PMOS_NOSF[454]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2179.305 187.44 2179.585 188.44 ;
    END
  END Data_PMOS_NOSF[454]
  PIN Data_PMOS_NOSF[461]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2178.745 187.44 2179.025 188.44 ;
    END
  END Data_PMOS_NOSF[461]
  PIN Data_PMOS_NOSF[455]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2178.185 187.44 2178.465 188.44 ;
    END
  END Data_PMOS_NOSF[455]
  PIN Data_PMOS_NOSF[448]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2177.625 187.44 2177.905 188.44 ;
    END
  END Data_PMOS_NOSF[448]
  PIN Data_PMOS_NOSF[447]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2177.065 187.44 2177.345 188.44 ;
    END
  END Data_PMOS_NOSF[447]
  PIN nTOK_PMOS_NOSF[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2174.825 187.44 2175.105 188.44 ;
    END
  END nTOK_PMOS_NOSF[21]
  PIN FREEZE_PMOS_NOSF[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2172.025 187.44 2172.305 188.44 ;
    END
  END FREEZE_PMOS_NOSF[21]
  PIN Read_PMOS_NOSF[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2171.465 187.44 2171.745 188.44 ;
    END
  END Read_PMOS_NOSF[21]
  PIN Data_PMOS_NOSF[444]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2159.145 187.44 2159.425 188.44 ;
    END
  END Data_PMOS_NOSF[444]
  PIN Data_PMOS_NOSF[443]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2158.585 187.44 2158.865 188.44 ;
    END
  END Data_PMOS_NOSF[443]
  PIN Data_PMOS_NOSF[456]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2157.465 187.44 2157.745 188.44 ;
    END
  END Data_PMOS_NOSF[456]
  PIN Data_PMOS_NOSF[450]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2158.025 187.44 2158.305 188.44 ;
    END
  END Data_PMOS_NOSF[450]
  PIN Data_PMOS_NOSF[451]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2156.905 187.44 2157.185 188.44 ;
    END
  END Data_PMOS_NOSF[451]
  PIN Data_PMOS_NOSF[445]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2156.345 187.44 2156.625 188.44 ;
    END
  END Data_PMOS_NOSF[445]
  PIN Data_PMOS_NOSF[457]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2155.785 187.44 2156.065 188.44 ;
    END
  END Data_PMOS_NOSF[457]
  PIN Data_PMOS_NOSF[452]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2155.225 187.44 2155.505 188.44 ;
    END
  END Data_PMOS_NOSF[452]
  PIN Data_PMOS_NOSF[442]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2154.665 187.44 2154.945 188.44 ;
    END
  END Data_PMOS_NOSF[442]
  PIN Data_PMOS_NOSF[441]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2154.105 187.44 2154.385 188.44 ;
    END
  END Data_PMOS_NOSF[441]
  PIN Data_PMOS_NOSF[458]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2153.545 187.44 2153.825 188.44 ;
    END
  END Data_PMOS_NOSF[458]
  PIN DIG_MON_PMOS_NOSF[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2148.785 187.44 2149.065 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[42]
  PIN FREEZE_PMOS_NOSF[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2401.625 187.44 2401.905 188.44 ;
    END
  END FREEZE_PMOS_NOSF[24]
  PIN DIG_MON_PMOS_NOSF[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3238.265 187.44 3238.545 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[69]
  PIN Data_PMOS_NOSF[732]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3236.025 187.44 3236.305 188.44 ;
    END
  END Data_PMOS_NOSF[732]
  PIN Data_PMOS_NOSF[722]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3235.465 187.44 3235.745 188.44 ;
    END
  END Data_PMOS_NOSF[722]
  PIN Data_PMOS_NOSF[726]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3234.905 187.44 3235.185 188.44 ;
    END
  END Data_PMOS_NOSF[726]
  PIN Data_PMOS_NOSF[733]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3234.345 187.44 3234.625 188.44 ;
    END
  END Data_PMOS_NOSF[733]
  PIN Data_PMOS_NOSF[719]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3233.785 187.44 3234.065 188.44 ;
    END
  END Data_PMOS_NOSF[719]
  PIN Data_PMOS_NOSF[727]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3233.225 187.44 3233.505 188.44 ;
    END
  END Data_PMOS_NOSF[727]
  PIN Data_PMOS_NOSF[734]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3232.665 187.44 3232.945 188.44 ;
    END
  END Data_PMOS_NOSF[734]
  PIN Data_PMOS_NOSF[728]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3232.105 187.44 3232.385 188.44 ;
    END
  END Data_PMOS_NOSF[728]
  PIN Data_PMOS_NOSF[721]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3231.545 187.44 3231.825 188.44 ;
    END
  END Data_PMOS_NOSF[721]
  PIN Data_PMOS_NOSF[720]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3230.985 187.44 3231.265 188.44 ;
    END
  END Data_PMOS_NOSF[720]
  PIN nTOK_PMOS_NOSF[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3228.745 187.44 3229.025 188.44 ;
    END
  END nTOK_PMOS_NOSF[34]
  PIN FREEZE_PMOS_NOSF[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3212.505 187.44 3212.785 188.44 ;
    END
  END FREEZE_PMOS_NOSF[34]
  PIN Read_PMOS_NOSF[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3211.945 187.44 3212.225 188.44 ;
    END
  END Read_PMOS_NOSF[34]
  PIN Data_PMOS_NOSF[717]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3208.025 187.44 3208.305 188.44 ;
    END
  END Data_PMOS_NOSF[717]
  PIN Data_PMOS_NOSF[716]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3207.465 187.44 3207.745 188.44 ;
    END
  END Data_PMOS_NOSF[716]
  PIN Data_PMOS_NOSF[723]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3206.905 187.44 3207.185 188.44 ;
    END
  END Data_PMOS_NOSF[723]
  PIN Data_PMOS_NOSF[729]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3206.345 187.44 3206.625 188.44 ;
    END
  END Data_PMOS_NOSF[729]
  PIN Data_PMOS_NOSF[724]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3205.785 187.44 3206.065 188.44 ;
    END
  END Data_PMOS_NOSF[724]
  PIN Data_PMOS_NOSF[718]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3205.225 187.44 3205.505 188.44 ;
    END
  END Data_PMOS_NOSF[718]
  PIN Data_PMOS_NOSF[730]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3204.665 187.44 3204.945 188.44 ;
    END
  END Data_PMOS_NOSF[730]
  PIN Data_PMOS_NOSF[725]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3204.105 187.44 3204.385 188.44 ;
    END
  END Data_PMOS_NOSF[725]
  PIN Data_PMOS_NOSF[715]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3203.545 187.44 3203.825 188.44 ;
    END
  END Data_PMOS_NOSF[715]
  PIN Data_PMOS_NOSF[714]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3202.985 187.44 3203.265 188.44 ;
    END
  END Data_PMOS_NOSF[714]
  PIN Data_PMOS_NOSF[731]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3202.425 187.44 3202.705 188.44 ;
    END
  END Data_PMOS_NOSF[731]
  PIN DIG_MON_PMOS_NOSF[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3160.985 187.44 3161.265 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[68]
  PIN DIG_MON_PMOS_NOSF[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3156.505 187.44 3156.785 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[67]
  PIN Data_PMOS_NOSF[711]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3154.265 187.44 3154.545 188.44 ;
    END
  END Data_PMOS_NOSF[711]
  PIN Data_PMOS_NOSF[701]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3153.705 187.44 3153.985 188.44 ;
    END
  END Data_PMOS_NOSF[701]
  PIN Data_PMOS_NOSF[705]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3153.145 187.44 3153.425 188.44 ;
    END
  END Data_PMOS_NOSF[705]
  PIN Data_PMOS_NOSF[712]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3152.585 187.44 3152.865 188.44 ;
    END
  END Data_PMOS_NOSF[712]
  PIN Data_PMOS_NOSF[698]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3152.025 187.44 3152.305 188.44 ;
    END
  END Data_PMOS_NOSF[698]
  PIN Data_PMOS_NOSF[706]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3151.465 187.44 3151.745 188.44 ;
    END
  END Data_PMOS_NOSF[706]
  PIN Data_PMOS_NOSF[713]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3150.905 187.44 3151.185 188.44 ;
    END
  END Data_PMOS_NOSF[713]
  PIN Data_PMOS_NOSF[707]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3150.345 187.44 3150.625 188.44 ;
    END
  END Data_PMOS_NOSF[707]
  PIN Data_PMOS_NOSF[700]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3149.785 187.44 3150.065 188.44 ;
    END
  END Data_PMOS_NOSF[700]
  PIN Data_PMOS_NOSF[699]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3140.825 187.44 3141.105 188.44 ;
    END
  END Data_PMOS_NOSF[699]
  PIN nTOK_PMOS_NOSF[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3138.585 187.44 3138.865 188.44 ;
    END
  END nTOK_PMOS_NOSF[33]
  PIN FREEZE_PMOS_NOSF[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3135.785 187.44 3136.065 188.44 ;
    END
  END FREEZE_PMOS_NOSF[33]
  PIN Read_PMOS_NOSF[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3135.225 187.44 3135.505 188.44 ;
    END
  END Read_PMOS_NOSF[33]
  PIN Data_PMOS_NOSF[696]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3129.345 187.44 3129.625 188.44 ;
    END
  END Data_PMOS_NOSF[696]
  PIN Data_PMOS_NOSF[695]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3128.785 187.44 3129.065 188.44 ;
    END
  END Data_PMOS_NOSF[695]
  PIN Data_PMOS_NOSF[702]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3128.225 187.44 3128.505 188.44 ;
    END
  END Data_PMOS_NOSF[702]
  PIN Data_PMOS_NOSF[708]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3127.665 187.44 3127.945 188.44 ;
    END
  END Data_PMOS_NOSF[708]
  PIN Data_PMOS_NOSF[703]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3127.105 187.44 3127.385 188.44 ;
    END
  END Data_PMOS_NOSF[703]
  PIN Data_PMOS_NOSF[697]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3101.065 187.44 3101.345 188.44 ;
    END
  END Data_PMOS_NOSF[697]
  PIN Data_PMOS_NOSF[709]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3100.505 187.44 3100.785 188.44 ;
    END
  END Data_PMOS_NOSF[709]
  PIN Data_PMOS_NOSF[704]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3099.945 187.44 3100.225 188.44 ;
    END
  END Data_PMOS_NOSF[704]
  PIN Data_PMOS_NOSF[694]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3099.385 187.44 3099.665 188.44 ;
    END
  END Data_PMOS_NOSF[694]
  PIN Data_PMOS_NOSF[693]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3098.825 187.44 3099.105 188.44 ;
    END
  END Data_PMOS_NOSF[693]
  PIN Data_PMOS_NOSF[710]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3098.265 187.44 3098.545 188.44 ;
    END
  END Data_PMOS_NOSF[710]
  PIN DIG_MON_PMOS_NOSF[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3095.465 187.44 3095.745 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[66]
  PIN DIG_MON_PMOS_NOSF[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3090.985 187.44 3091.265 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[65]
  PIN Data_PMOS_NOSF[690]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3088.745 187.44 3089.025 188.44 ;
    END
  END Data_PMOS_NOSF[690]
  PIN Data_PMOS_NOSF[680]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3088.185 187.44 3088.465 188.44 ;
    END
  END Data_PMOS_NOSF[680]
  PIN Data_PMOS_NOSF[684]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3074.745 187.44 3075.025 188.44 ;
    END
  END Data_PMOS_NOSF[684]
  PIN Data_PMOS_NOSF[691]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3074.185 187.44 3074.465 188.44 ;
    END
  END Data_PMOS_NOSF[691]
  PIN Data_PMOS_NOSF[677]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3073.625 187.44 3073.905 188.44 ;
    END
  END Data_PMOS_NOSF[677]
  PIN Data_PMOS_NOSF[685]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3073.065 187.44 3073.345 188.44 ;
    END
  END Data_PMOS_NOSF[685]
  PIN Data_PMOS_NOSF[692]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3072.505 187.44 3072.785 188.44 ;
    END
  END Data_PMOS_NOSF[692]
  PIN Data_PMOS_NOSF[686]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3071.945 187.44 3072.225 188.44 ;
    END
  END Data_PMOS_NOSF[686]
  PIN Data_PMOS_NOSF[679]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3071.385 187.44 3071.665 188.44 ;
    END
  END Data_PMOS_NOSF[679]
  PIN Data_PMOS_NOSF[678]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3070.825 187.44 3071.105 188.44 ;
    END
  END Data_PMOS_NOSF[678]
  PIN nTOK_PMOS_NOSF[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3068.585 187.44 3068.865 188.44 ;
    END
  END nTOK_PMOS_NOSF[32]
  PIN FREEZE_PMOS_NOSF[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3065.785 187.44 3066.065 188.44 ;
    END
  END FREEZE_PMOS_NOSF[32]
  PIN Read_PMOS_NOSF[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3065.225 187.44 3065.505 188.44 ;
    END
  END Read_PMOS_NOSF[32]
  PIN Data_PMOS_NOSF[675]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3022.665 187.44 3022.945 188.44 ;
    END
  END Data_PMOS_NOSF[675]
  PIN Data_PMOS_NOSF[674]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3022.105 187.44 3022.385 188.44 ;
    END
  END Data_PMOS_NOSF[674]
  PIN Data_PMOS_NOSF[681]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3021.545 187.44 3021.825 188.44 ;
    END
  END Data_PMOS_NOSF[681]
  PIN Data_PMOS_NOSF[687]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3020.985 187.44 3021.265 188.44 ;
    END
  END Data_PMOS_NOSF[687]
  PIN Data_PMOS_NOSF[682]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3020.425 187.44 3020.705 188.44 ;
    END
  END Data_PMOS_NOSF[682]
  PIN Data_PMOS_NOSF[676]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3019.865 187.44 3020.145 188.44 ;
    END
  END Data_PMOS_NOSF[676]
  PIN Data_PMOS_NOSF[688]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3019.305 187.44 3019.585 188.44 ;
    END
  END Data_PMOS_NOSF[688]
  PIN Data_PMOS_NOSF[683]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3018.745 187.44 3019.025 188.44 ;
    END
  END Data_PMOS_NOSF[683]
  PIN Data_PMOS_NOSF[673]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3018.185 187.44 3018.465 188.44 ;
    END
  END Data_PMOS_NOSF[673]
  PIN Data_PMOS_NOSF[672]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3017.625 187.44 3017.905 188.44 ;
    END
  END Data_PMOS_NOSF[672]
  PIN Data_PMOS_NOSF[689]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3017.065 187.44 3017.345 188.44 ;
    END
  END Data_PMOS_NOSF[689]
  PIN DIG_MON_PMOS_NOSF[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3014.265 187.44 3014.545 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[64]
  PIN DIG_MON_PMOS_NOSF[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3009.785 187.44 3010.065 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[63]
  PIN Data_PMOS_NOSF[669]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2999.145 187.44 2999.425 188.44 ;
    END
  END Data_PMOS_NOSF[669]
  PIN Data_PMOS_NOSF[659]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2998.585 187.44 2998.865 188.44 ;
    END
  END Data_PMOS_NOSF[659]
  PIN Data_PMOS_NOSF[663]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2998.025 187.44 2998.305 188.44 ;
    END
  END Data_PMOS_NOSF[663]
  PIN Data_PMOS_NOSF[670]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2997.465 187.44 2997.745 188.44 ;
    END
  END Data_PMOS_NOSF[670]
  PIN Data_PMOS_NOSF[656]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2996.905 187.44 2997.185 188.44 ;
    END
  END Data_PMOS_NOSF[656]
  PIN Data_PMOS_NOSF[664]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2996.345 187.44 2996.625 188.44 ;
    END
  END Data_PMOS_NOSF[664]
  PIN Data_PMOS_NOSF[671]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2995.785 187.44 2996.065 188.44 ;
    END
  END Data_PMOS_NOSF[671]
  PIN Data_PMOS_NOSF[665]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2995.225 187.44 2995.505 188.44 ;
    END
  END Data_PMOS_NOSF[665]
  PIN Data_PMOS_NOSF[658]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2994.665 187.44 2994.945 188.44 ;
    END
  END Data_PMOS_NOSF[658]
  PIN Data_PMOS_NOSF[657]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2994.105 187.44 2994.385 188.44 ;
    END
  END Data_PMOS_NOSF[657]
  PIN nTOK_PMOS_NOSF[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2989.905 187.44 2990.185 188.44 ;
    END
  END nTOK_PMOS_NOSF[31]
  PIN Read_PMOS_NOSF[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2961.065 187.44 2961.345 188.44 ;
    END
  END Read_PMOS_NOSF[31]
  PIN Data_PMOS_NOSF[654]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2957.145 187.44 2957.425 188.44 ;
    END
  END Data_PMOS_NOSF[654]
  PIN Data_PMOS_NOSF[653]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2956.585 187.44 2956.865 188.44 ;
    END
  END Data_PMOS_NOSF[653]
  PIN Data_PMOS_NOSF[660]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2956.025 187.44 2956.305 188.44 ;
    END
  END Data_PMOS_NOSF[660]
  PIN Data_PMOS_NOSF[666]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2955.465 187.44 2955.745 188.44 ;
    END
  END Data_PMOS_NOSF[666]
  PIN Data_PMOS_NOSF[661]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2954.905 187.44 2955.185 188.44 ;
    END
  END Data_PMOS_NOSF[661]
  PIN Data_PMOS_NOSF[655]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2954.345 187.44 2954.625 188.44 ;
    END
  END Data_PMOS_NOSF[655]
  PIN Data_PMOS_NOSF[667]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2953.785 187.44 2954.065 188.44 ;
    END
  END Data_PMOS_NOSF[667]
  PIN Data_PMOS_NOSF[662]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2953.225 187.44 2953.505 188.44 ;
    END
  END Data_PMOS_NOSF[662]
  PIN Data_PMOS_NOSF[652]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2952.665 187.44 2952.945 188.44 ;
    END
  END Data_PMOS_NOSF[652]
  PIN Data_PMOS_NOSF[651]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2952.105 187.44 2952.385 188.44 ;
    END
  END Data_PMOS_NOSF[651]
  PIN Data_PMOS_NOSF[668]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2951.545 187.44 2951.825 188.44 ;
    END
  END Data_PMOS_NOSF[668]
  PIN DIG_MON_PMOS_NOSF[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2948.745 187.44 2949.025 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[62]
  PIN DIG_MON_PMOS_NOSF[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2931.385 187.44 2931.665 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[61]
  PIN Data_PMOS_NOSF[648]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2929.145 187.44 2929.425 188.44 ;
    END
  END Data_PMOS_NOSF[648]
  PIN Data_PMOS_NOSF[638]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2928.585 187.44 2928.865 188.44 ;
    END
  END Data_PMOS_NOSF[638]
  PIN Data_PMOS_NOSF[642]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2928.025 187.44 2928.305 188.44 ;
    END
  END Data_PMOS_NOSF[642]
  PIN Data_PMOS_NOSF[649]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2927.465 187.44 2927.745 188.44 ;
    END
  END Data_PMOS_NOSF[649]
  PIN Data_PMOS_NOSF[635]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2926.905 187.44 2927.185 188.44 ;
    END
  END Data_PMOS_NOSF[635]
  PIN Data_PMOS_NOSF[643]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2926.345 187.44 2926.625 188.44 ;
    END
  END Data_PMOS_NOSF[643]
  PIN Data_PMOS_NOSF[650]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2925.785 187.44 2926.065 188.44 ;
    END
  END Data_PMOS_NOSF[650]
  PIN Data_PMOS_NOSF[644]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2925.225 187.44 2925.505 188.44 ;
    END
  END Data_PMOS_NOSF[644]
  PIN Data_PMOS_NOSF[637]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2924.665 187.44 2924.945 188.44 ;
    END
  END Data_PMOS_NOSF[637]
  PIN Data_PMOS_NOSF[636]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2924.105 187.44 2924.385 188.44 ;
    END
  END Data_PMOS_NOSF[636]
  PIN nTOK_PMOS_NOSF[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2882.665 187.44 2882.945 188.44 ;
    END
  END nTOK_PMOS_NOSF[30]
  PIN FREEZE_PMOS_NOSF[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2879.865 187.44 2880.145 188.44 ;
    END
  END FREEZE_PMOS_NOSF[30]
  PIN Read_PMOS_NOSF[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2879.305 187.44 2879.585 188.44 ;
    END
  END Read_PMOS_NOSF[30]
  PIN Data_PMOS_NOSF[633]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2875.385 187.44 2875.665 188.44 ;
    END
  END Data_PMOS_NOSF[633]
  PIN Data_PMOS_NOSF[632]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2874.825 187.44 2875.105 188.44 ;
    END
  END Data_PMOS_NOSF[632]
  PIN Data_PMOS_NOSF[639]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2874.265 187.44 2874.545 188.44 ;
    END
  END Data_PMOS_NOSF[639]
  PIN Data_PMOS_NOSF[645]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2873.705 187.44 2873.985 188.44 ;
    END
  END Data_PMOS_NOSF[645]
  PIN Data_PMOS_NOSF[640]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2873.145 187.44 2873.425 188.44 ;
    END
  END Data_PMOS_NOSF[640]
  PIN Data_PMOS_NOSF[634]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2872.585 187.44 2872.865 188.44 ;
    END
  END Data_PMOS_NOSF[634]
  PIN Data_PMOS_NOSF[646]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2872.025 187.44 2872.305 188.44 ;
    END
  END Data_PMOS_NOSF[646]
  PIN Data_PMOS_NOSF[641]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2871.465 187.44 2871.745 188.44 ;
    END
  END Data_PMOS_NOSF[641]
  PIN Data_PMOS_NOSF[631]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2870.905 187.44 2871.185 188.44 ;
    END
  END Data_PMOS_NOSF[631]
  PIN Data_PMOS_NOSF[630]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2870.345 187.44 2870.625 188.44 ;
    END
  END Data_PMOS_NOSF[630]
  PIN Data_PMOS_NOSF[647]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2869.785 187.44 2870.065 188.44 ;
    END
  END Data_PMOS_NOSF[647]
  PIN DIG_MON_PMOS_NOSF[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2858.585 187.44 2858.865 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[60]
  PIN DIG_MON_PMOS_NOSF[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2854.105 187.44 2854.385 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[59]
  PIN Data_PMOS_NOSF[627]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2849.905 187.44 2850.185 188.44 ;
    END
  END Data_PMOS_NOSF[627]
  PIN Data_PMOS_NOSF[617]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2849.345 187.44 2849.625 188.44 ;
    END
  END Data_PMOS_NOSF[617]
  PIN Data_PMOS_NOSF[621]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2848.785 187.44 2849.065 188.44 ;
    END
  END Data_PMOS_NOSF[621]
  PIN Data_PMOS_NOSF[628]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2848.225 187.44 2848.505 188.44 ;
    END
  END Data_PMOS_NOSF[628]
  PIN Data_PMOS_NOSF[614]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2847.665 187.44 2847.945 188.44 ;
    END
  END Data_PMOS_NOSF[614]
  PIN Data_PMOS_NOSF[622]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2821.625 187.44 2821.905 188.44 ;
    END
  END Data_PMOS_NOSF[622]
  PIN Data_PMOS_NOSF[629]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2821.065 187.44 2821.345 188.44 ;
    END
  END Data_PMOS_NOSF[629]
  PIN Data_PMOS_NOSF[623]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2820.505 187.44 2820.785 188.44 ;
    END
  END Data_PMOS_NOSF[623]
  PIN Data_PMOS_NOSF[616]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2819.945 187.44 2820.225 188.44 ;
    END
  END Data_PMOS_NOSF[616]
  PIN Data_PMOS_NOSF[615]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2819.385 187.44 2819.665 188.44 ;
    END
  END Data_PMOS_NOSF[615]
  PIN nTOK_PMOS_NOSF[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2817.145 187.44 2817.425 188.44 ;
    END
  END nTOK_PMOS_NOSF[29]
  PIN FREEZE_PMOS_NOSF[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2814.345 187.44 2814.625 188.44 ;
    END
  END FREEZE_PMOS_NOSF[29]
  PIN Read_PMOS_NOSF[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2813.785 187.44 2814.065 188.44 ;
    END
  END Read_PMOS_NOSF[29]
  PIN Data_PMOS_NOSF[612]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2809.865 187.44 2810.145 188.44 ;
    END
  END Data_PMOS_NOSF[612]
  PIN Data_PMOS_NOSF[611]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2809.305 187.44 2809.585 188.44 ;
    END
  END Data_PMOS_NOSF[611]
  PIN Data_PMOS_NOSF[618]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2808.745 187.44 2809.025 188.44 ;
    END
  END Data_PMOS_NOSF[618]
  PIN Data_PMOS_NOSF[624]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2795.305 187.44 2795.585 188.44 ;
    END
  END Data_PMOS_NOSF[624]
  PIN Data_PMOS_NOSF[619]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2794.745 187.44 2795.025 188.44 ;
    END
  END Data_PMOS_NOSF[619]
  PIN Data_PMOS_NOSF[613]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2794.185 187.44 2794.465 188.44 ;
    END
  END Data_PMOS_NOSF[613]
  PIN Data_PMOS_NOSF[625]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2793.625 187.44 2793.905 188.44 ;
    END
  END Data_PMOS_NOSF[625]
  PIN Data_PMOS_NOSF[620]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2793.065 187.44 2793.345 188.44 ;
    END
  END Data_PMOS_NOSF[620]
  PIN Data_PMOS_NOSF[610]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2792.505 187.44 2792.785 188.44 ;
    END
  END Data_PMOS_NOSF[610]
  PIN Data_PMOS_NOSF[609]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2791.945 187.44 2792.225 188.44 ;
    END
  END Data_PMOS_NOSF[609]
  PIN Data_PMOS_NOSF[626]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2791.385 187.44 2791.665 188.44 ;
    END
  END Data_PMOS_NOSF[626]
  PIN DIG_MON_PMOS_NOSF[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2788.585 187.44 2788.865 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[58]
  PIN DIG_MON_PMOS_NOSF[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2784.105 187.44 2784.385 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[57]
  PIN Data_PMOS_NOSF[606]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2742.105 187.44 2742.385 188.44 ;
    END
  END Data_PMOS_NOSF[606]
  PIN Data_PMOS_NOSF[596]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2741.545 187.44 2741.825 188.44 ;
    END
  END Data_PMOS_NOSF[596]
  PIN Data_PMOS_NOSF[600]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2740.985 187.44 2741.265 188.44 ;
    END
  END Data_PMOS_NOSF[600]
  PIN Data_PMOS_NOSF[607]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2740.425 187.44 2740.705 188.44 ;
    END
  END Data_PMOS_NOSF[607]
  PIN Data_PMOS_NOSF[593]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2739.865 187.44 2740.145 188.44 ;
    END
  END Data_PMOS_NOSF[593]
  PIN Data_PMOS_NOSF[601]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2739.305 187.44 2739.585 188.44 ;
    END
  END Data_PMOS_NOSF[601]
  PIN Data_PMOS_NOSF[608]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2738.745 187.44 2739.025 188.44 ;
    END
  END Data_PMOS_NOSF[608]
  PIN Data_PMOS_NOSF[602]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2738.185 187.44 2738.465 188.44 ;
    END
  END Data_PMOS_NOSF[602]
  PIN Data_PMOS_NOSF[595]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2737.625 187.44 2737.905 188.44 ;
    END
  END Data_PMOS_NOSF[595]
  PIN Data_PMOS_NOSF[594]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2737.065 187.44 2737.345 188.44 ;
    END
  END Data_PMOS_NOSF[594]
  PIN nTOK_PMOS_NOSF[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2734.825 187.44 2735.105 188.44 ;
    END
  END nTOK_PMOS_NOSF[28]
  PIN FREEZE_PMOS_NOSF[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2732.025 187.44 2732.305 188.44 ;
    END
  END FREEZE_PMOS_NOSF[28]
  PIN Read_PMOS_NOSF[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2731.465 187.44 2731.745 188.44 ;
    END
  END Read_PMOS_NOSF[28]
  PIN Data_PMOS_NOSF[591]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2719.145 187.44 2719.425 188.44 ;
    END
  END Data_PMOS_NOSF[591]
  PIN Data_PMOS_NOSF[590]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2718.585 187.44 2718.865 188.44 ;
    END
  END Data_PMOS_NOSF[590]
  PIN Data_PMOS_NOSF[603]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2717.465 187.44 2717.745 188.44 ;
    END
  END Data_PMOS_NOSF[603]
  PIN Data_PMOS_NOSF[597]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2718.025 187.44 2718.305 188.44 ;
    END
  END Data_PMOS_NOSF[597]
  PIN Data_PMOS_NOSF[598]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2716.905 187.44 2717.185 188.44 ;
    END
  END Data_PMOS_NOSF[598]
  PIN Data_PMOS_NOSF[592]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2716.345 187.44 2716.625 188.44 ;
    END
  END Data_PMOS_NOSF[592]
  PIN Data_PMOS_NOSF[604]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2715.785 187.44 2716.065 188.44 ;
    END
  END Data_PMOS_NOSF[604]
  PIN Data_PMOS_NOSF[599]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2715.225 187.44 2715.505 188.44 ;
    END
  END Data_PMOS_NOSF[599]
  PIN Data_PMOS_NOSF[589]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2714.665 187.44 2714.945 188.44 ;
    END
  END Data_PMOS_NOSF[589]
  PIN Data_PMOS_NOSF[588]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2714.105 187.44 2714.385 188.44 ;
    END
  END Data_PMOS_NOSF[588]
  PIN Data_PMOS_NOSF[605]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2713.545 187.44 2713.825 188.44 ;
    END
  END Data_PMOS_NOSF[605]
  PIN DIG_MON_PMOS_NOSF[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2708.785 187.44 2709.065 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[56]
  PIN FREEZE_PMOS_NOSF[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2961.625 187.44 2961.905 188.44 ;
    END
  END FREEZE_PMOS_NOSF[31]
  PIN DIG_MON_PMOS_NOSF[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3798.265 187.44 3798.545 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[83]
  PIN Data_PMOS_NOSF[879]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3796.025 187.44 3796.305 188.44 ;
    END
  END Data_PMOS_NOSF[879]
  PIN Data_PMOS_NOSF[869]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3795.465 187.44 3795.745 188.44 ;
    END
  END Data_PMOS_NOSF[869]
  PIN Data_PMOS_NOSF[873]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3794.905 187.44 3795.185 188.44 ;
    END
  END Data_PMOS_NOSF[873]
  PIN Data_PMOS_NOSF[880]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3794.345 187.44 3794.625 188.44 ;
    END
  END Data_PMOS_NOSF[880]
  PIN Data_PMOS_NOSF[866]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3793.785 187.44 3794.065 188.44 ;
    END
  END Data_PMOS_NOSF[866]
  PIN Data_PMOS_NOSF[874]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3793.225 187.44 3793.505 188.44 ;
    END
  END Data_PMOS_NOSF[874]
  PIN Data_PMOS_NOSF[881]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3792.665 187.44 3792.945 188.44 ;
    END
  END Data_PMOS_NOSF[881]
  PIN Data_PMOS_NOSF[875]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3792.105 187.44 3792.385 188.44 ;
    END
  END Data_PMOS_NOSF[875]
  PIN Data_PMOS_NOSF[868]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3791.545 187.44 3791.825 188.44 ;
    END
  END Data_PMOS_NOSF[868]
  PIN Data_PMOS_NOSF[867]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3790.985 187.44 3791.265 188.44 ;
    END
  END Data_PMOS_NOSF[867]
  PIN nTOK_PMOS_NOSF[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3788.745 187.44 3789.025 188.44 ;
    END
  END nTOK_PMOS_NOSF[41]
  PIN FREEZE_PMOS_NOSF[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3772.505 187.44 3772.785 188.44 ;
    END
  END FREEZE_PMOS_NOSF[41]
  PIN Read_PMOS_NOSF[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3771.945 187.44 3772.225 188.44 ;
    END
  END Read_PMOS_NOSF[41]
  PIN Data_PMOS_NOSF[864]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3768.025 187.44 3768.305 188.44 ;
    END
  END Data_PMOS_NOSF[864]
  PIN Data_PMOS_NOSF[863]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3767.465 187.44 3767.745 188.44 ;
    END
  END Data_PMOS_NOSF[863]
  PIN Data_PMOS_NOSF[870]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3766.905 187.44 3767.185 188.44 ;
    END
  END Data_PMOS_NOSF[870]
  PIN Data_PMOS_NOSF[876]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3766.345 187.44 3766.625 188.44 ;
    END
  END Data_PMOS_NOSF[876]
  PIN Data_PMOS_NOSF[871]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3765.785 187.44 3766.065 188.44 ;
    END
  END Data_PMOS_NOSF[871]
  PIN Data_PMOS_NOSF[865]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3765.225 187.44 3765.505 188.44 ;
    END
  END Data_PMOS_NOSF[865]
  PIN Data_PMOS_NOSF[877]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3764.665 187.44 3764.945 188.44 ;
    END
  END Data_PMOS_NOSF[877]
  PIN Data_PMOS_NOSF[872]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3764.105 187.44 3764.385 188.44 ;
    END
  END Data_PMOS_NOSF[872]
  PIN Data_PMOS_NOSF[862]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3763.545 187.44 3763.825 188.44 ;
    END
  END Data_PMOS_NOSF[862]
  PIN Data_PMOS_NOSF[861]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3762.985 187.44 3763.265 188.44 ;
    END
  END Data_PMOS_NOSF[861]
  PIN Data_PMOS_NOSF[878]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3762.425 187.44 3762.705 188.44 ;
    END
  END Data_PMOS_NOSF[878]
  PIN DIG_MON_PMOS_NOSF[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3720.985 187.44 3721.265 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[82]
  PIN DIG_MON_PMOS_NOSF[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3716.505 187.44 3716.785 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[81]
  PIN Data_PMOS_NOSF[858]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3714.265 187.44 3714.545 188.44 ;
    END
  END Data_PMOS_NOSF[858]
  PIN Data_PMOS_NOSF[848]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3713.705 187.44 3713.985 188.44 ;
    END
  END Data_PMOS_NOSF[848]
  PIN Data_PMOS_NOSF[852]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3713.145 187.44 3713.425 188.44 ;
    END
  END Data_PMOS_NOSF[852]
  PIN Data_PMOS_NOSF[859]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3712.585 187.44 3712.865 188.44 ;
    END
  END Data_PMOS_NOSF[859]
  PIN Data_PMOS_NOSF[845]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3712.025 187.44 3712.305 188.44 ;
    END
  END Data_PMOS_NOSF[845]
  PIN Data_PMOS_NOSF[853]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3711.465 187.44 3711.745 188.44 ;
    END
  END Data_PMOS_NOSF[853]
  PIN Data_PMOS_NOSF[860]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3710.905 187.44 3711.185 188.44 ;
    END
  END Data_PMOS_NOSF[860]
  PIN Data_PMOS_NOSF[854]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3710.345 187.44 3710.625 188.44 ;
    END
  END Data_PMOS_NOSF[854]
  PIN Data_PMOS_NOSF[847]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3709.785 187.44 3710.065 188.44 ;
    END
  END Data_PMOS_NOSF[847]
  PIN Data_PMOS_NOSF[846]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3700.825 187.44 3701.105 188.44 ;
    END
  END Data_PMOS_NOSF[846]
  PIN nTOK_PMOS_NOSF[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3698.585 187.44 3698.865 188.44 ;
    END
  END nTOK_PMOS_NOSF[40]
  PIN FREEZE_PMOS_NOSF[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3695.785 187.44 3696.065 188.44 ;
    END
  END FREEZE_PMOS_NOSF[40]
  PIN Read_PMOS_NOSF[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3695.225 187.44 3695.505 188.44 ;
    END
  END Read_PMOS_NOSF[40]
  PIN Data_PMOS_NOSF[843]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3689.345 187.44 3689.625 188.44 ;
    END
  END Data_PMOS_NOSF[843]
  PIN Data_PMOS_NOSF[842]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3688.785 187.44 3689.065 188.44 ;
    END
  END Data_PMOS_NOSF[842]
  PIN Data_PMOS_NOSF[849]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3688.225 187.44 3688.505 188.44 ;
    END
  END Data_PMOS_NOSF[849]
  PIN Data_PMOS_NOSF[855]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3687.665 187.44 3687.945 188.44 ;
    END
  END Data_PMOS_NOSF[855]
  PIN Data_PMOS_NOSF[850]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3687.105 187.44 3687.385 188.44 ;
    END
  END Data_PMOS_NOSF[850]
  PIN Data_PMOS_NOSF[844]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3661.065 187.44 3661.345 188.44 ;
    END
  END Data_PMOS_NOSF[844]
  PIN Data_PMOS_NOSF[856]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3660.505 187.44 3660.785 188.44 ;
    END
  END Data_PMOS_NOSF[856]
  PIN Data_PMOS_NOSF[851]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3659.945 187.44 3660.225 188.44 ;
    END
  END Data_PMOS_NOSF[851]
  PIN Data_PMOS_NOSF[841]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3659.385 187.44 3659.665 188.44 ;
    END
  END Data_PMOS_NOSF[841]
  PIN Data_PMOS_NOSF[840]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3658.825 187.44 3659.105 188.44 ;
    END
  END Data_PMOS_NOSF[840]
  PIN Data_PMOS_NOSF[857]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3658.265 187.44 3658.545 188.44 ;
    END
  END Data_PMOS_NOSF[857]
  PIN DIG_MON_PMOS_NOSF[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3655.465 187.44 3655.745 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[80]
  PIN DIG_MON_PMOS_NOSF[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3650.985 187.44 3651.265 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[79]
  PIN Data_PMOS_NOSF[837]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3648.745 187.44 3649.025 188.44 ;
    END
  END Data_PMOS_NOSF[837]
  PIN Data_PMOS_NOSF[827]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3648.185 187.44 3648.465 188.44 ;
    END
  END Data_PMOS_NOSF[827]
  PIN Data_PMOS_NOSF[831]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3634.745 187.44 3635.025 188.44 ;
    END
  END Data_PMOS_NOSF[831]
  PIN Data_PMOS_NOSF[838]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3634.185 187.44 3634.465 188.44 ;
    END
  END Data_PMOS_NOSF[838]
  PIN Data_PMOS_NOSF[824]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3633.625 187.44 3633.905 188.44 ;
    END
  END Data_PMOS_NOSF[824]
  PIN Data_PMOS_NOSF[832]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3633.065 187.44 3633.345 188.44 ;
    END
  END Data_PMOS_NOSF[832]
  PIN Data_PMOS_NOSF[839]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3632.505 187.44 3632.785 188.44 ;
    END
  END Data_PMOS_NOSF[839]
  PIN Data_PMOS_NOSF[833]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3631.945 187.44 3632.225 188.44 ;
    END
  END Data_PMOS_NOSF[833]
  PIN Data_PMOS_NOSF[826]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3631.385 187.44 3631.665 188.44 ;
    END
  END Data_PMOS_NOSF[826]
  PIN Data_PMOS_NOSF[825]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3630.825 187.44 3631.105 188.44 ;
    END
  END Data_PMOS_NOSF[825]
  PIN nTOK_PMOS_NOSF[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3628.585 187.44 3628.865 188.44 ;
    END
  END nTOK_PMOS_NOSF[39]
  PIN FREEZE_PMOS_NOSF[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3625.785 187.44 3626.065 188.44 ;
    END
  END FREEZE_PMOS_NOSF[39]
  PIN Read_PMOS_NOSF[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3625.225 187.44 3625.505 188.44 ;
    END
  END Read_PMOS_NOSF[39]
  PIN Data_PMOS_NOSF[822]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3582.665 187.44 3582.945 188.44 ;
    END
  END Data_PMOS_NOSF[822]
  PIN Data_PMOS_NOSF[821]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3582.105 187.44 3582.385 188.44 ;
    END
  END Data_PMOS_NOSF[821]
  PIN Data_PMOS_NOSF[828]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3581.545 187.44 3581.825 188.44 ;
    END
  END Data_PMOS_NOSF[828]
  PIN Data_PMOS_NOSF[834]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3580.985 187.44 3581.265 188.44 ;
    END
  END Data_PMOS_NOSF[834]
  PIN Data_PMOS_NOSF[829]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3580.425 187.44 3580.705 188.44 ;
    END
  END Data_PMOS_NOSF[829]
  PIN Data_PMOS_NOSF[823]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3579.865 187.44 3580.145 188.44 ;
    END
  END Data_PMOS_NOSF[823]
  PIN Data_PMOS_NOSF[835]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3579.305 187.44 3579.585 188.44 ;
    END
  END Data_PMOS_NOSF[835]
  PIN Data_PMOS_NOSF[830]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3578.745 187.44 3579.025 188.44 ;
    END
  END Data_PMOS_NOSF[830]
  PIN Data_PMOS_NOSF[820]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3578.185 187.44 3578.465 188.44 ;
    END
  END Data_PMOS_NOSF[820]
  PIN Data_PMOS_NOSF[819]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3577.625 187.44 3577.905 188.44 ;
    END
  END Data_PMOS_NOSF[819]
  PIN Data_PMOS_NOSF[836]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3577.065 187.44 3577.345 188.44 ;
    END
  END Data_PMOS_NOSF[836]
  PIN DIG_MON_PMOS_NOSF[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3574.265 187.44 3574.545 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[78]
  PIN DIG_MON_PMOS_NOSF[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3569.785 187.44 3570.065 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[77]
  PIN Data_PMOS_NOSF[816]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3559.145 187.44 3559.425 188.44 ;
    END
  END Data_PMOS_NOSF[816]
  PIN Data_PMOS_NOSF[806]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3558.585 187.44 3558.865 188.44 ;
    END
  END Data_PMOS_NOSF[806]
  PIN Data_PMOS_NOSF[810]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3558.025 187.44 3558.305 188.44 ;
    END
  END Data_PMOS_NOSF[810]
  PIN Data_PMOS_NOSF[817]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3557.465 187.44 3557.745 188.44 ;
    END
  END Data_PMOS_NOSF[817]
  PIN Data_PMOS_NOSF[803]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3556.905 187.44 3557.185 188.44 ;
    END
  END Data_PMOS_NOSF[803]
  PIN Data_PMOS_NOSF[811]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3556.345 187.44 3556.625 188.44 ;
    END
  END Data_PMOS_NOSF[811]
  PIN Data_PMOS_NOSF[818]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3555.785 187.44 3556.065 188.44 ;
    END
  END Data_PMOS_NOSF[818]
  PIN Data_PMOS_NOSF[812]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3555.225 187.44 3555.505 188.44 ;
    END
  END Data_PMOS_NOSF[812]
  PIN Data_PMOS_NOSF[805]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3554.665 187.44 3554.945 188.44 ;
    END
  END Data_PMOS_NOSF[805]
  PIN Data_PMOS_NOSF[804]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3554.105 187.44 3554.385 188.44 ;
    END
  END Data_PMOS_NOSF[804]
  PIN nTOK_PMOS_NOSF[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3549.905 187.44 3550.185 188.44 ;
    END
  END nTOK_PMOS_NOSF[38]
  PIN Read_PMOS_NOSF[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3521.065 187.44 3521.345 188.44 ;
    END
  END Read_PMOS_NOSF[38]
  PIN Data_PMOS_NOSF[801]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3517.145 187.44 3517.425 188.44 ;
    END
  END Data_PMOS_NOSF[801]
  PIN Data_PMOS_NOSF[800]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3516.585 187.44 3516.865 188.44 ;
    END
  END Data_PMOS_NOSF[800]
  PIN Data_PMOS_NOSF[807]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3516.025 187.44 3516.305 188.44 ;
    END
  END Data_PMOS_NOSF[807]
  PIN Data_PMOS_NOSF[813]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3515.465 187.44 3515.745 188.44 ;
    END
  END Data_PMOS_NOSF[813]
  PIN Data_PMOS_NOSF[808]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3514.905 187.44 3515.185 188.44 ;
    END
  END Data_PMOS_NOSF[808]
  PIN Data_PMOS_NOSF[802]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3514.345 187.44 3514.625 188.44 ;
    END
  END Data_PMOS_NOSF[802]
  PIN Data_PMOS_NOSF[814]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3513.785 187.44 3514.065 188.44 ;
    END
  END Data_PMOS_NOSF[814]
  PIN Data_PMOS_NOSF[809]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3513.225 187.44 3513.505 188.44 ;
    END
  END Data_PMOS_NOSF[809]
  PIN Data_PMOS_NOSF[799]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3512.665 187.44 3512.945 188.44 ;
    END
  END Data_PMOS_NOSF[799]
  PIN Data_PMOS_NOSF[798]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3512.105 187.44 3512.385 188.44 ;
    END
  END Data_PMOS_NOSF[798]
  PIN Data_PMOS_NOSF[815]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3511.545 187.44 3511.825 188.44 ;
    END
  END Data_PMOS_NOSF[815]
  PIN DIG_MON_PMOS_NOSF[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3508.745 187.44 3509.025 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[76]
  PIN DIG_MON_PMOS_NOSF[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3491.385 187.44 3491.665 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[75]
  PIN Data_PMOS_NOSF[795]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3489.145 187.44 3489.425 188.44 ;
    END
  END Data_PMOS_NOSF[795]
  PIN Data_PMOS_NOSF[785]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3488.585 187.44 3488.865 188.44 ;
    END
  END Data_PMOS_NOSF[785]
  PIN Data_PMOS_NOSF[789]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3488.025 187.44 3488.305 188.44 ;
    END
  END Data_PMOS_NOSF[789]
  PIN Data_PMOS_NOSF[796]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3487.465 187.44 3487.745 188.44 ;
    END
  END Data_PMOS_NOSF[796]
  PIN Data_PMOS_NOSF[782]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3486.905 187.44 3487.185 188.44 ;
    END
  END Data_PMOS_NOSF[782]
  PIN Data_PMOS_NOSF[790]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3486.345 187.44 3486.625 188.44 ;
    END
  END Data_PMOS_NOSF[790]
  PIN Data_PMOS_NOSF[797]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3485.785 187.44 3486.065 188.44 ;
    END
  END Data_PMOS_NOSF[797]
  PIN Data_PMOS_NOSF[791]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3485.225 187.44 3485.505 188.44 ;
    END
  END Data_PMOS_NOSF[791]
  PIN Data_PMOS_NOSF[784]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3484.665 187.44 3484.945 188.44 ;
    END
  END Data_PMOS_NOSF[784]
  PIN Data_PMOS_NOSF[783]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3484.105 187.44 3484.385 188.44 ;
    END
  END Data_PMOS_NOSF[783]
  PIN nTOK_PMOS_NOSF[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3442.665 187.44 3442.945 188.44 ;
    END
  END nTOK_PMOS_NOSF[37]
  PIN FREEZE_PMOS_NOSF[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3439.865 187.44 3440.145 188.44 ;
    END
  END FREEZE_PMOS_NOSF[37]
  PIN Read_PMOS_NOSF[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3439.305 187.44 3439.585 188.44 ;
    END
  END Read_PMOS_NOSF[37]
  PIN Data_PMOS_NOSF[780]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3435.385 187.44 3435.665 188.44 ;
    END
  END Data_PMOS_NOSF[780]
  PIN Data_PMOS_NOSF[779]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3434.825 187.44 3435.105 188.44 ;
    END
  END Data_PMOS_NOSF[779]
  PIN Data_PMOS_NOSF[786]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3434.265 187.44 3434.545 188.44 ;
    END
  END Data_PMOS_NOSF[786]
  PIN Data_PMOS_NOSF[792]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3433.705 187.44 3433.985 188.44 ;
    END
  END Data_PMOS_NOSF[792]
  PIN Data_PMOS_NOSF[787]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3433.145 187.44 3433.425 188.44 ;
    END
  END Data_PMOS_NOSF[787]
  PIN Data_PMOS_NOSF[781]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3432.585 187.44 3432.865 188.44 ;
    END
  END Data_PMOS_NOSF[781]
  PIN Data_PMOS_NOSF[793]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3432.025 187.44 3432.305 188.44 ;
    END
  END Data_PMOS_NOSF[793]
  PIN Data_PMOS_NOSF[788]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3431.465 187.44 3431.745 188.44 ;
    END
  END Data_PMOS_NOSF[788]
  PIN Data_PMOS_NOSF[778]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3430.905 187.44 3431.185 188.44 ;
    END
  END Data_PMOS_NOSF[778]
  PIN Data_PMOS_NOSF[777]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3430.345 187.44 3430.625 188.44 ;
    END
  END Data_PMOS_NOSF[777]
  PIN Data_PMOS_NOSF[794]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3429.785 187.44 3430.065 188.44 ;
    END
  END Data_PMOS_NOSF[794]
  PIN DIG_MON_PMOS_NOSF[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3418.585 187.44 3418.865 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[74]
  PIN DIG_MON_PMOS_NOSF[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3414.105 187.44 3414.385 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[73]
  PIN Data_PMOS_NOSF[774]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3409.905 187.44 3410.185 188.44 ;
    END
  END Data_PMOS_NOSF[774]
  PIN Data_PMOS_NOSF[764]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3409.345 187.44 3409.625 188.44 ;
    END
  END Data_PMOS_NOSF[764]
  PIN Data_PMOS_NOSF[768]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3408.785 187.44 3409.065 188.44 ;
    END
  END Data_PMOS_NOSF[768]
  PIN Data_PMOS_NOSF[775]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3408.225 187.44 3408.505 188.44 ;
    END
  END Data_PMOS_NOSF[775]
  PIN Data_PMOS_NOSF[761]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3407.665 187.44 3407.945 188.44 ;
    END
  END Data_PMOS_NOSF[761]
  PIN Data_PMOS_NOSF[769]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3381.625 187.44 3381.905 188.44 ;
    END
  END Data_PMOS_NOSF[769]
  PIN Data_PMOS_NOSF[776]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3381.065 187.44 3381.345 188.44 ;
    END
  END Data_PMOS_NOSF[776]
  PIN Data_PMOS_NOSF[770]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3380.505 187.44 3380.785 188.44 ;
    END
  END Data_PMOS_NOSF[770]
  PIN Data_PMOS_NOSF[763]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3379.945 187.44 3380.225 188.44 ;
    END
  END Data_PMOS_NOSF[763]
  PIN Data_PMOS_NOSF[762]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3379.385 187.44 3379.665 188.44 ;
    END
  END Data_PMOS_NOSF[762]
  PIN nTOK_PMOS_NOSF[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3377.145 187.44 3377.425 188.44 ;
    END
  END nTOK_PMOS_NOSF[36]
  PIN FREEZE_PMOS_NOSF[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3374.345 187.44 3374.625 188.44 ;
    END
  END FREEZE_PMOS_NOSF[36]
  PIN Read_PMOS_NOSF[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3373.785 187.44 3374.065 188.44 ;
    END
  END Read_PMOS_NOSF[36]
  PIN Data_PMOS_NOSF[759]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3369.865 187.44 3370.145 188.44 ;
    END
  END Data_PMOS_NOSF[759]
  PIN Data_PMOS_NOSF[758]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3369.305 187.44 3369.585 188.44 ;
    END
  END Data_PMOS_NOSF[758]
  PIN Data_PMOS_NOSF[765]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3368.745 187.44 3369.025 188.44 ;
    END
  END Data_PMOS_NOSF[765]
  PIN Data_PMOS_NOSF[771]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3355.305 187.44 3355.585 188.44 ;
    END
  END Data_PMOS_NOSF[771]
  PIN Data_PMOS_NOSF[766]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3354.745 187.44 3355.025 188.44 ;
    END
  END Data_PMOS_NOSF[766]
  PIN Data_PMOS_NOSF[760]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3354.185 187.44 3354.465 188.44 ;
    END
  END Data_PMOS_NOSF[760]
  PIN Data_PMOS_NOSF[772]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3353.625 187.44 3353.905 188.44 ;
    END
  END Data_PMOS_NOSF[772]
  PIN Data_PMOS_NOSF[767]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3353.065 187.44 3353.345 188.44 ;
    END
  END Data_PMOS_NOSF[767]
  PIN Data_PMOS_NOSF[757]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3352.505 187.44 3352.785 188.44 ;
    END
  END Data_PMOS_NOSF[757]
  PIN Data_PMOS_NOSF[756]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3351.945 187.44 3352.225 188.44 ;
    END
  END Data_PMOS_NOSF[756]
  PIN Data_PMOS_NOSF[773]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3351.385 187.44 3351.665 188.44 ;
    END
  END Data_PMOS_NOSF[773]
  PIN DIG_MON_PMOS_NOSF[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3348.585 187.44 3348.865 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[72]
  PIN DIG_MON_PMOS_NOSF[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3344.105 187.44 3344.385 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[71]
  PIN Data_PMOS_NOSF[753]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3302.105 187.44 3302.385 188.44 ;
    END
  END Data_PMOS_NOSF[753]
  PIN Data_PMOS_NOSF[743]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3301.545 187.44 3301.825 188.44 ;
    END
  END Data_PMOS_NOSF[743]
  PIN Data_PMOS_NOSF[747]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3300.985 187.44 3301.265 188.44 ;
    END
  END Data_PMOS_NOSF[747]
  PIN Data_PMOS_NOSF[754]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3300.425 187.44 3300.705 188.44 ;
    END
  END Data_PMOS_NOSF[754]
  PIN Data_PMOS_NOSF[740]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3299.865 187.44 3300.145 188.44 ;
    END
  END Data_PMOS_NOSF[740]
  PIN Data_PMOS_NOSF[748]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3299.305 187.44 3299.585 188.44 ;
    END
  END Data_PMOS_NOSF[748]
  PIN Data_PMOS_NOSF[755]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3298.745 187.44 3299.025 188.44 ;
    END
  END Data_PMOS_NOSF[755]
  PIN Data_PMOS_NOSF[749]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3298.185 187.44 3298.465 188.44 ;
    END
  END Data_PMOS_NOSF[749]
  PIN Data_PMOS_NOSF[742]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3297.625 187.44 3297.905 188.44 ;
    END
  END Data_PMOS_NOSF[742]
  PIN Data_PMOS_NOSF[741]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3297.065 187.44 3297.345 188.44 ;
    END
  END Data_PMOS_NOSF[741]
  PIN nTOK_PMOS_NOSF[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3294.825 187.44 3295.105 188.44 ;
    END
  END nTOK_PMOS_NOSF[35]
  PIN FREEZE_PMOS_NOSF[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3292.025 187.44 3292.305 188.44 ;
    END
  END FREEZE_PMOS_NOSF[35]
  PIN Read_PMOS_NOSF[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3291.465 187.44 3291.745 188.44 ;
    END
  END Read_PMOS_NOSF[35]
  PIN Data_PMOS_NOSF[738]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3279.145 187.44 3279.425 188.44 ;
    END
  END Data_PMOS_NOSF[738]
  PIN Data_PMOS_NOSF[737]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3278.585 187.44 3278.865 188.44 ;
    END
  END Data_PMOS_NOSF[737]
  PIN Data_PMOS_NOSF[750]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3277.465 187.44 3277.745 188.44 ;
    END
  END Data_PMOS_NOSF[750]
  PIN Data_PMOS_NOSF[744]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3278.025 187.44 3278.305 188.44 ;
    END
  END Data_PMOS_NOSF[744]
  PIN Data_PMOS_NOSF[745]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3276.905 187.44 3277.185 188.44 ;
    END
  END Data_PMOS_NOSF[745]
  PIN Data_PMOS_NOSF[739]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3276.345 187.44 3276.625 188.44 ;
    END
  END Data_PMOS_NOSF[739]
  PIN Data_PMOS_NOSF[751]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3275.785 187.44 3276.065 188.44 ;
    END
  END Data_PMOS_NOSF[751]
  PIN Data_PMOS_NOSF[746]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3275.225 187.44 3275.505 188.44 ;
    END
  END Data_PMOS_NOSF[746]
  PIN Data_PMOS_NOSF[736]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3274.665 187.44 3274.945 188.44 ;
    END
  END Data_PMOS_NOSF[736]
  PIN Data_PMOS_NOSF[735]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3274.105 187.44 3274.385 188.44 ;
    END
  END Data_PMOS_NOSF[735]
  PIN Data_PMOS_NOSF[752]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3273.545 187.44 3273.825 188.44 ;
    END
  END Data_PMOS_NOSF[752]
  PIN DIG_MON_PMOS_NOSF[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3268.785 187.44 3269.065 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[70]
  PIN FREEZE_PMOS_NOSF[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3521.625 187.44 3521.905 188.44 ;
    END
  END FREEZE_PMOS_NOSF[38]
  PIN DIG_MON_PMOS_NOSF[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4358.265 187.44 4358.545 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[97]
  PIN Data_PMOS_NOSF[1026]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4356.025 187.44 4356.305 188.44 ;
    END
  END Data_PMOS_NOSF[1026]
  PIN Data_PMOS_NOSF[1016]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4355.465 187.44 4355.745 188.44 ;
    END
  END Data_PMOS_NOSF[1016]
  PIN Data_PMOS_NOSF[1020]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4354.905 187.44 4355.185 188.44 ;
    END
  END Data_PMOS_NOSF[1020]
  PIN Data_PMOS_NOSF[1027]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4354.345 187.44 4354.625 188.44 ;
    END
  END Data_PMOS_NOSF[1027]
  PIN Data_PMOS_NOSF[1013]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4353.785 187.44 4354.065 188.44 ;
    END
  END Data_PMOS_NOSF[1013]
  PIN Data_PMOS_NOSF[1021]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4353.225 187.44 4353.505 188.44 ;
    END
  END Data_PMOS_NOSF[1021]
  PIN Data_PMOS_NOSF[1028]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4352.665 187.44 4352.945 188.44 ;
    END
  END Data_PMOS_NOSF[1028]
  PIN Data_PMOS_NOSF[1022]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4352.105 187.44 4352.385 188.44 ;
    END
  END Data_PMOS_NOSF[1022]
  PIN Data_PMOS_NOSF[1015]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4351.545 187.44 4351.825 188.44 ;
    END
  END Data_PMOS_NOSF[1015]
  PIN Data_PMOS_NOSF[1014]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4350.985 187.44 4351.265 188.44 ;
    END
  END Data_PMOS_NOSF[1014]
  PIN nTOK_PMOS_NOSF[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4348.745 187.44 4349.025 188.44 ;
    END
  END nTOK_PMOS_NOSF[48]
  PIN FREEZE_PMOS_NOSF[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4332.505 187.44 4332.785 188.44 ;
    END
  END FREEZE_PMOS_NOSF[48]
  PIN Read_PMOS_NOSF[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4331.945 187.44 4332.225 188.44 ;
    END
  END Read_PMOS_NOSF[48]
  PIN Data_PMOS_NOSF[1011]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4328.025 187.44 4328.305 188.44 ;
    END
  END Data_PMOS_NOSF[1011]
  PIN Data_PMOS_NOSF[1010]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4327.465 187.44 4327.745 188.44 ;
    END
  END Data_PMOS_NOSF[1010]
  PIN Data_PMOS_NOSF[1017]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4326.905 187.44 4327.185 188.44 ;
    END
  END Data_PMOS_NOSF[1017]
  PIN Data_PMOS_NOSF[1023]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4326.345 187.44 4326.625 188.44 ;
    END
  END Data_PMOS_NOSF[1023]
  PIN Data_PMOS_NOSF[1018]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4325.785 187.44 4326.065 188.44 ;
    END
  END Data_PMOS_NOSF[1018]
  PIN Data_PMOS_NOSF[1012]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4325.225 187.44 4325.505 188.44 ;
    END
  END Data_PMOS_NOSF[1012]
  PIN Data_PMOS_NOSF[1024]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4324.665 187.44 4324.945 188.44 ;
    END
  END Data_PMOS_NOSF[1024]
  PIN Data_PMOS_NOSF[1019]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4324.105 187.44 4324.385 188.44 ;
    END
  END Data_PMOS_NOSF[1019]
  PIN Data_PMOS_NOSF[1009]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4323.545 187.44 4323.825 188.44 ;
    END
  END Data_PMOS_NOSF[1009]
  PIN Data_PMOS_NOSF[1008]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4322.985 187.44 4323.265 188.44 ;
    END
  END Data_PMOS_NOSF[1008]
  PIN Data_PMOS_NOSF[1025]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4322.425 187.44 4322.705 188.44 ;
    END
  END Data_PMOS_NOSF[1025]
  PIN DIG_MON_PMOS_NOSF[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4280.985 187.44 4281.265 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[96]
  PIN DIG_MON_PMOS_NOSF[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4276.505 187.44 4276.785 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[95]
  PIN Data_PMOS_NOSF[1005]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4274.265 187.44 4274.545 188.44 ;
    END
  END Data_PMOS_NOSF[1005]
  PIN Data_PMOS_NOSF[995]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4273.705 187.44 4273.985 188.44 ;
    END
  END Data_PMOS_NOSF[995]
  PIN Data_PMOS_NOSF[999]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4273.145 187.44 4273.425 188.44 ;
    END
  END Data_PMOS_NOSF[999]
  PIN Data_PMOS_NOSF[1006]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4272.585 187.44 4272.865 188.44 ;
    END
  END Data_PMOS_NOSF[1006]
  PIN Data_PMOS_NOSF[992]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4272.025 187.44 4272.305 188.44 ;
    END
  END Data_PMOS_NOSF[992]
  PIN Data_PMOS_NOSF[1000]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4271.465 187.44 4271.745 188.44 ;
    END
  END Data_PMOS_NOSF[1000]
  PIN Data_PMOS_NOSF[1007]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4270.905 187.44 4271.185 188.44 ;
    END
  END Data_PMOS_NOSF[1007]
  PIN Data_PMOS_NOSF[1001]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4270.345 187.44 4270.625 188.44 ;
    END
  END Data_PMOS_NOSF[1001]
  PIN Data_PMOS_NOSF[994]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4269.785 187.44 4270.065 188.44 ;
    END
  END Data_PMOS_NOSF[994]
  PIN Data_PMOS_NOSF[993]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4260.825 187.44 4261.105 188.44 ;
    END
  END Data_PMOS_NOSF[993]
  PIN nTOK_PMOS_NOSF[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4258.585 187.44 4258.865 188.44 ;
    END
  END nTOK_PMOS_NOSF[47]
  PIN FREEZE_PMOS_NOSF[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4255.785 187.44 4256.065 188.44 ;
    END
  END FREEZE_PMOS_NOSF[47]
  PIN Read_PMOS_NOSF[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4255.225 187.44 4255.505 188.44 ;
    END
  END Read_PMOS_NOSF[47]
  PIN Data_PMOS_NOSF[990]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4249.345 187.44 4249.625 188.44 ;
    END
  END Data_PMOS_NOSF[990]
  PIN Data_PMOS_NOSF[989]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4248.785 187.44 4249.065 188.44 ;
    END
  END Data_PMOS_NOSF[989]
  PIN Data_PMOS_NOSF[996]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4248.225 187.44 4248.505 188.44 ;
    END
  END Data_PMOS_NOSF[996]
  PIN Data_PMOS_NOSF[1002]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4247.665 187.44 4247.945 188.44 ;
    END
  END Data_PMOS_NOSF[1002]
  PIN Data_PMOS_NOSF[997]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4247.105 187.44 4247.385 188.44 ;
    END
  END Data_PMOS_NOSF[997]
  PIN Data_PMOS_NOSF[991]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4221.065 187.44 4221.345 188.44 ;
    END
  END Data_PMOS_NOSF[991]
  PIN Data_PMOS_NOSF[1003]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4220.505 187.44 4220.785 188.44 ;
    END
  END Data_PMOS_NOSF[1003]
  PIN Data_PMOS_NOSF[998]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4219.945 187.44 4220.225 188.44 ;
    END
  END Data_PMOS_NOSF[998]
  PIN Data_PMOS_NOSF[988]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4219.385 187.44 4219.665 188.44 ;
    END
  END Data_PMOS_NOSF[988]
  PIN Data_PMOS_NOSF[987]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4218.825 187.44 4219.105 188.44 ;
    END
  END Data_PMOS_NOSF[987]
  PIN Data_PMOS_NOSF[1004]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4218.265 187.44 4218.545 188.44 ;
    END
  END Data_PMOS_NOSF[1004]
  PIN DIG_MON_PMOS_NOSF[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4215.465 187.44 4215.745 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[94]
  PIN DIG_MON_PMOS_NOSF[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4210.985 187.44 4211.265 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[93]
  PIN Data_PMOS_NOSF[984]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4208.745 187.44 4209.025 188.44 ;
    END
  END Data_PMOS_NOSF[984]
  PIN Data_PMOS_NOSF[974]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4208.185 187.44 4208.465 188.44 ;
    END
  END Data_PMOS_NOSF[974]
  PIN Data_PMOS_NOSF[978]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4194.745 187.44 4195.025 188.44 ;
    END
  END Data_PMOS_NOSF[978]
  PIN Data_PMOS_NOSF[985]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4194.185 187.44 4194.465 188.44 ;
    END
  END Data_PMOS_NOSF[985]
  PIN Data_PMOS_NOSF[971]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4193.625 187.44 4193.905 188.44 ;
    END
  END Data_PMOS_NOSF[971]
  PIN Data_PMOS_NOSF[979]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4193.065 187.44 4193.345 188.44 ;
    END
  END Data_PMOS_NOSF[979]
  PIN Data_PMOS_NOSF[986]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4192.505 187.44 4192.785 188.44 ;
    END
  END Data_PMOS_NOSF[986]
  PIN Data_PMOS_NOSF[980]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4191.945 187.44 4192.225 188.44 ;
    END
  END Data_PMOS_NOSF[980]
  PIN Data_PMOS_NOSF[973]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4191.385 187.44 4191.665 188.44 ;
    END
  END Data_PMOS_NOSF[973]
  PIN Data_PMOS_NOSF[972]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4190.825 187.44 4191.105 188.44 ;
    END
  END Data_PMOS_NOSF[972]
  PIN nTOK_PMOS_NOSF[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4188.585 187.44 4188.865 188.44 ;
    END
  END nTOK_PMOS_NOSF[46]
  PIN FREEZE_PMOS_NOSF[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4185.785 187.44 4186.065 188.44 ;
    END
  END FREEZE_PMOS_NOSF[46]
  PIN Read_PMOS_NOSF[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4185.225 187.44 4185.505 188.44 ;
    END
  END Read_PMOS_NOSF[46]
  PIN Data_PMOS_NOSF[969]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4142.665 187.44 4142.945 188.44 ;
    END
  END Data_PMOS_NOSF[969]
  PIN Data_PMOS_NOSF[968]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4142.105 187.44 4142.385 188.44 ;
    END
  END Data_PMOS_NOSF[968]
  PIN Data_PMOS_NOSF[975]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4141.545 187.44 4141.825 188.44 ;
    END
  END Data_PMOS_NOSF[975]
  PIN Data_PMOS_NOSF[981]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4140.985 187.44 4141.265 188.44 ;
    END
  END Data_PMOS_NOSF[981]
  PIN Data_PMOS_NOSF[976]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4140.425 187.44 4140.705 188.44 ;
    END
  END Data_PMOS_NOSF[976]
  PIN Data_PMOS_NOSF[970]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4139.865 187.44 4140.145 188.44 ;
    END
  END Data_PMOS_NOSF[970]
  PIN Data_PMOS_NOSF[982]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4139.305 187.44 4139.585 188.44 ;
    END
  END Data_PMOS_NOSF[982]
  PIN Data_PMOS_NOSF[977]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4138.745 187.44 4139.025 188.44 ;
    END
  END Data_PMOS_NOSF[977]
  PIN Data_PMOS_NOSF[967]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4138.185 187.44 4138.465 188.44 ;
    END
  END Data_PMOS_NOSF[967]
  PIN Data_PMOS_NOSF[966]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4137.625 187.44 4137.905 188.44 ;
    END
  END Data_PMOS_NOSF[966]
  PIN Data_PMOS_NOSF[983]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4137.065 187.44 4137.345 188.44 ;
    END
  END Data_PMOS_NOSF[983]
  PIN DIG_MON_PMOS_NOSF[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4134.265 187.44 4134.545 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[92]
  PIN DIG_MON_PMOS_NOSF[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4129.785 187.44 4130.065 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[91]
  PIN Data_PMOS_NOSF[963]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4119.145 187.44 4119.425 188.44 ;
    END
  END Data_PMOS_NOSF[963]
  PIN Data_PMOS_NOSF[953]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4118.585 187.44 4118.865 188.44 ;
    END
  END Data_PMOS_NOSF[953]
  PIN Data_PMOS_NOSF[957]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4118.025 187.44 4118.305 188.44 ;
    END
  END Data_PMOS_NOSF[957]
  PIN Data_PMOS_NOSF[964]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4117.465 187.44 4117.745 188.44 ;
    END
  END Data_PMOS_NOSF[964]
  PIN Data_PMOS_NOSF[950]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4116.905 187.44 4117.185 188.44 ;
    END
  END Data_PMOS_NOSF[950]
  PIN Data_PMOS_NOSF[958]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4116.345 187.44 4116.625 188.44 ;
    END
  END Data_PMOS_NOSF[958]
  PIN Data_PMOS_NOSF[965]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4115.785 187.44 4116.065 188.44 ;
    END
  END Data_PMOS_NOSF[965]
  PIN Data_PMOS_NOSF[959]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4115.225 187.44 4115.505 188.44 ;
    END
  END Data_PMOS_NOSF[959]
  PIN Data_PMOS_NOSF[952]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4114.665 187.44 4114.945 188.44 ;
    END
  END Data_PMOS_NOSF[952]
  PIN Data_PMOS_NOSF[951]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4114.105 187.44 4114.385 188.44 ;
    END
  END Data_PMOS_NOSF[951]
  PIN nTOK_PMOS_NOSF[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4109.905 187.44 4110.185 188.44 ;
    END
  END nTOK_PMOS_NOSF[45]
  PIN Read_PMOS_NOSF[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4081.065 187.44 4081.345 188.44 ;
    END
  END Read_PMOS_NOSF[45]
  PIN Data_PMOS_NOSF[948]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4077.145 187.44 4077.425 188.44 ;
    END
  END Data_PMOS_NOSF[948]
  PIN Data_PMOS_NOSF[947]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4076.585 187.44 4076.865 188.44 ;
    END
  END Data_PMOS_NOSF[947]
  PIN Data_PMOS_NOSF[954]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4076.025 187.44 4076.305 188.44 ;
    END
  END Data_PMOS_NOSF[954]
  PIN Data_PMOS_NOSF[960]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4075.465 187.44 4075.745 188.44 ;
    END
  END Data_PMOS_NOSF[960]
  PIN Data_PMOS_NOSF[955]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4074.905 187.44 4075.185 188.44 ;
    END
  END Data_PMOS_NOSF[955]
  PIN Data_PMOS_NOSF[949]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4074.345 187.44 4074.625 188.44 ;
    END
  END Data_PMOS_NOSF[949]
  PIN Data_PMOS_NOSF[961]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4073.785 187.44 4074.065 188.44 ;
    END
  END Data_PMOS_NOSF[961]
  PIN Data_PMOS_NOSF[956]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4073.225 187.44 4073.505 188.44 ;
    END
  END Data_PMOS_NOSF[956]
  PIN Data_PMOS_NOSF[946]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4072.665 187.44 4072.945 188.44 ;
    END
  END Data_PMOS_NOSF[946]
  PIN Data_PMOS_NOSF[945]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4072.105 187.44 4072.385 188.44 ;
    END
  END Data_PMOS_NOSF[945]
  PIN Data_PMOS_NOSF[962]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4071.545 187.44 4071.825 188.44 ;
    END
  END Data_PMOS_NOSF[962]
  PIN DIG_MON_PMOS_NOSF[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4068.745 187.44 4069.025 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[90]
  PIN DIG_MON_PMOS_NOSF[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4051.385 187.44 4051.665 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[89]
  PIN Data_PMOS_NOSF[942]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4049.145 187.44 4049.425 188.44 ;
    END
  END Data_PMOS_NOSF[942]
  PIN Data_PMOS_NOSF[932]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4048.585 187.44 4048.865 188.44 ;
    END
  END Data_PMOS_NOSF[932]
  PIN Data_PMOS_NOSF[936]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4048.025 187.44 4048.305 188.44 ;
    END
  END Data_PMOS_NOSF[936]
  PIN Data_PMOS_NOSF[943]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4047.465 187.44 4047.745 188.44 ;
    END
  END Data_PMOS_NOSF[943]
  PIN Data_PMOS_NOSF[929]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4046.905 187.44 4047.185 188.44 ;
    END
  END Data_PMOS_NOSF[929]
  PIN Data_PMOS_NOSF[937]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4046.345 187.44 4046.625 188.44 ;
    END
  END Data_PMOS_NOSF[937]
  PIN Data_PMOS_NOSF[944]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4045.785 187.44 4046.065 188.44 ;
    END
  END Data_PMOS_NOSF[944]
  PIN Data_PMOS_NOSF[938]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4045.225 187.44 4045.505 188.44 ;
    END
  END Data_PMOS_NOSF[938]
  PIN Data_PMOS_NOSF[931]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4044.665 187.44 4044.945 188.44 ;
    END
  END Data_PMOS_NOSF[931]
  PIN Data_PMOS_NOSF[930]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4044.105 187.44 4044.385 188.44 ;
    END
  END Data_PMOS_NOSF[930]
  PIN nTOK_PMOS_NOSF[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4002.665 187.44 4002.945 188.44 ;
    END
  END nTOK_PMOS_NOSF[44]
  PIN FREEZE_PMOS_NOSF[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3999.865 187.44 4000.145 188.44 ;
    END
  END FREEZE_PMOS_NOSF[44]
  PIN Read_PMOS_NOSF[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3999.305 187.44 3999.585 188.44 ;
    END
  END Read_PMOS_NOSF[44]
  PIN Data_PMOS_NOSF[927]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3995.385 187.44 3995.665 188.44 ;
    END
  END Data_PMOS_NOSF[927]
  PIN Data_PMOS_NOSF[926]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3994.825 187.44 3995.105 188.44 ;
    END
  END Data_PMOS_NOSF[926]
  PIN Data_PMOS_NOSF[933]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3994.265 187.44 3994.545 188.44 ;
    END
  END Data_PMOS_NOSF[933]
  PIN Data_PMOS_NOSF[939]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3993.705 187.44 3993.985 188.44 ;
    END
  END Data_PMOS_NOSF[939]
  PIN Data_PMOS_NOSF[934]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3993.145 187.44 3993.425 188.44 ;
    END
  END Data_PMOS_NOSF[934]
  PIN Data_PMOS_NOSF[928]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3992.585 187.44 3992.865 188.44 ;
    END
  END Data_PMOS_NOSF[928]
  PIN Data_PMOS_NOSF[940]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3992.025 187.44 3992.305 188.44 ;
    END
  END Data_PMOS_NOSF[940]
  PIN Data_PMOS_NOSF[935]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3991.465 187.44 3991.745 188.44 ;
    END
  END Data_PMOS_NOSF[935]
  PIN Data_PMOS_NOSF[925]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3990.905 187.44 3991.185 188.44 ;
    END
  END Data_PMOS_NOSF[925]
  PIN Data_PMOS_NOSF[924]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3990.345 187.44 3990.625 188.44 ;
    END
  END Data_PMOS_NOSF[924]
  PIN Data_PMOS_NOSF[941]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3989.785 187.44 3990.065 188.44 ;
    END
  END Data_PMOS_NOSF[941]
  PIN DIG_MON_PMOS_NOSF[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3978.585 187.44 3978.865 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[88]
  PIN DIG_MON_PMOS_NOSF[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3974.105 187.44 3974.385 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[87]
  PIN Data_PMOS_NOSF[921]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3969.905 187.44 3970.185 188.44 ;
    END
  END Data_PMOS_NOSF[921]
  PIN Data_PMOS_NOSF[911]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3969.345 187.44 3969.625 188.44 ;
    END
  END Data_PMOS_NOSF[911]
  PIN Data_PMOS_NOSF[915]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3968.785 187.44 3969.065 188.44 ;
    END
  END Data_PMOS_NOSF[915]
  PIN Data_PMOS_NOSF[922]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3968.225 187.44 3968.505 188.44 ;
    END
  END Data_PMOS_NOSF[922]
  PIN Data_PMOS_NOSF[908]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3967.665 187.44 3967.945 188.44 ;
    END
  END Data_PMOS_NOSF[908]
  PIN Data_PMOS_NOSF[916]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3941.625 187.44 3941.905 188.44 ;
    END
  END Data_PMOS_NOSF[916]
  PIN Data_PMOS_NOSF[923]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3941.065 187.44 3941.345 188.44 ;
    END
  END Data_PMOS_NOSF[923]
  PIN Data_PMOS_NOSF[917]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3940.505 187.44 3940.785 188.44 ;
    END
  END Data_PMOS_NOSF[917]
  PIN Data_PMOS_NOSF[910]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3939.945 187.44 3940.225 188.44 ;
    END
  END Data_PMOS_NOSF[910]
  PIN Data_PMOS_NOSF[909]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3939.385 187.44 3939.665 188.44 ;
    END
  END Data_PMOS_NOSF[909]
  PIN nTOK_PMOS_NOSF[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3937.145 187.44 3937.425 188.44 ;
    END
  END nTOK_PMOS_NOSF[43]
  PIN FREEZE_PMOS_NOSF[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3934.345 187.44 3934.625 188.44 ;
    END
  END FREEZE_PMOS_NOSF[43]
  PIN Read_PMOS_NOSF[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3933.785 187.44 3934.065 188.44 ;
    END
  END Read_PMOS_NOSF[43]
  PIN Data_PMOS_NOSF[906]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3929.865 187.44 3930.145 188.44 ;
    END
  END Data_PMOS_NOSF[906]
  PIN Data_PMOS_NOSF[905]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3929.305 187.44 3929.585 188.44 ;
    END
  END Data_PMOS_NOSF[905]
  PIN Data_PMOS_NOSF[912]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3928.745 187.44 3929.025 188.44 ;
    END
  END Data_PMOS_NOSF[912]
  PIN Data_PMOS_NOSF[918]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3915.305 187.44 3915.585 188.44 ;
    END
  END Data_PMOS_NOSF[918]
  PIN Data_PMOS_NOSF[913]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3914.745 187.44 3915.025 188.44 ;
    END
  END Data_PMOS_NOSF[913]
  PIN Data_PMOS_NOSF[907]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3914.185 187.44 3914.465 188.44 ;
    END
  END Data_PMOS_NOSF[907]
  PIN Data_PMOS_NOSF[919]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3913.625 187.44 3913.905 188.44 ;
    END
  END Data_PMOS_NOSF[919]
  PIN Data_PMOS_NOSF[914]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3913.065 187.44 3913.345 188.44 ;
    END
  END Data_PMOS_NOSF[914]
  PIN Data_PMOS_NOSF[904]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3912.505 187.44 3912.785 188.44 ;
    END
  END Data_PMOS_NOSF[904]
  PIN Data_PMOS_NOSF[903]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3911.945 187.44 3912.225 188.44 ;
    END
  END Data_PMOS_NOSF[903]
  PIN Data_PMOS_NOSF[920]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3911.385 187.44 3911.665 188.44 ;
    END
  END Data_PMOS_NOSF[920]
  PIN DIG_MON_PMOS_NOSF[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3908.585 187.44 3908.865 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[86]
  PIN DIG_MON_PMOS_NOSF[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3904.105 187.44 3904.385 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[85]
  PIN Data_PMOS_NOSF[900]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3862.105 187.44 3862.385 188.44 ;
    END
  END Data_PMOS_NOSF[900]
  PIN Data_PMOS_NOSF[890]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3861.545 187.44 3861.825 188.44 ;
    END
  END Data_PMOS_NOSF[890]
  PIN Data_PMOS_NOSF[894]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3860.985 187.44 3861.265 188.44 ;
    END
  END Data_PMOS_NOSF[894]
  PIN Data_PMOS_NOSF[901]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3860.425 187.44 3860.705 188.44 ;
    END
  END Data_PMOS_NOSF[901]
  PIN Data_PMOS_NOSF[887]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3859.865 187.44 3860.145 188.44 ;
    END
  END Data_PMOS_NOSF[887]
  PIN Data_PMOS_NOSF[895]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3859.305 187.44 3859.585 188.44 ;
    END
  END Data_PMOS_NOSF[895]
  PIN Data_PMOS_NOSF[902]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3858.745 187.44 3859.025 188.44 ;
    END
  END Data_PMOS_NOSF[902]
  PIN Data_PMOS_NOSF[896]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3858.185 187.44 3858.465 188.44 ;
    END
  END Data_PMOS_NOSF[896]
  PIN Data_PMOS_NOSF[889]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3857.625 187.44 3857.905 188.44 ;
    END
  END Data_PMOS_NOSF[889]
  PIN Data_PMOS_NOSF[888]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3857.065 187.44 3857.345 188.44 ;
    END
  END Data_PMOS_NOSF[888]
  PIN nTOK_PMOS_NOSF[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3854.825 187.44 3855.105 188.44 ;
    END
  END nTOK_PMOS_NOSF[42]
  PIN FREEZE_PMOS_NOSF[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3852.025 187.44 3852.305 188.44 ;
    END
  END FREEZE_PMOS_NOSF[42]
  PIN Read_PMOS_NOSF[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3851.465 187.44 3851.745 188.44 ;
    END
  END Read_PMOS_NOSF[42]
  PIN Data_PMOS_NOSF[885]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3839.145 187.44 3839.425 188.44 ;
    END
  END Data_PMOS_NOSF[885]
  PIN Data_PMOS_NOSF[884]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3838.585 187.44 3838.865 188.44 ;
    END
  END Data_PMOS_NOSF[884]
  PIN Data_PMOS_NOSF[897]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3837.465 187.44 3837.745 188.44 ;
    END
  END Data_PMOS_NOSF[897]
  PIN Data_PMOS_NOSF[891]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3838.025 187.44 3838.305 188.44 ;
    END
  END Data_PMOS_NOSF[891]
  PIN Data_PMOS_NOSF[892]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3836.905 187.44 3837.185 188.44 ;
    END
  END Data_PMOS_NOSF[892]
  PIN Data_PMOS_NOSF[886]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3836.345 187.44 3836.625 188.44 ;
    END
  END Data_PMOS_NOSF[886]
  PIN Data_PMOS_NOSF[898]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3835.785 187.44 3836.065 188.44 ;
    END
  END Data_PMOS_NOSF[898]
  PIN Data_PMOS_NOSF[893]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3835.225 187.44 3835.505 188.44 ;
    END
  END Data_PMOS_NOSF[893]
  PIN Data_PMOS_NOSF[883]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3834.665 187.44 3834.945 188.44 ;
    END
  END Data_PMOS_NOSF[883]
  PIN Data_PMOS_NOSF[882]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3834.105 187.44 3834.385 188.44 ;
    END
  END Data_PMOS_NOSF[882]
  PIN Data_PMOS_NOSF[899]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3833.545 187.44 3833.825 188.44 ;
    END
  END Data_PMOS_NOSF[899]
  PIN DIG_MON_PMOS_NOSF[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3828.785 187.44 3829.065 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[84]
  PIN FREEZE_PMOS_NOSF[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4081.625 187.44 4081.905 188.44 ;
    END
  END FREEZE_PMOS_NOSF[45]
  PIN DIG_MON_PMOS_NOSF[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4918.265 187.44 4918.545 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[111]
  PIN Data_PMOS_NOSF[1173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4916.025 187.44 4916.305 188.44 ;
    END
  END Data_PMOS_NOSF[1173]
  PIN Data_PMOS_NOSF[1163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4915.465 187.44 4915.745 188.44 ;
    END
  END Data_PMOS_NOSF[1163]
  PIN Data_PMOS_NOSF[1167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4914.905 187.44 4915.185 188.44 ;
    END
  END Data_PMOS_NOSF[1167]
  PIN Data_PMOS_NOSF[1174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4914.345 187.44 4914.625 188.44 ;
    END
  END Data_PMOS_NOSF[1174]
  PIN Data_PMOS_NOSF[1160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4913.785 187.44 4914.065 188.44 ;
    END
  END Data_PMOS_NOSF[1160]
  PIN Data_PMOS_NOSF[1168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4913.225 187.44 4913.505 188.44 ;
    END
  END Data_PMOS_NOSF[1168]
  PIN Data_PMOS_NOSF[1175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4912.665 187.44 4912.945 188.44 ;
    END
  END Data_PMOS_NOSF[1175]
  PIN Data_PMOS_NOSF[1169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4912.105 187.44 4912.385 188.44 ;
    END
  END Data_PMOS_NOSF[1169]
  PIN Data_PMOS_NOSF[1162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4911.545 187.44 4911.825 188.44 ;
    END
  END Data_PMOS_NOSF[1162]
  PIN Data_PMOS_NOSF[1161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4910.985 187.44 4911.265 188.44 ;
    END
  END Data_PMOS_NOSF[1161]
  PIN nTOK_PMOS_NOSF[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4908.745 187.44 4909.025 188.44 ;
    END
  END nTOK_PMOS_NOSF[55]
  PIN FREEZE_PMOS_NOSF[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4892.505 187.44 4892.785 188.44 ;
    END
  END FREEZE_PMOS_NOSF[55]
  PIN Read_PMOS_NOSF[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4891.945 187.44 4892.225 188.44 ;
    END
  END Read_PMOS_NOSF[55]
  PIN Data_PMOS_NOSF[1158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4888.025 187.44 4888.305 188.44 ;
    END
  END Data_PMOS_NOSF[1158]
  PIN Data_PMOS_NOSF[1157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4887.465 187.44 4887.745 188.44 ;
    END
  END Data_PMOS_NOSF[1157]
  PIN Data_PMOS_NOSF[1164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4886.905 187.44 4887.185 188.44 ;
    END
  END Data_PMOS_NOSF[1164]
  PIN Data_PMOS_NOSF[1170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4886.345 187.44 4886.625 188.44 ;
    END
  END Data_PMOS_NOSF[1170]
  PIN Data_PMOS_NOSF[1165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4885.785 187.44 4886.065 188.44 ;
    END
  END Data_PMOS_NOSF[1165]
  PIN Data_PMOS_NOSF[1159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4885.225 187.44 4885.505 188.44 ;
    END
  END Data_PMOS_NOSF[1159]
  PIN Data_PMOS_NOSF[1171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4884.665 187.44 4884.945 188.44 ;
    END
  END Data_PMOS_NOSF[1171]
  PIN Data_PMOS_NOSF[1166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4884.105 187.44 4884.385 188.44 ;
    END
  END Data_PMOS_NOSF[1166]
  PIN Data_PMOS_NOSF[1156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4883.545 187.44 4883.825 188.44 ;
    END
  END Data_PMOS_NOSF[1156]
  PIN Data_PMOS_NOSF[1155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4882.985 187.44 4883.265 188.44 ;
    END
  END Data_PMOS_NOSF[1155]
  PIN Data_PMOS_NOSF[1172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4882.425 187.44 4882.705 188.44 ;
    END
  END Data_PMOS_NOSF[1172]
  PIN DIG_MON_PMOS_NOSF[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4840.985 187.44 4841.265 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[110]
  PIN DIG_MON_PMOS_NOSF[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4836.505 187.44 4836.785 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[109]
  PIN Data_PMOS_NOSF[1152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4834.265 187.44 4834.545 188.44 ;
    END
  END Data_PMOS_NOSF[1152]
  PIN Data_PMOS_NOSF[1142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4833.705 187.44 4833.985 188.44 ;
    END
  END Data_PMOS_NOSF[1142]
  PIN Data_PMOS_NOSF[1146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4833.145 187.44 4833.425 188.44 ;
    END
  END Data_PMOS_NOSF[1146]
  PIN Data_PMOS_NOSF[1153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4832.585 187.44 4832.865 188.44 ;
    END
  END Data_PMOS_NOSF[1153]
  PIN Data_PMOS_NOSF[1139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4832.025 187.44 4832.305 188.44 ;
    END
  END Data_PMOS_NOSF[1139]
  PIN Data_PMOS_NOSF[1147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4831.465 187.44 4831.745 188.44 ;
    END
  END Data_PMOS_NOSF[1147]
  PIN Data_PMOS_NOSF[1154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4830.905 187.44 4831.185 188.44 ;
    END
  END Data_PMOS_NOSF[1154]
  PIN Data_PMOS_NOSF[1148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4830.345 187.44 4830.625 188.44 ;
    END
  END Data_PMOS_NOSF[1148]
  PIN Data_PMOS_NOSF[1141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4829.785 187.44 4830.065 188.44 ;
    END
  END Data_PMOS_NOSF[1141]
  PIN Data_PMOS_NOSF[1140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4820.825 187.44 4821.105 188.44 ;
    END
  END Data_PMOS_NOSF[1140]
  PIN nTOK_PMOS_NOSF[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4818.585 187.44 4818.865 188.44 ;
    END
  END nTOK_PMOS_NOSF[54]
  PIN FREEZE_PMOS_NOSF[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4815.785 187.44 4816.065 188.44 ;
    END
  END FREEZE_PMOS_NOSF[54]
  PIN Read_PMOS_NOSF[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4815.225 187.44 4815.505 188.44 ;
    END
  END Read_PMOS_NOSF[54]
  PIN Data_PMOS_NOSF[1137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4809.345 187.44 4809.625 188.44 ;
    END
  END Data_PMOS_NOSF[1137]
  PIN Data_PMOS_NOSF[1136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4808.785 187.44 4809.065 188.44 ;
    END
  END Data_PMOS_NOSF[1136]
  PIN Data_PMOS_NOSF[1143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4808.225 187.44 4808.505 188.44 ;
    END
  END Data_PMOS_NOSF[1143]
  PIN Data_PMOS_NOSF[1149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4807.665 187.44 4807.945 188.44 ;
    END
  END Data_PMOS_NOSF[1149]
  PIN Data_PMOS_NOSF[1144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4807.105 187.44 4807.385 188.44 ;
    END
  END Data_PMOS_NOSF[1144]
  PIN Data_PMOS_NOSF[1138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4781.065 187.44 4781.345 188.44 ;
    END
  END Data_PMOS_NOSF[1138]
  PIN Data_PMOS_NOSF[1150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4780.505 187.44 4780.785 188.44 ;
    END
  END Data_PMOS_NOSF[1150]
  PIN Data_PMOS_NOSF[1145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4779.945 187.44 4780.225 188.44 ;
    END
  END Data_PMOS_NOSF[1145]
  PIN Data_PMOS_NOSF[1135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4779.385 187.44 4779.665 188.44 ;
    END
  END Data_PMOS_NOSF[1135]
  PIN Data_PMOS_NOSF[1134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4778.825 187.44 4779.105 188.44 ;
    END
  END Data_PMOS_NOSF[1134]
  PIN Data_PMOS_NOSF[1151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4778.265 187.44 4778.545 188.44 ;
    END
  END Data_PMOS_NOSF[1151]
  PIN DIG_MON_PMOS_NOSF[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4775.465 187.44 4775.745 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[108]
  PIN DIG_MON_PMOS_NOSF[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4770.985 187.44 4771.265 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[107]
  PIN Data_PMOS_NOSF[1131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4768.745 187.44 4769.025 188.44 ;
    END
  END Data_PMOS_NOSF[1131]
  PIN Data_PMOS_NOSF[1121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4768.185 187.44 4768.465 188.44 ;
    END
  END Data_PMOS_NOSF[1121]
  PIN Data_PMOS_NOSF[1125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4754.745 187.44 4755.025 188.44 ;
    END
  END Data_PMOS_NOSF[1125]
  PIN Data_PMOS_NOSF[1132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4754.185 187.44 4754.465 188.44 ;
    END
  END Data_PMOS_NOSF[1132]
  PIN Data_PMOS_NOSF[1118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4753.625 187.44 4753.905 188.44 ;
    END
  END Data_PMOS_NOSF[1118]
  PIN Data_PMOS_NOSF[1126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4753.065 187.44 4753.345 188.44 ;
    END
  END Data_PMOS_NOSF[1126]
  PIN Data_PMOS_NOSF[1133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4752.505 187.44 4752.785 188.44 ;
    END
  END Data_PMOS_NOSF[1133]
  PIN Data_PMOS_NOSF[1127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4751.945 187.44 4752.225 188.44 ;
    END
  END Data_PMOS_NOSF[1127]
  PIN Data_PMOS_NOSF[1120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4751.385 187.44 4751.665 188.44 ;
    END
  END Data_PMOS_NOSF[1120]
  PIN Data_PMOS_NOSF[1119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4750.825 187.44 4751.105 188.44 ;
    END
  END Data_PMOS_NOSF[1119]
  PIN nTOK_PMOS_NOSF[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4748.585 187.44 4748.865 188.44 ;
    END
  END nTOK_PMOS_NOSF[53]
  PIN FREEZE_PMOS_NOSF[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4745.785 187.44 4746.065 188.44 ;
    END
  END FREEZE_PMOS_NOSF[53]
  PIN Read_PMOS_NOSF[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4745.225 187.44 4745.505 188.44 ;
    END
  END Read_PMOS_NOSF[53]
  PIN Data_PMOS_NOSF[1116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4702.665 187.44 4702.945 188.44 ;
    END
  END Data_PMOS_NOSF[1116]
  PIN Data_PMOS_NOSF[1115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4702.105 187.44 4702.385 188.44 ;
    END
  END Data_PMOS_NOSF[1115]
  PIN Data_PMOS_NOSF[1122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4701.545 187.44 4701.825 188.44 ;
    END
  END Data_PMOS_NOSF[1122]
  PIN Data_PMOS_NOSF[1128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4700.985 187.44 4701.265 188.44 ;
    END
  END Data_PMOS_NOSF[1128]
  PIN Data_PMOS_NOSF[1123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4700.425 187.44 4700.705 188.44 ;
    END
  END Data_PMOS_NOSF[1123]
  PIN Data_PMOS_NOSF[1117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4699.865 187.44 4700.145 188.44 ;
    END
  END Data_PMOS_NOSF[1117]
  PIN Data_PMOS_NOSF[1129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4699.305 187.44 4699.585 188.44 ;
    END
  END Data_PMOS_NOSF[1129]
  PIN Data_PMOS_NOSF[1124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4698.745 187.44 4699.025 188.44 ;
    END
  END Data_PMOS_NOSF[1124]
  PIN Data_PMOS_NOSF[1114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4698.185 187.44 4698.465 188.44 ;
    END
  END Data_PMOS_NOSF[1114]
  PIN Data_PMOS_NOSF[1113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4697.625 187.44 4697.905 188.44 ;
    END
  END Data_PMOS_NOSF[1113]
  PIN Data_PMOS_NOSF[1130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4697.065 187.44 4697.345 188.44 ;
    END
  END Data_PMOS_NOSF[1130]
  PIN DIG_MON_PMOS_NOSF[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4694.265 187.44 4694.545 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[106]
  PIN DIG_MON_PMOS_NOSF[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4689.785 187.44 4690.065 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[105]
  PIN Data_PMOS_NOSF[1110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4679.145 187.44 4679.425 188.44 ;
    END
  END Data_PMOS_NOSF[1110]
  PIN Data_PMOS_NOSF[1100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4678.585 187.44 4678.865 188.44 ;
    END
  END Data_PMOS_NOSF[1100]
  PIN Data_PMOS_NOSF[1104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4678.025 187.44 4678.305 188.44 ;
    END
  END Data_PMOS_NOSF[1104]
  PIN Data_PMOS_NOSF[1111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4677.465 187.44 4677.745 188.44 ;
    END
  END Data_PMOS_NOSF[1111]
  PIN Data_PMOS_NOSF[1097]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4676.905 187.44 4677.185 188.44 ;
    END
  END Data_PMOS_NOSF[1097]
  PIN Data_PMOS_NOSF[1105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4676.345 187.44 4676.625 188.44 ;
    END
  END Data_PMOS_NOSF[1105]
  PIN Data_PMOS_NOSF[1112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4675.785 187.44 4676.065 188.44 ;
    END
  END Data_PMOS_NOSF[1112]
  PIN Data_PMOS_NOSF[1106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4675.225 187.44 4675.505 188.44 ;
    END
  END Data_PMOS_NOSF[1106]
  PIN Data_PMOS_NOSF[1099]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4674.665 187.44 4674.945 188.44 ;
    END
  END Data_PMOS_NOSF[1099]
  PIN Data_PMOS_NOSF[1098]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4674.105 187.44 4674.385 188.44 ;
    END
  END Data_PMOS_NOSF[1098]
  PIN nTOK_PMOS_NOSF[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4669.905 187.44 4670.185 188.44 ;
    END
  END nTOK_PMOS_NOSF[52]
  PIN Read_PMOS_NOSF[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4641.065 187.44 4641.345 188.44 ;
    END
  END Read_PMOS_NOSF[52]
  PIN Data_PMOS_NOSF[1095]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4637.145 187.44 4637.425 188.44 ;
    END
  END Data_PMOS_NOSF[1095]
  PIN Data_PMOS_NOSF[1094]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4636.585 187.44 4636.865 188.44 ;
    END
  END Data_PMOS_NOSF[1094]
  PIN Data_PMOS_NOSF[1101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4636.025 187.44 4636.305 188.44 ;
    END
  END Data_PMOS_NOSF[1101]
  PIN Data_PMOS_NOSF[1107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4635.465 187.44 4635.745 188.44 ;
    END
  END Data_PMOS_NOSF[1107]
  PIN Data_PMOS_NOSF[1102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4634.905 187.44 4635.185 188.44 ;
    END
  END Data_PMOS_NOSF[1102]
  PIN Data_PMOS_NOSF[1096]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4634.345 187.44 4634.625 188.44 ;
    END
  END Data_PMOS_NOSF[1096]
  PIN Data_PMOS_NOSF[1108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4633.785 187.44 4634.065 188.44 ;
    END
  END Data_PMOS_NOSF[1108]
  PIN Data_PMOS_NOSF[1103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4633.225 187.44 4633.505 188.44 ;
    END
  END Data_PMOS_NOSF[1103]
  PIN Data_PMOS_NOSF[1093]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4632.665 187.44 4632.945 188.44 ;
    END
  END Data_PMOS_NOSF[1093]
  PIN Data_PMOS_NOSF[1092]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4632.105 187.44 4632.385 188.44 ;
    END
  END Data_PMOS_NOSF[1092]
  PIN Data_PMOS_NOSF[1109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4631.545 187.44 4631.825 188.44 ;
    END
  END Data_PMOS_NOSF[1109]
  PIN DIG_MON_PMOS_NOSF[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4628.745 187.44 4629.025 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[104]
  PIN DIG_MON_PMOS_NOSF[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4611.385 187.44 4611.665 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[103]
  PIN Data_PMOS_NOSF[1089]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4609.145 187.44 4609.425 188.44 ;
    END
  END Data_PMOS_NOSF[1089]
  PIN Data_PMOS_NOSF[1079]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4608.585 187.44 4608.865 188.44 ;
    END
  END Data_PMOS_NOSF[1079]
  PIN Data_PMOS_NOSF[1083]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4608.025 187.44 4608.305 188.44 ;
    END
  END Data_PMOS_NOSF[1083]
  PIN Data_PMOS_NOSF[1090]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4607.465 187.44 4607.745 188.44 ;
    END
  END Data_PMOS_NOSF[1090]
  PIN Data_PMOS_NOSF[1076]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4606.905 187.44 4607.185 188.44 ;
    END
  END Data_PMOS_NOSF[1076]
  PIN Data_PMOS_NOSF[1084]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4606.345 187.44 4606.625 188.44 ;
    END
  END Data_PMOS_NOSF[1084]
  PIN Data_PMOS_NOSF[1091]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4605.785 187.44 4606.065 188.44 ;
    END
  END Data_PMOS_NOSF[1091]
  PIN Data_PMOS_NOSF[1085]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4605.225 187.44 4605.505 188.44 ;
    END
  END Data_PMOS_NOSF[1085]
  PIN Data_PMOS_NOSF[1078]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4604.665 187.44 4604.945 188.44 ;
    END
  END Data_PMOS_NOSF[1078]
  PIN Data_PMOS_NOSF[1077]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4604.105 187.44 4604.385 188.44 ;
    END
  END Data_PMOS_NOSF[1077]
  PIN nTOK_PMOS_NOSF[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4562.665 187.44 4562.945 188.44 ;
    END
  END nTOK_PMOS_NOSF[51]
  PIN FREEZE_PMOS_NOSF[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4559.865 187.44 4560.145 188.44 ;
    END
  END FREEZE_PMOS_NOSF[51]
  PIN Read_PMOS_NOSF[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4559.305 187.44 4559.585 188.44 ;
    END
  END Read_PMOS_NOSF[51]
  PIN Data_PMOS_NOSF[1074]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4555.385 187.44 4555.665 188.44 ;
    END
  END Data_PMOS_NOSF[1074]
  PIN Data_PMOS_NOSF[1073]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4554.825 187.44 4555.105 188.44 ;
    END
  END Data_PMOS_NOSF[1073]
  PIN Data_PMOS_NOSF[1080]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4554.265 187.44 4554.545 188.44 ;
    END
  END Data_PMOS_NOSF[1080]
  PIN Data_PMOS_NOSF[1086]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4553.705 187.44 4553.985 188.44 ;
    END
  END Data_PMOS_NOSF[1086]
  PIN Data_PMOS_NOSF[1081]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4553.145 187.44 4553.425 188.44 ;
    END
  END Data_PMOS_NOSF[1081]
  PIN Data_PMOS_NOSF[1075]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4552.585 187.44 4552.865 188.44 ;
    END
  END Data_PMOS_NOSF[1075]
  PIN Data_PMOS_NOSF[1087]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4552.025 187.44 4552.305 188.44 ;
    END
  END Data_PMOS_NOSF[1087]
  PIN Data_PMOS_NOSF[1082]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4551.465 187.44 4551.745 188.44 ;
    END
  END Data_PMOS_NOSF[1082]
  PIN Data_PMOS_NOSF[1072]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4550.905 187.44 4551.185 188.44 ;
    END
  END Data_PMOS_NOSF[1072]
  PIN Data_PMOS_NOSF[1071]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4550.345 187.44 4550.625 188.44 ;
    END
  END Data_PMOS_NOSF[1071]
  PIN Data_PMOS_NOSF[1088]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4549.785 187.44 4550.065 188.44 ;
    END
  END Data_PMOS_NOSF[1088]
  PIN DIG_MON_PMOS_NOSF[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4538.585 187.44 4538.865 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[102]
  PIN DIG_MON_PMOS_NOSF[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4534.105 187.44 4534.385 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[101]
  PIN Data_PMOS_NOSF[1068]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4529.905 187.44 4530.185 188.44 ;
    END
  END Data_PMOS_NOSF[1068]
  PIN Data_PMOS_NOSF[1058]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4529.345 187.44 4529.625 188.44 ;
    END
  END Data_PMOS_NOSF[1058]
  PIN Data_PMOS_NOSF[1062]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4528.785 187.44 4529.065 188.44 ;
    END
  END Data_PMOS_NOSF[1062]
  PIN Data_PMOS_NOSF[1069]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4528.225 187.44 4528.505 188.44 ;
    END
  END Data_PMOS_NOSF[1069]
  PIN Data_PMOS_NOSF[1055]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4527.665 187.44 4527.945 188.44 ;
    END
  END Data_PMOS_NOSF[1055]
  PIN Data_PMOS_NOSF[1063]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4501.625 187.44 4501.905 188.44 ;
    END
  END Data_PMOS_NOSF[1063]
  PIN Data_PMOS_NOSF[1070]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4501.065 187.44 4501.345 188.44 ;
    END
  END Data_PMOS_NOSF[1070]
  PIN Data_PMOS_NOSF[1064]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4500.505 187.44 4500.785 188.44 ;
    END
  END Data_PMOS_NOSF[1064]
  PIN Data_PMOS_NOSF[1057]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4499.945 187.44 4500.225 188.44 ;
    END
  END Data_PMOS_NOSF[1057]
  PIN Data_PMOS_NOSF[1056]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4499.385 187.44 4499.665 188.44 ;
    END
  END Data_PMOS_NOSF[1056]
  PIN nTOK_PMOS_NOSF[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4497.145 187.44 4497.425 188.44 ;
    END
  END nTOK_PMOS_NOSF[50]
  PIN FREEZE_PMOS_NOSF[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4494.345 187.44 4494.625 188.44 ;
    END
  END FREEZE_PMOS_NOSF[50]
  PIN Read_PMOS_NOSF[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4493.785 187.44 4494.065 188.44 ;
    END
  END Read_PMOS_NOSF[50]
  PIN Data_PMOS_NOSF[1053]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4489.865 187.44 4490.145 188.44 ;
    END
  END Data_PMOS_NOSF[1053]
  PIN Data_PMOS_NOSF[1052]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4489.305 187.44 4489.585 188.44 ;
    END
  END Data_PMOS_NOSF[1052]
  PIN Data_PMOS_NOSF[1059]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4488.745 187.44 4489.025 188.44 ;
    END
  END Data_PMOS_NOSF[1059]
  PIN Data_PMOS_NOSF[1065]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4475.305 187.44 4475.585 188.44 ;
    END
  END Data_PMOS_NOSF[1065]
  PIN Data_PMOS_NOSF[1060]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4474.745 187.44 4475.025 188.44 ;
    END
  END Data_PMOS_NOSF[1060]
  PIN Data_PMOS_NOSF[1054]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4474.185 187.44 4474.465 188.44 ;
    END
  END Data_PMOS_NOSF[1054]
  PIN Data_PMOS_NOSF[1066]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4473.625 187.44 4473.905 188.44 ;
    END
  END Data_PMOS_NOSF[1066]
  PIN Data_PMOS_NOSF[1061]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4473.065 187.44 4473.345 188.44 ;
    END
  END Data_PMOS_NOSF[1061]
  PIN Data_PMOS_NOSF[1051]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4472.505 187.44 4472.785 188.44 ;
    END
  END Data_PMOS_NOSF[1051]
  PIN Data_PMOS_NOSF[1050]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4471.945 187.44 4472.225 188.44 ;
    END
  END Data_PMOS_NOSF[1050]
  PIN Data_PMOS_NOSF[1067]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4471.385 187.44 4471.665 188.44 ;
    END
  END Data_PMOS_NOSF[1067]
  PIN DIG_MON_PMOS_NOSF[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4468.585 187.44 4468.865 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[100]
  PIN DIG_MON_PMOS_NOSF[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4464.105 187.44 4464.385 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[99]
  PIN Data_PMOS_NOSF[1047]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4422.105 187.44 4422.385 188.44 ;
    END
  END Data_PMOS_NOSF[1047]
  PIN Data_PMOS_NOSF[1037]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4421.545 187.44 4421.825 188.44 ;
    END
  END Data_PMOS_NOSF[1037]
  PIN Data_PMOS_NOSF[1041]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4420.985 187.44 4421.265 188.44 ;
    END
  END Data_PMOS_NOSF[1041]
  PIN Data_PMOS_NOSF[1048]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4420.425 187.44 4420.705 188.44 ;
    END
  END Data_PMOS_NOSF[1048]
  PIN Data_PMOS_NOSF[1034]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4419.865 187.44 4420.145 188.44 ;
    END
  END Data_PMOS_NOSF[1034]
  PIN Data_PMOS_NOSF[1042]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4419.305 187.44 4419.585 188.44 ;
    END
  END Data_PMOS_NOSF[1042]
  PIN Data_PMOS_NOSF[1049]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4418.745 187.44 4419.025 188.44 ;
    END
  END Data_PMOS_NOSF[1049]
  PIN Data_PMOS_NOSF[1043]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4418.185 187.44 4418.465 188.44 ;
    END
  END Data_PMOS_NOSF[1043]
  PIN Data_PMOS_NOSF[1036]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4417.625 187.44 4417.905 188.44 ;
    END
  END Data_PMOS_NOSF[1036]
  PIN Data_PMOS_NOSF[1035]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4417.065 187.44 4417.345 188.44 ;
    END
  END Data_PMOS_NOSF[1035]
  PIN nTOK_PMOS_NOSF[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4414.825 187.44 4415.105 188.44 ;
    END
  END nTOK_PMOS_NOSF[49]
  PIN FREEZE_PMOS_NOSF[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4412.025 187.44 4412.305 188.44 ;
    END
  END FREEZE_PMOS_NOSF[49]
  PIN Read_PMOS_NOSF[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4411.465 187.44 4411.745 188.44 ;
    END
  END Read_PMOS_NOSF[49]
  PIN Data_PMOS_NOSF[1032]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4399.145 187.44 4399.425 188.44 ;
    END
  END Data_PMOS_NOSF[1032]
  PIN Data_PMOS_NOSF[1031]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4398.585 187.44 4398.865 188.44 ;
    END
  END Data_PMOS_NOSF[1031]
  PIN Data_PMOS_NOSF[1044]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4397.465 187.44 4397.745 188.44 ;
    END
  END Data_PMOS_NOSF[1044]
  PIN Data_PMOS_NOSF[1038]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4398.025 187.44 4398.305 188.44 ;
    END
  END Data_PMOS_NOSF[1038]
  PIN Data_PMOS_NOSF[1039]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4396.905 187.44 4397.185 188.44 ;
    END
  END Data_PMOS_NOSF[1039]
  PIN Data_PMOS_NOSF[1033]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4396.345 187.44 4396.625 188.44 ;
    END
  END Data_PMOS_NOSF[1033]
  PIN Data_PMOS_NOSF[1045]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4395.785 187.44 4396.065 188.44 ;
    END
  END Data_PMOS_NOSF[1045]
  PIN Data_PMOS_NOSF[1040]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4395.225 187.44 4395.505 188.44 ;
    END
  END Data_PMOS_NOSF[1040]
  PIN Data_PMOS_NOSF[1030]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4394.665 187.44 4394.945 188.44 ;
    END
  END Data_PMOS_NOSF[1030]
  PIN Data_PMOS_NOSF[1029]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4394.105 187.44 4394.385 188.44 ;
    END
  END Data_PMOS_NOSF[1029]
  PIN Data_PMOS_NOSF[1046]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4393.545 187.44 4393.825 188.44 ;
    END
  END Data_PMOS_NOSF[1046]
  PIN DIG_MON_PMOS_NOSF[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4388.785 187.44 4389.065 188.44 ;
    END
  END DIG_MON_PMOS_NOSF[98]
  PIN FREEZE_PMOS_NOSF[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4641.625 187.44 4641.905 188.44 ;
    END
  END FREEZE_PMOS_NOSF[52]
  OBS
    LAYER M1 SPACING 0.23 ;
      RECT 326.66 187.44 18490.46 8613.565 ;
    LAYER M2 ;
      RECT 9429.265 189.04 9431.205 189.225 ;
      RECT 9431.115 188.945 9431.205 189.225 ;
      RECT 9429.265 188.945 9429.355 189.225 ;
      RECT 18484.435 189.04 18484.715 252.385 ;
      RECT 18483.875 189.04 18484.155 252.385 ;
      RECT 18483.315 189.04 18483.595 252.385 ;
      RECT 18482.755 189.04 18483.035 252.385 ;
      RECT 18482.195 189.04 18482.475 252.385 ;
      RECT 18481.635 189.04 18481.915 252.385 ;
      RECT 18481.075 189.04 18481.355 252.385 ;
      RECT 18480.515 189.04 18480.795 252.385 ;
      RECT 18356.515 189.04 18356.795 190.305 ;
      RECT 18352.875 189.04 18353.155 190.27 ;
      RECT 18349.235 189.04 18349.515 190.325 ;
      RECT 18345.595 189.04 18345.875 190.365 ;
      RECT 18341.955 189.04 18342.235 190.35 ;
      RECT 18338.315 189.04 18338.595 190.26 ;
      RECT 18279.235 189.04 18279.515 190.16 ;
      RECT 18275.315 189.04 18275.595 190.205 ;
      RECT 18271.395 189.04 18271.675 189.935 ;
      RECT 18267.475 189.04 18267.755 190.16 ;
      RECT 18263.555 189.04 18263.835 205.605 ;
      RECT 18216.515 189.04 18216.795 190.305 ;
      RECT 18212.875 189.04 18213.155 190.27 ;
      RECT 18209.235 189.04 18209.515 190.325 ;
      RECT 18205.595 189.04 18205.875 190.365 ;
      RECT 18201.955 189.04 18202.235 190.35 ;
      RECT 18198.315 189.04 18198.595 190.26 ;
      RECT 18139.235 189.04 18139.515 190.16 ;
      RECT 18135.315 189.04 18135.595 190.205 ;
      RECT 18131.395 189.04 18131.675 189.935 ;
      RECT 18127.475 189.04 18127.755 190.16 ;
      RECT 18123.555 189.04 18123.835 205.605 ;
      RECT 18076.515 189.04 18076.795 190.305 ;
      RECT 18072.875 189.04 18073.155 190.27 ;
      RECT 18069.235 189.04 18069.515 190.325 ;
      RECT 18065.595 189.04 18065.875 190.365 ;
      RECT 18061.955 189.04 18062.235 190.35 ;
      RECT 18058.315 189.04 18058.595 190.26 ;
      RECT 17999.235 189.04 17999.515 190.16 ;
      RECT 17995.315 189.04 17995.595 190.205 ;
      RECT 17991.395 189.04 17991.675 189.935 ;
      RECT 17987.475 189.04 17987.755 190.16 ;
      RECT 17983.555 189.04 17983.835 205.605 ;
      RECT 17936.515 189.04 17936.795 190.305 ;
      RECT 17932.875 189.04 17933.155 190.27 ;
      RECT 17929.235 189.04 17929.515 190.325 ;
      RECT 17925.595 189.04 17925.875 190.365 ;
      RECT 17921.955 189.04 17922.235 190.35 ;
      RECT 17918.315 189.04 17918.595 190.26 ;
      RECT 17859.235 189.04 17859.515 190.16 ;
      RECT 17855.315 189.04 17855.595 190.205 ;
      RECT 17851.395 189.04 17851.675 189.935 ;
      RECT 17847.475 189.04 17847.755 190.16 ;
      RECT 17843.555 189.04 17843.835 205.605 ;
      RECT 17796.515 189.04 17796.795 190.305 ;
      RECT 17792.875 189.04 17793.155 190.27 ;
      RECT 17789.235 189.04 17789.515 190.325 ;
      RECT 17785.595 189.04 17785.875 190.365 ;
      RECT 17781.955 189.04 17782.235 190.35 ;
      RECT 17778.315 189.04 17778.595 190.26 ;
      RECT 17719.235 189.04 17719.515 190.16 ;
      RECT 17715.315 189.04 17715.595 190.205 ;
      RECT 17711.395 189.04 17711.675 189.935 ;
      RECT 17707.475 189.04 17707.755 190.16 ;
      RECT 17703.555 189.04 17703.835 205.605 ;
      RECT 17656.515 189.04 17656.795 190.305 ;
      RECT 17652.875 189.04 17653.155 190.27 ;
      RECT 17649.235 189.04 17649.515 190.325 ;
      RECT 17645.595 189.04 17645.875 190.365 ;
      RECT 17641.955 189.04 17642.235 190.35 ;
      RECT 17638.315 189.04 17638.595 190.26 ;
      RECT 17579.235 189.04 17579.515 190.16 ;
      RECT 17575.315 189.04 17575.595 190.205 ;
      RECT 17571.395 189.04 17571.675 189.935 ;
      RECT 17567.475 189.04 17567.755 190.16 ;
      RECT 17563.555 189.04 17563.835 205.605 ;
      RECT 17516.515 189.04 17516.795 190.305 ;
      RECT 17512.875 189.04 17513.155 190.27 ;
      RECT 17509.235 189.04 17509.515 190.325 ;
      RECT 17505.595 189.04 17505.875 190.365 ;
      RECT 17501.955 189.04 17502.235 190.35 ;
      RECT 17498.315 189.04 17498.595 190.26 ;
      RECT 17439.235 189.04 17439.515 190.16 ;
      RECT 17435.315 189.04 17435.595 190.205 ;
      RECT 17431.395 189.04 17431.675 189.935 ;
      RECT 17427.475 189.04 17427.755 190.16 ;
      RECT 17423.555 189.04 17423.835 205.605 ;
      RECT 17376.515 189.04 17376.795 190.305 ;
      RECT 17372.875 189.04 17373.155 190.27 ;
      RECT 17369.235 189.04 17369.515 190.325 ;
      RECT 17365.595 189.04 17365.875 190.365 ;
      RECT 17361.955 189.04 17362.235 190.35 ;
      RECT 17358.315 189.04 17358.595 190.26 ;
      RECT 17299.235 189.04 17299.515 190.16 ;
      RECT 17295.315 189.04 17295.595 190.205 ;
      RECT 17291.395 189.04 17291.675 189.935 ;
      RECT 17287.475 189.04 17287.755 190.16 ;
      RECT 17283.555 189.04 17283.835 205.605 ;
      RECT 17236.515 189.04 17236.795 190.305 ;
      RECT 17232.875 189.04 17233.155 190.27 ;
      RECT 17229.235 189.04 17229.515 190.325 ;
      RECT 17225.595 189.04 17225.875 190.365 ;
      RECT 17221.955 189.04 17222.235 190.35 ;
      RECT 17218.315 189.04 17218.595 190.26 ;
      RECT 17159.235 189.04 17159.515 190.16 ;
      RECT 17155.315 189.04 17155.595 190.205 ;
      RECT 17151.395 189.04 17151.675 189.935 ;
      RECT 17147.475 189.04 17147.755 190.16 ;
      RECT 17143.555 189.04 17143.835 205.605 ;
      RECT 17096.515 189.04 17096.795 190.305 ;
      RECT 17092.875 189.04 17093.155 190.27 ;
      RECT 17089.235 189.04 17089.515 190.325 ;
      RECT 17085.595 189.04 17085.875 190.365 ;
      RECT 17081.955 189.04 17082.235 190.35 ;
      RECT 17078.315 189.04 17078.595 190.26 ;
      RECT 17019.235 189.04 17019.515 190.16 ;
      RECT 17015.315 189.04 17015.595 190.205 ;
      RECT 17011.395 189.04 17011.675 189.935 ;
      RECT 17007.475 189.04 17007.755 190.16 ;
      RECT 17003.555 189.04 17003.835 205.605 ;
      RECT 16956.515 189.04 16956.795 190.305 ;
      RECT 16952.875 189.04 16953.155 190.27 ;
      RECT 16949.235 189.04 16949.515 190.325 ;
      RECT 16945.595 189.04 16945.875 190.365 ;
      RECT 16941.955 189.04 16942.235 190.35 ;
      RECT 16938.315 189.04 16938.595 190.26 ;
      RECT 16879.235 189.04 16879.515 190.16 ;
      RECT 16875.315 189.04 16875.595 190.205 ;
      RECT 16871.395 189.04 16871.675 189.935 ;
      RECT 16867.475 189.04 16867.755 190.16 ;
      RECT 16863.555 189.04 16863.835 205.605 ;
      RECT 16816.515 189.04 16816.795 190.305 ;
      RECT 16812.875 189.04 16813.155 190.27 ;
      RECT 16809.235 189.04 16809.515 190.325 ;
      RECT 16805.595 189.04 16805.875 190.365 ;
      RECT 16801.955 189.04 16802.235 190.35 ;
      RECT 16798.315 189.04 16798.595 190.26 ;
      RECT 16739.235 189.04 16739.515 190.16 ;
      RECT 16735.315 189.04 16735.595 190.205 ;
      RECT 16731.395 189.04 16731.675 189.935 ;
      RECT 16727.475 189.04 16727.755 190.16 ;
      RECT 16723.555 189.04 16723.835 205.605 ;
      RECT 16676.515 189.04 16676.795 190.305 ;
      RECT 16672.875 189.04 16673.155 190.27 ;
      RECT 16669.235 189.04 16669.515 190.325 ;
      RECT 16665.595 189.04 16665.875 190.365 ;
      RECT 16661.955 189.04 16662.235 190.35 ;
      RECT 16658.315 189.04 16658.595 190.26 ;
      RECT 16599.235 189.04 16599.515 190.16 ;
      RECT 16595.315 189.04 16595.595 190.205 ;
      RECT 16591.395 189.04 16591.675 189.935 ;
      RECT 16587.475 189.04 16587.755 190.16 ;
      RECT 16583.555 189.04 16583.835 205.605 ;
      RECT 16536.515 189.04 16536.795 190.305 ;
      RECT 16532.875 189.04 16533.155 190.27 ;
      RECT 16529.235 189.04 16529.515 190.325 ;
      RECT 16525.595 189.04 16525.875 190.365 ;
      RECT 16521.955 189.04 16522.235 190.35 ;
      RECT 16518.315 189.04 16518.595 190.26 ;
      RECT 16459.235 189.04 16459.515 190.16 ;
      RECT 16455.315 189.04 16455.595 190.205 ;
      RECT 16451.395 189.04 16451.675 189.935 ;
      RECT 16447.475 189.04 16447.755 190.16 ;
      RECT 16443.555 189.04 16443.835 205.605 ;
      RECT 16396.515 189.04 16396.795 190.305 ;
      RECT 16392.875 189.04 16393.155 190.27 ;
      RECT 16389.235 189.04 16389.515 190.325 ;
      RECT 16385.595 189.04 16385.875 190.365 ;
      RECT 16381.955 189.04 16382.235 190.35 ;
      RECT 16378.315 189.04 16378.595 190.26 ;
      RECT 16319.235 189.04 16319.515 190.16 ;
      RECT 16315.315 189.04 16315.595 190.205 ;
      RECT 16311.395 189.04 16311.675 189.935 ;
      RECT 16307.475 189.04 16307.755 190.16 ;
      RECT 16303.555 189.04 16303.835 205.605 ;
      RECT 16256.515 189.04 16256.795 190.305 ;
      RECT 16252.875 189.04 16253.155 190.27 ;
      RECT 16249.235 189.04 16249.515 190.325 ;
      RECT 16245.595 189.04 16245.875 190.365 ;
      RECT 16241.955 189.04 16242.235 190.35 ;
      RECT 16238.315 189.04 16238.595 190.26 ;
      RECT 16179.235 189.04 16179.515 190.16 ;
      RECT 16175.315 189.04 16175.595 190.205 ;
      RECT 16171.395 189.04 16171.675 189.935 ;
      RECT 16167.475 189.04 16167.755 190.16 ;
      RECT 16163.555 189.04 16163.835 205.605 ;
      RECT 16116.515 189.04 16116.795 190.305 ;
      RECT 16112.875 189.04 16113.155 190.27 ;
      RECT 16109.235 189.04 16109.515 190.325 ;
      RECT 16105.595 189.04 16105.875 190.365 ;
      RECT 16101.955 189.04 16102.235 190.35 ;
      RECT 16098.315 189.04 16098.595 190.26 ;
      RECT 16039.235 189.04 16039.515 190.16 ;
      RECT 16035.315 189.04 16035.595 190.205 ;
      RECT 16031.395 189.04 16031.675 189.935 ;
      RECT 16027.475 189.04 16027.755 190.16 ;
      RECT 16023.555 189.04 16023.835 205.605 ;
      RECT 15976.515 189.04 15976.795 190.305 ;
      RECT 15972.875 189.04 15973.155 190.27 ;
      RECT 15969.235 189.04 15969.515 190.325 ;
      RECT 15965.595 189.04 15965.875 190.365 ;
      RECT 15961.955 189.04 15962.235 190.35 ;
      RECT 15958.315 189.04 15958.595 190.26 ;
      RECT 15899.235 189.04 15899.515 190.16 ;
      RECT 15895.315 189.04 15895.595 190.205 ;
      RECT 15891.395 189.04 15891.675 189.935 ;
      RECT 15887.475 189.04 15887.755 190.16 ;
      RECT 15883.555 189.04 15883.835 205.605 ;
      RECT 15836.515 189.04 15836.795 190.305 ;
      RECT 15832.875 189.04 15833.155 190.27 ;
      RECT 15829.235 189.04 15829.515 190.325 ;
      RECT 15825.595 189.04 15825.875 190.365 ;
      RECT 15821.955 189.04 15822.235 190.35 ;
      RECT 15818.315 189.04 15818.595 190.26 ;
      RECT 15759.235 189.04 15759.515 190.16 ;
      RECT 15755.315 189.04 15755.595 190.205 ;
      RECT 15751.395 189.04 15751.675 189.935 ;
      RECT 15747.475 189.04 15747.755 190.16 ;
      RECT 15743.555 189.04 15743.835 205.605 ;
      RECT 15696.515 189.04 15696.795 190.305 ;
      RECT 15692.875 189.04 15693.155 190.27 ;
      RECT 15689.235 189.04 15689.515 190.325 ;
      RECT 15685.595 189.04 15685.875 190.365 ;
      RECT 15681.955 189.04 15682.235 190.35 ;
      RECT 15678.315 189.04 15678.595 190.26 ;
      RECT 15619.235 189.04 15619.515 190.16 ;
      RECT 15615.315 189.04 15615.595 190.205 ;
      RECT 15611.395 189.04 15611.675 189.935 ;
      RECT 15607.475 189.04 15607.755 190.16 ;
      RECT 15603.555 189.04 15603.835 205.605 ;
      RECT 15556.515 189.04 15556.795 190.305 ;
      RECT 15552.875 189.04 15553.155 190.27 ;
      RECT 15549.235 189.04 15549.515 190.325 ;
      RECT 15545.595 189.04 15545.875 190.365 ;
      RECT 15541.955 189.04 15542.235 190.35 ;
      RECT 15538.315 189.04 15538.595 190.26 ;
      RECT 15479.235 189.04 15479.515 190.16 ;
      RECT 15475.315 189.04 15475.595 190.205 ;
      RECT 15471.395 189.04 15471.675 189.935 ;
      RECT 15467.475 189.04 15467.755 190.16 ;
      RECT 15463.555 189.04 15463.835 205.605 ;
      RECT 15416.515 189.04 15416.795 190.305 ;
      RECT 15412.875 189.04 15413.155 190.27 ;
      RECT 15409.235 189.04 15409.515 190.325 ;
      RECT 15405.595 189.04 15405.875 190.365 ;
      RECT 15401.955 189.04 15402.235 190.35 ;
      RECT 15398.315 189.04 15398.595 190.26 ;
      RECT 15339.235 189.04 15339.515 190.16 ;
      RECT 15335.315 189.04 15335.595 190.205 ;
      RECT 15331.395 189.04 15331.675 189.935 ;
      RECT 15327.475 189.04 15327.755 190.16 ;
      RECT 15323.555 189.04 15323.835 205.605 ;
      RECT 15276.515 189.04 15276.795 190.305 ;
      RECT 15272.875 189.04 15273.155 190.27 ;
      RECT 15269.235 189.04 15269.515 190.325 ;
      RECT 15265.595 189.04 15265.875 190.365 ;
      RECT 15261.955 189.04 15262.235 190.35 ;
      RECT 15258.315 189.04 15258.595 190.26 ;
      RECT 15199.235 189.04 15199.515 190.16 ;
      RECT 15195.315 189.04 15195.595 190.205 ;
      RECT 15191.395 189.04 15191.675 189.935 ;
      RECT 15187.475 189.04 15187.755 190.16 ;
      RECT 15183.555 189.04 15183.835 205.605 ;
      RECT 15136.515 189.04 15136.795 190.305 ;
      RECT 15132.875 189.04 15133.155 190.27 ;
      RECT 15129.235 189.04 15129.515 190.325 ;
      RECT 15125.595 189.04 15125.875 190.365 ;
      RECT 15121.955 189.04 15122.235 190.35 ;
      RECT 15118.315 189.04 15118.595 190.26 ;
      RECT 15059.235 189.04 15059.515 190.16 ;
      RECT 15055.315 189.04 15055.595 190.205 ;
      RECT 15051.395 189.04 15051.675 189.935 ;
      RECT 15047.475 189.04 15047.755 190.16 ;
      RECT 15043.555 189.04 15043.835 205.605 ;
      RECT 14996.515 189.04 14996.795 190.305 ;
      RECT 14992.875 189.04 14993.155 190.27 ;
      RECT 14989.235 189.04 14989.515 190.325 ;
      RECT 14985.595 189.04 14985.875 190.365 ;
      RECT 14981.955 189.04 14982.235 190.35 ;
      RECT 14978.315 189.04 14978.595 190.26 ;
      RECT 14919.235 189.04 14919.515 190.16 ;
      RECT 14915.315 189.04 14915.595 190.205 ;
      RECT 14911.395 189.04 14911.675 189.935 ;
      RECT 14907.475 189.04 14907.755 190.16 ;
      RECT 14903.555 189.04 14903.835 205.605 ;
      RECT 14856.515 189.04 14856.795 190.305 ;
      RECT 14852.875 189.04 14853.155 190.27 ;
      RECT 14849.235 189.04 14849.515 190.325 ;
      RECT 14845.595 189.04 14845.875 190.365 ;
      RECT 14841.955 189.04 14842.235 190.35 ;
      RECT 14838.315 189.04 14838.595 190.26 ;
      RECT 14779.235 189.04 14779.515 190.16 ;
      RECT 14775.315 189.04 14775.595 190.205 ;
      RECT 14771.395 189.04 14771.675 189.935 ;
      RECT 14767.475 189.04 14767.755 190.16 ;
      RECT 14763.555 189.04 14763.835 205.605 ;
      RECT 14716.515 189.04 14716.795 190.305 ;
      RECT 14712.875 189.04 14713.155 190.27 ;
      RECT 14709.235 189.04 14709.515 190.325 ;
      RECT 14705.595 189.04 14705.875 190.365 ;
      RECT 14701.955 189.04 14702.235 190.35 ;
      RECT 14698.315 189.04 14698.595 190.26 ;
      RECT 14639.235 189.04 14639.515 190.16 ;
      RECT 14635.315 189.04 14635.595 190.205 ;
      RECT 14631.395 189.04 14631.675 189.935 ;
      RECT 14627.475 189.04 14627.755 190.16 ;
      RECT 14623.555 189.04 14623.835 205.605 ;
      RECT 14576.515 189.04 14576.795 190.305 ;
      RECT 14572.875 189.04 14573.155 190.27 ;
      RECT 14569.235 189.04 14569.515 190.325 ;
      RECT 14565.595 189.04 14565.875 190.365 ;
      RECT 14561.955 189.04 14562.235 190.35 ;
      RECT 14558.315 189.04 14558.595 190.26 ;
      RECT 14499.235 189.04 14499.515 190.16 ;
      RECT 14495.315 189.04 14495.595 190.205 ;
      RECT 14491.395 189.04 14491.675 189.935 ;
      RECT 14487.475 189.04 14487.755 190.16 ;
      RECT 14483.555 189.04 14483.835 205.605 ;
      RECT 14436.515 189.04 14436.795 190.305 ;
      RECT 14432.875 189.04 14433.155 190.27 ;
      RECT 14429.235 189.04 14429.515 190.325 ;
      RECT 14425.595 189.04 14425.875 190.365 ;
      RECT 14421.955 189.04 14422.235 190.35 ;
      RECT 14418.315 189.04 14418.595 190.26 ;
      RECT 14359.235 189.04 14359.515 190.16 ;
      RECT 14355.315 189.04 14355.595 190.205 ;
      RECT 14351.395 189.04 14351.675 189.935 ;
      RECT 14347.475 189.04 14347.755 190.16 ;
      RECT 14343.555 189.04 14343.835 205.605 ;
      RECT 14296.515 189.04 14296.795 190.305 ;
      RECT 14292.875 189.04 14293.155 190.27 ;
      RECT 14289.235 189.04 14289.515 190.325 ;
      RECT 14285.595 189.04 14285.875 190.365 ;
      RECT 14281.955 189.04 14282.235 190.35 ;
      RECT 14278.315 189.04 14278.595 190.26 ;
      RECT 14219.235 189.04 14219.515 190.16 ;
      RECT 14215.315 189.04 14215.595 190.205 ;
      RECT 14211.395 189.04 14211.675 189.935 ;
      RECT 14207.475 189.04 14207.755 190.16 ;
      RECT 14203.555 189.04 14203.835 205.605 ;
      RECT 14156.515 189.04 14156.795 190.305 ;
      RECT 14152.875 189.04 14153.155 190.27 ;
      RECT 14149.235 189.04 14149.515 190.325 ;
      RECT 14145.595 189.04 14145.875 190.365 ;
      RECT 14141.955 189.04 14142.235 190.35 ;
      RECT 14138.315 189.04 14138.595 190.26 ;
      RECT 14079.235 189.04 14079.515 190.16 ;
      RECT 14075.315 189.04 14075.595 190.205 ;
      RECT 14071.395 189.04 14071.675 189.935 ;
      RECT 14067.475 189.04 14067.755 190.16 ;
      RECT 14063.555 189.04 14063.835 205.605 ;
      RECT 14016.515 189.04 14016.795 190.305 ;
      RECT 14012.875 189.04 14013.155 190.27 ;
      RECT 14009.235 189.04 14009.515 190.325 ;
      RECT 14005.595 189.04 14005.875 190.365 ;
      RECT 14001.955 189.04 14002.235 190.35 ;
      RECT 13998.315 189.04 13998.595 190.26 ;
      RECT 13939.235 189.04 13939.515 190.16 ;
      RECT 13935.315 189.04 13935.595 190.205 ;
      RECT 13931.395 189.04 13931.675 189.935 ;
      RECT 13927.475 189.04 13927.755 190.16 ;
      RECT 13923.555 189.04 13923.835 205.605 ;
      RECT 13876.515 189.04 13876.795 190.305 ;
      RECT 13872.875 189.04 13873.155 190.27 ;
      RECT 13869.235 189.04 13869.515 190.325 ;
      RECT 13865.595 189.04 13865.875 190.365 ;
      RECT 13861.955 189.04 13862.235 190.35 ;
      RECT 13858.315 189.04 13858.595 190.26 ;
      RECT 13799.235 189.04 13799.515 190.16 ;
      RECT 13795.315 189.04 13795.595 190.205 ;
      RECT 13791.395 189.04 13791.675 189.935 ;
      RECT 13787.475 189.04 13787.755 190.16 ;
      RECT 13783.555 189.04 13783.835 205.605 ;
      RECT 13736.515 189.04 13736.795 190.305 ;
      RECT 13732.875 189.04 13733.155 190.27 ;
      RECT 13729.235 189.04 13729.515 190.325 ;
      RECT 13725.595 189.04 13725.875 190.365 ;
      RECT 13721.955 189.04 13722.235 190.35 ;
      RECT 13718.315 189.04 13718.595 190.26 ;
      RECT 13659.235 189.04 13659.515 190.16 ;
      RECT 13655.315 189.04 13655.595 190.205 ;
      RECT 13651.395 189.04 13651.675 189.935 ;
      RECT 13647.475 189.04 13647.755 190.16 ;
      RECT 13643.555 189.04 13643.835 205.605 ;
      RECT 13596.515 189.04 13596.795 190.305 ;
      RECT 13592.875 189.04 13593.155 190.27 ;
      RECT 13589.235 189.04 13589.515 190.325 ;
      RECT 13585.595 189.04 13585.875 190.365 ;
      RECT 13581.955 189.04 13582.235 190.35 ;
      RECT 13578.315 189.04 13578.595 190.26 ;
      RECT 13519.235 189.04 13519.515 190.16 ;
      RECT 13515.315 189.04 13515.595 190.205 ;
      RECT 13511.395 189.04 13511.675 189.935 ;
      RECT 13507.475 189.04 13507.755 190.16 ;
      RECT 13503.555 189.04 13503.835 205.605 ;
      RECT 13456.515 189.04 13456.795 190.305 ;
      RECT 13452.875 189.04 13453.155 190.27 ;
      RECT 13449.235 189.04 13449.515 190.325 ;
      RECT 13445.595 189.04 13445.875 190.365 ;
      RECT 13441.955 189.04 13442.235 190.35 ;
      RECT 13438.315 189.04 13438.595 190.26 ;
      RECT 13379.235 189.04 13379.515 190.16 ;
      RECT 13375.315 189.04 13375.595 190.205 ;
      RECT 13371.395 189.04 13371.675 189.935 ;
      RECT 13367.475 189.04 13367.755 190.16 ;
      RECT 13363.555 189.04 13363.835 205.605 ;
      RECT 13316.515 189.04 13316.795 190.305 ;
      RECT 13312.875 189.04 13313.155 190.27 ;
      RECT 13309.235 189.04 13309.515 190.325 ;
      RECT 13305.595 189.04 13305.875 190.365 ;
      RECT 13301.955 189.04 13302.235 190.35 ;
      RECT 13298.315 189.04 13298.595 190.26 ;
      RECT 13239.235 189.04 13239.515 190.16 ;
      RECT 13235.315 189.04 13235.595 190.205 ;
      RECT 13231.395 189.04 13231.675 189.935 ;
      RECT 13227.475 189.04 13227.755 190.16 ;
      RECT 13223.555 189.04 13223.835 205.605 ;
      RECT 13176.515 189.04 13176.795 190.305 ;
      RECT 13172.875 189.04 13173.155 190.27 ;
      RECT 13169.235 189.04 13169.515 190.325 ;
      RECT 13165.595 189.04 13165.875 190.365 ;
      RECT 13161.955 189.04 13162.235 190.35 ;
      RECT 13158.315 189.04 13158.595 190.26 ;
      RECT 13099.235 189.04 13099.515 190.16 ;
      RECT 13095.315 189.04 13095.595 190.205 ;
      RECT 13091.395 189.04 13091.675 189.935 ;
      RECT 13087.475 189.04 13087.755 190.16 ;
      RECT 13083.555 189.04 13083.835 205.605 ;
      RECT 13036.515 189.04 13036.795 190.305 ;
      RECT 13032.875 189.04 13033.155 190.27 ;
      RECT 13029.235 189.04 13029.515 190.325 ;
      RECT 13025.595 189.04 13025.875 190.365 ;
      RECT 13021.955 189.04 13022.235 190.35 ;
      RECT 13018.315 189.04 13018.595 190.26 ;
      RECT 12959.235 189.04 12959.515 190.16 ;
      RECT 12955.315 189.04 12955.595 190.205 ;
      RECT 12951.395 189.04 12951.675 189.935 ;
      RECT 12947.475 189.04 12947.755 190.16 ;
      RECT 12943.555 189.04 12943.835 205.605 ;
      RECT 12896.515 189.04 12896.795 190.305 ;
      RECT 12892.875 189.04 12893.155 190.27 ;
      RECT 12889.235 189.04 12889.515 190.325 ;
      RECT 12885.595 189.04 12885.875 190.365 ;
      RECT 12881.955 189.04 12882.235 190.35 ;
      RECT 12878.315 189.04 12878.595 190.26 ;
      RECT 12819.235 189.04 12819.515 190.16 ;
      RECT 12815.315 189.04 12815.595 190.205 ;
      RECT 12811.395 189.04 12811.675 189.935 ;
      RECT 12807.475 189.04 12807.755 190.16 ;
      RECT 12803.555 189.04 12803.835 205.605 ;
      RECT 12756.515 189.04 12756.795 190.305 ;
      RECT 12752.875 189.04 12753.155 190.27 ;
      RECT 12749.235 189.04 12749.515 190.325 ;
      RECT 12745.595 189.04 12745.875 190.365 ;
      RECT 12741.955 189.04 12742.235 190.35 ;
      RECT 12738.315 189.04 12738.595 190.26 ;
      RECT 12679.235 189.04 12679.515 190.16 ;
      RECT 12675.315 189.04 12675.595 190.205 ;
      RECT 12671.395 189.04 12671.675 189.935 ;
      RECT 12667.475 189.04 12667.755 190.16 ;
      RECT 12663.555 189.04 12663.835 205.605 ;
      RECT 12616.515 189.04 12616.795 190.305 ;
      RECT 12612.875 189.04 12613.155 190.27 ;
      RECT 12609.235 189.04 12609.515 190.325 ;
      RECT 12605.595 189.04 12605.875 190.365 ;
      RECT 12601.955 189.04 12602.235 190.35 ;
      RECT 12598.315 189.04 12598.595 190.26 ;
      RECT 12539.235 189.04 12539.515 190.16 ;
      RECT 12535.315 189.04 12535.595 190.205 ;
      RECT 12531.395 189.04 12531.675 189.935 ;
      RECT 12527.475 189.04 12527.755 190.16 ;
      RECT 12523.555 189.04 12523.835 205.605 ;
      RECT 12476.515 189.04 12476.795 190.305 ;
      RECT 12472.875 189.04 12473.155 190.27 ;
      RECT 12469.235 189.04 12469.515 190.325 ;
      RECT 12465.595 189.04 12465.875 190.365 ;
      RECT 12461.955 189.04 12462.235 190.35 ;
      RECT 12458.315 189.04 12458.595 190.26 ;
      RECT 12399.235 189.04 12399.515 190.16 ;
      RECT 12395.315 189.04 12395.595 190.205 ;
      RECT 12391.395 189.04 12391.675 189.935 ;
      RECT 12387.475 189.04 12387.755 190.16 ;
      RECT 12383.555 189.04 12383.835 205.605 ;
      RECT 12336.515 189.04 12336.795 190.305 ;
      RECT 12332.875 189.04 12333.155 190.27 ;
      RECT 12329.235 189.04 12329.515 190.325 ;
      RECT 12325.595 189.04 12325.875 190.365 ;
      RECT 12321.955 189.04 12322.235 190.35 ;
      RECT 12318.315 189.04 12318.595 190.26 ;
      RECT 12259.235 189.04 12259.515 190.16 ;
      RECT 12255.315 189.04 12255.595 190.205 ;
      RECT 12251.395 189.04 12251.675 189.935 ;
      RECT 12247.475 189.04 12247.755 190.16 ;
      RECT 12243.555 189.04 12243.835 205.605 ;
      RECT 12196.515 189.04 12196.795 190.305 ;
      RECT 12192.875 189.04 12193.155 190.27 ;
      RECT 12189.235 189.04 12189.515 190.325 ;
      RECT 12185.595 189.04 12185.875 190.365 ;
      RECT 12181.955 189.04 12182.235 190.35 ;
      RECT 12178.315 189.04 12178.595 190.26 ;
      RECT 12119.235 189.04 12119.515 190.16 ;
      RECT 12115.315 189.04 12115.595 190.205 ;
      RECT 12111.395 189.04 12111.675 189.935 ;
      RECT 12107.475 189.04 12107.755 190.16 ;
      RECT 12103.555 189.04 12103.835 205.605 ;
      RECT 12056.515 189.04 12056.795 190.305 ;
      RECT 12052.875 189.04 12053.155 190.27 ;
      RECT 12049.235 189.04 12049.515 190.325 ;
      RECT 12045.595 189.04 12045.875 190.365 ;
      RECT 12041.955 189.04 12042.235 190.35 ;
      RECT 12038.315 189.04 12038.595 190.26 ;
      RECT 11979.235 189.04 11979.515 190.16 ;
      RECT 11975.315 189.04 11975.595 190.205 ;
      RECT 11971.395 189.04 11971.675 189.935 ;
      RECT 11967.475 189.04 11967.755 190.16 ;
      RECT 11963.555 189.04 11963.835 205.605 ;
      RECT 11916.515 189.04 11916.795 190.305 ;
      RECT 11912.875 189.04 11913.155 190.27 ;
      RECT 11909.235 189.04 11909.515 190.325 ;
      RECT 11905.595 189.04 11905.875 190.365 ;
      RECT 11901.955 189.04 11902.235 190.35 ;
      RECT 11898.315 189.04 11898.595 190.26 ;
      RECT 11839.235 189.04 11839.515 190.16 ;
      RECT 11835.315 189.04 11835.595 190.205 ;
      RECT 11831.395 189.04 11831.675 189.935 ;
      RECT 11827.475 189.04 11827.755 190.16 ;
      RECT 11823.555 189.04 11823.835 205.605 ;
      RECT 11776.515 189.04 11776.795 190.305 ;
      RECT 11772.875 189.04 11773.155 190.27 ;
      RECT 11769.235 189.04 11769.515 190.325 ;
      RECT 11765.595 189.04 11765.875 190.365 ;
      RECT 11761.955 189.04 11762.235 190.35 ;
      RECT 11758.315 189.04 11758.595 190.26 ;
      RECT 11699.235 189.04 11699.515 190.16 ;
      RECT 11695.315 189.04 11695.595 190.205 ;
      RECT 11691.395 189.04 11691.675 189.935 ;
      RECT 11687.475 189.04 11687.755 190.16 ;
      RECT 11683.555 189.04 11683.835 205.605 ;
      RECT 11636.515 189.04 11636.795 190.305 ;
      RECT 11632.875 189.04 11633.155 190.27 ;
      RECT 11629.235 189.04 11629.515 190.325 ;
      RECT 11625.595 189.04 11625.875 190.365 ;
      RECT 11621.955 189.04 11622.235 190.35 ;
      RECT 11618.315 189.04 11618.595 190.26 ;
      RECT 11559.235 189.04 11559.515 190.16 ;
      RECT 11555.315 189.04 11555.595 190.205 ;
      RECT 11551.395 189.04 11551.675 189.935 ;
      RECT 11547.475 189.04 11547.755 190.16 ;
      RECT 11543.555 189.04 11543.835 205.605 ;
      RECT 11496.515 189.04 11496.795 190.305 ;
      RECT 11492.875 189.04 11493.155 190.27 ;
      RECT 11489.235 189.04 11489.515 190.325 ;
      RECT 11485.595 189.04 11485.875 190.365 ;
      RECT 11481.955 189.04 11482.235 190.35 ;
      RECT 11478.315 189.04 11478.595 190.26 ;
      RECT 11419.235 189.04 11419.515 190.16 ;
      RECT 11415.315 189.04 11415.595 190.205 ;
      RECT 11411.395 189.04 11411.675 189.935 ;
      RECT 11407.475 189.04 11407.755 190.16 ;
      RECT 11403.555 189.04 11403.835 205.605 ;
      RECT 11356.515 189.04 11356.795 190.305 ;
      RECT 11352.875 189.04 11353.155 190.27 ;
      RECT 11349.235 189.04 11349.515 190.325 ;
      RECT 11345.595 189.04 11345.875 190.365 ;
      RECT 11341.955 189.04 11342.235 190.35 ;
      RECT 11338.315 189.04 11338.595 190.26 ;
      RECT 11279.235 189.04 11279.515 190.16 ;
      RECT 11275.315 189.04 11275.595 190.205 ;
      RECT 11271.395 189.04 11271.675 189.935 ;
      RECT 11267.475 189.04 11267.755 190.16 ;
      RECT 11263.555 189.04 11263.835 205.605 ;
      RECT 11216.515 189.04 11216.795 190.305 ;
      RECT 11212.875 189.04 11213.155 190.27 ;
      RECT 11209.235 189.04 11209.515 190.325 ;
      RECT 11205.595 189.04 11205.875 190.365 ;
      RECT 11201.955 189.04 11202.235 190.35 ;
      RECT 11198.315 189.04 11198.595 190.26 ;
      RECT 11139.235 189.04 11139.515 190.16 ;
      RECT 11135.315 189.04 11135.595 190.205 ;
      RECT 11131.395 189.04 11131.675 189.935 ;
      RECT 11127.475 189.04 11127.755 190.16 ;
      RECT 11123.555 189.04 11123.835 205.605 ;
      RECT 11076.515 189.04 11076.795 190.305 ;
      RECT 11072.875 189.04 11073.155 190.27 ;
      RECT 11069.235 189.04 11069.515 190.325 ;
      RECT 11065.595 189.04 11065.875 190.365 ;
      RECT 11061.955 189.04 11062.235 190.35 ;
      RECT 11058.315 189.04 11058.595 190.26 ;
      RECT 10999.235 189.04 10999.515 190.16 ;
      RECT 10995.315 189.04 10995.595 190.205 ;
      RECT 10991.395 189.04 10991.675 189.935 ;
      RECT 10987.475 189.04 10987.755 190.16 ;
      RECT 10983.555 189.04 10983.835 205.605 ;
      RECT 10936.515 189.04 10936.795 190.305 ;
      RECT 10932.875 189.04 10933.155 190.27 ;
      RECT 10929.235 189.04 10929.515 190.325 ;
      RECT 10925.595 189.04 10925.875 190.365 ;
      RECT 10921.955 189.04 10922.235 190.35 ;
      RECT 10918.315 189.04 10918.595 190.26 ;
      RECT 10859.235 189.04 10859.515 190.16 ;
      RECT 10855.315 189.04 10855.595 190.205 ;
      RECT 10851.395 189.04 10851.675 189.935 ;
      RECT 10847.475 189.04 10847.755 190.16 ;
      RECT 10843.555 189.04 10843.835 205.605 ;
      RECT 10796.515 189.04 10796.795 190.305 ;
      RECT 10792.875 189.04 10793.155 190.27 ;
      RECT 10789.235 189.04 10789.515 190.325 ;
      RECT 10785.595 189.04 10785.875 190.365 ;
      RECT 10781.955 189.04 10782.235 190.35 ;
      RECT 10778.315 189.04 10778.595 190.26 ;
      RECT 10719.235 189.04 10719.515 190.16 ;
      RECT 10715.315 189.04 10715.595 190.205 ;
      RECT 10711.395 189.04 10711.675 189.935 ;
      RECT 10707.475 189.04 10707.755 190.16 ;
      RECT 10703.555 189.04 10703.835 205.605 ;
      RECT 10656.515 189.04 10656.795 190.305 ;
      RECT 10652.875 189.04 10653.155 190.27 ;
      RECT 10649.235 189.04 10649.515 190.325 ;
      RECT 10645.595 189.04 10645.875 190.365 ;
      RECT 10641.955 189.04 10642.235 190.35 ;
      RECT 10638.315 189.04 10638.595 190.26 ;
      RECT 10579.235 189.04 10579.515 190.16 ;
      RECT 10575.315 189.04 10575.595 190.205 ;
      RECT 10571.395 189.04 10571.675 189.935 ;
      RECT 10567.475 189.04 10567.755 190.16 ;
      RECT 10563.555 189.04 10563.835 205.605 ;
      RECT 10516.515 189.04 10516.795 190.305 ;
      RECT 10512.875 189.04 10513.155 190.27 ;
      RECT 10509.235 189.04 10509.515 190.325 ;
      RECT 10505.595 189.04 10505.875 190.365 ;
      RECT 10501.955 189.04 10502.235 190.35 ;
      RECT 10498.315 189.04 10498.595 190.26 ;
      RECT 10439.235 189.04 10439.515 190.16 ;
      RECT 10435.315 189.04 10435.595 190.205 ;
      RECT 10431.395 189.04 10431.675 189.935 ;
      RECT 10427.475 189.04 10427.755 190.16 ;
      RECT 10423.555 189.04 10423.835 205.605 ;
      RECT 10376.515 189.04 10376.795 190.305 ;
      RECT 10372.875 189.04 10373.155 190.27 ;
      RECT 10369.235 189.04 10369.515 190.325 ;
      RECT 10365.595 189.04 10365.875 190.365 ;
      RECT 10361.955 189.04 10362.235 190.35 ;
      RECT 10358.315 189.04 10358.595 190.26 ;
      RECT 10299.235 189.04 10299.515 190.16 ;
      RECT 10295.315 189.04 10295.595 190.205 ;
      RECT 10291.395 189.04 10291.675 189.935 ;
      RECT 10287.475 189.04 10287.755 190.16 ;
      RECT 10283.555 189.04 10283.835 205.605 ;
      RECT 10236.515 189.04 10236.795 190.305 ;
      RECT 10232.875 189.04 10233.155 190.27 ;
      RECT 10229.235 189.04 10229.515 190.325 ;
      RECT 10225.595 189.04 10225.875 190.365 ;
      RECT 10221.955 189.04 10222.235 190.35 ;
      RECT 10218.315 189.04 10218.595 190.26 ;
      RECT 10159.235 189.04 10159.515 190.16 ;
      RECT 10155.315 189.04 10155.595 190.205 ;
      RECT 10151.395 189.04 10151.675 189.935 ;
      RECT 10147.475 189.04 10147.755 190.16 ;
      RECT 10143.555 189.04 10143.835 205.605 ;
      RECT 10096.515 189.04 10096.795 190.305 ;
      RECT 10092.875 189.04 10093.155 190.27 ;
      RECT 10089.235 189.04 10089.515 190.325 ;
      RECT 10085.595 189.04 10085.875 190.365 ;
      RECT 10081.955 189.04 10082.235 190.35 ;
      RECT 10078.315 189.04 10078.595 190.26 ;
      RECT 10019.235 189.04 10019.515 190.16 ;
      RECT 10015.315 189.04 10015.595 190.205 ;
      RECT 10011.395 189.04 10011.675 189.935 ;
      RECT 10007.475 189.04 10007.755 190.16 ;
      RECT 10003.555 189.04 10003.835 205.605 ;
      RECT 9956.515 189.04 9956.795 190.305 ;
      RECT 9952.875 189.04 9953.155 190.27 ;
      RECT 9949.235 189.04 9949.515 190.325 ;
      RECT 9945.595 189.04 9945.875 190.365 ;
      RECT 9941.955 189.04 9942.235 190.35 ;
      RECT 9938.315 189.04 9938.595 190.26 ;
      RECT 9879.235 189.04 9879.515 190.16 ;
      RECT 9875.315 189.04 9875.595 190.205 ;
      RECT 9871.395 189.04 9871.675 189.935 ;
      RECT 9867.475 189.04 9867.755 190.16 ;
      RECT 9863.555 189.04 9863.835 205.605 ;
      RECT 9816.515 189.04 9816.795 190.305 ;
      RECT 9812.875 189.04 9813.155 190.27 ;
      RECT 9809.235 189.04 9809.515 190.325 ;
      RECT 9805.595 189.04 9805.875 190.365 ;
      RECT 9801.955 189.04 9802.235 190.35 ;
      RECT 9798.315 189.04 9798.595 190.26 ;
      RECT 9739.235 189.04 9739.515 190.16 ;
      RECT 9735.315 189.04 9735.595 190.205 ;
      RECT 9731.395 189.04 9731.675 189.935 ;
      RECT 9727.475 189.04 9727.755 190.16 ;
      RECT 9723.555 189.04 9723.835 205.605 ;
      RECT 9676.515 189.04 9676.795 190.305 ;
      RECT 9672.875 189.04 9673.155 190.27 ;
      RECT 9669.235 189.04 9669.515 190.325 ;
      RECT 9665.595 189.04 9665.875 190.365 ;
      RECT 9661.955 189.04 9662.235 190.35 ;
      RECT 9658.315 189.04 9658.595 190.26 ;
      RECT 9599.235 189.04 9599.515 190.16 ;
      RECT 9595.315 189.04 9595.595 190.205 ;
      RECT 9591.395 189.04 9591.675 189.935 ;
      RECT 9587.475 189.04 9587.755 190.16 ;
      RECT 9583.555 189.04 9583.835 205.605 ;
      RECT 9536.515 189.04 9536.795 190.305 ;
      RECT 9532.875 189.04 9533.155 190.27 ;
      RECT 9529.235 189.04 9529.515 190.325 ;
      RECT 9525.595 189.04 9525.875 190.365 ;
      RECT 9521.955 189.04 9522.235 190.35 ;
      RECT 9518.315 189.04 9518.595 190.26 ;
      RECT 9459.235 189.04 9459.515 190.16 ;
      RECT 9455.315 189.04 9455.595 190.205 ;
      RECT 9451.395 189.04 9451.675 189.935 ;
      RECT 9447.475 189.04 9447.755 190.16 ;
      RECT 9443.555 189.04 9443.835 205.605 ;
      RECT 9432.795 188.015 9432.885 188.295 ;
      RECT 9430.945 188.015 9431.035 188.295 ;
      RECT 9428.275 189.04 9428.835 190.015 ;
      RECT 9426.595 189.04 9427.155 190.945 ;
      RECT 9424.915 189.04 9425.475 191.875 ;
      RECT 9423.235 189.04 9423.795 192.805 ;
      RECT 9421.555 189.04 9422.115 193.735 ;
      RECT 9419.875 189.04 9420.435 194.665 ;
      RECT 9418.195 189.04 9418.755 195.595 ;
      RECT 9416.515 189.04 9417.075 196.515 ;
      RECT 9414.835 189.04 9415.395 197.445 ;
      RECT 9413.155 189.04 9413.715 198.375 ;
      RECT 9411.475 189.04 9412.035 199.305 ;
      RECT 9409.795 189.04 9410.355 200.235 ;
      RECT 9408.115 189.04 9408.675 201.165 ;
      RECT 9396.515 189.04 9396.795 190.305 ;
      RECT 9392.875 189.04 9393.155 190.27 ;
      RECT 9389.235 189.04 9389.515 190.325 ;
      RECT 9385.595 189.04 9385.875 190.365 ;
      RECT 9381.955 189.04 9382.235 190.35 ;
      RECT 9378.315 189.04 9378.595 190.26 ;
      RECT 9319.235 189.04 9319.515 190.16 ;
      RECT 9315.315 189.04 9315.595 190.205 ;
      RECT 9311.395 189.04 9311.675 189.935 ;
      RECT 9307.475 189.04 9307.755 190.16 ;
      RECT 9303.555 189.04 9303.835 205.605 ;
      RECT 9256.515 189.04 9256.795 190.305 ;
      RECT 9252.875 189.04 9253.155 190.27 ;
      RECT 9249.235 189.04 9249.515 190.325 ;
      RECT 9245.595 189.04 9245.875 190.365 ;
      RECT 9241.955 189.04 9242.235 190.35 ;
      RECT 9238.315 189.04 9238.595 190.26 ;
      RECT 9179.235 189.04 9179.515 190.16 ;
      RECT 9175.315 189.04 9175.595 190.205 ;
      RECT 9171.395 189.04 9171.675 189.935 ;
      RECT 9167.475 189.04 9167.755 190.16 ;
      RECT 9163.555 189.04 9163.835 205.605 ;
      RECT 9116.515 189.04 9116.795 190.305 ;
      RECT 9112.875 189.04 9113.155 190.27 ;
      RECT 9109.235 189.04 9109.515 190.325 ;
      RECT 9105.595 189.04 9105.875 190.365 ;
      RECT 9101.955 189.04 9102.235 190.35 ;
      RECT 9098.315 189.04 9098.595 190.26 ;
      RECT 9039.235 189.04 9039.515 190.16 ;
      RECT 9035.315 189.04 9035.595 190.205 ;
      RECT 9031.395 189.04 9031.675 189.935 ;
      RECT 9027.475 189.04 9027.755 190.16 ;
      RECT 9023.555 189.04 9023.835 205.605 ;
      RECT 8976.515 189.04 8976.795 190.305 ;
      RECT 8972.875 189.04 8973.155 190.27 ;
      RECT 8969.235 189.04 8969.515 190.325 ;
      RECT 8965.595 189.04 8965.875 190.365 ;
      RECT 8961.955 189.04 8962.235 190.35 ;
      RECT 8958.315 189.04 8958.595 190.26 ;
      RECT 8899.235 189.04 8899.515 190.16 ;
      RECT 8895.315 189.04 8895.595 190.205 ;
      RECT 8891.395 189.04 8891.675 189.935 ;
      RECT 8887.475 189.04 8887.755 190.16 ;
      RECT 8883.555 189.04 8883.835 205.605 ;
      RECT 8836.515 189.04 8836.795 190.305 ;
      RECT 8832.875 189.04 8833.155 190.27 ;
      RECT 8829.235 189.04 8829.515 190.325 ;
      RECT 8825.595 189.04 8825.875 190.365 ;
      RECT 8821.955 189.04 8822.235 190.35 ;
      RECT 8818.315 189.04 8818.595 190.26 ;
      RECT 8759.235 189.04 8759.515 190.16 ;
      RECT 8755.315 189.04 8755.595 190.205 ;
      RECT 8751.395 189.04 8751.675 189.935 ;
      RECT 8747.475 189.04 8747.755 190.16 ;
      RECT 8743.555 189.04 8743.835 205.605 ;
      RECT 8696.515 189.04 8696.795 190.305 ;
      RECT 8692.875 189.04 8693.155 190.27 ;
      RECT 8689.235 189.04 8689.515 190.325 ;
      RECT 8685.595 189.04 8685.875 190.365 ;
      RECT 8681.955 189.04 8682.235 190.35 ;
      RECT 8678.315 189.04 8678.595 190.26 ;
      RECT 8619.235 189.04 8619.515 190.16 ;
      RECT 8615.315 189.04 8615.595 190.205 ;
      RECT 8611.395 189.04 8611.675 189.935 ;
      RECT 8607.475 189.04 8607.755 190.16 ;
      RECT 8603.555 189.04 8603.835 205.605 ;
      RECT 8556.515 189.04 8556.795 190.305 ;
      RECT 8552.875 189.04 8553.155 190.27 ;
      RECT 8549.235 189.04 8549.515 190.325 ;
      RECT 8545.595 189.04 8545.875 190.365 ;
      RECT 8541.955 189.04 8542.235 190.35 ;
      RECT 8538.315 189.04 8538.595 190.26 ;
      RECT 8479.235 189.04 8479.515 190.16 ;
      RECT 8475.315 189.04 8475.595 190.205 ;
      RECT 8471.395 189.04 8471.675 189.935 ;
      RECT 8467.475 189.04 8467.755 190.16 ;
      RECT 8463.555 189.04 8463.835 205.605 ;
      RECT 8416.515 189.04 8416.795 190.305 ;
      RECT 8412.875 189.04 8413.155 190.27 ;
      RECT 8409.235 189.04 8409.515 190.325 ;
      RECT 8405.595 189.04 8405.875 190.365 ;
      RECT 8401.955 189.04 8402.235 190.35 ;
      RECT 8398.315 189.04 8398.595 190.26 ;
      RECT 8339.235 189.04 8339.515 190.16 ;
      RECT 8335.315 189.04 8335.595 190.205 ;
      RECT 8331.395 189.04 8331.675 189.935 ;
      RECT 8327.475 189.04 8327.755 190.16 ;
      RECT 8323.555 189.04 8323.835 205.605 ;
      RECT 8276.515 189.04 8276.795 190.305 ;
      RECT 8272.875 189.04 8273.155 190.27 ;
      RECT 8269.235 189.04 8269.515 190.325 ;
      RECT 8265.595 189.04 8265.875 190.365 ;
      RECT 8261.955 189.04 8262.235 190.35 ;
      RECT 8258.315 189.04 8258.595 190.26 ;
      RECT 8199.235 189.04 8199.515 190.16 ;
      RECT 8195.315 189.04 8195.595 190.205 ;
      RECT 8191.395 189.04 8191.675 189.935 ;
      RECT 8187.475 189.04 8187.755 190.16 ;
      RECT 8183.555 189.04 8183.835 205.605 ;
      RECT 8136.515 189.04 8136.795 190.305 ;
      RECT 8132.875 189.04 8133.155 190.27 ;
      RECT 8129.235 189.04 8129.515 190.325 ;
      RECT 8125.595 189.04 8125.875 190.365 ;
      RECT 8121.955 189.04 8122.235 190.35 ;
      RECT 8118.315 189.04 8118.595 190.26 ;
      RECT 8059.235 189.04 8059.515 190.16 ;
      RECT 8055.315 189.04 8055.595 190.205 ;
      RECT 8051.395 189.04 8051.675 189.935 ;
      RECT 8047.475 189.04 8047.755 190.16 ;
      RECT 8043.555 189.04 8043.835 205.605 ;
      RECT 7996.515 189.04 7996.795 190.305 ;
      RECT 7992.875 189.04 7993.155 190.27 ;
      RECT 7989.235 189.04 7989.515 190.325 ;
      RECT 7985.595 189.04 7985.875 190.365 ;
      RECT 7981.955 189.04 7982.235 190.35 ;
      RECT 7978.315 189.04 7978.595 190.26 ;
      RECT 7919.235 189.04 7919.515 190.16 ;
      RECT 7915.315 189.04 7915.595 190.205 ;
      RECT 7911.395 189.04 7911.675 189.935 ;
      RECT 7907.475 189.04 7907.755 190.16 ;
      RECT 7903.555 189.04 7903.835 205.605 ;
      RECT 7856.515 189.04 7856.795 190.305 ;
      RECT 7852.875 189.04 7853.155 190.27 ;
      RECT 7849.235 189.04 7849.515 190.325 ;
      RECT 7845.595 189.04 7845.875 190.365 ;
      RECT 7841.955 189.04 7842.235 190.35 ;
      RECT 7838.315 189.04 7838.595 190.26 ;
      RECT 7779.235 189.04 7779.515 190.16 ;
      RECT 7775.315 189.04 7775.595 190.205 ;
      RECT 7771.395 189.04 7771.675 189.935 ;
      RECT 7767.475 189.04 7767.755 190.16 ;
      RECT 7763.555 189.04 7763.835 205.605 ;
      RECT 7716.515 189.04 7716.795 190.305 ;
      RECT 7712.875 189.04 7713.155 190.27 ;
      RECT 7709.235 189.04 7709.515 190.325 ;
      RECT 7705.595 189.04 7705.875 190.365 ;
      RECT 7701.955 189.04 7702.235 190.35 ;
      RECT 7698.315 189.04 7698.595 190.26 ;
      RECT 7639.235 189.04 7639.515 190.16 ;
      RECT 7635.315 189.04 7635.595 190.205 ;
      RECT 7631.395 189.04 7631.675 189.935 ;
      RECT 7627.475 189.04 7627.755 190.16 ;
      RECT 7623.555 189.04 7623.835 205.605 ;
      RECT 7576.515 189.04 7576.795 190.305 ;
      RECT 7572.875 189.04 7573.155 190.27 ;
      RECT 7569.235 189.04 7569.515 190.325 ;
      RECT 7565.595 189.04 7565.875 190.365 ;
      RECT 7561.955 189.04 7562.235 190.35 ;
      RECT 7558.315 189.04 7558.595 190.26 ;
      RECT 7499.235 189.04 7499.515 190.16 ;
      RECT 7495.315 189.04 7495.595 190.205 ;
      RECT 7491.395 189.04 7491.675 189.935 ;
      RECT 7487.475 189.04 7487.755 190.16 ;
      RECT 7483.555 189.04 7483.835 205.605 ;
      RECT 7436.515 189.04 7436.795 190.305 ;
      RECT 7432.875 189.04 7433.155 190.27 ;
      RECT 7429.235 189.04 7429.515 190.325 ;
      RECT 7425.595 189.04 7425.875 190.365 ;
      RECT 7421.955 189.04 7422.235 190.35 ;
      RECT 7418.315 189.04 7418.595 190.26 ;
      RECT 7359.235 189.04 7359.515 190.16 ;
      RECT 7355.315 189.04 7355.595 190.205 ;
      RECT 7351.395 189.04 7351.675 189.935 ;
      RECT 7347.475 189.04 7347.755 190.16 ;
      RECT 7343.555 189.04 7343.835 205.605 ;
      RECT 7296.515 189.04 7296.795 190.305 ;
      RECT 7292.875 189.04 7293.155 190.27 ;
      RECT 7289.235 189.04 7289.515 190.325 ;
      RECT 7285.595 189.04 7285.875 190.365 ;
      RECT 7281.955 189.04 7282.235 190.35 ;
      RECT 7278.315 189.04 7278.595 190.26 ;
      RECT 7219.235 189.04 7219.515 190.16 ;
      RECT 7215.315 189.04 7215.595 190.205 ;
      RECT 7211.395 189.04 7211.675 189.935 ;
      RECT 7207.475 189.04 7207.755 190.16 ;
      RECT 7203.555 189.04 7203.835 205.605 ;
      RECT 7156.515 189.04 7156.795 190.305 ;
      RECT 7152.875 189.04 7153.155 190.27 ;
      RECT 7149.235 189.04 7149.515 190.325 ;
      RECT 7145.595 189.04 7145.875 190.365 ;
      RECT 7141.955 189.04 7142.235 190.35 ;
      RECT 7138.315 189.04 7138.595 190.26 ;
      RECT 7079.235 189.04 7079.515 190.16 ;
      RECT 7075.315 189.04 7075.595 190.205 ;
      RECT 7071.395 189.04 7071.675 189.935 ;
      RECT 7067.475 189.04 7067.755 190.16 ;
      RECT 7063.555 189.04 7063.835 205.605 ;
      RECT 7016.515 189.04 7016.795 190.305 ;
      RECT 7012.875 189.04 7013.155 190.27 ;
      RECT 7009.235 189.04 7009.515 190.325 ;
      RECT 7005.595 189.04 7005.875 190.365 ;
      RECT 7001.955 189.04 7002.235 190.35 ;
      RECT 6998.315 189.04 6998.595 190.26 ;
      RECT 6939.235 189.04 6939.515 190.16 ;
      RECT 6935.315 189.04 6935.595 190.205 ;
      RECT 6931.395 189.04 6931.675 189.935 ;
      RECT 6927.475 189.04 6927.755 190.16 ;
      RECT 6923.555 189.04 6923.835 205.605 ;
      RECT 6876.515 189.04 6876.795 190.305 ;
      RECT 6872.875 189.04 6873.155 190.27 ;
      RECT 6869.235 189.04 6869.515 190.325 ;
      RECT 6865.595 189.04 6865.875 190.365 ;
      RECT 6861.955 189.04 6862.235 190.35 ;
      RECT 6858.315 189.04 6858.595 190.26 ;
      RECT 6799.235 189.04 6799.515 190.16 ;
      RECT 6795.315 189.04 6795.595 190.205 ;
      RECT 6791.395 189.04 6791.675 189.935 ;
      RECT 6787.475 189.04 6787.755 190.16 ;
      RECT 6783.555 189.04 6783.835 205.605 ;
      RECT 6736.515 189.04 6736.795 190.305 ;
      RECT 6732.875 189.04 6733.155 190.27 ;
      RECT 6729.235 189.04 6729.515 190.325 ;
      RECT 6725.595 189.04 6725.875 190.365 ;
      RECT 6721.955 189.04 6722.235 190.35 ;
      RECT 6718.315 189.04 6718.595 190.26 ;
      RECT 6659.235 189.04 6659.515 190.16 ;
      RECT 6655.315 189.04 6655.595 190.205 ;
      RECT 6651.395 189.04 6651.675 189.935 ;
      RECT 6647.475 189.04 6647.755 190.16 ;
      RECT 6643.555 189.04 6643.835 205.605 ;
      RECT 6596.515 189.04 6596.795 190.305 ;
      RECT 6592.875 189.04 6593.155 190.27 ;
      RECT 6589.235 189.04 6589.515 190.325 ;
      RECT 6585.595 189.04 6585.875 190.365 ;
      RECT 6581.955 189.04 6582.235 190.35 ;
      RECT 6578.315 189.04 6578.595 190.26 ;
      RECT 6519.235 189.04 6519.515 190.16 ;
      RECT 6515.315 189.04 6515.595 190.205 ;
      RECT 6511.395 189.04 6511.675 189.935 ;
      RECT 6507.475 189.04 6507.755 190.16 ;
      RECT 6503.555 189.04 6503.835 205.605 ;
      RECT 6456.515 189.04 6456.795 190.305 ;
      RECT 6452.875 189.04 6453.155 190.27 ;
      RECT 6449.235 189.04 6449.515 190.325 ;
      RECT 6445.595 189.04 6445.875 190.365 ;
      RECT 6441.955 189.04 6442.235 190.35 ;
      RECT 6438.315 189.04 6438.595 190.26 ;
      RECT 6379.235 189.04 6379.515 190.16 ;
      RECT 6375.315 189.04 6375.595 190.205 ;
      RECT 6371.395 189.04 6371.675 189.935 ;
      RECT 6367.475 189.04 6367.755 190.16 ;
      RECT 6363.555 189.04 6363.835 205.605 ;
      RECT 6316.515 189.04 6316.795 190.305 ;
      RECT 6312.875 189.04 6313.155 190.27 ;
      RECT 6309.235 189.04 6309.515 190.325 ;
      RECT 6305.595 189.04 6305.875 190.365 ;
      RECT 6301.955 189.04 6302.235 190.35 ;
      RECT 6298.315 189.04 6298.595 190.26 ;
      RECT 6239.235 189.04 6239.515 190.16 ;
      RECT 6235.315 189.04 6235.595 190.205 ;
      RECT 6231.395 189.04 6231.675 189.935 ;
      RECT 6227.475 189.04 6227.755 190.16 ;
      RECT 6223.555 189.04 6223.835 205.605 ;
      RECT 6176.515 189.04 6176.795 190.305 ;
      RECT 6172.875 189.04 6173.155 190.27 ;
      RECT 6169.235 189.04 6169.515 190.325 ;
      RECT 6165.595 189.04 6165.875 190.365 ;
      RECT 6161.955 189.04 6162.235 190.35 ;
      RECT 6158.315 189.04 6158.595 190.26 ;
      RECT 6099.235 189.04 6099.515 190.16 ;
      RECT 6095.315 189.04 6095.595 190.205 ;
      RECT 6091.395 189.04 6091.675 189.935 ;
      RECT 6087.475 189.04 6087.755 190.16 ;
      RECT 6083.555 189.04 6083.835 205.605 ;
      RECT 6036.515 189.04 6036.795 190.305 ;
      RECT 6032.875 189.04 6033.155 190.27 ;
      RECT 6029.235 189.04 6029.515 190.325 ;
      RECT 6025.595 189.04 6025.875 190.365 ;
      RECT 6021.955 189.04 6022.235 190.35 ;
      RECT 6018.315 189.04 6018.595 190.26 ;
      RECT 5959.235 189.04 5959.515 190.16 ;
      RECT 5955.315 189.04 5955.595 190.205 ;
      RECT 5951.395 189.04 5951.675 189.935 ;
      RECT 5947.475 189.04 5947.755 190.16 ;
      RECT 5943.555 189.04 5943.835 205.605 ;
      RECT 5896.515 189.04 5896.795 190.305 ;
      RECT 5892.875 189.04 5893.155 190.27 ;
      RECT 5889.235 189.04 5889.515 190.325 ;
      RECT 5885.595 189.04 5885.875 190.365 ;
      RECT 5881.955 189.04 5882.235 190.35 ;
      RECT 5878.315 189.04 5878.595 190.26 ;
      RECT 5819.235 189.04 5819.515 190.16 ;
      RECT 5815.315 189.04 5815.595 190.205 ;
      RECT 5811.395 189.04 5811.675 189.935 ;
      RECT 5807.475 189.04 5807.755 190.16 ;
      RECT 5803.555 189.04 5803.835 205.605 ;
      RECT 5756.515 189.04 5756.795 190.305 ;
      RECT 5752.875 189.04 5753.155 190.27 ;
      RECT 5749.235 189.04 5749.515 190.325 ;
      RECT 5745.595 189.04 5745.875 190.365 ;
      RECT 5741.955 189.04 5742.235 190.35 ;
      RECT 5738.315 189.04 5738.595 190.26 ;
      RECT 5679.235 189.04 5679.515 190.16 ;
      RECT 5675.315 189.04 5675.595 190.205 ;
      RECT 5671.395 189.04 5671.675 189.935 ;
      RECT 5667.475 189.04 5667.755 190.16 ;
      RECT 5663.555 189.04 5663.835 205.605 ;
      RECT 5616.515 189.04 5616.795 190.305 ;
      RECT 5612.875 189.04 5613.155 190.27 ;
      RECT 5609.235 189.04 5609.515 190.325 ;
      RECT 5605.595 189.04 5605.875 190.365 ;
      RECT 5601.955 189.04 5602.235 190.35 ;
      RECT 5598.315 189.04 5598.595 190.26 ;
      RECT 5539.235 189.04 5539.515 190.16 ;
      RECT 5535.315 189.04 5535.595 190.205 ;
      RECT 5531.395 189.04 5531.675 189.935 ;
      RECT 5527.475 189.04 5527.755 190.16 ;
      RECT 5523.555 189.04 5523.835 205.605 ;
      RECT 5476.515 189.04 5476.795 190.305 ;
      RECT 5472.875 189.04 5473.155 190.27 ;
      RECT 5469.235 189.04 5469.515 190.325 ;
      RECT 5465.595 189.04 5465.875 190.365 ;
      RECT 5461.955 189.04 5462.235 190.35 ;
      RECT 5458.315 189.04 5458.595 190.26 ;
      RECT 5399.235 189.04 5399.515 190.16 ;
      RECT 5395.315 189.04 5395.595 190.205 ;
      RECT 5391.395 189.04 5391.675 189.935 ;
      RECT 5387.475 189.04 5387.755 190.16 ;
      RECT 5383.555 189.04 5383.835 205.605 ;
      RECT 5336.515 189.04 5336.795 190.305 ;
      RECT 5332.875 189.04 5333.155 190.27 ;
      RECT 5329.235 189.04 5329.515 190.325 ;
      RECT 5325.595 189.04 5325.875 190.365 ;
      RECT 5321.955 189.04 5322.235 190.35 ;
      RECT 5318.315 189.04 5318.595 190.26 ;
      RECT 5259.235 189.04 5259.515 190.16 ;
      RECT 5255.315 189.04 5255.595 190.205 ;
      RECT 5251.395 189.04 5251.675 189.935 ;
      RECT 5247.475 189.04 5247.755 190.16 ;
      RECT 5243.555 189.04 5243.835 205.605 ;
      RECT 5196.515 189.04 5196.795 190.305 ;
      RECT 5192.875 189.04 5193.155 190.27 ;
      RECT 5189.235 189.04 5189.515 190.325 ;
      RECT 5185.595 189.04 5185.875 190.365 ;
      RECT 5181.955 189.04 5182.235 190.35 ;
      RECT 5178.315 189.04 5178.595 190.26 ;
      RECT 5119.235 189.04 5119.515 190.16 ;
      RECT 5115.315 189.04 5115.595 190.205 ;
      RECT 5111.395 189.04 5111.675 189.935 ;
      RECT 5107.475 189.04 5107.755 190.16 ;
      RECT 5103.555 189.04 5103.835 205.605 ;
      RECT 5056.515 189.04 5056.795 190.305 ;
      RECT 5052.875 189.04 5053.155 190.27 ;
      RECT 5049.235 189.04 5049.515 190.325 ;
      RECT 5045.595 189.04 5045.875 190.365 ;
      RECT 5041.955 189.04 5042.235 190.35 ;
      RECT 5038.315 189.04 5038.595 190.26 ;
      RECT 4979.235 189.04 4979.515 190.16 ;
      RECT 4975.315 189.04 4975.595 190.205 ;
      RECT 4971.395 189.04 4971.675 189.935 ;
      RECT 4967.475 189.04 4967.755 190.16 ;
      RECT 4963.555 189.04 4963.835 205.605 ;
      RECT 4916.515 189.04 4916.795 190.305 ;
      RECT 4912.875 189.04 4913.155 190.27 ;
      RECT 4909.235 189.04 4909.515 190.325 ;
      RECT 4905.595 189.04 4905.875 190.365 ;
      RECT 4901.955 189.04 4902.235 190.35 ;
      RECT 4898.315 189.04 4898.595 190.26 ;
      RECT 4839.235 189.04 4839.515 190.16 ;
      RECT 4835.315 189.04 4835.595 190.205 ;
      RECT 4831.395 189.04 4831.675 189.935 ;
      RECT 4827.475 189.04 4827.755 190.16 ;
      RECT 4823.555 189.04 4823.835 205.605 ;
      RECT 4776.515 189.04 4776.795 190.305 ;
      RECT 4772.875 189.04 4773.155 190.27 ;
      RECT 4769.235 189.04 4769.515 190.325 ;
      RECT 4765.595 189.04 4765.875 190.365 ;
      RECT 4761.955 189.04 4762.235 190.35 ;
      RECT 4758.315 189.04 4758.595 190.26 ;
      RECT 4699.235 189.04 4699.515 190.16 ;
      RECT 4695.315 189.04 4695.595 190.205 ;
      RECT 4691.395 189.04 4691.675 189.935 ;
      RECT 4687.475 189.04 4687.755 190.16 ;
      RECT 4683.555 189.04 4683.835 205.605 ;
      RECT 4636.515 189.04 4636.795 190.305 ;
      RECT 4632.875 189.04 4633.155 190.27 ;
      RECT 4629.235 189.04 4629.515 190.325 ;
      RECT 4625.595 189.04 4625.875 190.365 ;
      RECT 4621.955 189.04 4622.235 190.35 ;
      RECT 4618.315 189.04 4618.595 190.26 ;
      RECT 4559.235 189.04 4559.515 190.16 ;
      RECT 4555.315 189.04 4555.595 190.205 ;
      RECT 4551.395 189.04 4551.675 189.935 ;
      RECT 4547.475 189.04 4547.755 190.16 ;
      RECT 4543.555 189.04 4543.835 205.605 ;
      RECT 4496.515 189.04 4496.795 190.305 ;
      RECT 4492.875 189.04 4493.155 190.27 ;
      RECT 4489.235 189.04 4489.515 190.325 ;
      RECT 4485.595 189.04 4485.875 190.365 ;
      RECT 4481.955 189.04 4482.235 190.35 ;
      RECT 4478.315 189.04 4478.595 190.26 ;
      RECT 4419.235 189.04 4419.515 190.16 ;
      RECT 4415.315 189.04 4415.595 190.205 ;
      RECT 4411.395 189.04 4411.675 189.935 ;
      RECT 4407.475 189.04 4407.755 190.16 ;
      RECT 4403.555 189.04 4403.835 205.605 ;
      RECT 4356.515 189.04 4356.795 190.305 ;
      RECT 4352.875 189.04 4353.155 190.27 ;
      RECT 4349.235 189.04 4349.515 190.325 ;
      RECT 4345.595 189.04 4345.875 190.365 ;
      RECT 4341.955 189.04 4342.235 190.35 ;
      RECT 4338.315 189.04 4338.595 190.26 ;
      RECT 4279.235 189.04 4279.515 190.16 ;
      RECT 4275.315 189.04 4275.595 190.205 ;
      RECT 4271.395 189.04 4271.675 189.935 ;
      RECT 4267.475 189.04 4267.755 190.16 ;
      RECT 4263.555 189.04 4263.835 205.605 ;
      RECT 4216.515 189.04 4216.795 190.305 ;
      RECT 4212.875 189.04 4213.155 190.27 ;
      RECT 4209.235 189.04 4209.515 190.325 ;
      RECT 4205.595 189.04 4205.875 190.365 ;
      RECT 4201.955 189.04 4202.235 190.35 ;
      RECT 4198.315 189.04 4198.595 190.26 ;
      RECT 4139.235 189.04 4139.515 190.16 ;
      RECT 4135.315 189.04 4135.595 190.205 ;
      RECT 4131.395 189.04 4131.675 189.935 ;
      RECT 4127.475 189.04 4127.755 190.16 ;
      RECT 4123.555 189.04 4123.835 205.605 ;
      RECT 4076.515 189.04 4076.795 190.305 ;
      RECT 4072.875 189.04 4073.155 190.27 ;
      RECT 4069.235 189.04 4069.515 190.325 ;
      RECT 4065.595 189.04 4065.875 190.365 ;
      RECT 4061.955 189.04 4062.235 190.35 ;
      RECT 4058.315 189.04 4058.595 190.26 ;
      RECT 3999.235 189.04 3999.515 190.16 ;
      RECT 3995.315 189.04 3995.595 190.205 ;
      RECT 3991.395 189.04 3991.675 189.935 ;
      RECT 3987.475 189.04 3987.755 190.16 ;
      RECT 3983.555 189.04 3983.835 205.605 ;
      RECT 3936.515 189.04 3936.795 190.305 ;
      RECT 3932.875 189.04 3933.155 190.27 ;
      RECT 3929.235 189.04 3929.515 190.325 ;
      RECT 3925.595 189.04 3925.875 190.365 ;
      RECT 3921.955 189.04 3922.235 190.35 ;
      RECT 3918.315 189.04 3918.595 190.26 ;
      RECT 3859.235 189.04 3859.515 190.16 ;
      RECT 3855.315 189.04 3855.595 190.205 ;
      RECT 3851.395 189.04 3851.675 189.935 ;
      RECT 3847.475 189.04 3847.755 190.16 ;
      RECT 3843.555 189.04 3843.835 205.605 ;
      RECT 3796.515 189.04 3796.795 190.305 ;
      RECT 3792.875 189.04 3793.155 190.27 ;
      RECT 3789.235 189.04 3789.515 190.325 ;
      RECT 3785.595 189.04 3785.875 190.365 ;
      RECT 3781.955 189.04 3782.235 190.35 ;
      RECT 3778.315 189.04 3778.595 190.26 ;
      RECT 3719.235 189.04 3719.515 190.16 ;
      RECT 3715.315 189.04 3715.595 190.205 ;
      RECT 3711.395 189.04 3711.675 189.935 ;
      RECT 3707.475 189.04 3707.755 190.16 ;
      RECT 3703.555 189.04 3703.835 205.605 ;
      RECT 3656.515 189.04 3656.795 190.305 ;
      RECT 3652.875 189.04 3653.155 190.27 ;
      RECT 3649.235 189.04 3649.515 190.325 ;
      RECT 3645.595 189.04 3645.875 190.365 ;
      RECT 3641.955 189.04 3642.235 190.35 ;
      RECT 3638.315 189.04 3638.595 190.26 ;
      RECT 3579.235 189.04 3579.515 190.16 ;
      RECT 3575.315 189.04 3575.595 190.205 ;
      RECT 3571.395 189.04 3571.675 189.935 ;
      RECT 3567.475 189.04 3567.755 190.16 ;
      RECT 3563.555 189.04 3563.835 205.605 ;
      RECT 3516.515 189.04 3516.795 190.305 ;
      RECT 3512.875 189.04 3513.155 190.27 ;
      RECT 3509.235 189.04 3509.515 190.325 ;
      RECT 3505.595 189.04 3505.875 190.365 ;
      RECT 3501.955 189.04 3502.235 190.35 ;
      RECT 3498.315 189.04 3498.595 190.26 ;
      RECT 3439.235 189.04 3439.515 190.16 ;
      RECT 3435.315 189.04 3435.595 190.205 ;
      RECT 3431.395 189.04 3431.675 189.935 ;
      RECT 3427.475 189.04 3427.755 190.16 ;
      RECT 3423.555 189.04 3423.835 205.605 ;
      RECT 3376.515 189.04 3376.795 190.305 ;
      RECT 3372.875 189.04 3373.155 190.27 ;
      RECT 3369.235 189.04 3369.515 190.325 ;
      RECT 3365.595 189.04 3365.875 190.365 ;
      RECT 3361.955 189.04 3362.235 190.35 ;
      RECT 3358.315 189.04 3358.595 190.26 ;
      RECT 3299.235 189.04 3299.515 190.16 ;
      RECT 3295.315 189.04 3295.595 190.205 ;
      RECT 3291.395 189.04 3291.675 189.935 ;
      RECT 3287.475 189.04 3287.755 190.16 ;
      RECT 3283.555 189.04 3283.835 205.605 ;
      RECT 3236.515 189.04 3236.795 190.305 ;
      RECT 3232.875 189.04 3233.155 190.27 ;
      RECT 3229.235 189.04 3229.515 190.325 ;
      RECT 3225.595 189.04 3225.875 190.365 ;
      RECT 3221.955 189.04 3222.235 190.35 ;
      RECT 3218.315 189.04 3218.595 190.26 ;
      RECT 3159.235 189.04 3159.515 190.16 ;
      RECT 3155.315 189.04 3155.595 190.205 ;
      RECT 3151.395 189.04 3151.675 189.935 ;
      RECT 3147.475 189.04 3147.755 190.16 ;
      RECT 3143.555 189.04 3143.835 205.605 ;
      RECT 3096.515 189.04 3096.795 190.305 ;
      RECT 3092.875 189.04 3093.155 190.27 ;
      RECT 3089.235 189.04 3089.515 190.325 ;
      RECT 3085.595 189.04 3085.875 190.365 ;
      RECT 3081.955 189.04 3082.235 190.35 ;
      RECT 3078.315 189.04 3078.595 190.26 ;
      RECT 3019.235 189.04 3019.515 190.16 ;
      RECT 3015.315 189.04 3015.595 190.205 ;
      RECT 3011.395 189.04 3011.675 189.935 ;
      RECT 3007.475 189.04 3007.755 190.16 ;
      RECT 3003.555 189.04 3003.835 205.605 ;
      RECT 2956.515 189.04 2956.795 190.305 ;
      RECT 2952.875 189.04 2953.155 190.27 ;
      RECT 2949.235 189.04 2949.515 190.325 ;
      RECT 2945.595 189.04 2945.875 190.365 ;
      RECT 2941.955 189.04 2942.235 190.35 ;
      RECT 2938.315 189.04 2938.595 190.26 ;
      RECT 2879.235 189.04 2879.515 190.16 ;
      RECT 2875.315 189.04 2875.595 190.205 ;
      RECT 2871.395 189.04 2871.675 189.935 ;
      RECT 2867.475 189.04 2867.755 190.16 ;
      RECT 2863.555 189.04 2863.835 205.605 ;
      RECT 2816.515 189.04 2816.795 190.305 ;
      RECT 2812.875 189.04 2813.155 190.27 ;
      RECT 2809.235 189.04 2809.515 190.325 ;
      RECT 2805.595 189.04 2805.875 190.365 ;
      RECT 2801.955 189.04 2802.235 190.35 ;
      RECT 2798.315 189.04 2798.595 190.26 ;
      RECT 2739.235 189.04 2739.515 190.16 ;
      RECT 2735.315 189.04 2735.595 190.205 ;
      RECT 2731.395 189.04 2731.675 189.935 ;
      RECT 2727.475 189.04 2727.755 190.16 ;
      RECT 2723.555 189.04 2723.835 205.605 ;
      RECT 2676.515 189.04 2676.795 190.305 ;
      RECT 2672.875 189.04 2673.155 190.27 ;
      RECT 2669.235 189.04 2669.515 190.325 ;
      RECT 2665.595 189.04 2665.875 190.365 ;
      RECT 2661.955 189.04 2662.235 190.35 ;
      RECT 2658.315 189.04 2658.595 190.26 ;
      RECT 2599.235 189.04 2599.515 190.16 ;
      RECT 2595.315 189.04 2595.595 190.205 ;
      RECT 2591.395 189.04 2591.675 189.935 ;
      RECT 2587.475 189.04 2587.755 190.16 ;
      RECT 2583.555 189.04 2583.835 205.605 ;
      RECT 2536.515 189.04 2536.795 190.305 ;
      RECT 2532.875 189.04 2533.155 190.27 ;
      RECT 2529.235 189.04 2529.515 190.325 ;
      RECT 2525.595 189.04 2525.875 190.365 ;
      RECT 2521.955 189.04 2522.235 190.35 ;
      RECT 2518.315 189.04 2518.595 190.26 ;
      RECT 2459.235 189.04 2459.515 190.16 ;
      RECT 2455.315 189.04 2455.595 190.205 ;
      RECT 2451.395 189.04 2451.675 189.935 ;
      RECT 2447.475 189.04 2447.755 190.16 ;
      RECT 2443.555 189.04 2443.835 205.605 ;
      RECT 2396.515 189.04 2396.795 190.305 ;
      RECT 2392.875 189.04 2393.155 190.27 ;
      RECT 2389.235 189.04 2389.515 190.325 ;
      RECT 2385.595 189.04 2385.875 190.365 ;
      RECT 2381.955 189.04 2382.235 190.35 ;
      RECT 2378.315 189.04 2378.595 190.26 ;
      RECT 2319.235 189.04 2319.515 190.16 ;
      RECT 2315.315 189.04 2315.595 190.205 ;
      RECT 2311.395 189.04 2311.675 189.935 ;
      RECT 2307.475 189.04 2307.755 190.16 ;
      RECT 2303.555 189.04 2303.835 205.605 ;
      RECT 2256.515 189.04 2256.795 190.305 ;
      RECT 2252.875 189.04 2253.155 190.27 ;
      RECT 2249.235 189.04 2249.515 190.325 ;
      RECT 2245.595 189.04 2245.875 190.365 ;
      RECT 2241.955 189.04 2242.235 190.35 ;
      RECT 2238.315 189.04 2238.595 190.26 ;
      RECT 2179.235 189.04 2179.515 190.16 ;
      RECT 2175.315 189.04 2175.595 190.205 ;
      RECT 2171.395 189.04 2171.675 189.935 ;
      RECT 2167.475 189.04 2167.755 190.16 ;
      RECT 2163.555 189.04 2163.835 205.605 ;
      RECT 2116.515 189.04 2116.795 190.305 ;
      RECT 2112.875 189.04 2113.155 190.27 ;
      RECT 2109.235 189.04 2109.515 190.325 ;
      RECT 2105.595 189.04 2105.875 190.365 ;
      RECT 2101.955 189.04 2102.235 190.35 ;
      RECT 2098.315 189.04 2098.595 190.26 ;
      RECT 2039.235 189.04 2039.515 190.16 ;
      RECT 2035.315 189.04 2035.595 190.205 ;
      RECT 2031.395 189.04 2031.675 189.935 ;
      RECT 2027.475 189.04 2027.755 190.16 ;
      RECT 2023.555 189.04 2023.835 205.605 ;
      RECT 1976.515 189.04 1976.795 190.305 ;
      RECT 1972.875 189.04 1973.155 190.27 ;
      RECT 1969.235 189.04 1969.515 190.325 ;
      RECT 1965.595 189.04 1965.875 190.365 ;
      RECT 1961.955 189.04 1962.235 190.35 ;
      RECT 1958.315 189.04 1958.595 190.26 ;
      RECT 1899.235 189.04 1899.515 190.16 ;
      RECT 1895.315 189.04 1895.595 190.205 ;
      RECT 1891.395 189.04 1891.675 189.935 ;
      RECT 1887.475 189.04 1887.755 190.16 ;
      RECT 1883.555 189.04 1883.835 205.605 ;
      RECT 1836.515 189.04 1836.795 190.305 ;
      RECT 1832.875 189.04 1833.155 190.27 ;
      RECT 1829.235 189.04 1829.515 190.325 ;
      RECT 1825.595 189.04 1825.875 190.365 ;
      RECT 1821.955 189.04 1822.235 190.35 ;
      RECT 1818.315 189.04 1818.595 190.26 ;
      RECT 1759.235 189.04 1759.515 190.16 ;
      RECT 1755.315 189.04 1755.595 190.205 ;
      RECT 1751.395 189.04 1751.675 189.935 ;
      RECT 1747.475 189.04 1747.755 190.16 ;
      RECT 1743.555 189.04 1743.835 205.605 ;
      RECT 1696.515 189.04 1696.795 190.305 ;
      RECT 1692.875 189.04 1693.155 190.27 ;
      RECT 1689.235 189.04 1689.515 190.325 ;
      RECT 1685.595 189.04 1685.875 190.365 ;
      RECT 1681.955 189.04 1682.235 190.35 ;
      RECT 1678.315 189.04 1678.595 190.26 ;
      RECT 1619.235 189.04 1619.515 190.16 ;
      RECT 1615.315 189.04 1615.595 190.205 ;
      RECT 1611.395 189.04 1611.675 189.935 ;
      RECT 1607.475 189.04 1607.755 190.16 ;
      RECT 1603.555 189.04 1603.835 205.605 ;
      RECT 1556.515 189.04 1556.795 190.305 ;
      RECT 1552.875 189.04 1553.155 190.27 ;
      RECT 1549.235 189.04 1549.515 190.325 ;
      RECT 1545.595 189.04 1545.875 190.365 ;
      RECT 1541.955 189.04 1542.235 190.35 ;
      RECT 1538.315 189.04 1538.595 190.26 ;
      RECT 1479.235 189.04 1479.515 190.16 ;
      RECT 1475.315 189.04 1475.595 190.205 ;
      RECT 1471.395 189.04 1471.675 189.935 ;
      RECT 1467.475 189.04 1467.755 190.16 ;
      RECT 1463.555 189.04 1463.835 205.605 ;
      RECT 1416.515 189.04 1416.795 190.305 ;
      RECT 1412.875 189.04 1413.155 190.27 ;
      RECT 1409.235 189.04 1409.515 190.325 ;
      RECT 1405.595 189.04 1405.875 190.365 ;
      RECT 1401.955 189.04 1402.235 190.35 ;
      RECT 1398.315 189.04 1398.595 190.26 ;
      RECT 1339.235 189.04 1339.515 190.16 ;
      RECT 1335.315 189.04 1335.595 190.205 ;
      RECT 1331.395 189.04 1331.675 189.935 ;
      RECT 1327.475 189.04 1327.755 190.16 ;
      RECT 1323.555 189.04 1323.835 205.605 ;
      RECT 1276.515 189.04 1276.795 190.305 ;
      RECT 1272.875 189.04 1273.155 190.27 ;
      RECT 1269.235 189.04 1269.515 190.325 ;
      RECT 1265.595 189.04 1265.875 190.365 ;
      RECT 1261.955 189.04 1262.235 190.35 ;
      RECT 1258.315 189.04 1258.595 190.26 ;
      RECT 1199.235 189.04 1199.515 190.16 ;
      RECT 1195.315 189.04 1195.595 190.205 ;
      RECT 1191.395 189.04 1191.675 189.935 ;
      RECT 1187.475 189.04 1187.755 190.16 ;
      RECT 1183.555 189.04 1183.835 205.605 ;
      RECT 1136.515 189.04 1136.795 190.305 ;
      RECT 1132.875 189.04 1133.155 190.27 ;
      RECT 1129.235 189.04 1129.515 190.325 ;
      RECT 1125.595 189.04 1125.875 190.365 ;
      RECT 1121.955 189.04 1122.235 190.35 ;
      RECT 1118.315 189.04 1118.595 190.26 ;
      RECT 1059.235 189.04 1059.515 190.16 ;
      RECT 1055.315 189.04 1055.595 190.205 ;
      RECT 1051.395 189.04 1051.675 189.935 ;
      RECT 1047.475 189.04 1047.755 190.16 ;
      RECT 1043.555 189.04 1043.835 205.605 ;
      RECT 996.515 189.04 996.795 190.305 ;
      RECT 992.875 189.04 993.155 190.27 ;
      RECT 989.235 189.04 989.515 190.325 ;
      RECT 985.595 189.04 985.875 190.365 ;
      RECT 981.955 189.04 982.235 190.35 ;
      RECT 978.315 189.04 978.595 190.26 ;
      RECT 919.235 189.04 919.515 190.16 ;
      RECT 915.315 189.04 915.595 190.205 ;
      RECT 911.395 189.04 911.675 189.935 ;
      RECT 907.475 189.04 907.755 190.16 ;
      RECT 903.555 189.04 903.835 205.605 ;
      RECT 856.515 189.04 856.795 190.305 ;
      RECT 852.875 189.04 853.155 190.27 ;
      RECT 849.235 189.04 849.515 190.325 ;
      RECT 845.595 189.04 845.875 190.365 ;
      RECT 841.955 189.04 842.235 190.35 ;
      RECT 838.315 189.04 838.595 190.26 ;
      RECT 779.235 189.04 779.515 190.16 ;
      RECT 775.315 189.04 775.595 190.205 ;
      RECT 771.395 189.04 771.675 189.935 ;
      RECT 767.475 189.04 767.755 190.16 ;
      RECT 763.555 189.04 763.835 205.605 ;
      RECT 716.515 189.04 716.795 190.305 ;
      RECT 712.875 189.04 713.155 190.27 ;
      RECT 709.235 189.04 709.515 190.325 ;
      RECT 705.595 189.04 705.875 190.365 ;
      RECT 701.955 189.04 702.235 190.35 ;
      RECT 698.315 189.04 698.595 190.26 ;
      RECT 639.235 189.04 639.515 190.16 ;
      RECT 635.315 189.04 635.595 190.205 ;
      RECT 631.395 189.04 631.675 189.935 ;
      RECT 627.475 189.04 627.755 190.16 ;
      RECT 623.555 189.04 623.835 205.605 ;
      RECT 576.515 189.04 576.795 190.305 ;
      RECT 572.875 189.04 573.155 190.27 ;
      RECT 569.235 189.04 569.515 190.325 ;
      RECT 565.595 189.04 565.875 190.365 ;
      RECT 561.955 189.04 562.235 190.35 ;
      RECT 558.315 189.04 558.595 190.26 ;
      RECT 499.235 189.04 499.515 190.16 ;
      RECT 495.315 189.04 495.595 190.205 ;
      RECT 491.395 189.04 491.675 189.935 ;
      RECT 487.475 189.04 487.755 190.16 ;
      RECT 483.555 189.04 483.835 205.605 ;
      RECT 336.325 189.04 336.605 252.385 ;
      RECT 335.765 189.04 336.045 252.385 ;
      RECT 335.205 189.04 335.485 252.385 ;
      RECT 334.645 189.04 334.925 252.385 ;
      RECT 334.085 189.04 334.365 252.385 ;
      RECT 333.525 189.04 333.805 252.385 ;
      RECT 332.965 189.04 333.245 252.385 ;
      RECT 332.405 189.04 332.685 252.385 ;
    LAYER M2 SPACING 0.28 ;
      RECT 12958.815 188.86 18490.46 8613.565 ;
      RECT 18485.135 187.44 18490.46 8613.565 ;
      RECT 18357.215 187.44 18480.095 8613.565 ;
      RECT 18353.575 187.44 18356.095 8613.565 ;
      RECT 18349.935 187.44 18352.455 8613.565 ;
      RECT 18346.295 187.44 18348.815 8613.565 ;
      RECT 18342.655 187.44 18345.175 8613.565 ;
      RECT 18339.015 187.44 18341.535 8613.565 ;
      RECT 18279.935 187.44 18337.895 8613.565 ;
      RECT 18276.015 187.44 18278.815 8613.565 ;
      RECT 18272.095 187.44 18274.895 8613.565 ;
      RECT 18268.175 187.44 18270.975 8613.565 ;
      RECT 18264.255 187.44 18267.055 8613.565 ;
      RECT 18217.215 187.44 18263.135 8613.565 ;
      RECT 18213.575 187.44 18216.095 8613.565 ;
      RECT 18209.935 187.44 18212.455 8613.565 ;
      RECT 18206.295 187.44 18208.815 8613.565 ;
      RECT 18202.655 187.44 18205.175 8613.565 ;
      RECT 18199.015 187.44 18201.535 8613.565 ;
      RECT 18139.935 187.44 18197.895 8613.565 ;
      RECT 18136.015 187.44 18138.815 8613.565 ;
      RECT 18132.095 187.44 18134.895 8613.565 ;
      RECT 18128.175 187.44 18130.975 8613.565 ;
      RECT 18124.255 187.44 18127.055 8613.565 ;
      RECT 18077.215 187.44 18123.135 8613.565 ;
      RECT 18073.575 187.44 18076.095 8613.565 ;
      RECT 18069.935 187.44 18072.455 8613.565 ;
      RECT 18066.295 187.44 18068.815 8613.565 ;
      RECT 18062.655 187.44 18065.175 8613.565 ;
      RECT 18059.015 187.44 18061.535 8613.565 ;
      RECT 17999.935 187.44 18057.895 8613.565 ;
      RECT 17996.015 187.44 17998.815 8613.565 ;
      RECT 17992.095 187.44 17994.895 8613.565 ;
      RECT 17988.175 187.44 17990.975 8613.565 ;
      RECT 17984.255 187.44 17987.055 8613.565 ;
      RECT 17937.215 187.44 17983.135 8613.565 ;
      RECT 17933.575 187.44 17936.095 8613.565 ;
      RECT 17929.935 187.44 17932.455 8613.565 ;
      RECT 17926.295 187.44 17928.815 8613.565 ;
      RECT 17922.655 187.44 17925.175 8613.565 ;
      RECT 17919.015 187.44 17921.535 8613.565 ;
      RECT 17859.935 187.44 17917.895 8613.565 ;
      RECT 17856.015 187.44 17858.815 8613.565 ;
      RECT 17852.095 187.44 17854.895 8613.565 ;
      RECT 17848.175 187.44 17850.975 8613.565 ;
      RECT 17844.255 187.44 17847.055 8613.565 ;
      RECT 17797.215 187.44 17843.135 8613.565 ;
      RECT 17793.575 187.44 17796.095 8613.565 ;
      RECT 17789.935 187.44 17792.455 8613.565 ;
      RECT 17786.295 187.44 17788.815 8613.565 ;
      RECT 17782.655 187.44 17785.175 8613.565 ;
      RECT 17779.015 187.44 17781.535 8613.565 ;
      RECT 17719.935 187.44 17777.895 8613.565 ;
      RECT 17716.015 187.44 17718.815 8613.565 ;
      RECT 17712.095 187.44 17714.895 8613.565 ;
      RECT 17708.175 187.44 17710.975 8613.565 ;
      RECT 17704.255 187.44 17707.055 8613.565 ;
      RECT 17657.215 187.44 17703.135 8613.565 ;
      RECT 17653.575 187.44 17656.095 8613.565 ;
      RECT 17649.935 187.44 17652.455 8613.565 ;
      RECT 17646.295 187.44 17648.815 8613.565 ;
      RECT 17642.655 187.44 17645.175 8613.565 ;
      RECT 17639.015 187.44 17641.535 8613.565 ;
      RECT 17579.935 187.44 17637.895 8613.565 ;
      RECT 17576.015 187.44 17578.815 8613.565 ;
      RECT 17572.095 187.44 17574.895 8613.565 ;
      RECT 17568.175 187.44 17570.975 8613.565 ;
      RECT 17564.255 187.44 17567.055 8613.565 ;
      RECT 17517.215 187.44 17563.135 8613.565 ;
      RECT 17513.575 187.44 17516.095 8613.565 ;
      RECT 17509.935 187.44 17512.455 8613.565 ;
      RECT 17506.295 187.44 17508.815 8613.565 ;
      RECT 17502.655 187.44 17505.175 8613.565 ;
      RECT 17499.015 187.44 17501.535 8613.565 ;
      RECT 17439.935 187.44 17497.895 8613.565 ;
      RECT 17436.015 187.44 17438.815 8613.565 ;
      RECT 17432.095 187.44 17434.895 8613.565 ;
      RECT 17428.175 187.44 17430.975 8613.565 ;
      RECT 17424.255 187.44 17427.055 8613.565 ;
      RECT 17377.215 187.44 17423.135 8613.565 ;
      RECT 17373.575 187.44 17376.095 8613.565 ;
      RECT 17369.935 187.44 17372.455 8613.565 ;
      RECT 17366.295 187.44 17368.815 8613.565 ;
      RECT 17362.655 187.44 17365.175 8613.565 ;
      RECT 17359.015 187.44 17361.535 8613.565 ;
      RECT 17299.935 187.44 17357.895 8613.565 ;
      RECT 17296.015 187.44 17298.815 8613.565 ;
      RECT 17292.095 187.44 17294.895 8613.565 ;
      RECT 17288.175 187.44 17290.975 8613.565 ;
      RECT 17284.255 187.44 17287.055 8613.565 ;
      RECT 17237.215 187.44 17283.135 8613.565 ;
      RECT 17233.575 187.44 17236.095 8613.565 ;
      RECT 17229.935 187.44 17232.455 8613.565 ;
      RECT 17226.295 187.44 17228.815 8613.565 ;
      RECT 17222.655 187.44 17225.175 8613.565 ;
      RECT 17219.015 187.44 17221.535 8613.565 ;
      RECT 17159.935 187.44 17217.895 8613.565 ;
      RECT 17156.015 187.44 17158.815 8613.565 ;
      RECT 17152.095 187.44 17154.895 8613.565 ;
      RECT 17148.175 187.44 17150.975 8613.565 ;
      RECT 17144.255 187.44 17147.055 8613.565 ;
      RECT 17097.215 187.44 17143.135 8613.565 ;
      RECT 17093.575 187.44 17096.095 8613.565 ;
      RECT 17089.935 187.44 17092.455 8613.565 ;
      RECT 17086.295 187.44 17088.815 8613.565 ;
      RECT 17082.655 187.44 17085.175 8613.565 ;
      RECT 17079.015 187.44 17081.535 8613.565 ;
      RECT 17019.935 187.44 17077.895 8613.565 ;
      RECT 17016.015 187.44 17018.815 8613.565 ;
      RECT 17012.095 187.44 17014.895 8613.565 ;
      RECT 17008.175 187.44 17010.975 8613.565 ;
      RECT 17004.255 187.44 17007.055 8613.565 ;
      RECT 16957.215 187.44 17003.135 8613.565 ;
      RECT 16953.575 187.44 16956.095 8613.565 ;
      RECT 16949.935 187.44 16952.455 8613.565 ;
      RECT 16946.295 187.44 16948.815 8613.565 ;
      RECT 16942.655 187.44 16945.175 8613.565 ;
      RECT 16939.015 187.44 16941.535 8613.565 ;
      RECT 16879.935 187.44 16937.895 8613.565 ;
      RECT 16876.015 187.44 16878.815 8613.565 ;
      RECT 16872.095 187.44 16874.895 8613.565 ;
      RECT 16868.175 187.44 16870.975 8613.565 ;
      RECT 16864.255 187.44 16867.055 8613.565 ;
      RECT 16817.215 187.44 16863.135 8613.565 ;
      RECT 16813.575 187.44 16816.095 8613.565 ;
      RECT 16809.935 187.44 16812.455 8613.565 ;
      RECT 16806.295 187.44 16808.815 8613.565 ;
      RECT 16802.655 187.44 16805.175 8613.565 ;
      RECT 16799.015 187.44 16801.535 8613.565 ;
      RECT 16739.935 187.44 16797.895 8613.565 ;
      RECT 16736.015 187.44 16738.815 8613.565 ;
      RECT 16732.095 187.44 16734.895 8613.565 ;
      RECT 16728.175 187.44 16730.975 8613.565 ;
      RECT 16724.255 187.44 16727.055 8613.565 ;
      RECT 16677.215 187.44 16723.135 8613.565 ;
      RECT 16673.575 187.44 16676.095 8613.565 ;
      RECT 16669.935 187.44 16672.455 8613.565 ;
      RECT 16666.295 187.44 16668.815 8613.565 ;
      RECT 16662.655 187.44 16665.175 8613.565 ;
      RECT 16659.015 187.44 16661.535 8613.565 ;
      RECT 16599.935 187.44 16657.895 8613.565 ;
      RECT 16596.015 187.44 16598.815 8613.565 ;
      RECT 16592.095 187.44 16594.895 8613.565 ;
      RECT 16588.175 187.44 16590.975 8613.565 ;
      RECT 16584.255 187.44 16587.055 8613.565 ;
      RECT 16537.215 187.44 16583.135 8613.565 ;
      RECT 16533.575 187.44 16536.095 8613.565 ;
      RECT 16529.935 187.44 16532.455 8613.565 ;
      RECT 16526.295 187.44 16528.815 8613.565 ;
      RECT 16522.655 187.44 16525.175 8613.565 ;
      RECT 16519.015 187.44 16521.535 8613.565 ;
      RECT 16459.935 187.44 16517.895 8613.565 ;
      RECT 16456.015 187.44 16458.815 8613.565 ;
      RECT 16452.095 187.44 16454.895 8613.565 ;
      RECT 16448.175 187.44 16450.975 8613.565 ;
      RECT 16444.255 187.44 16447.055 8613.565 ;
      RECT 16397.215 187.44 16443.135 8613.565 ;
      RECT 16393.575 187.44 16396.095 8613.565 ;
      RECT 16389.935 187.44 16392.455 8613.565 ;
      RECT 16386.295 187.44 16388.815 8613.565 ;
      RECT 16382.655 187.44 16385.175 8613.565 ;
      RECT 16379.015 187.44 16381.535 8613.565 ;
      RECT 16319.935 187.44 16377.895 8613.565 ;
      RECT 16316.015 187.44 16318.815 8613.565 ;
      RECT 16312.095 187.44 16314.895 8613.565 ;
      RECT 16308.175 187.44 16310.975 8613.565 ;
      RECT 16304.255 187.44 16307.055 8613.565 ;
      RECT 16257.215 187.44 16303.135 8613.565 ;
      RECT 16253.575 187.44 16256.095 8613.565 ;
      RECT 16249.935 187.44 16252.455 8613.565 ;
      RECT 16246.295 187.44 16248.815 8613.565 ;
      RECT 16242.655 187.44 16245.175 8613.565 ;
      RECT 16239.015 187.44 16241.535 8613.565 ;
      RECT 16179.935 187.44 16237.895 8613.565 ;
      RECT 16176.015 187.44 16178.815 8613.565 ;
      RECT 16172.095 187.44 16174.895 8613.565 ;
      RECT 16168.175 187.44 16170.975 8613.565 ;
      RECT 16164.255 187.44 16167.055 8613.565 ;
      RECT 16117.215 187.44 16163.135 8613.565 ;
      RECT 16113.575 187.44 16116.095 8613.565 ;
      RECT 16109.935 187.44 16112.455 8613.565 ;
      RECT 16106.295 187.44 16108.815 8613.565 ;
      RECT 16102.655 187.44 16105.175 8613.565 ;
      RECT 16099.015 187.44 16101.535 8613.565 ;
      RECT 16039.935 187.44 16097.895 8613.565 ;
      RECT 16036.015 187.44 16038.815 8613.565 ;
      RECT 16032.095 187.44 16034.895 8613.565 ;
      RECT 16028.175 187.44 16030.975 8613.565 ;
      RECT 16024.255 187.44 16027.055 8613.565 ;
      RECT 15977.215 187.44 16023.135 8613.565 ;
      RECT 15973.575 187.44 15976.095 8613.565 ;
      RECT 15969.935 187.44 15972.455 8613.565 ;
      RECT 15966.295 187.44 15968.815 8613.565 ;
      RECT 15962.655 187.44 15965.175 8613.565 ;
      RECT 15959.015 187.44 15961.535 8613.565 ;
      RECT 15899.935 187.44 15957.895 8613.565 ;
      RECT 15896.015 187.44 15898.815 8613.565 ;
      RECT 15892.095 187.44 15894.895 8613.565 ;
      RECT 15888.175 187.44 15890.975 8613.565 ;
      RECT 15884.255 187.44 15887.055 8613.565 ;
      RECT 15837.215 187.44 15883.135 8613.565 ;
      RECT 15833.575 187.44 15836.095 8613.565 ;
      RECT 15829.935 187.44 15832.455 8613.565 ;
      RECT 15826.295 187.44 15828.815 8613.565 ;
      RECT 15822.655 187.44 15825.175 8613.565 ;
      RECT 15819.015 187.44 15821.535 8613.565 ;
      RECT 15759.935 187.44 15817.895 8613.565 ;
      RECT 15756.015 187.44 15758.815 8613.565 ;
      RECT 15752.095 187.44 15754.895 8613.565 ;
      RECT 15748.175 187.44 15750.975 8613.565 ;
      RECT 15744.255 187.44 15747.055 8613.565 ;
      RECT 15697.215 187.44 15743.135 8613.565 ;
      RECT 15693.575 187.44 15696.095 8613.565 ;
      RECT 15689.935 187.44 15692.455 8613.565 ;
      RECT 15686.295 187.44 15688.815 8613.565 ;
      RECT 15682.655 187.44 15685.175 8613.565 ;
      RECT 15679.015 187.44 15681.535 8613.565 ;
      RECT 15619.935 187.44 15677.895 8613.565 ;
      RECT 15616.015 187.44 15618.815 8613.565 ;
      RECT 15612.095 187.44 15614.895 8613.565 ;
      RECT 15608.175 187.44 15610.975 8613.565 ;
      RECT 15604.255 187.44 15607.055 8613.565 ;
      RECT 15557.215 187.44 15603.135 8613.565 ;
      RECT 15553.575 187.44 15556.095 8613.565 ;
      RECT 15549.935 187.44 15552.455 8613.565 ;
      RECT 15546.295 187.44 15548.815 8613.565 ;
      RECT 15542.655 187.44 15545.175 8613.565 ;
      RECT 15539.015 187.44 15541.535 8613.565 ;
      RECT 15479.935 187.44 15537.895 8613.565 ;
      RECT 15476.015 187.44 15478.815 8613.565 ;
      RECT 15472.095 187.44 15474.895 8613.565 ;
      RECT 15468.175 187.44 15470.975 8613.565 ;
      RECT 15464.255 187.44 15467.055 8613.565 ;
      RECT 15417.215 187.44 15463.135 8613.565 ;
      RECT 15413.575 187.44 15416.095 8613.565 ;
      RECT 15409.935 187.44 15412.455 8613.565 ;
      RECT 15406.295 187.44 15408.815 8613.565 ;
      RECT 15402.655 187.44 15405.175 8613.565 ;
      RECT 15399.015 187.44 15401.535 8613.565 ;
      RECT 15339.935 187.44 15397.895 8613.565 ;
      RECT 15336.015 187.44 15338.815 8613.565 ;
      RECT 15332.095 187.44 15334.895 8613.565 ;
      RECT 15328.175 187.44 15330.975 8613.565 ;
      RECT 15324.255 187.44 15327.055 8613.565 ;
      RECT 15277.215 187.44 15323.135 8613.565 ;
      RECT 15273.575 187.44 15276.095 8613.565 ;
      RECT 15269.935 187.44 15272.455 8613.565 ;
      RECT 15266.295 187.44 15268.815 8613.565 ;
      RECT 15262.655 187.44 15265.175 8613.565 ;
      RECT 15259.015 187.44 15261.535 8613.565 ;
      RECT 15199.935 187.44 15257.895 8613.565 ;
      RECT 15196.015 187.44 15198.815 8613.565 ;
      RECT 15192.095 187.44 15194.895 8613.565 ;
      RECT 15188.175 187.44 15190.975 8613.565 ;
      RECT 15184.255 187.44 15187.055 8613.565 ;
      RECT 15137.215 187.44 15183.135 8613.565 ;
      RECT 15133.575 187.44 15136.095 8613.565 ;
      RECT 15129.935 187.44 15132.455 8613.565 ;
      RECT 15126.295 187.44 15128.815 8613.565 ;
      RECT 15122.655 187.44 15125.175 8613.565 ;
      RECT 15119.015 187.44 15121.535 8613.565 ;
      RECT 15059.935 187.44 15117.895 8613.565 ;
      RECT 15056.015 187.44 15058.815 8613.565 ;
      RECT 15052.095 187.44 15054.895 8613.565 ;
      RECT 15048.175 187.44 15050.975 8613.565 ;
      RECT 15044.255 187.44 15047.055 8613.565 ;
      RECT 14997.215 187.44 15043.135 8613.565 ;
      RECT 14993.575 187.44 14996.095 8613.565 ;
      RECT 14989.935 187.44 14992.455 8613.565 ;
      RECT 14986.295 187.44 14988.815 8613.565 ;
      RECT 14982.655 187.44 14985.175 8613.565 ;
      RECT 14979.015 187.44 14981.535 8613.565 ;
      RECT 14919.935 187.44 14977.895 8613.565 ;
      RECT 14916.015 187.44 14918.815 8613.565 ;
      RECT 14912.095 187.44 14914.895 8613.565 ;
      RECT 14908.175 187.44 14910.975 8613.565 ;
      RECT 14904.255 187.44 14907.055 8613.565 ;
      RECT 14857.215 187.44 14903.135 8613.565 ;
      RECT 14853.575 187.44 14856.095 8613.565 ;
      RECT 14849.935 187.44 14852.455 8613.565 ;
      RECT 14846.295 187.44 14848.815 8613.565 ;
      RECT 14842.655 187.44 14845.175 8613.565 ;
      RECT 14839.015 187.44 14841.535 8613.565 ;
      RECT 14779.935 187.44 14837.895 8613.565 ;
      RECT 14776.015 187.44 14778.815 8613.565 ;
      RECT 14772.095 187.44 14774.895 8613.565 ;
      RECT 14768.175 187.44 14770.975 8613.565 ;
      RECT 14764.255 187.44 14767.055 8613.565 ;
      RECT 14717.215 187.44 14763.135 8613.565 ;
      RECT 14713.575 187.44 14716.095 8613.565 ;
      RECT 14709.935 187.44 14712.455 8613.565 ;
      RECT 14706.295 187.44 14708.815 8613.565 ;
      RECT 14702.655 187.44 14705.175 8613.565 ;
      RECT 14699.015 187.44 14701.535 8613.565 ;
      RECT 14639.935 187.44 14697.895 8613.565 ;
      RECT 14636.015 187.44 14638.815 8613.565 ;
      RECT 14632.095 187.44 14634.895 8613.565 ;
      RECT 14628.175 187.44 14630.975 8613.565 ;
      RECT 14624.255 187.44 14627.055 8613.565 ;
      RECT 14577.215 187.44 14623.135 8613.565 ;
      RECT 14573.575 187.44 14576.095 8613.565 ;
      RECT 14569.935 187.44 14572.455 8613.565 ;
      RECT 14566.295 187.44 14568.815 8613.565 ;
      RECT 14562.655 187.44 14565.175 8613.565 ;
      RECT 14559.015 187.44 14561.535 8613.565 ;
      RECT 14499.935 187.44 14557.895 8613.565 ;
      RECT 14496.015 187.44 14498.815 8613.565 ;
      RECT 14492.095 187.44 14494.895 8613.565 ;
      RECT 14488.175 187.44 14490.975 8613.565 ;
      RECT 14484.255 187.44 14487.055 8613.565 ;
      RECT 14437.215 187.44 14483.135 8613.565 ;
      RECT 14433.575 187.44 14436.095 8613.565 ;
      RECT 14429.935 187.44 14432.455 8613.565 ;
      RECT 14426.295 187.44 14428.815 8613.565 ;
      RECT 14422.655 187.44 14425.175 8613.565 ;
      RECT 14419.015 187.44 14421.535 8613.565 ;
      RECT 14359.935 187.44 14417.895 8613.565 ;
      RECT 14356.015 187.44 14358.815 8613.565 ;
      RECT 14352.095 187.44 14354.895 8613.565 ;
      RECT 14348.175 187.44 14350.975 8613.565 ;
      RECT 14344.255 187.44 14347.055 8613.565 ;
      RECT 14297.215 187.44 14343.135 8613.565 ;
      RECT 14293.575 187.44 14296.095 8613.565 ;
      RECT 14289.935 187.44 14292.455 8613.565 ;
      RECT 14286.295 187.44 14288.815 8613.565 ;
      RECT 14282.655 187.44 14285.175 8613.565 ;
      RECT 14279.015 187.44 14281.535 8613.565 ;
      RECT 14219.935 187.44 14277.895 8613.565 ;
      RECT 14216.015 187.44 14218.815 8613.565 ;
      RECT 14212.095 187.44 14214.895 8613.565 ;
      RECT 14208.175 187.44 14210.975 8613.565 ;
      RECT 14204.255 187.44 14207.055 8613.565 ;
      RECT 14157.215 187.44 14203.135 8613.565 ;
      RECT 14153.575 187.44 14156.095 8613.565 ;
      RECT 14149.935 187.44 14152.455 8613.565 ;
      RECT 14146.295 187.44 14148.815 8613.565 ;
      RECT 14142.655 187.44 14145.175 8613.565 ;
      RECT 14139.015 187.44 14141.535 8613.565 ;
      RECT 14079.935 187.44 14137.895 8613.565 ;
      RECT 14076.015 187.44 14078.815 8613.565 ;
      RECT 14072.095 187.44 14074.895 8613.565 ;
      RECT 14068.175 187.44 14070.975 8613.565 ;
      RECT 14064.255 187.44 14067.055 8613.565 ;
      RECT 14017.215 187.44 14063.135 8613.565 ;
      RECT 14013.575 187.44 14016.095 8613.565 ;
      RECT 14009.935 187.44 14012.455 8613.565 ;
      RECT 14006.295 187.44 14008.815 8613.565 ;
      RECT 14002.655 187.44 14005.175 8613.565 ;
      RECT 13999.015 187.44 14001.535 8613.565 ;
      RECT 13939.935 187.44 13997.895 8613.565 ;
      RECT 13936.015 187.44 13938.815 8613.565 ;
      RECT 13932.095 187.44 13934.895 8613.565 ;
      RECT 13928.175 187.44 13930.975 8613.565 ;
      RECT 13924.255 187.44 13927.055 8613.565 ;
      RECT 13877.215 187.44 13923.135 8613.565 ;
      RECT 13873.575 187.44 13876.095 8613.565 ;
      RECT 13869.935 187.44 13872.455 8613.565 ;
      RECT 13866.295 187.44 13868.815 8613.565 ;
      RECT 13862.655 187.44 13865.175 8613.565 ;
      RECT 13859.015 187.44 13861.535 8613.565 ;
      RECT 13799.935 187.44 13857.895 8613.565 ;
      RECT 13796.015 187.44 13798.815 8613.565 ;
      RECT 13792.095 187.44 13794.895 8613.565 ;
      RECT 13788.175 187.44 13790.975 8613.565 ;
      RECT 13784.255 187.44 13787.055 8613.565 ;
      RECT 13737.215 187.44 13783.135 8613.565 ;
      RECT 13733.575 187.44 13736.095 8613.565 ;
      RECT 13729.935 187.44 13732.455 8613.565 ;
      RECT 13726.295 187.44 13728.815 8613.565 ;
      RECT 13722.655 187.44 13725.175 8613.565 ;
      RECT 13719.015 187.44 13721.535 8613.565 ;
      RECT 13659.935 187.44 13717.895 8613.565 ;
      RECT 13656.015 187.44 13658.815 8613.565 ;
      RECT 13652.095 187.44 13654.895 8613.565 ;
      RECT 13648.175 187.44 13650.975 8613.565 ;
      RECT 13644.255 187.44 13647.055 8613.565 ;
      RECT 13597.215 187.44 13643.135 8613.565 ;
      RECT 13593.575 187.44 13596.095 8613.565 ;
      RECT 13589.935 187.44 13592.455 8613.565 ;
      RECT 13586.295 187.44 13588.815 8613.565 ;
      RECT 13582.655 187.44 13585.175 8613.565 ;
      RECT 13579.015 187.44 13581.535 8613.565 ;
      RECT 13519.935 187.44 13577.895 8613.565 ;
      RECT 13516.015 187.44 13518.815 8613.565 ;
      RECT 13512.095 187.44 13514.895 8613.565 ;
      RECT 13508.175 187.44 13510.975 8613.565 ;
      RECT 13504.255 187.44 13507.055 8613.565 ;
      RECT 13457.215 187.44 13503.135 8613.565 ;
      RECT 13453.575 187.44 13456.095 8613.565 ;
      RECT 13449.935 187.44 13452.455 8613.565 ;
      RECT 13446.295 187.44 13448.815 8613.565 ;
      RECT 13442.655 187.44 13445.175 8613.565 ;
      RECT 13439.015 187.44 13441.535 8613.565 ;
      RECT 13379.935 187.44 13437.895 8613.565 ;
      RECT 13376.015 187.44 13378.815 8613.565 ;
      RECT 13372.095 187.44 13374.895 8613.565 ;
      RECT 13368.175 187.44 13370.975 8613.565 ;
      RECT 13364.255 187.44 13367.055 8613.565 ;
      RECT 13317.215 187.44 13363.135 8613.565 ;
      RECT 13313.575 187.44 13316.095 8613.565 ;
      RECT 13309.935 187.44 13312.455 8613.565 ;
      RECT 13306.295 187.44 13308.815 8613.565 ;
      RECT 13302.655 187.44 13305.175 8613.565 ;
      RECT 13299.015 187.44 13301.535 8613.565 ;
      RECT 13239.935 187.44 13297.895 8613.565 ;
      RECT 13236.015 187.44 13238.815 8613.565 ;
      RECT 13232.095 187.44 13234.895 8613.565 ;
      RECT 13228.175 187.44 13230.975 8613.565 ;
      RECT 13224.255 187.44 13227.055 8613.565 ;
      RECT 13177.215 187.44 13223.135 8613.565 ;
      RECT 13173.575 187.44 13176.095 8613.565 ;
      RECT 13169.935 187.44 13172.455 8613.565 ;
      RECT 13166.295 187.44 13168.815 8613.565 ;
      RECT 13162.655 187.44 13165.175 8613.565 ;
      RECT 13159.015 187.44 13161.535 8613.565 ;
      RECT 13099.935 187.44 13157.895 8613.565 ;
      RECT 13096.015 187.44 13098.815 8613.565 ;
      RECT 13092.095 187.44 13094.895 8613.565 ;
      RECT 13088.175 187.44 13090.975 8613.565 ;
      RECT 13084.255 187.44 13087.055 8613.565 ;
      RECT 13037.215 187.44 13083.135 8613.565 ;
      RECT 13033.575 187.44 13036.095 8613.565 ;
      RECT 13029.935 187.44 13032.455 8613.565 ;
      RECT 13026.295 187.44 13028.815 8613.565 ;
      RECT 13022.655 187.44 13025.175 8613.565 ;
      RECT 13019.015 187.44 13021.535 8613.565 ;
      RECT 12959.935 187.44 13017.895 8613.565 ;
      RECT 326.66 188.86 12958.815 8613.565 ;
      RECT 12956.015 187.44 12958.815 8613.565 ;
      RECT 12952.095 187.44 12954.895 8613.565 ;
      RECT 12948.175 187.44 12950.975 8613.565 ;
      RECT 12944.255 187.44 12947.055 8613.565 ;
      RECT 12897.215 187.44 12943.135 8613.565 ;
      RECT 12893.575 187.44 12896.095 8613.565 ;
      RECT 12889.935 187.44 12892.455 8613.565 ;
      RECT 12886.295 187.44 12888.815 8613.565 ;
      RECT 12882.655 187.44 12885.175 8613.565 ;
      RECT 12879.015 187.44 12881.535 8613.565 ;
      RECT 12819.935 187.44 12877.895 8613.565 ;
      RECT 12816.015 187.44 12818.815 8613.565 ;
      RECT 12812.095 187.44 12814.895 8613.565 ;
      RECT 12808.175 187.44 12810.975 8613.565 ;
      RECT 12804.255 187.44 12807.055 8613.565 ;
      RECT 12757.215 187.44 12803.135 8613.565 ;
      RECT 12753.575 187.44 12756.095 8613.565 ;
      RECT 12749.935 187.44 12752.455 8613.565 ;
      RECT 12746.295 187.44 12748.815 8613.565 ;
      RECT 12742.655 187.44 12745.175 8613.565 ;
      RECT 12739.015 187.44 12741.535 8613.565 ;
      RECT 12679.935 187.44 12737.895 8613.565 ;
      RECT 12676.015 187.44 12678.815 8613.565 ;
      RECT 12672.095 187.44 12674.895 8613.565 ;
      RECT 12668.175 187.44 12670.975 8613.565 ;
      RECT 12664.255 187.44 12667.055 8613.565 ;
      RECT 12617.215 187.44 12663.135 8613.565 ;
      RECT 12613.575 187.44 12616.095 8613.565 ;
      RECT 12609.935 187.44 12612.455 8613.565 ;
      RECT 12606.295 187.44 12608.815 8613.565 ;
      RECT 12602.655 187.44 12605.175 8613.565 ;
      RECT 12599.015 187.44 12601.535 8613.565 ;
      RECT 12539.935 187.44 12597.895 8613.565 ;
      RECT 12536.015 187.44 12538.815 8613.565 ;
      RECT 12532.095 187.44 12534.895 8613.565 ;
      RECT 12528.175 187.44 12530.975 8613.565 ;
      RECT 12524.255 187.44 12527.055 8613.565 ;
      RECT 12477.215 187.44 12523.135 8613.565 ;
      RECT 12473.575 187.44 12476.095 8613.565 ;
      RECT 12469.935 187.44 12472.455 8613.565 ;
      RECT 12466.295 187.44 12468.815 8613.565 ;
      RECT 12462.655 187.44 12465.175 8613.565 ;
      RECT 12459.015 187.44 12461.535 8613.565 ;
      RECT 12399.935 187.44 12457.895 8613.565 ;
      RECT 12396.015 187.44 12398.815 8613.565 ;
      RECT 12392.095 187.44 12394.895 8613.565 ;
      RECT 12388.175 187.44 12390.975 8613.565 ;
      RECT 12384.255 187.44 12387.055 8613.565 ;
      RECT 12337.215 187.44 12383.135 8613.565 ;
      RECT 12333.575 187.44 12336.095 8613.565 ;
      RECT 12329.935 187.44 12332.455 8613.565 ;
      RECT 12326.295 187.44 12328.815 8613.565 ;
      RECT 12322.655 187.44 12325.175 8613.565 ;
      RECT 12319.015 187.44 12321.535 8613.565 ;
      RECT 12259.935 187.44 12317.895 8613.565 ;
      RECT 12256.015 187.44 12258.815 8613.565 ;
      RECT 12252.095 187.44 12254.895 8613.565 ;
      RECT 12248.175 187.44 12250.975 8613.565 ;
      RECT 12244.255 187.44 12247.055 8613.565 ;
      RECT 12197.215 187.44 12243.135 8613.565 ;
      RECT 12193.575 187.44 12196.095 8613.565 ;
      RECT 12189.935 187.44 12192.455 8613.565 ;
      RECT 12186.295 187.44 12188.815 8613.565 ;
      RECT 12182.655 187.44 12185.175 8613.565 ;
      RECT 12179.015 187.44 12181.535 8613.565 ;
      RECT 12119.935 187.44 12177.895 8613.565 ;
      RECT 12116.015 187.44 12118.815 8613.565 ;
      RECT 12112.095 187.44 12114.895 8613.565 ;
      RECT 12108.175 187.44 12110.975 8613.565 ;
      RECT 12104.255 187.44 12107.055 8613.565 ;
      RECT 12057.215 187.44 12103.135 8613.565 ;
      RECT 12053.575 187.44 12056.095 8613.565 ;
      RECT 12049.935 187.44 12052.455 8613.565 ;
      RECT 12046.295 187.44 12048.815 8613.565 ;
      RECT 12042.655 187.44 12045.175 8613.565 ;
      RECT 12039.015 187.44 12041.535 8613.565 ;
      RECT 11979.935 187.44 12037.895 8613.565 ;
      RECT 11976.015 187.44 11978.815 8613.565 ;
      RECT 11972.095 187.44 11974.895 8613.565 ;
      RECT 11968.175 187.44 11970.975 8613.565 ;
      RECT 11964.255 187.44 11967.055 8613.565 ;
      RECT 11917.215 187.44 11963.135 8613.565 ;
      RECT 11913.575 187.44 11916.095 8613.565 ;
      RECT 11909.935 187.44 11912.455 8613.565 ;
      RECT 11906.295 187.44 11908.815 8613.565 ;
      RECT 11902.655 187.44 11905.175 8613.565 ;
      RECT 11899.015 187.44 11901.535 8613.565 ;
      RECT 11839.935 187.44 11897.895 8613.565 ;
      RECT 11836.015 187.44 11838.815 8613.565 ;
      RECT 11832.095 187.44 11834.895 8613.565 ;
      RECT 11828.175 187.44 11830.975 8613.565 ;
      RECT 11824.255 187.44 11827.055 8613.565 ;
      RECT 11777.215 187.44 11823.135 8613.565 ;
      RECT 11773.575 187.44 11776.095 8613.565 ;
      RECT 11769.935 187.44 11772.455 8613.565 ;
      RECT 11766.295 187.44 11768.815 8613.565 ;
      RECT 11762.655 187.44 11765.175 8613.565 ;
      RECT 11759.015 187.44 11761.535 8613.565 ;
      RECT 11699.935 187.44 11757.895 8613.565 ;
      RECT 11696.015 187.44 11698.815 8613.565 ;
      RECT 11692.095 187.44 11694.895 8613.565 ;
      RECT 11688.175 187.44 11690.975 8613.565 ;
      RECT 11684.255 187.44 11687.055 8613.565 ;
      RECT 11637.215 187.44 11683.135 8613.565 ;
      RECT 11633.575 187.44 11636.095 8613.565 ;
      RECT 11629.935 187.44 11632.455 8613.565 ;
      RECT 11626.295 187.44 11628.815 8613.565 ;
      RECT 11622.655 187.44 11625.175 8613.565 ;
      RECT 11619.015 187.44 11621.535 8613.565 ;
      RECT 11559.935 187.44 11617.895 8613.565 ;
      RECT 11556.015 187.44 11558.815 8613.565 ;
      RECT 11552.095 187.44 11554.895 8613.565 ;
      RECT 11548.175 187.44 11550.975 8613.565 ;
      RECT 11544.255 187.44 11547.055 8613.565 ;
      RECT 11497.215 187.44 11543.135 8613.565 ;
      RECT 11493.575 187.44 11496.095 8613.565 ;
      RECT 11489.935 187.44 11492.455 8613.565 ;
      RECT 11486.295 187.44 11488.815 8613.565 ;
      RECT 11482.655 187.44 11485.175 8613.565 ;
      RECT 11479.015 187.44 11481.535 8613.565 ;
      RECT 11419.935 187.44 11477.895 8613.565 ;
      RECT 11416.015 187.44 11418.815 8613.565 ;
      RECT 11412.095 187.44 11414.895 8613.565 ;
      RECT 11408.175 187.44 11410.975 8613.565 ;
      RECT 11404.255 187.44 11407.055 8613.565 ;
      RECT 11357.215 187.44 11403.135 8613.565 ;
      RECT 11353.575 187.44 11356.095 8613.565 ;
      RECT 11349.935 187.44 11352.455 8613.565 ;
      RECT 11346.295 187.44 11348.815 8613.565 ;
      RECT 11342.655 187.44 11345.175 8613.565 ;
      RECT 11339.015 187.44 11341.535 8613.565 ;
      RECT 11279.935 187.44 11337.895 8613.565 ;
      RECT 11276.015 187.44 11278.815 8613.565 ;
      RECT 11272.095 187.44 11274.895 8613.565 ;
      RECT 11268.175 187.44 11270.975 8613.565 ;
      RECT 11264.255 187.44 11267.055 8613.565 ;
      RECT 11217.215 187.44 11263.135 8613.565 ;
      RECT 11213.575 187.44 11216.095 8613.565 ;
      RECT 11209.935 187.44 11212.455 8613.565 ;
      RECT 11206.295 187.44 11208.815 8613.565 ;
      RECT 11202.655 187.44 11205.175 8613.565 ;
      RECT 11199.015 187.44 11201.535 8613.565 ;
      RECT 11139.935 187.44 11197.895 8613.565 ;
      RECT 11136.015 187.44 11138.815 8613.565 ;
      RECT 11132.095 187.44 11134.895 8613.565 ;
      RECT 11128.175 187.44 11130.975 8613.565 ;
      RECT 11124.255 187.44 11127.055 8613.565 ;
      RECT 11077.215 187.44 11123.135 8613.565 ;
      RECT 11073.575 187.44 11076.095 8613.565 ;
      RECT 11069.935 187.44 11072.455 8613.565 ;
      RECT 11066.295 187.44 11068.815 8613.565 ;
      RECT 11062.655 187.44 11065.175 8613.565 ;
      RECT 11059.015 187.44 11061.535 8613.565 ;
      RECT 10999.935 187.44 11057.895 8613.565 ;
      RECT 10996.015 187.44 10998.815 8613.565 ;
      RECT 10992.095 187.44 10994.895 8613.565 ;
      RECT 10988.175 187.44 10990.975 8613.565 ;
      RECT 10984.255 187.44 10987.055 8613.565 ;
      RECT 10937.215 187.44 10983.135 8613.565 ;
      RECT 10933.575 187.44 10936.095 8613.565 ;
      RECT 10929.935 187.44 10932.455 8613.565 ;
      RECT 10926.295 187.44 10928.815 8613.565 ;
      RECT 10922.655 187.44 10925.175 8613.565 ;
      RECT 10919.015 187.44 10921.535 8613.565 ;
      RECT 10859.935 187.44 10917.895 8613.565 ;
      RECT 10856.015 187.44 10858.815 8613.565 ;
      RECT 10852.095 187.44 10854.895 8613.565 ;
      RECT 10848.175 187.44 10850.975 8613.565 ;
      RECT 10844.255 187.44 10847.055 8613.565 ;
      RECT 10797.215 187.44 10843.135 8613.565 ;
      RECT 10793.575 187.44 10796.095 8613.565 ;
      RECT 10789.935 187.44 10792.455 8613.565 ;
      RECT 10786.295 187.44 10788.815 8613.565 ;
      RECT 10782.655 187.44 10785.175 8613.565 ;
      RECT 10779.015 187.44 10781.535 8613.565 ;
      RECT 10719.935 187.44 10777.895 8613.565 ;
      RECT 10716.015 187.44 10718.815 8613.565 ;
      RECT 10712.095 187.44 10714.895 8613.565 ;
      RECT 10708.175 187.44 10710.975 8613.565 ;
      RECT 10704.255 187.44 10707.055 8613.565 ;
      RECT 10657.215 187.44 10703.135 8613.565 ;
      RECT 10653.575 187.44 10656.095 8613.565 ;
      RECT 10649.935 187.44 10652.455 8613.565 ;
      RECT 10646.295 187.44 10648.815 8613.565 ;
      RECT 10642.655 187.44 10645.175 8613.565 ;
      RECT 10639.015 187.44 10641.535 8613.565 ;
      RECT 10579.935 187.44 10637.895 8613.565 ;
      RECT 10576.015 187.44 10578.815 8613.565 ;
      RECT 10572.095 187.44 10574.895 8613.565 ;
      RECT 10568.175 187.44 10570.975 8613.565 ;
      RECT 10564.255 187.44 10567.055 8613.565 ;
      RECT 10517.215 187.44 10563.135 8613.565 ;
      RECT 10513.575 187.44 10516.095 8613.565 ;
      RECT 10509.935 187.44 10512.455 8613.565 ;
      RECT 10506.295 187.44 10508.815 8613.565 ;
      RECT 10502.655 187.44 10505.175 8613.565 ;
      RECT 10499.015 187.44 10501.535 8613.565 ;
      RECT 10439.935 187.44 10497.895 8613.565 ;
      RECT 10436.015 187.44 10438.815 8613.565 ;
      RECT 10432.095 187.44 10434.895 8613.565 ;
      RECT 10428.175 187.44 10430.975 8613.565 ;
      RECT 10424.255 187.44 10427.055 8613.565 ;
      RECT 10377.215 187.44 10423.135 8613.565 ;
      RECT 10373.575 187.44 10376.095 8613.565 ;
      RECT 10369.935 187.44 10372.455 8613.565 ;
      RECT 10366.295 187.44 10368.815 8613.565 ;
      RECT 10362.655 187.44 10365.175 8613.565 ;
      RECT 10359.015 187.44 10361.535 8613.565 ;
      RECT 10299.935 187.44 10357.895 8613.565 ;
      RECT 10296.015 187.44 10298.815 8613.565 ;
      RECT 10292.095 187.44 10294.895 8613.565 ;
      RECT 10288.175 187.44 10290.975 8613.565 ;
      RECT 10284.255 187.44 10287.055 8613.565 ;
      RECT 10237.215 187.44 10283.135 8613.565 ;
      RECT 10233.575 187.44 10236.095 8613.565 ;
      RECT 10229.935 187.44 10232.455 8613.565 ;
      RECT 10226.295 187.44 10228.815 8613.565 ;
      RECT 10222.655 187.44 10225.175 8613.565 ;
      RECT 10219.015 187.44 10221.535 8613.565 ;
      RECT 10159.935 187.44 10217.895 8613.565 ;
      RECT 10156.015 187.44 10158.815 8613.565 ;
      RECT 10152.095 187.44 10154.895 8613.565 ;
      RECT 10148.175 187.44 10150.975 8613.565 ;
      RECT 10144.255 187.44 10147.055 8613.565 ;
      RECT 10097.215 187.44 10143.135 8613.565 ;
      RECT 10093.575 187.44 10096.095 8613.565 ;
      RECT 10089.935 187.44 10092.455 8613.565 ;
      RECT 10086.295 187.44 10088.815 8613.565 ;
      RECT 10082.655 187.44 10085.175 8613.565 ;
      RECT 10079.015 187.44 10081.535 8613.565 ;
      RECT 10019.935 187.44 10077.895 8613.565 ;
      RECT 10016.015 187.44 10018.815 8613.565 ;
      RECT 10012.095 187.44 10014.895 8613.565 ;
      RECT 10008.175 187.44 10010.975 8613.565 ;
      RECT 10004.255 187.44 10007.055 8613.565 ;
      RECT 9957.215 187.44 10003.135 8613.565 ;
      RECT 9953.575 187.44 9956.095 8613.565 ;
      RECT 9949.935 187.44 9952.455 8613.565 ;
      RECT 9946.295 187.44 9948.815 8613.565 ;
      RECT 9942.655 187.44 9945.175 8613.565 ;
      RECT 9939.015 187.44 9941.535 8613.565 ;
      RECT 9879.935 187.44 9937.895 8613.565 ;
      RECT 9876.015 187.44 9878.815 8613.565 ;
      RECT 9872.095 187.44 9874.895 8613.565 ;
      RECT 9868.175 187.44 9870.975 8613.565 ;
      RECT 9864.255 187.44 9867.055 8613.565 ;
      RECT 9817.215 187.44 9863.135 8613.565 ;
      RECT 9813.575 187.44 9816.095 8613.565 ;
      RECT 9809.935 187.44 9812.455 8613.565 ;
      RECT 9806.295 187.44 9808.815 8613.565 ;
      RECT 9802.655 187.44 9805.175 8613.565 ;
      RECT 9799.015 187.44 9801.535 8613.565 ;
      RECT 9739.935 187.44 9797.895 8613.565 ;
      RECT 9736.015 187.44 9738.815 8613.565 ;
      RECT 9732.095 187.44 9734.895 8613.565 ;
      RECT 9728.175 187.44 9730.975 8613.565 ;
      RECT 9724.255 187.44 9727.055 8613.565 ;
      RECT 9677.215 187.44 9723.135 8613.565 ;
      RECT 9673.575 187.44 9676.095 8613.565 ;
      RECT 9669.935 187.44 9672.455 8613.565 ;
      RECT 9666.295 187.44 9668.815 8613.565 ;
      RECT 9662.655 187.44 9665.175 8613.565 ;
      RECT 9659.015 187.44 9661.535 8613.565 ;
      RECT 9599.935 187.44 9657.895 8613.565 ;
      RECT 9596.015 187.44 9598.815 8613.565 ;
      RECT 9592.095 187.44 9594.895 8613.565 ;
      RECT 9588.175 187.44 9590.975 8613.565 ;
      RECT 9584.255 187.44 9587.055 8613.565 ;
      RECT 9537.215 187.44 9583.135 8613.565 ;
      RECT 9533.575 187.44 9536.095 8613.565 ;
      RECT 9529.935 187.44 9532.455 8613.565 ;
      RECT 9526.295 187.44 9528.815 8613.565 ;
      RECT 9522.655 187.44 9525.175 8613.565 ;
      RECT 9519.015 187.44 9521.535 8613.565 ;
      RECT 9459.935 187.44 9517.895 8613.565 ;
      RECT 9456.015 187.44 9458.815 8613.565 ;
      RECT 9452.095 187.44 9454.895 8613.565 ;
      RECT 9448.175 187.44 9450.975 8613.565 ;
      RECT 9444.255 187.44 9447.055 8613.565 ;
      RECT 9430.935 188.715 9443.135 8613.565 ;
      RECT 9432.615 187.44 9443.135 8613.565 ;
      RECT 9429.255 187.44 9429.535 8613.565 ;
      RECT 9427.575 187.44 9427.855 8613.565 ;
      RECT 9425.895 187.44 9426.175 8613.565 ;
      RECT 9424.215 187.44 9424.495 8613.565 ;
      RECT 9422.535 187.44 9422.815 8613.565 ;
      RECT 9420.855 187.44 9421.135 8613.565 ;
      RECT 9419.175 187.44 9419.455 8613.565 ;
      RECT 9417.495 187.44 9417.775 8613.565 ;
      RECT 9415.815 187.44 9416.095 8613.565 ;
      RECT 9414.135 187.44 9414.415 8613.565 ;
      RECT 9412.455 187.44 9412.735 8613.565 ;
      RECT 9410.775 187.44 9411.055 8613.565 ;
      RECT 9409.095 187.44 9409.375 8613.565 ;
      RECT 9397.215 187.44 9407.695 8613.565 ;
      RECT 9393.575 187.44 9396.095 8613.565 ;
      RECT 9389.935 187.44 9392.455 8613.565 ;
      RECT 9386.295 187.44 9388.815 8613.565 ;
      RECT 9382.655 187.44 9385.175 8613.565 ;
      RECT 9379.015 187.44 9381.535 8613.565 ;
      RECT 9319.935 187.44 9377.895 8613.565 ;
      RECT 9316.015 187.44 9318.815 8613.565 ;
      RECT 9312.095 187.44 9314.895 8613.565 ;
      RECT 9308.175 187.44 9310.975 8613.565 ;
      RECT 9304.255 187.44 9307.055 8613.565 ;
      RECT 9257.215 187.44 9303.135 8613.565 ;
      RECT 9253.575 187.44 9256.095 8613.565 ;
      RECT 9249.935 187.44 9252.455 8613.565 ;
      RECT 9246.295 187.44 9248.815 8613.565 ;
      RECT 9242.655 187.44 9245.175 8613.565 ;
      RECT 9239.015 187.44 9241.535 8613.565 ;
      RECT 9179.935 187.44 9237.895 8613.565 ;
      RECT 9176.015 187.44 9178.815 8613.565 ;
      RECT 9172.095 187.44 9174.895 8613.565 ;
      RECT 9168.175 187.44 9170.975 8613.565 ;
      RECT 9164.255 187.44 9167.055 8613.565 ;
      RECT 9117.215 187.44 9163.135 8613.565 ;
      RECT 9113.575 187.44 9116.095 8613.565 ;
      RECT 9109.935 187.44 9112.455 8613.565 ;
      RECT 9106.295 187.44 9108.815 8613.565 ;
      RECT 9102.655 187.44 9105.175 8613.565 ;
      RECT 9099.015 187.44 9101.535 8613.565 ;
      RECT 9039.935 187.44 9097.895 8613.565 ;
      RECT 9036.015 187.44 9038.815 8613.565 ;
      RECT 9032.095 187.44 9034.895 8613.565 ;
      RECT 9028.175 187.44 9030.975 8613.565 ;
      RECT 9024.255 187.44 9027.055 8613.565 ;
      RECT 8977.215 187.44 9023.135 8613.565 ;
      RECT 8973.575 187.44 8976.095 8613.565 ;
      RECT 8969.935 187.44 8972.455 8613.565 ;
      RECT 8966.295 187.44 8968.815 8613.565 ;
      RECT 8962.655 187.44 8965.175 8613.565 ;
      RECT 8959.015 187.44 8961.535 8613.565 ;
      RECT 8899.935 187.44 8957.895 8613.565 ;
      RECT 8896.015 187.44 8898.815 8613.565 ;
      RECT 8892.095 187.44 8894.895 8613.565 ;
      RECT 8888.175 187.44 8890.975 8613.565 ;
      RECT 8884.255 187.44 8887.055 8613.565 ;
      RECT 8837.215 187.44 8883.135 8613.565 ;
      RECT 8833.575 187.44 8836.095 8613.565 ;
      RECT 8829.935 187.44 8832.455 8613.565 ;
      RECT 8826.295 187.44 8828.815 8613.565 ;
      RECT 8822.655 187.44 8825.175 8613.565 ;
      RECT 8819.015 187.44 8821.535 8613.565 ;
      RECT 8759.935 187.44 8817.895 8613.565 ;
      RECT 8756.015 187.44 8758.815 8613.565 ;
      RECT 8752.095 187.44 8754.895 8613.565 ;
      RECT 8748.175 187.44 8750.975 8613.565 ;
      RECT 8744.255 187.44 8747.055 8613.565 ;
      RECT 8697.215 187.44 8743.135 8613.565 ;
      RECT 8693.575 187.44 8696.095 8613.565 ;
      RECT 8689.935 187.44 8692.455 8613.565 ;
      RECT 8686.295 187.44 8688.815 8613.565 ;
      RECT 8682.655 187.44 8685.175 8613.565 ;
      RECT 8679.015 187.44 8681.535 8613.565 ;
      RECT 8619.935 187.44 8677.895 8613.565 ;
      RECT 8616.015 187.44 8618.815 8613.565 ;
      RECT 8612.095 187.44 8614.895 8613.565 ;
      RECT 8608.175 187.44 8610.975 8613.565 ;
      RECT 8604.255 187.44 8607.055 8613.565 ;
      RECT 8557.215 187.44 8603.135 8613.565 ;
      RECT 8553.575 187.44 8556.095 8613.565 ;
      RECT 8549.935 187.44 8552.455 8613.565 ;
      RECT 8546.295 187.44 8548.815 8613.565 ;
      RECT 8542.655 187.44 8545.175 8613.565 ;
      RECT 8539.015 187.44 8541.535 8613.565 ;
      RECT 8479.935 187.44 8537.895 8613.565 ;
      RECT 8476.015 187.44 8478.815 8613.565 ;
      RECT 8472.095 187.44 8474.895 8613.565 ;
      RECT 8468.175 187.44 8470.975 8613.565 ;
      RECT 8464.255 187.44 8467.055 8613.565 ;
      RECT 8417.215 187.44 8463.135 8613.565 ;
      RECT 8413.575 187.44 8416.095 8613.565 ;
      RECT 8409.935 187.44 8412.455 8613.565 ;
      RECT 8406.295 187.44 8408.815 8613.565 ;
      RECT 8402.655 187.44 8405.175 8613.565 ;
      RECT 8399.015 187.44 8401.535 8613.565 ;
      RECT 8339.935 187.44 8397.895 8613.565 ;
      RECT 8336.015 187.44 8338.815 8613.565 ;
      RECT 8332.095 187.44 8334.895 8613.565 ;
      RECT 8328.175 187.44 8330.975 8613.565 ;
      RECT 8324.255 187.44 8327.055 8613.565 ;
      RECT 8277.215 187.44 8323.135 8613.565 ;
      RECT 8273.575 187.44 8276.095 8613.565 ;
      RECT 8269.935 187.44 8272.455 8613.565 ;
      RECT 8266.295 187.44 8268.815 8613.565 ;
      RECT 8262.655 187.44 8265.175 8613.565 ;
      RECT 8259.015 187.44 8261.535 8613.565 ;
      RECT 8199.935 187.44 8257.895 8613.565 ;
      RECT 8196.015 187.44 8198.815 8613.565 ;
      RECT 8192.095 187.44 8194.895 8613.565 ;
      RECT 8188.175 187.44 8190.975 8613.565 ;
      RECT 8184.255 187.44 8187.055 8613.565 ;
      RECT 8137.215 187.44 8183.135 8613.565 ;
      RECT 8133.575 187.44 8136.095 8613.565 ;
      RECT 8129.935 187.44 8132.455 8613.565 ;
      RECT 8126.295 187.44 8128.815 8613.565 ;
      RECT 8122.655 187.44 8125.175 8613.565 ;
      RECT 8119.015 187.44 8121.535 8613.565 ;
      RECT 8059.935 187.44 8117.895 8613.565 ;
      RECT 8056.015 187.44 8058.815 8613.565 ;
      RECT 8052.095 187.44 8054.895 8613.565 ;
      RECT 8048.175 187.44 8050.975 8613.565 ;
      RECT 8044.255 187.44 8047.055 8613.565 ;
      RECT 7997.215 187.44 8043.135 8613.565 ;
      RECT 7993.575 187.44 7996.095 8613.565 ;
      RECT 7989.935 187.44 7992.455 8613.565 ;
      RECT 7986.295 187.44 7988.815 8613.565 ;
      RECT 7982.655 187.44 7985.175 8613.565 ;
      RECT 7979.015 187.44 7981.535 8613.565 ;
      RECT 7919.935 187.44 7977.895 8613.565 ;
      RECT 7916.015 187.44 7918.815 8613.565 ;
      RECT 7912.095 187.44 7914.895 8613.565 ;
      RECT 7908.175 187.44 7910.975 8613.565 ;
      RECT 7904.255 187.44 7907.055 8613.565 ;
      RECT 7857.215 187.44 7903.135 8613.565 ;
      RECT 7853.575 187.44 7856.095 8613.565 ;
      RECT 7849.935 187.44 7852.455 8613.565 ;
      RECT 7846.295 187.44 7848.815 8613.565 ;
      RECT 7842.655 187.44 7845.175 8613.565 ;
      RECT 7839.015 187.44 7841.535 8613.565 ;
      RECT 7779.935 187.44 7837.895 8613.565 ;
      RECT 7776.015 187.44 7778.815 8613.565 ;
      RECT 7772.095 187.44 7774.895 8613.565 ;
      RECT 7768.175 187.44 7770.975 8613.565 ;
      RECT 7764.255 187.44 7767.055 8613.565 ;
      RECT 7717.215 187.44 7763.135 8613.565 ;
      RECT 7713.575 187.44 7716.095 8613.565 ;
      RECT 7709.935 187.44 7712.455 8613.565 ;
      RECT 7706.295 187.44 7708.815 8613.565 ;
      RECT 7702.655 187.44 7705.175 8613.565 ;
      RECT 7699.015 187.44 7701.535 8613.565 ;
      RECT 7639.935 187.44 7697.895 8613.565 ;
      RECT 7636.015 187.44 7638.815 8613.565 ;
      RECT 7632.095 187.44 7634.895 8613.565 ;
      RECT 7628.175 187.44 7630.975 8613.565 ;
      RECT 7624.255 187.44 7627.055 8613.565 ;
      RECT 7577.215 187.44 7623.135 8613.565 ;
      RECT 7573.575 187.44 7576.095 8613.565 ;
      RECT 7569.935 187.44 7572.455 8613.565 ;
      RECT 7566.295 187.44 7568.815 8613.565 ;
      RECT 7562.655 187.44 7565.175 8613.565 ;
      RECT 7559.015 187.44 7561.535 8613.565 ;
      RECT 7499.935 187.44 7557.895 8613.565 ;
      RECT 7496.015 187.44 7498.815 8613.565 ;
      RECT 7492.095 187.44 7494.895 8613.565 ;
      RECT 7488.175 187.44 7490.975 8613.565 ;
      RECT 7484.255 187.44 7487.055 8613.565 ;
      RECT 7437.215 187.44 7483.135 8613.565 ;
      RECT 7433.575 187.44 7436.095 8613.565 ;
      RECT 7429.935 187.44 7432.455 8613.565 ;
      RECT 7426.295 187.44 7428.815 8613.565 ;
      RECT 7422.655 187.44 7425.175 8613.565 ;
      RECT 7419.015 187.44 7421.535 8613.565 ;
      RECT 7359.935 187.44 7417.895 8613.565 ;
      RECT 7356.015 187.44 7358.815 8613.565 ;
      RECT 7352.095 187.44 7354.895 8613.565 ;
      RECT 7348.175 187.44 7350.975 8613.565 ;
      RECT 7344.255 187.44 7347.055 8613.565 ;
      RECT 7297.215 187.44 7343.135 8613.565 ;
      RECT 7293.575 187.44 7296.095 8613.565 ;
      RECT 7289.935 187.44 7292.455 8613.565 ;
      RECT 7286.295 187.44 7288.815 8613.565 ;
      RECT 7282.655 187.44 7285.175 8613.565 ;
      RECT 7279.015 187.44 7281.535 8613.565 ;
      RECT 7219.935 187.44 7277.895 8613.565 ;
      RECT 7216.015 187.44 7218.815 8613.565 ;
      RECT 7212.095 187.44 7214.895 8613.565 ;
      RECT 7208.175 187.44 7210.975 8613.565 ;
      RECT 7204.255 187.44 7207.055 8613.565 ;
      RECT 7157.215 187.44 7203.135 8613.565 ;
      RECT 7153.575 187.44 7156.095 8613.565 ;
      RECT 7149.935 187.44 7152.455 8613.565 ;
      RECT 7146.295 187.44 7148.815 8613.565 ;
      RECT 7142.655 187.44 7145.175 8613.565 ;
      RECT 7139.015 187.44 7141.535 8613.565 ;
      RECT 7079.935 187.44 7137.895 8613.565 ;
      RECT 7076.015 187.44 7078.815 8613.565 ;
      RECT 7072.095 187.44 7074.895 8613.565 ;
      RECT 7068.175 187.44 7070.975 8613.565 ;
      RECT 7064.255 187.44 7067.055 8613.565 ;
      RECT 7017.215 187.44 7063.135 8613.565 ;
      RECT 7013.575 187.44 7016.095 8613.565 ;
      RECT 7009.935 187.44 7012.455 8613.565 ;
      RECT 7006.295 187.44 7008.815 8613.565 ;
      RECT 7002.655 187.44 7005.175 8613.565 ;
      RECT 6999.015 187.44 7001.535 8613.565 ;
      RECT 6939.935 187.44 6997.895 8613.565 ;
      RECT 6936.015 187.44 6938.815 8613.565 ;
      RECT 6932.095 187.44 6934.895 8613.565 ;
      RECT 6928.175 187.44 6930.975 8613.565 ;
      RECT 6924.255 187.44 6927.055 8613.565 ;
      RECT 6877.215 187.44 6923.135 8613.565 ;
      RECT 6873.575 187.44 6876.095 8613.565 ;
      RECT 6869.935 187.44 6872.455 8613.565 ;
      RECT 6866.295 187.44 6868.815 8613.565 ;
      RECT 6862.655 187.44 6865.175 8613.565 ;
      RECT 6859.015 187.44 6861.535 8613.565 ;
      RECT 6799.935 187.44 6857.895 8613.565 ;
      RECT 6796.015 187.44 6798.815 8613.565 ;
      RECT 6792.095 187.44 6794.895 8613.565 ;
      RECT 6788.175 187.44 6790.975 8613.565 ;
      RECT 6784.255 187.44 6787.055 8613.565 ;
      RECT 6737.215 187.44 6783.135 8613.565 ;
      RECT 6733.575 187.44 6736.095 8613.565 ;
      RECT 6729.935 187.44 6732.455 8613.565 ;
      RECT 6726.295 187.44 6728.815 8613.565 ;
      RECT 6722.655 187.44 6725.175 8613.565 ;
      RECT 6719.015 187.44 6721.535 8613.565 ;
      RECT 6659.935 187.44 6717.895 8613.565 ;
      RECT 6656.015 187.44 6658.815 8613.565 ;
      RECT 6652.095 187.44 6654.895 8613.565 ;
      RECT 6648.175 187.44 6650.975 8613.565 ;
      RECT 6644.255 187.44 6647.055 8613.565 ;
      RECT 6597.215 187.44 6643.135 8613.565 ;
      RECT 6593.575 187.44 6596.095 8613.565 ;
      RECT 6589.935 187.44 6592.455 8613.565 ;
      RECT 6586.295 187.44 6588.815 8613.565 ;
      RECT 6582.655 187.44 6585.175 8613.565 ;
      RECT 6579.015 187.44 6581.535 8613.565 ;
      RECT 6519.935 187.44 6577.895 8613.565 ;
      RECT 6516.015 187.44 6518.815 8613.565 ;
      RECT 6512.095 187.44 6514.895 8613.565 ;
      RECT 6508.175 187.44 6510.975 8613.565 ;
      RECT 6504.255 187.44 6507.055 8613.565 ;
      RECT 6457.215 187.44 6503.135 8613.565 ;
      RECT 6453.575 187.44 6456.095 8613.565 ;
      RECT 6449.935 187.44 6452.455 8613.565 ;
      RECT 6446.295 187.44 6448.815 8613.565 ;
      RECT 6442.655 187.44 6445.175 8613.565 ;
      RECT 6439.015 187.44 6441.535 8613.565 ;
      RECT 6379.935 187.44 6437.895 8613.565 ;
      RECT 6376.015 187.44 6378.815 8613.565 ;
      RECT 6372.095 187.44 6374.895 8613.565 ;
      RECT 6368.175 187.44 6370.975 8613.565 ;
      RECT 6364.255 187.44 6367.055 8613.565 ;
      RECT 6317.215 187.44 6363.135 8613.565 ;
      RECT 6313.575 187.44 6316.095 8613.565 ;
      RECT 6309.935 187.44 6312.455 8613.565 ;
      RECT 6306.295 187.44 6308.815 8613.565 ;
      RECT 6302.655 187.44 6305.175 8613.565 ;
      RECT 6299.015 187.44 6301.535 8613.565 ;
      RECT 6239.935 187.44 6297.895 8613.565 ;
      RECT 6236.015 187.44 6238.815 8613.565 ;
      RECT 6232.095 187.44 6234.895 8613.565 ;
      RECT 6228.175 187.44 6230.975 8613.565 ;
      RECT 6224.255 187.44 6227.055 8613.565 ;
      RECT 6177.215 187.44 6223.135 8613.565 ;
      RECT 6173.575 187.44 6176.095 8613.565 ;
      RECT 6169.935 187.44 6172.455 8613.565 ;
      RECT 6166.295 187.44 6168.815 8613.565 ;
      RECT 6162.655 187.44 6165.175 8613.565 ;
      RECT 6159.015 187.44 6161.535 8613.565 ;
      RECT 6099.935 187.44 6157.895 8613.565 ;
      RECT 6096.015 187.44 6098.815 8613.565 ;
      RECT 6092.095 187.44 6094.895 8613.565 ;
      RECT 6088.175 187.44 6090.975 8613.565 ;
      RECT 6084.255 187.44 6087.055 8613.565 ;
      RECT 6037.215 187.44 6083.135 8613.565 ;
      RECT 6033.575 187.44 6036.095 8613.565 ;
      RECT 6029.935 187.44 6032.455 8613.565 ;
      RECT 6026.295 187.44 6028.815 8613.565 ;
      RECT 6022.655 187.44 6025.175 8613.565 ;
      RECT 6019.015 187.44 6021.535 8613.565 ;
      RECT 5959.935 187.44 6017.895 8613.565 ;
      RECT 5956.015 187.44 5958.815 8613.565 ;
      RECT 5952.095 187.44 5954.895 8613.565 ;
      RECT 5948.175 187.44 5950.975 8613.565 ;
      RECT 5944.255 187.44 5947.055 8613.565 ;
      RECT 5897.215 187.44 5943.135 8613.565 ;
      RECT 5893.575 187.44 5896.095 8613.565 ;
      RECT 5889.935 187.44 5892.455 8613.565 ;
      RECT 5886.295 187.44 5888.815 8613.565 ;
      RECT 5882.655 187.44 5885.175 8613.565 ;
      RECT 5879.015 187.44 5881.535 8613.565 ;
      RECT 5819.935 187.44 5877.895 8613.565 ;
      RECT 5816.015 187.44 5818.815 8613.565 ;
      RECT 5812.095 187.44 5814.895 8613.565 ;
      RECT 5808.175 187.44 5810.975 8613.565 ;
      RECT 5804.255 187.44 5807.055 8613.565 ;
      RECT 5757.215 187.44 5803.135 8613.565 ;
      RECT 5753.575 187.44 5756.095 8613.565 ;
      RECT 5749.935 187.44 5752.455 8613.565 ;
      RECT 5746.295 187.44 5748.815 8613.565 ;
      RECT 5742.655 187.44 5745.175 8613.565 ;
      RECT 5739.015 187.44 5741.535 8613.565 ;
      RECT 5679.935 187.44 5737.895 8613.565 ;
      RECT 5676.015 187.44 5678.815 8613.565 ;
      RECT 5672.095 187.44 5674.895 8613.565 ;
      RECT 5668.175 187.44 5670.975 8613.565 ;
      RECT 5664.255 187.44 5667.055 8613.565 ;
      RECT 5617.215 187.44 5663.135 8613.565 ;
      RECT 5613.575 187.44 5616.095 8613.565 ;
      RECT 5609.935 187.44 5612.455 8613.565 ;
      RECT 5606.295 187.44 5608.815 8613.565 ;
      RECT 5602.655 187.44 5605.175 8613.565 ;
      RECT 5599.015 187.44 5601.535 8613.565 ;
      RECT 5539.935 187.44 5597.895 8613.565 ;
      RECT 5536.015 187.44 5538.815 8613.565 ;
      RECT 5532.095 187.44 5534.895 8613.565 ;
      RECT 5528.175 187.44 5530.975 8613.565 ;
      RECT 5524.255 187.44 5527.055 8613.565 ;
      RECT 5477.215 187.44 5523.135 8613.565 ;
      RECT 5473.575 187.44 5476.095 8613.565 ;
      RECT 5469.935 187.44 5472.455 8613.565 ;
      RECT 5466.295 187.44 5468.815 8613.565 ;
      RECT 5462.655 187.44 5465.175 8613.565 ;
      RECT 5459.015 187.44 5461.535 8613.565 ;
      RECT 5399.935 187.44 5457.895 8613.565 ;
      RECT 5396.015 187.44 5398.815 8613.565 ;
      RECT 5392.095 187.44 5394.895 8613.565 ;
      RECT 5388.175 187.44 5390.975 8613.565 ;
      RECT 5384.255 187.44 5387.055 8613.565 ;
      RECT 5337.215 187.44 5383.135 8613.565 ;
      RECT 5333.575 187.44 5336.095 8613.565 ;
      RECT 5329.935 187.44 5332.455 8613.565 ;
      RECT 5326.295 187.44 5328.815 8613.565 ;
      RECT 5322.655 187.44 5325.175 8613.565 ;
      RECT 5319.015 187.44 5321.535 8613.565 ;
      RECT 5259.935 187.44 5317.895 8613.565 ;
      RECT 5256.015 187.44 5258.815 8613.565 ;
      RECT 5252.095 187.44 5254.895 8613.565 ;
      RECT 5248.175 187.44 5250.975 8613.565 ;
      RECT 5244.255 187.44 5247.055 8613.565 ;
      RECT 5197.215 187.44 5243.135 8613.565 ;
      RECT 5193.575 187.44 5196.095 8613.565 ;
      RECT 5189.935 187.44 5192.455 8613.565 ;
      RECT 5186.295 187.44 5188.815 8613.565 ;
      RECT 5182.655 187.44 5185.175 8613.565 ;
      RECT 5179.015 187.44 5181.535 8613.565 ;
      RECT 5119.935 187.44 5177.895 8613.565 ;
      RECT 5116.015 187.44 5118.815 8613.565 ;
      RECT 5112.095 187.44 5114.895 8613.565 ;
      RECT 5108.175 187.44 5110.975 8613.565 ;
      RECT 5104.255 187.44 5107.055 8613.565 ;
      RECT 5057.215 187.44 5103.135 8613.565 ;
      RECT 5053.575 187.44 5056.095 8613.565 ;
      RECT 5049.935 187.44 5052.455 8613.565 ;
      RECT 5046.295 187.44 5048.815 8613.565 ;
      RECT 5042.655 187.44 5045.175 8613.565 ;
      RECT 5039.015 187.44 5041.535 8613.565 ;
      RECT 4979.935 187.44 5037.895 8613.565 ;
      RECT 4976.015 187.44 4978.815 8613.565 ;
      RECT 4972.095 187.44 4974.895 8613.565 ;
      RECT 4968.175 187.44 4970.975 8613.565 ;
      RECT 4964.255 187.44 4967.055 8613.565 ;
      RECT 4917.215 187.44 4963.135 8613.565 ;
      RECT 4913.575 187.44 4916.095 8613.565 ;
      RECT 4909.935 187.44 4912.455 8613.565 ;
      RECT 4906.295 187.44 4908.815 8613.565 ;
      RECT 4902.655 187.44 4905.175 8613.565 ;
      RECT 4899.015 187.44 4901.535 8613.565 ;
      RECT 4839.935 187.44 4897.895 8613.565 ;
      RECT 4836.015 187.44 4838.815 8613.565 ;
      RECT 4832.095 187.44 4834.895 8613.565 ;
      RECT 4828.175 187.44 4830.975 8613.565 ;
      RECT 4824.255 187.44 4827.055 8613.565 ;
      RECT 4777.215 187.44 4823.135 8613.565 ;
      RECT 4773.575 187.44 4776.095 8613.565 ;
      RECT 4769.935 187.44 4772.455 8613.565 ;
      RECT 4766.295 187.44 4768.815 8613.565 ;
      RECT 4762.655 187.44 4765.175 8613.565 ;
      RECT 4759.015 187.44 4761.535 8613.565 ;
      RECT 4699.935 187.44 4757.895 8613.565 ;
      RECT 4696.015 187.44 4698.815 8613.565 ;
      RECT 4692.095 187.44 4694.895 8613.565 ;
      RECT 4688.175 187.44 4690.975 8613.565 ;
      RECT 4684.255 187.44 4687.055 8613.565 ;
      RECT 4637.215 187.44 4683.135 8613.565 ;
      RECT 4633.575 187.44 4636.095 8613.565 ;
      RECT 4629.935 187.44 4632.455 8613.565 ;
      RECT 4626.295 187.44 4628.815 8613.565 ;
      RECT 4622.655 187.44 4625.175 8613.565 ;
      RECT 4619.015 187.44 4621.535 8613.565 ;
      RECT 4559.935 187.44 4617.895 8613.565 ;
      RECT 4556.015 187.44 4558.815 8613.565 ;
      RECT 4552.095 187.44 4554.895 8613.565 ;
      RECT 4548.175 187.44 4550.975 8613.565 ;
      RECT 4544.255 187.44 4547.055 8613.565 ;
      RECT 4497.215 187.44 4543.135 8613.565 ;
      RECT 4493.575 187.44 4496.095 8613.565 ;
      RECT 4489.935 187.44 4492.455 8613.565 ;
      RECT 4486.295 187.44 4488.815 8613.565 ;
      RECT 4482.655 187.44 4485.175 8613.565 ;
      RECT 4479.015 187.44 4481.535 8613.565 ;
      RECT 4419.935 187.44 4477.895 8613.565 ;
      RECT 4416.015 187.44 4418.815 8613.565 ;
      RECT 4412.095 187.44 4414.895 8613.565 ;
      RECT 4408.175 187.44 4410.975 8613.565 ;
      RECT 4404.255 187.44 4407.055 8613.565 ;
      RECT 4357.215 187.44 4403.135 8613.565 ;
      RECT 4353.575 187.44 4356.095 8613.565 ;
      RECT 4349.935 187.44 4352.455 8613.565 ;
      RECT 4346.295 187.44 4348.815 8613.565 ;
      RECT 4342.655 187.44 4345.175 8613.565 ;
      RECT 4339.015 187.44 4341.535 8613.565 ;
      RECT 4279.935 187.44 4337.895 8613.565 ;
      RECT 4276.015 187.44 4278.815 8613.565 ;
      RECT 4272.095 187.44 4274.895 8613.565 ;
      RECT 4268.175 187.44 4270.975 8613.565 ;
      RECT 4264.255 187.44 4267.055 8613.565 ;
      RECT 4217.215 187.44 4263.135 8613.565 ;
      RECT 4213.575 187.44 4216.095 8613.565 ;
      RECT 4209.935 187.44 4212.455 8613.565 ;
      RECT 4206.295 187.44 4208.815 8613.565 ;
      RECT 4202.655 187.44 4205.175 8613.565 ;
      RECT 4199.015 187.44 4201.535 8613.565 ;
      RECT 4139.935 187.44 4197.895 8613.565 ;
      RECT 4136.015 187.44 4138.815 8613.565 ;
      RECT 4132.095 187.44 4134.895 8613.565 ;
      RECT 4128.175 187.44 4130.975 8613.565 ;
      RECT 4124.255 187.44 4127.055 8613.565 ;
      RECT 4077.215 187.44 4123.135 8613.565 ;
      RECT 4073.575 187.44 4076.095 8613.565 ;
      RECT 4069.935 187.44 4072.455 8613.565 ;
      RECT 4066.295 187.44 4068.815 8613.565 ;
      RECT 4062.655 187.44 4065.175 8613.565 ;
      RECT 4059.015 187.44 4061.535 8613.565 ;
      RECT 3999.935 187.44 4057.895 8613.565 ;
      RECT 3996.015 187.44 3998.815 8613.565 ;
      RECT 3992.095 187.44 3994.895 8613.565 ;
      RECT 3988.175 187.44 3990.975 8613.565 ;
      RECT 3984.255 187.44 3987.055 8613.565 ;
      RECT 3937.215 187.44 3983.135 8613.565 ;
      RECT 3933.575 187.44 3936.095 8613.565 ;
      RECT 3929.935 187.44 3932.455 8613.565 ;
      RECT 3926.295 187.44 3928.815 8613.565 ;
      RECT 3922.655 187.44 3925.175 8613.565 ;
      RECT 3919.015 187.44 3921.535 8613.565 ;
      RECT 3859.935 187.44 3917.895 8613.565 ;
      RECT 3856.015 187.44 3858.815 8613.565 ;
      RECT 3852.095 187.44 3854.895 8613.565 ;
      RECT 3848.175 187.44 3850.975 8613.565 ;
      RECT 3844.255 187.44 3847.055 8613.565 ;
      RECT 3797.215 187.44 3843.135 8613.565 ;
      RECT 3793.575 187.44 3796.095 8613.565 ;
      RECT 3789.935 187.44 3792.455 8613.565 ;
      RECT 3786.295 187.44 3788.815 8613.565 ;
      RECT 3782.655 187.44 3785.175 8613.565 ;
      RECT 3779.015 187.44 3781.535 8613.565 ;
      RECT 3719.935 187.44 3777.895 8613.565 ;
      RECT 3716.015 187.44 3718.815 8613.565 ;
      RECT 3712.095 187.44 3714.895 8613.565 ;
      RECT 3708.175 187.44 3710.975 8613.565 ;
      RECT 3704.255 187.44 3707.055 8613.565 ;
      RECT 3657.215 187.44 3703.135 8613.565 ;
      RECT 3653.575 187.44 3656.095 8613.565 ;
      RECT 3649.935 187.44 3652.455 8613.565 ;
      RECT 3646.295 187.44 3648.815 8613.565 ;
      RECT 3642.655 187.44 3645.175 8613.565 ;
      RECT 3639.015 187.44 3641.535 8613.565 ;
      RECT 3579.935 187.44 3637.895 8613.565 ;
      RECT 3576.015 187.44 3578.815 8613.565 ;
      RECT 3572.095 187.44 3574.895 8613.565 ;
      RECT 3568.175 187.44 3570.975 8613.565 ;
      RECT 3564.255 187.44 3567.055 8613.565 ;
      RECT 3517.215 187.44 3563.135 8613.565 ;
      RECT 3513.575 187.44 3516.095 8613.565 ;
      RECT 3509.935 187.44 3512.455 8613.565 ;
      RECT 3506.295 187.44 3508.815 8613.565 ;
      RECT 3502.655 187.44 3505.175 8613.565 ;
      RECT 3499.015 187.44 3501.535 8613.565 ;
      RECT 3439.935 187.44 3497.895 8613.565 ;
      RECT 3436.015 187.44 3438.815 8613.565 ;
      RECT 3432.095 187.44 3434.895 8613.565 ;
      RECT 3428.175 187.44 3430.975 8613.565 ;
      RECT 3424.255 187.44 3427.055 8613.565 ;
      RECT 3377.215 187.44 3423.135 8613.565 ;
      RECT 3373.575 187.44 3376.095 8613.565 ;
      RECT 3369.935 187.44 3372.455 8613.565 ;
      RECT 3366.295 187.44 3368.815 8613.565 ;
      RECT 3362.655 187.44 3365.175 8613.565 ;
      RECT 3359.015 187.44 3361.535 8613.565 ;
      RECT 3299.935 187.44 3357.895 8613.565 ;
      RECT 3296.015 187.44 3298.815 8613.565 ;
      RECT 3292.095 187.44 3294.895 8613.565 ;
      RECT 3288.175 187.44 3290.975 8613.565 ;
      RECT 3284.255 187.44 3287.055 8613.565 ;
      RECT 3237.215 187.44 3283.135 8613.565 ;
      RECT 3233.575 187.44 3236.095 8613.565 ;
      RECT 3229.935 187.44 3232.455 8613.565 ;
      RECT 3226.295 187.44 3228.815 8613.565 ;
      RECT 3222.655 187.44 3225.175 8613.565 ;
      RECT 3219.015 187.44 3221.535 8613.565 ;
      RECT 3159.935 187.44 3217.895 8613.565 ;
      RECT 3156.015 187.44 3158.815 8613.565 ;
      RECT 3152.095 187.44 3154.895 8613.565 ;
      RECT 3148.175 187.44 3150.975 8613.565 ;
      RECT 3144.255 187.44 3147.055 8613.565 ;
      RECT 3097.215 187.44 3143.135 8613.565 ;
      RECT 3093.575 187.44 3096.095 8613.565 ;
      RECT 3089.935 187.44 3092.455 8613.565 ;
      RECT 3086.295 187.44 3088.815 8613.565 ;
      RECT 3082.655 187.44 3085.175 8613.565 ;
      RECT 3079.015 187.44 3081.535 8613.565 ;
      RECT 3019.935 187.44 3077.895 8613.565 ;
      RECT 3016.015 187.44 3018.815 8613.565 ;
      RECT 3012.095 187.44 3014.895 8613.565 ;
      RECT 3008.175 187.44 3010.975 8613.565 ;
      RECT 3004.255 187.44 3007.055 8613.565 ;
      RECT 2957.215 187.44 3003.135 8613.565 ;
      RECT 2953.575 187.44 2956.095 8613.565 ;
      RECT 2949.935 187.44 2952.455 8613.565 ;
      RECT 2946.295 187.44 2948.815 8613.565 ;
      RECT 2942.655 187.44 2945.175 8613.565 ;
      RECT 2939.015 187.44 2941.535 8613.565 ;
      RECT 2879.935 187.44 2937.895 8613.565 ;
      RECT 2876.015 187.44 2878.815 8613.565 ;
      RECT 2872.095 187.44 2874.895 8613.565 ;
      RECT 2868.175 187.44 2870.975 8613.565 ;
      RECT 2864.255 187.44 2867.055 8613.565 ;
      RECT 2817.215 187.44 2863.135 8613.565 ;
      RECT 2813.575 187.44 2816.095 8613.565 ;
      RECT 2809.935 187.44 2812.455 8613.565 ;
      RECT 2806.295 187.44 2808.815 8613.565 ;
      RECT 2802.655 187.44 2805.175 8613.565 ;
      RECT 2799.015 187.44 2801.535 8613.565 ;
      RECT 2739.935 187.44 2797.895 8613.565 ;
      RECT 2736.015 187.44 2738.815 8613.565 ;
      RECT 2732.095 187.44 2734.895 8613.565 ;
      RECT 2728.175 187.44 2730.975 8613.565 ;
      RECT 2724.255 187.44 2727.055 8613.565 ;
      RECT 2677.215 187.44 2723.135 8613.565 ;
      RECT 2673.575 187.44 2676.095 8613.565 ;
      RECT 2669.935 187.44 2672.455 8613.565 ;
      RECT 2666.295 187.44 2668.815 8613.565 ;
      RECT 2662.655 187.44 2665.175 8613.565 ;
      RECT 2659.015 187.44 2661.535 8613.565 ;
      RECT 2599.935 187.44 2657.895 8613.565 ;
      RECT 2596.015 187.44 2598.815 8613.565 ;
      RECT 2592.095 187.44 2594.895 8613.565 ;
      RECT 2588.175 187.44 2590.975 8613.565 ;
      RECT 2584.255 187.44 2587.055 8613.565 ;
      RECT 2537.215 187.44 2583.135 8613.565 ;
      RECT 2533.575 187.44 2536.095 8613.565 ;
      RECT 2529.935 187.44 2532.455 8613.565 ;
      RECT 2526.295 187.44 2528.815 8613.565 ;
      RECT 2522.655 187.44 2525.175 8613.565 ;
      RECT 2519.015 187.44 2521.535 8613.565 ;
      RECT 2459.935 187.44 2517.895 8613.565 ;
      RECT 2456.015 187.44 2458.815 8613.565 ;
      RECT 2452.095 187.44 2454.895 8613.565 ;
      RECT 2448.175 187.44 2450.975 8613.565 ;
      RECT 2444.255 187.44 2447.055 8613.565 ;
      RECT 2397.215 187.44 2443.135 8613.565 ;
      RECT 2393.575 187.44 2396.095 8613.565 ;
      RECT 2389.935 187.44 2392.455 8613.565 ;
      RECT 2386.295 187.44 2388.815 8613.565 ;
      RECT 2382.655 187.44 2385.175 8613.565 ;
      RECT 2379.015 187.44 2381.535 8613.565 ;
      RECT 2319.935 187.44 2377.895 8613.565 ;
      RECT 2316.015 187.44 2318.815 8613.565 ;
      RECT 2312.095 187.44 2314.895 8613.565 ;
      RECT 2308.175 187.44 2310.975 8613.565 ;
      RECT 2304.255 187.44 2307.055 8613.565 ;
      RECT 2257.215 187.44 2303.135 8613.565 ;
      RECT 2253.575 187.44 2256.095 8613.565 ;
      RECT 2249.935 187.44 2252.455 8613.565 ;
      RECT 2246.295 187.44 2248.815 8613.565 ;
      RECT 2242.655 187.44 2245.175 8613.565 ;
      RECT 2239.015 187.44 2241.535 8613.565 ;
      RECT 2179.935 187.44 2237.895 8613.565 ;
      RECT 2176.015 187.44 2178.815 8613.565 ;
      RECT 2172.095 187.44 2174.895 8613.565 ;
      RECT 2168.175 187.44 2170.975 8613.565 ;
      RECT 2164.255 187.44 2167.055 8613.565 ;
      RECT 2117.215 187.44 2163.135 8613.565 ;
      RECT 2113.575 187.44 2116.095 8613.565 ;
      RECT 2109.935 187.44 2112.455 8613.565 ;
      RECT 2106.295 187.44 2108.815 8613.565 ;
      RECT 2102.655 187.44 2105.175 8613.565 ;
      RECT 2099.015 187.44 2101.535 8613.565 ;
      RECT 2039.935 187.44 2097.895 8613.565 ;
      RECT 2036.015 187.44 2038.815 8613.565 ;
      RECT 2032.095 187.44 2034.895 8613.565 ;
      RECT 2028.175 187.44 2030.975 8613.565 ;
      RECT 2024.255 187.44 2027.055 8613.565 ;
      RECT 1977.215 187.44 2023.135 8613.565 ;
      RECT 1973.575 187.44 1976.095 8613.565 ;
      RECT 1969.935 187.44 1972.455 8613.565 ;
      RECT 1966.295 187.44 1968.815 8613.565 ;
      RECT 1962.655 187.44 1965.175 8613.565 ;
      RECT 1959.015 187.44 1961.535 8613.565 ;
      RECT 1899.935 187.44 1957.895 8613.565 ;
      RECT 1896.015 187.44 1898.815 8613.565 ;
      RECT 1892.095 187.44 1894.895 8613.565 ;
      RECT 1888.175 187.44 1890.975 8613.565 ;
      RECT 1884.255 187.44 1887.055 8613.565 ;
      RECT 1837.215 187.44 1883.135 8613.565 ;
      RECT 1833.575 187.44 1836.095 8613.565 ;
      RECT 1829.935 187.44 1832.455 8613.565 ;
      RECT 1826.295 187.44 1828.815 8613.565 ;
      RECT 1822.655 187.44 1825.175 8613.565 ;
      RECT 1819.015 187.44 1821.535 8613.565 ;
      RECT 1759.935 187.44 1817.895 8613.565 ;
      RECT 1756.015 187.44 1758.815 8613.565 ;
      RECT 1752.095 187.44 1754.895 8613.565 ;
      RECT 1748.175 187.44 1750.975 8613.565 ;
      RECT 1744.255 187.44 1747.055 8613.565 ;
      RECT 1697.215 187.44 1743.135 8613.565 ;
      RECT 1693.575 187.44 1696.095 8613.565 ;
      RECT 1689.935 187.44 1692.455 8613.565 ;
      RECT 1686.295 187.44 1688.815 8613.565 ;
      RECT 1682.655 187.44 1685.175 8613.565 ;
      RECT 1679.015 187.44 1681.535 8613.565 ;
      RECT 1619.935 187.44 1677.895 8613.565 ;
      RECT 1616.015 187.44 1618.815 8613.565 ;
      RECT 1612.095 187.44 1614.895 8613.565 ;
      RECT 1608.175 187.44 1610.975 8613.565 ;
      RECT 1604.255 187.44 1607.055 8613.565 ;
      RECT 1557.215 187.44 1603.135 8613.565 ;
      RECT 1553.575 187.44 1556.095 8613.565 ;
      RECT 1549.935 187.44 1552.455 8613.565 ;
      RECT 1546.295 187.44 1548.815 8613.565 ;
      RECT 1542.655 187.44 1545.175 8613.565 ;
      RECT 1539.015 187.44 1541.535 8613.565 ;
      RECT 1479.935 187.44 1537.895 8613.565 ;
      RECT 1476.015 187.44 1478.815 8613.565 ;
      RECT 1472.095 187.44 1474.895 8613.565 ;
      RECT 1468.175 187.44 1470.975 8613.565 ;
      RECT 1464.255 187.44 1467.055 8613.565 ;
      RECT 1417.215 187.44 1463.135 8613.565 ;
      RECT 1413.575 187.44 1416.095 8613.565 ;
      RECT 1409.935 187.44 1412.455 8613.565 ;
      RECT 1406.295 187.44 1408.815 8613.565 ;
      RECT 1402.655 187.44 1405.175 8613.565 ;
      RECT 1399.015 187.44 1401.535 8613.565 ;
      RECT 1339.935 187.44 1397.895 8613.565 ;
      RECT 1336.015 187.44 1338.815 8613.565 ;
      RECT 1332.095 187.44 1334.895 8613.565 ;
      RECT 1328.175 187.44 1330.975 8613.565 ;
      RECT 1324.255 187.44 1327.055 8613.565 ;
      RECT 1277.215 187.44 1323.135 8613.565 ;
      RECT 1273.575 187.44 1276.095 8613.565 ;
      RECT 1269.935 187.44 1272.455 8613.565 ;
      RECT 1266.295 187.44 1268.815 8613.565 ;
      RECT 1262.655 187.44 1265.175 8613.565 ;
      RECT 1259.015 187.44 1261.535 8613.565 ;
      RECT 1199.935 187.44 1257.895 8613.565 ;
      RECT 1196.015 187.44 1198.815 8613.565 ;
      RECT 1192.095 187.44 1194.895 8613.565 ;
      RECT 1188.175 187.44 1190.975 8613.565 ;
      RECT 1184.255 187.44 1187.055 8613.565 ;
      RECT 1137.215 187.44 1183.135 8613.565 ;
      RECT 1133.575 187.44 1136.095 8613.565 ;
      RECT 1129.935 187.44 1132.455 8613.565 ;
      RECT 1126.295 187.44 1128.815 8613.565 ;
      RECT 1122.655 187.44 1125.175 8613.565 ;
      RECT 1119.015 187.44 1121.535 8613.565 ;
      RECT 1059.935 187.44 1117.895 8613.565 ;
      RECT 1056.015 187.44 1058.815 8613.565 ;
      RECT 1052.095 187.44 1054.895 8613.565 ;
      RECT 1048.175 187.44 1050.975 8613.565 ;
      RECT 1044.255 187.44 1047.055 8613.565 ;
      RECT 997.215 187.44 1043.135 8613.565 ;
      RECT 993.575 187.44 996.095 8613.565 ;
      RECT 989.935 187.44 992.455 8613.565 ;
      RECT 986.295 187.44 988.815 8613.565 ;
      RECT 982.655 187.44 985.175 8613.565 ;
      RECT 979.015 187.44 981.535 8613.565 ;
      RECT 919.935 187.44 977.895 8613.565 ;
      RECT 916.015 187.44 918.815 8613.565 ;
      RECT 912.095 187.44 914.895 8613.565 ;
      RECT 908.175 187.44 910.975 8613.565 ;
      RECT 904.255 187.44 907.055 8613.565 ;
      RECT 857.215 187.44 903.135 8613.565 ;
      RECT 853.575 187.44 856.095 8613.565 ;
      RECT 849.935 187.44 852.455 8613.565 ;
      RECT 846.295 187.44 848.815 8613.565 ;
      RECT 842.655 187.44 845.175 8613.565 ;
      RECT 839.015 187.44 841.535 8613.565 ;
      RECT 779.935 187.44 837.895 8613.565 ;
      RECT 776.015 187.44 778.815 8613.565 ;
      RECT 772.095 187.44 774.895 8613.565 ;
      RECT 768.175 187.44 770.975 8613.565 ;
      RECT 764.255 187.44 767.055 8613.565 ;
      RECT 717.215 187.44 763.135 8613.565 ;
      RECT 713.575 187.44 716.095 8613.565 ;
      RECT 709.935 187.44 712.455 8613.565 ;
      RECT 706.295 187.44 708.815 8613.565 ;
      RECT 702.655 187.44 705.175 8613.565 ;
      RECT 699.015 187.44 701.535 8613.565 ;
      RECT 639.935 187.44 697.895 8613.565 ;
      RECT 636.015 187.44 638.815 8613.565 ;
      RECT 632.095 187.44 634.895 8613.565 ;
      RECT 628.175 187.44 630.975 8613.565 ;
      RECT 624.255 187.44 627.055 8613.565 ;
      RECT 577.215 187.44 623.135 8613.565 ;
      RECT 573.575 187.44 576.095 8613.565 ;
      RECT 569.935 187.44 572.455 8613.565 ;
      RECT 566.295 187.44 568.815 8613.565 ;
      RECT 562.655 187.44 565.175 8613.565 ;
      RECT 559.015 187.44 561.535 8613.565 ;
      RECT 499.935 187.44 557.895 8613.565 ;
      RECT 496.015 187.44 498.815 8613.565 ;
      RECT 492.095 187.44 494.895 8613.565 ;
      RECT 488.175 187.44 490.975 8613.565 ;
      RECT 484.255 187.44 487.055 8613.565 ;
      RECT 337.025 187.44 483.135 8613.565 ;
      RECT 326.66 187.44 331.985 8613.565 ;
      RECT 9430.935 187.44 9431.215 8613.565 ;
    LAYER M3 ;
      RECT 18342.915 187.94 18367.915 330.165 ;
      RECT 18316.915 187.94 18340.915 330.165 ;
      RECT 18266.305 187.94 18290.305 259.845 ;
      RECT 18253.305 187.94 18264.305 259.845 ;
      RECT 18202.915 187.94 18227.915 330.165 ;
      RECT 18176.915 187.94 18200.915 330.165 ;
      RECT 18126.305 187.94 18150.305 259.845 ;
      RECT 18113.305 187.94 18124.305 259.845 ;
      RECT 18062.915 187.94 18087.915 330.165 ;
      RECT 18036.915 187.94 18060.915 330.165 ;
      RECT 17986.305 187.94 18010.305 259.845 ;
      RECT 17973.305 187.94 17984.305 259.845 ;
      RECT 17922.915 187.94 17947.915 330.165 ;
      RECT 17896.915 187.94 17920.915 330.165 ;
      RECT 17846.305 187.94 17870.305 259.845 ;
      RECT 17833.305 187.94 17844.305 259.845 ;
      RECT 17782.915 187.94 17807.915 330.165 ;
      RECT 17756.915 187.94 17780.915 330.165 ;
      RECT 17706.305 187.94 17730.305 259.845 ;
      RECT 17693.305 187.94 17704.305 259.845 ;
      RECT 17642.915 187.94 17667.915 330.165 ;
      RECT 17616.915 187.94 17640.915 330.165 ;
      RECT 17566.305 187.94 17590.305 259.845 ;
      RECT 17553.305 187.94 17564.305 259.845 ;
      RECT 17502.915 187.94 17527.915 330.165 ;
      RECT 17476.915 187.94 17500.915 330.165 ;
      RECT 17426.305 187.94 17450.305 259.845 ;
      RECT 17413.305 187.94 17424.305 259.845 ;
      RECT 17362.915 187.94 17387.915 330.165 ;
      RECT 17336.915 187.94 17360.915 330.165 ;
      RECT 17286.305 187.94 17310.305 259.845 ;
      RECT 17273.305 187.94 17284.305 259.845 ;
      RECT 17222.915 187.94 17247.915 330.165 ;
      RECT 17196.915 187.94 17220.915 330.165 ;
      RECT 17146.305 187.94 17170.305 259.845 ;
      RECT 17133.305 187.94 17144.305 259.845 ;
      RECT 17082.915 187.94 17107.915 330.165 ;
      RECT 17056.915 187.94 17080.915 330.165 ;
      RECT 17006.305 187.94 17030.305 259.845 ;
      RECT 16993.305 187.94 17004.305 259.845 ;
      RECT 16942.915 187.94 16967.915 330.165 ;
      RECT 16916.915 187.94 16940.915 330.165 ;
      RECT 16866.305 187.94 16890.305 259.845 ;
      RECT 16853.305 187.94 16864.305 259.845 ;
      RECT 16802.915 187.94 16827.915 330.165 ;
      RECT 16776.915 187.94 16800.915 330.165 ;
      RECT 16726.305 187.94 16750.305 259.845 ;
      RECT 16713.305 187.94 16724.305 259.845 ;
      RECT 16662.915 187.94 16687.915 330.165 ;
      RECT 16636.915 187.94 16660.915 330.165 ;
      RECT 16586.305 187.94 16610.305 259.845 ;
      RECT 16573.305 187.94 16584.305 259.845 ;
      RECT 16522.915 187.94 16547.915 330.165 ;
      RECT 16496.915 187.94 16520.915 330.165 ;
      RECT 16446.305 187.94 16470.305 259.845 ;
      RECT 16433.305 187.94 16444.305 259.845 ;
      RECT 16382.915 187.94 16407.915 330.165 ;
      RECT 16356.915 187.94 16380.915 330.165 ;
      RECT 16306.305 187.94 16330.305 259.845 ;
      RECT 16293.305 187.94 16304.305 259.845 ;
      RECT 16242.915 187.94 16267.915 330.165 ;
      RECT 16216.915 187.94 16240.915 330.165 ;
      RECT 16166.305 187.94 16190.305 259.845 ;
      RECT 16153.305 187.94 16164.305 259.845 ;
      RECT 16102.915 187.94 16127.915 330.165 ;
      RECT 16076.915 187.94 16100.915 330.165 ;
      RECT 16026.305 187.94 16050.305 259.845 ;
      RECT 16013.305 187.94 16024.305 259.845 ;
      RECT 15962.915 187.94 15987.915 330.165 ;
      RECT 15936.915 187.94 15960.915 330.165 ;
      RECT 15886.305 187.94 15910.305 259.845 ;
      RECT 15873.305 187.94 15884.305 259.845 ;
      RECT 15822.915 187.94 15847.915 330.165 ;
      RECT 15796.915 187.94 15820.915 330.165 ;
      RECT 15746.305 187.94 15770.305 259.845 ;
      RECT 15733.305 187.94 15744.305 259.845 ;
      RECT 15682.915 187.94 15707.915 330.165 ;
      RECT 15656.915 187.94 15680.915 330.165 ;
      RECT 15606.305 187.94 15630.305 259.845 ;
      RECT 15593.305 187.94 15604.305 259.845 ;
      RECT 15542.915 187.94 15567.915 330.165 ;
      RECT 15516.915 187.94 15540.915 330.165 ;
      RECT 15466.305 187.94 15490.305 259.845 ;
      RECT 15453.305 187.94 15464.305 259.845 ;
      RECT 15402.915 187.94 15427.915 330.165 ;
      RECT 15376.915 187.94 15400.915 330.165 ;
      RECT 15326.305 187.94 15350.305 259.845 ;
      RECT 15313.305 187.94 15324.305 259.845 ;
      RECT 15262.915 187.94 15287.915 330.165 ;
      RECT 15236.915 187.94 15260.915 330.165 ;
      RECT 15186.305 187.94 15210.305 259.845 ;
      RECT 15173.305 187.94 15184.305 259.845 ;
      RECT 15122.915 187.94 15147.915 330.165 ;
      RECT 15096.915 187.94 15120.915 330.165 ;
      RECT 15046.305 187.94 15070.305 259.845 ;
      RECT 15033.305 187.94 15044.305 259.845 ;
      RECT 14982.915 187.94 15007.915 330.165 ;
      RECT 14956.915 187.94 14980.915 330.165 ;
      RECT 14906.305 187.94 14930.305 259.845 ;
      RECT 14893.305 187.94 14904.305 259.845 ;
      RECT 14842.915 187.94 14867.915 330.165 ;
      RECT 14816.915 187.94 14840.915 330.165 ;
      RECT 14766.305 187.94 14790.305 259.845 ;
      RECT 14753.305 187.94 14764.305 259.845 ;
      RECT 14702.915 187.94 14727.915 330.165 ;
      RECT 14676.915 187.94 14700.915 330.165 ;
      RECT 14626.305 187.94 14650.305 259.845 ;
      RECT 14613.305 187.94 14624.305 259.845 ;
      RECT 14562.915 187.94 14587.915 330.165 ;
      RECT 14536.915 187.94 14560.915 330.165 ;
      RECT 14486.305 187.94 14510.305 259.845 ;
      RECT 14473.305 187.94 14484.305 259.845 ;
      RECT 14422.915 187.94 14447.915 330.165 ;
      RECT 14396.915 187.94 14420.915 330.165 ;
      RECT 14346.305 187.94 14370.305 259.845 ;
      RECT 14333.305 187.94 14344.305 259.845 ;
      RECT 14282.915 187.94 14307.915 330.165 ;
      RECT 14256.915 187.94 14280.915 330.165 ;
      RECT 14206.305 187.94 14230.305 259.845 ;
      RECT 14193.305 187.94 14204.305 259.845 ;
      RECT 14142.915 187.94 14167.915 330.165 ;
      RECT 14116.915 187.94 14140.915 330.165 ;
      RECT 14066.305 187.94 14090.305 259.845 ;
      RECT 14053.305 187.94 14064.305 259.845 ;
      RECT 14002.915 187.94 14027.915 330.165 ;
      RECT 13976.915 187.94 14000.915 330.165 ;
      RECT 13926.305 187.94 13950.305 259.845 ;
      RECT 13913.305 187.94 13924.305 259.845 ;
      RECT 13862.915 187.94 13887.915 330.165 ;
      RECT 13836.915 187.94 13860.915 330.165 ;
      RECT 13786.305 187.94 13810.305 259.845 ;
      RECT 13773.305 187.94 13784.305 259.845 ;
      RECT 13722.915 187.94 13747.915 330.165 ;
      RECT 13696.915 187.94 13720.915 330.165 ;
      RECT 13646.305 187.94 13670.305 259.845 ;
      RECT 13633.305 187.94 13644.305 259.845 ;
      RECT 13582.915 187.94 13607.915 330.165 ;
      RECT 13556.915 187.94 13580.915 330.165 ;
      RECT 13506.305 187.94 13530.305 259.845 ;
      RECT 13493.305 187.94 13504.305 259.845 ;
      RECT 13442.915 187.94 13467.915 330.165 ;
      RECT 13416.915 187.94 13440.915 330.165 ;
      RECT 13366.305 187.94 13390.305 259.845 ;
      RECT 13353.305 187.94 13364.305 259.845 ;
      RECT 13302.915 187.94 13327.915 330.165 ;
      RECT 13276.915 187.94 13300.915 330.165 ;
      RECT 13226.305 187.94 13250.305 259.845 ;
      RECT 13213.305 187.94 13224.305 259.845 ;
      RECT 13162.915 187.94 13187.915 330.165 ;
      RECT 13136.915 187.94 13160.915 330.165 ;
      RECT 13086.305 187.94 13110.305 259.845 ;
      RECT 13073.305 187.94 13084.305 259.845 ;
      RECT 13022.915 187.94 13047.915 330.165 ;
      RECT 12996.915 187.94 13020.915 330.165 ;
      RECT 12946.305 187.94 12970.305 259.845 ;
      RECT 12933.305 187.94 12944.305 259.845 ;
      RECT 12882.915 187.94 12907.915 330.165 ;
      RECT 12856.915 187.94 12880.915 330.165 ;
      RECT 12806.305 187.94 12830.305 259.845 ;
      RECT 12793.305 187.94 12804.305 259.845 ;
      RECT 12742.915 187.94 12767.915 330.165 ;
      RECT 12716.915 187.94 12740.915 330.165 ;
      RECT 12666.305 187.94 12690.305 259.845 ;
      RECT 12653.305 187.94 12664.305 259.845 ;
      RECT 12602.915 187.94 12627.915 330.165 ;
      RECT 12576.915 187.94 12600.915 330.165 ;
      RECT 12526.305 187.94 12550.305 259.845 ;
      RECT 12513.305 187.94 12524.305 259.845 ;
      RECT 12462.915 187.94 12487.915 330.165 ;
      RECT 12436.915 187.94 12460.915 330.165 ;
      RECT 12386.305 187.94 12410.305 259.845 ;
      RECT 12373.305 187.94 12384.305 259.845 ;
      RECT 12322.915 187.94 12347.915 330.165 ;
      RECT 12296.915 187.94 12320.915 330.165 ;
      RECT 12246.305 187.94 12270.305 259.845 ;
      RECT 12233.305 187.94 12244.305 259.845 ;
      RECT 12182.915 187.94 12207.915 330.165 ;
      RECT 12156.915 187.94 12180.915 330.165 ;
      RECT 12106.305 187.94 12130.305 259.845 ;
      RECT 12093.305 187.94 12104.305 259.845 ;
      RECT 12042.915 187.94 12067.915 330.165 ;
      RECT 12016.915 187.94 12040.915 330.165 ;
      RECT 11966.305 187.94 11990.305 259.845 ;
      RECT 11953.305 187.94 11964.305 259.845 ;
      RECT 11902.915 187.94 11927.915 330.165 ;
      RECT 11876.915 187.94 11900.915 330.165 ;
      RECT 11826.305 187.94 11850.305 259.845 ;
      RECT 11813.305 187.94 11824.305 259.845 ;
      RECT 11762.915 187.94 11787.915 330.165 ;
      RECT 11736.915 187.94 11760.915 330.165 ;
      RECT 11686.305 187.94 11710.305 259.845 ;
      RECT 11673.305 187.94 11684.305 259.845 ;
      RECT 11622.915 187.94 11647.915 330.165 ;
      RECT 11596.915 187.94 11620.915 330.165 ;
      RECT 11546.305 187.94 11570.305 259.845 ;
      RECT 11533.305 187.94 11544.305 259.845 ;
      RECT 11482.915 187.94 11507.915 330.165 ;
      RECT 11456.915 187.94 11480.915 330.165 ;
      RECT 11406.305 187.94 11430.305 259.845 ;
      RECT 11393.305 187.94 11404.305 259.845 ;
      RECT 11342.915 187.94 11367.915 330.165 ;
      RECT 11316.915 187.94 11340.915 330.165 ;
      RECT 11266.305 187.94 11290.305 259.845 ;
      RECT 11253.305 187.94 11264.305 259.845 ;
      RECT 11202.915 187.94 11227.915 330.165 ;
      RECT 11176.915 187.94 11200.915 330.165 ;
      RECT 11126.305 187.94 11150.305 259.845 ;
      RECT 11113.305 187.94 11124.305 259.845 ;
      RECT 11062.915 187.94 11087.915 330.165 ;
      RECT 11036.915 187.94 11060.915 330.165 ;
      RECT 10986.305 187.94 11010.305 259.845 ;
      RECT 10973.305 187.94 10984.305 259.845 ;
      RECT 10922.915 187.94 10947.915 330.165 ;
      RECT 10896.915 187.94 10920.915 330.165 ;
      RECT 10846.305 187.94 10870.305 259.845 ;
      RECT 10833.305 187.94 10844.305 259.845 ;
      RECT 10782.915 187.94 10807.915 330.165 ;
      RECT 10756.915 187.94 10780.915 330.165 ;
      RECT 10706.305 187.94 10730.305 259.845 ;
      RECT 10693.305 187.94 10704.305 259.845 ;
      RECT 10642.915 187.94 10667.915 330.165 ;
      RECT 10616.915 187.94 10640.915 330.165 ;
      RECT 10566.305 187.94 10590.305 259.845 ;
      RECT 10553.305 187.94 10564.305 259.845 ;
      RECT 10502.915 187.94 10527.915 330.165 ;
      RECT 10476.915 187.94 10500.915 330.165 ;
      RECT 10426.305 187.94 10450.305 259.845 ;
      RECT 10413.305 187.94 10424.305 259.845 ;
      RECT 10362.915 187.94 10387.915 330.165 ;
      RECT 10336.915 187.94 10360.915 330.165 ;
      RECT 10286.305 187.94 10310.305 259.845 ;
      RECT 10273.305 187.94 10284.305 259.845 ;
      RECT 10222.915 187.94 10247.915 330.165 ;
      RECT 10196.915 187.94 10220.915 330.165 ;
      RECT 10146.305 187.94 10170.305 259.845 ;
      RECT 10133.305 187.94 10144.305 259.845 ;
      RECT 10082.915 187.94 10107.915 330.165 ;
      RECT 10056.915 187.94 10080.915 330.165 ;
      RECT 10006.305 187.94 10030.305 259.845 ;
      RECT 9993.305 187.94 10004.305 259.845 ;
      RECT 9942.915 187.94 9967.915 330.165 ;
      RECT 9916.915 187.94 9940.915 330.165 ;
      RECT 9866.305 187.94 9890.305 259.845 ;
      RECT 9853.305 187.94 9864.305 259.845 ;
      RECT 9802.915 187.94 9827.915 330.165 ;
      RECT 9776.915 187.94 9800.915 330.165 ;
      RECT 9726.305 187.94 9750.305 259.845 ;
      RECT 9713.305 187.94 9724.305 259.845 ;
      RECT 9662.915 187.94 9687.915 330.165 ;
      RECT 9636.915 187.94 9660.915 330.165 ;
      RECT 9586.305 187.94 9610.305 259.845 ;
      RECT 9573.305 187.94 9584.305 259.845 ;
      RECT 9522.915 187.94 9547.915 330.165 ;
      RECT 9496.915 187.94 9520.915 330.165 ;
      RECT 9446.305 187.94 9470.305 259.845 ;
      RECT 9433.305 187.94 9444.305 259.845 ;
      RECT 9420.305 187.94 9431.305 297.965 ;
      RECT 9382.915 187.94 9407.915 330.165 ;
      RECT 9356.915 187.94 9380.915 330.165 ;
      RECT 9306.305 187.94 9330.305 259.845 ;
      RECT 9293.305 187.94 9304.305 259.845 ;
      RECT 9242.915 187.94 9267.915 330.165 ;
      RECT 9216.915 187.94 9240.915 330.165 ;
      RECT 9166.305 187.94 9190.305 259.845 ;
      RECT 9153.305 187.94 9164.305 259.845 ;
      RECT 9102.915 187.94 9127.915 330.165 ;
      RECT 9076.915 187.94 9100.915 330.165 ;
      RECT 9026.305 187.94 9050.305 259.845 ;
      RECT 9013.305 187.94 9024.305 259.845 ;
      RECT 8962.915 187.94 8987.915 330.165 ;
      RECT 8936.915 187.94 8960.915 330.165 ;
      RECT 8886.305 187.94 8910.305 259.845 ;
      RECT 8873.305 187.94 8884.305 259.845 ;
      RECT 8822.915 187.94 8847.915 330.165 ;
      RECT 8796.915 187.94 8820.915 330.165 ;
      RECT 8746.305 187.94 8770.305 259.845 ;
      RECT 8733.305 187.94 8744.305 259.845 ;
      RECT 8682.915 187.94 8707.915 330.165 ;
      RECT 8656.915 187.94 8680.915 330.165 ;
      RECT 8606.305 187.94 8630.305 259.845 ;
      RECT 8593.305 187.94 8604.305 259.845 ;
      RECT 8542.915 187.94 8567.915 330.165 ;
      RECT 8516.915 187.94 8540.915 330.165 ;
      RECT 8466.305 187.94 8490.305 259.845 ;
      RECT 8453.305 187.94 8464.305 259.845 ;
      RECT 8402.915 187.94 8427.915 330.165 ;
      RECT 8376.915 187.94 8400.915 330.165 ;
      RECT 8326.305 187.94 8350.305 259.845 ;
      RECT 8313.305 187.94 8324.305 259.845 ;
      RECT 8262.915 187.94 8287.915 330.165 ;
      RECT 8236.915 187.94 8260.915 330.165 ;
      RECT 8186.305 187.94 8210.305 259.845 ;
      RECT 8173.305 187.94 8184.305 259.845 ;
      RECT 8122.915 187.94 8147.915 330.165 ;
      RECT 8096.915 187.94 8120.915 330.165 ;
      RECT 8046.305 187.94 8070.305 259.845 ;
      RECT 8033.305 187.94 8044.305 259.845 ;
      RECT 7982.915 187.94 8007.915 330.165 ;
      RECT 7956.915 187.94 7980.915 330.165 ;
      RECT 7906.305 187.94 7930.305 259.845 ;
      RECT 7893.305 187.94 7904.305 259.845 ;
      RECT 7842.915 187.94 7867.915 330.165 ;
      RECT 7816.915 187.94 7840.915 330.165 ;
      RECT 7766.305 187.94 7790.305 259.845 ;
      RECT 7753.305 187.94 7764.305 259.845 ;
      RECT 7702.915 187.94 7727.915 330.165 ;
      RECT 7676.915 187.94 7700.915 330.165 ;
      RECT 7626.305 187.94 7650.305 259.845 ;
      RECT 7613.305 187.94 7624.305 259.845 ;
      RECT 7562.915 187.94 7587.915 330.165 ;
      RECT 7536.915 187.94 7560.915 330.165 ;
      RECT 7486.305 187.94 7510.305 259.845 ;
      RECT 7473.305 187.94 7484.305 259.845 ;
      RECT 7422.915 187.94 7447.915 330.165 ;
      RECT 7396.915 187.94 7420.915 330.165 ;
      RECT 7346.305 187.94 7370.305 259.845 ;
      RECT 7333.305 187.94 7344.305 259.845 ;
      RECT 7282.915 187.94 7307.915 330.165 ;
      RECT 7256.915 187.94 7280.915 330.165 ;
      RECT 7206.305 187.94 7230.305 259.845 ;
      RECT 7193.305 187.94 7204.305 259.845 ;
      RECT 7142.915 187.94 7167.915 330.165 ;
      RECT 7116.915 187.94 7140.915 330.165 ;
      RECT 7066.305 187.94 7090.305 259.845 ;
      RECT 7053.305 187.94 7064.305 259.845 ;
      RECT 7002.915 187.94 7027.915 330.165 ;
      RECT 6976.915 187.94 7000.915 330.165 ;
      RECT 6926.305 187.94 6950.305 259.845 ;
      RECT 6913.305 187.94 6924.305 259.845 ;
      RECT 6862.915 187.94 6887.915 330.165 ;
      RECT 6836.915 187.94 6860.915 330.165 ;
      RECT 6786.305 187.94 6810.305 259.845 ;
      RECT 6773.305 187.94 6784.305 259.845 ;
      RECT 6722.915 187.94 6747.915 330.165 ;
      RECT 6696.915 187.94 6720.915 330.165 ;
      RECT 6646.305 187.94 6670.305 259.845 ;
      RECT 6633.305 187.94 6644.305 259.845 ;
      RECT 6582.915 187.94 6607.915 330.165 ;
      RECT 6556.915 187.94 6580.915 330.165 ;
      RECT 6506.305 187.94 6530.305 259.845 ;
      RECT 6493.305 187.94 6504.305 259.845 ;
      RECT 6442.915 187.94 6467.915 330.165 ;
      RECT 6416.915 187.94 6440.915 330.165 ;
      RECT 6366.305 187.94 6390.305 259.845 ;
      RECT 6353.305 187.94 6364.305 259.845 ;
      RECT 6302.915 187.94 6327.915 330.165 ;
      RECT 6276.915 187.94 6300.915 330.165 ;
      RECT 6226.305 187.94 6250.305 259.845 ;
      RECT 6213.305 187.94 6224.305 259.845 ;
      RECT 6162.915 187.94 6187.915 330.165 ;
      RECT 6136.915 187.94 6160.915 330.165 ;
      RECT 6086.305 187.94 6110.305 259.845 ;
      RECT 6073.305 187.94 6084.305 259.845 ;
      RECT 6022.915 187.94 6047.915 330.165 ;
      RECT 5996.915 187.94 6020.915 330.165 ;
      RECT 5946.305 187.94 5970.305 259.845 ;
      RECT 5933.305 187.94 5944.305 259.845 ;
      RECT 5882.915 187.94 5907.915 330.165 ;
      RECT 5856.915 187.94 5880.915 330.165 ;
      RECT 5806.305 187.94 5830.305 259.845 ;
      RECT 5793.305 187.94 5804.305 259.845 ;
      RECT 5742.915 187.94 5767.915 330.165 ;
      RECT 5716.915 187.94 5740.915 330.165 ;
      RECT 5666.305 187.94 5690.305 259.845 ;
      RECT 5653.305 187.94 5664.305 259.845 ;
      RECT 5602.915 187.94 5627.915 330.165 ;
      RECT 5576.915 187.94 5600.915 330.165 ;
      RECT 5526.305 187.94 5550.305 259.845 ;
      RECT 5513.305 187.94 5524.305 259.845 ;
      RECT 5462.915 187.94 5487.915 330.165 ;
      RECT 5436.915 187.94 5460.915 330.165 ;
      RECT 5386.305 187.94 5410.305 259.845 ;
      RECT 5373.305 187.94 5384.305 259.845 ;
      RECT 5322.915 187.94 5347.915 330.165 ;
      RECT 5296.915 187.94 5320.915 330.165 ;
      RECT 5246.305 187.94 5270.305 259.845 ;
      RECT 5233.305 187.94 5244.305 259.845 ;
      RECT 5182.915 187.94 5207.915 330.165 ;
      RECT 5156.915 187.94 5180.915 330.165 ;
      RECT 5106.305 187.94 5130.305 259.845 ;
      RECT 5093.305 187.94 5104.305 259.845 ;
      RECT 5042.915 187.94 5067.915 330.165 ;
      RECT 5016.915 187.94 5040.915 330.165 ;
      RECT 4966.305 187.94 4990.305 259.845 ;
      RECT 4953.305 187.94 4964.305 259.845 ;
      RECT 4902.915 187.94 4927.915 330.165 ;
      RECT 4876.915 187.94 4900.915 330.165 ;
      RECT 4826.305 187.94 4850.305 259.845 ;
      RECT 4813.305 187.94 4824.305 259.845 ;
      RECT 4762.915 187.94 4787.915 330.165 ;
      RECT 4736.915 187.94 4760.915 330.165 ;
      RECT 4686.305 187.94 4710.305 259.845 ;
      RECT 4673.305 187.94 4684.305 259.845 ;
      RECT 4622.915 187.94 4647.915 330.165 ;
      RECT 4596.915 187.94 4620.915 330.165 ;
      RECT 4546.305 187.94 4570.305 259.845 ;
      RECT 4533.305 187.94 4544.305 259.845 ;
      RECT 4482.915 187.94 4507.915 330.165 ;
      RECT 4456.915 187.94 4480.915 330.165 ;
      RECT 4406.305 187.94 4430.305 259.845 ;
      RECT 4393.305 187.94 4404.305 259.845 ;
      RECT 4342.915 187.94 4367.915 330.165 ;
      RECT 4316.915 187.94 4340.915 330.165 ;
      RECT 4266.305 187.94 4290.305 259.845 ;
      RECT 4253.305 187.94 4264.305 259.845 ;
      RECT 4202.915 187.94 4227.915 330.165 ;
      RECT 4176.915 187.94 4200.915 330.165 ;
      RECT 4126.305 187.94 4150.305 259.845 ;
      RECT 4113.305 187.94 4124.305 259.845 ;
      RECT 4062.915 187.94 4087.915 330.165 ;
      RECT 4036.915 187.94 4060.915 330.165 ;
      RECT 3986.305 187.94 4010.305 259.845 ;
      RECT 3973.305 187.94 3984.305 259.845 ;
      RECT 3922.915 187.94 3947.915 330.165 ;
      RECT 3896.915 187.94 3920.915 330.165 ;
      RECT 3846.305 187.94 3870.305 259.845 ;
      RECT 3833.305 187.94 3844.305 259.845 ;
      RECT 3782.915 187.94 3807.915 330.165 ;
      RECT 3756.915 187.94 3780.915 330.165 ;
      RECT 3706.305 187.94 3730.305 259.845 ;
      RECT 3693.305 187.94 3704.305 259.845 ;
      RECT 3642.915 187.94 3667.915 330.165 ;
      RECT 3616.915 187.94 3640.915 330.165 ;
      RECT 3566.305 187.94 3590.305 259.845 ;
      RECT 3553.305 187.94 3564.305 259.845 ;
      RECT 3502.915 187.94 3527.915 330.165 ;
      RECT 3476.915 187.94 3500.915 330.165 ;
      RECT 3426.305 187.94 3450.305 259.845 ;
      RECT 3413.305 187.94 3424.305 259.845 ;
      RECT 3362.915 187.94 3387.915 330.165 ;
      RECT 3336.915 187.94 3360.915 330.165 ;
      RECT 3286.305 187.94 3310.305 259.845 ;
      RECT 3273.305 187.94 3284.305 259.845 ;
      RECT 3222.915 187.94 3247.915 330.165 ;
      RECT 3196.915 187.94 3220.915 330.165 ;
      RECT 3146.305 187.94 3170.305 259.845 ;
      RECT 3133.305 187.94 3144.305 259.845 ;
      RECT 3082.915 187.94 3107.915 330.165 ;
      RECT 3056.915 187.94 3080.915 330.165 ;
      RECT 3006.305 187.94 3030.305 259.845 ;
      RECT 2993.305 187.94 3004.305 259.845 ;
      RECT 2942.915 187.94 2967.915 330.165 ;
      RECT 2916.915 187.94 2940.915 330.165 ;
      RECT 2866.305 187.94 2890.305 259.845 ;
      RECT 2853.305 187.94 2864.305 259.845 ;
      RECT 2802.915 187.94 2827.915 330.165 ;
      RECT 2776.915 187.94 2800.915 330.165 ;
      RECT 2726.305 187.94 2750.305 259.845 ;
      RECT 2713.305 187.94 2724.305 259.845 ;
      RECT 2662.915 187.94 2687.915 330.165 ;
      RECT 2636.915 187.94 2660.915 330.165 ;
      RECT 2586.305 187.94 2610.305 259.845 ;
      RECT 2573.305 187.94 2584.305 259.845 ;
      RECT 2522.915 187.94 2547.915 330.165 ;
      RECT 2496.915 187.94 2520.915 330.165 ;
      RECT 2446.305 187.94 2470.305 259.845 ;
      RECT 2433.305 187.94 2444.305 259.845 ;
      RECT 2382.915 187.94 2407.915 330.165 ;
      RECT 2356.915 187.94 2380.915 330.165 ;
      RECT 2306.305 187.94 2330.305 259.845 ;
      RECT 2293.305 187.94 2304.305 259.845 ;
      RECT 2242.915 187.94 2267.915 330.165 ;
      RECT 2216.915 187.94 2240.915 330.165 ;
      RECT 2166.305 187.94 2190.305 259.845 ;
      RECT 2153.305 187.94 2164.305 259.845 ;
      RECT 2102.915 187.94 2127.915 330.165 ;
      RECT 2076.915 187.94 2100.915 330.165 ;
      RECT 2026.305 187.94 2050.305 259.845 ;
      RECT 2013.305 187.94 2024.305 259.845 ;
      RECT 1962.915 187.94 1987.915 330.165 ;
      RECT 1936.915 187.94 1960.915 330.165 ;
      RECT 1886.305 187.94 1910.305 259.845 ;
      RECT 1873.305 187.94 1884.305 259.845 ;
      RECT 1822.915 187.94 1847.915 330.165 ;
      RECT 1796.915 187.94 1820.915 330.165 ;
      RECT 1746.305 187.94 1770.305 259.845 ;
      RECT 1733.305 187.94 1744.305 259.845 ;
      RECT 1682.915 187.94 1707.915 330.165 ;
      RECT 1656.915 187.94 1680.915 330.165 ;
      RECT 1606.305 187.94 1630.305 259.845 ;
      RECT 1593.305 187.94 1604.305 259.845 ;
      RECT 1542.915 187.94 1567.915 330.165 ;
      RECT 1516.915 187.94 1540.915 330.165 ;
      RECT 1466.305 187.94 1490.305 259.845 ;
      RECT 1453.305 187.94 1464.305 259.845 ;
      RECT 1402.915 187.94 1427.915 330.165 ;
      RECT 1376.915 187.94 1400.915 330.165 ;
      RECT 1326.305 187.94 1350.305 259.845 ;
      RECT 1313.305 187.94 1324.305 259.845 ;
      RECT 1262.915 187.94 1287.915 330.165 ;
      RECT 1236.915 187.94 1260.915 330.165 ;
      RECT 1186.305 187.94 1210.305 259.845 ;
      RECT 1173.305 187.94 1184.305 259.845 ;
      RECT 1122.915 187.94 1147.915 330.165 ;
      RECT 1096.915 187.94 1120.915 330.165 ;
      RECT 1046.305 187.94 1070.305 259.845 ;
      RECT 1033.305 187.94 1044.305 259.845 ;
      RECT 982.915 187.94 1007.915 330.165 ;
      RECT 956.915 187.94 980.915 330.165 ;
      RECT 906.305 187.94 930.305 259.845 ;
      RECT 893.305 187.94 904.305 259.845 ;
      RECT 842.915 187.94 867.915 330.165 ;
      RECT 816.915 187.94 840.915 330.165 ;
      RECT 766.305 187.94 790.305 259.845 ;
      RECT 753.305 187.94 764.305 259.845 ;
      RECT 702.915 187.94 727.915 330.165 ;
      RECT 676.915 187.94 700.915 330.165 ;
      RECT 626.305 187.94 650.305 259.845 ;
      RECT 613.305 187.94 624.305 259.845 ;
      RECT 562.915 187.94 587.915 330.165 ;
      RECT 536.915 187.94 560.915 330.165 ;
      RECT 486.305 187.94 510.305 259.845 ;
      RECT 473.305 187.94 484.305 259.845 ;
    LAYER M3 SPACING 0.28 ;
      RECT 12952.095 188.86 18490.46 8613.565 ;
      RECT 18485.135 187.44 18490.46 8613.565 ;
      RECT 18342.655 187.94 18480.095 8613.565 ;
      RECT 18357.215 187.44 18480.095 8613.565 ;
      RECT 18202.655 187.94 18341.535 8613.565 ;
      RECT 18339.015 187.44 18341.535 8613.565 ;
      RECT 18062.655 187.94 18201.535 8613.565 ;
      RECT 18199.015 187.44 18201.535 8613.565 ;
      RECT 17922.655 187.94 18061.535 8613.565 ;
      RECT 18059.015 187.44 18061.535 8613.565 ;
      RECT 17782.655 187.94 17921.535 8613.565 ;
      RECT 17919.015 187.44 17921.535 8613.565 ;
      RECT 17642.655 187.94 17781.535 8613.565 ;
      RECT 17779.015 187.44 17781.535 8613.565 ;
      RECT 17502.655 187.94 17641.535 8613.565 ;
      RECT 17639.015 187.44 17641.535 8613.565 ;
      RECT 17362.655 187.94 17501.535 8613.565 ;
      RECT 17499.015 187.44 17501.535 8613.565 ;
      RECT 17222.655 187.94 17361.535 8613.565 ;
      RECT 17359.015 187.44 17361.535 8613.565 ;
      RECT 17082.655 187.94 17221.535 8613.565 ;
      RECT 17219.015 187.44 17221.535 8613.565 ;
      RECT 16942.655 187.94 17081.535 8613.565 ;
      RECT 17079.015 187.44 17081.535 8613.565 ;
      RECT 16802.655 187.94 16941.535 8613.565 ;
      RECT 16939.015 187.44 16941.535 8613.565 ;
      RECT 16662.655 187.94 16801.535 8613.565 ;
      RECT 16799.015 187.44 16801.535 8613.565 ;
      RECT 16522.655 187.94 16661.535 8613.565 ;
      RECT 16659.015 187.44 16661.535 8613.565 ;
      RECT 16382.655 187.94 16521.535 8613.565 ;
      RECT 16519.015 187.44 16521.535 8613.565 ;
      RECT 16242.655 187.94 16381.535 8613.565 ;
      RECT 16379.015 187.44 16381.535 8613.565 ;
      RECT 16102.655 187.94 16241.535 8613.565 ;
      RECT 16239.015 187.44 16241.535 8613.565 ;
      RECT 15962.655 187.94 16101.535 8613.565 ;
      RECT 16099.015 187.44 16101.535 8613.565 ;
      RECT 15822.655 187.94 15961.535 8613.565 ;
      RECT 15959.015 187.44 15961.535 8613.565 ;
      RECT 15682.655 187.94 15821.535 8613.565 ;
      RECT 15819.015 187.44 15821.535 8613.565 ;
      RECT 15542.655 187.94 15681.535 8613.565 ;
      RECT 15679.015 187.44 15681.535 8613.565 ;
      RECT 15402.655 187.94 15541.535 8613.565 ;
      RECT 15539.015 187.44 15541.535 8613.565 ;
      RECT 15262.655 187.94 15401.535 8613.565 ;
      RECT 15399.015 187.44 15401.535 8613.565 ;
      RECT 15122.655 187.94 15261.535 8613.565 ;
      RECT 15259.015 187.44 15261.535 8613.565 ;
      RECT 14982.655 187.94 15121.535 8613.565 ;
      RECT 15119.015 187.44 15121.535 8613.565 ;
      RECT 14842.655 187.94 14981.535 8613.565 ;
      RECT 14979.015 187.44 14981.535 8613.565 ;
      RECT 14702.655 187.94 14841.535 8613.565 ;
      RECT 14839.015 187.44 14841.535 8613.565 ;
      RECT 14562.655 187.94 14701.535 8613.565 ;
      RECT 14699.015 187.44 14701.535 8613.565 ;
      RECT 14422.655 187.94 14561.535 8613.565 ;
      RECT 14559.015 187.44 14561.535 8613.565 ;
      RECT 14282.655 187.94 14421.535 8613.565 ;
      RECT 14419.015 187.44 14421.535 8613.565 ;
      RECT 14142.655 187.94 14281.535 8613.565 ;
      RECT 14279.015 187.44 14281.535 8613.565 ;
      RECT 14002.655 187.94 14141.535 8613.565 ;
      RECT 14139.015 187.44 14141.535 8613.565 ;
      RECT 13862.655 187.94 14001.535 8613.565 ;
      RECT 13999.015 187.44 14001.535 8613.565 ;
      RECT 13722.655 187.94 13861.535 8613.565 ;
      RECT 13859.015 187.44 13861.535 8613.565 ;
      RECT 13582.655 187.94 13721.535 8613.565 ;
      RECT 13719.015 187.44 13721.535 8613.565 ;
      RECT 13442.655 187.94 13581.535 8613.565 ;
      RECT 13579.015 187.44 13581.535 8613.565 ;
      RECT 13302.655 187.94 13441.535 8613.565 ;
      RECT 13439.015 187.44 13441.535 8613.565 ;
      RECT 13162.655 187.94 13301.535 8613.565 ;
      RECT 13299.015 187.44 13301.535 8613.565 ;
      RECT 13022.655 187.94 13161.535 8613.565 ;
      RECT 13159.015 187.44 13161.535 8613.565 ;
      RECT 12952.095 187.94 13021.535 8613.565 ;
      RECT 13019.015 187.44 13021.535 8613.565 ;
      RECT 18353.575 187.44 18356.095 8613.565 ;
      RECT 18349.935 187.44 18352.455 8613.565 ;
      RECT 18346.295 187.44 18348.815 8613.565 ;
      RECT 18342.655 187.44 18345.175 8613.565 ;
      RECT 18279.935 187.44 18337.895 8613.565 ;
      RECT 18276.015 187.44 18278.815 8613.565 ;
      RECT 18272.095 187.44 18274.895 8613.565 ;
      RECT 18268.175 187.44 18270.975 8613.565 ;
      RECT 18264.255 187.44 18267.055 8613.565 ;
      RECT 18217.215 187.44 18263.135 8613.565 ;
      RECT 18213.575 187.44 18216.095 8613.565 ;
      RECT 18209.935 187.44 18212.455 8613.565 ;
      RECT 18206.295 187.44 18208.815 8613.565 ;
      RECT 18202.655 187.44 18205.175 8613.565 ;
      RECT 18139.935 187.44 18197.895 8613.565 ;
      RECT 18136.015 187.44 18138.815 8613.565 ;
      RECT 18132.095 187.44 18134.895 8613.565 ;
      RECT 18128.175 187.44 18130.975 8613.565 ;
      RECT 18124.255 187.44 18127.055 8613.565 ;
      RECT 18077.215 187.44 18123.135 8613.565 ;
      RECT 18073.575 187.44 18076.095 8613.565 ;
      RECT 18069.935 187.44 18072.455 8613.565 ;
      RECT 18066.295 187.44 18068.815 8613.565 ;
      RECT 18062.655 187.44 18065.175 8613.565 ;
      RECT 17999.935 187.44 18057.895 8613.565 ;
      RECT 17996.015 187.44 17998.815 8613.565 ;
      RECT 17992.095 187.44 17994.895 8613.565 ;
      RECT 17988.175 187.44 17990.975 8613.565 ;
      RECT 17984.255 187.44 17987.055 8613.565 ;
      RECT 17937.215 187.44 17983.135 8613.565 ;
      RECT 17933.575 187.44 17936.095 8613.565 ;
      RECT 17929.935 187.44 17932.455 8613.565 ;
      RECT 17926.295 187.44 17928.815 8613.565 ;
      RECT 17922.655 187.44 17925.175 8613.565 ;
      RECT 17859.935 187.44 17917.895 8613.565 ;
      RECT 17856.015 187.44 17858.815 8613.565 ;
      RECT 17852.095 187.44 17854.895 8613.565 ;
      RECT 17848.175 187.44 17850.975 8613.565 ;
      RECT 17844.255 187.44 17847.055 8613.565 ;
      RECT 17797.215 187.44 17843.135 8613.565 ;
      RECT 17793.575 187.44 17796.095 8613.565 ;
      RECT 17789.935 187.44 17792.455 8613.565 ;
      RECT 17786.295 187.44 17788.815 8613.565 ;
      RECT 17782.655 187.44 17785.175 8613.565 ;
      RECT 17719.935 187.44 17777.895 8613.565 ;
      RECT 17716.015 187.44 17718.815 8613.565 ;
      RECT 17712.095 187.44 17714.895 8613.565 ;
      RECT 17708.175 187.44 17710.975 8613.565 ;
      RECT 17704.255 187.44 17707.055 8613.565 ;
      RECT 17657.215 187.44 17703.135 8613.565 ;
      RECT 17653.575 187.44 17656.095 8613.565 ;
      RECT 17649.935 187.44 17652.455 8613.565 ;
      RECT 17646.295 187.44 17648.815 8613.565 ;
      RECT 17642.655 187.44 17645.175 8613.565 ;
      RECT 17579.935 187.44 17637.895 8613.565 ;
      RECT 17576.015 187.44 17578.815 8613.565 ;
      RECT 17572.095 187.44 17574.895 8613.565 ;
      RECT 17568.175 187.44 17570.975 8613.565 ;
      RECT 17564.255 187.44 17567.055 8613.565 ;
      RECT 17517.215 187.44 17563.135 8613.565 ;
      RECT 17513.575 187.44 17516.095 8613.565 ;
      RECT 17509.935 187.44 17512.455 8613.565 ;
      RECT 17506.295 187.44 17508.815 8613.565 ;
      RECT 17502.655 187.44 17505.175 8613.565 ;
      RECT 17439.935 187.44 17497.895 8613.565 ;
      RECT 17436.015 187.44 17438.815 8613.565 ;
      RECT 17432.095 187.44 17434.895 8613.565 ;
      RECT 17428.175 187.44 17430.975 8613.565 ;
      RECT 17424.255 187.44 17427.055 8613.565 ;
      RECT 17377.215 187.44 17423.135 8613.565 ;
      RECT 17373.575 187.44 17376.095 8613.565 ;
      RECT 17369.935 187.44 17372.455 8613.565 ;
      RECT 17366.295 187.44 17368.815 8613.565 ;
      RECT 17362.655 187.44 17365.175 8613.565 ;
      RECT 17299.935 187.44 17357.895 8613.565 ;
      RECT 17296.015 187.44 17298.815 8613.565 ;
      RECT 17292.095 187.44 17294.895 8613.565 ;
      RECT 17288.175 187.44 17290.975 8613.565 ;
      RECT 17284.255 187.44 17287.055 8613.565 ;
      RECT 17237.215 187.44 17283.135 8613.565 ;
      RECT 17233.575 187.44 17236.095 8613.565 ;
      RECT 17229.935 187.44 17232.455 8613.565 ;
      RECT 17226.295 187.44 17228.815 8613.565 ;
      RECT 17222.655 187.44 17225.175 8613.565 ;
      RECT 17159.935 187.44 17217.895 8613.565 ;
      RECT 17156.015 187.44 17158.815 8613.565 ;
      RECT 17152.095 187.44 17154.895 8613.565 ;
      RECT 17148.175 187.44 17150.975 8613.565 ;
      RECT 17144.255 187.44 17147.055 8613.565 ;
      RECT 17097.215 187.44 17143.135 8613.565 ;
      RECT 17093.575 187.44 17096.095 8613.565 ;
      RECT 17089.935 187.44 17092.455 8613.565 ;
      RECT 17086.295 187.44 17088.815 8613.565 ;
      RECT 17082.655 187.44 17085.175 8613.565 ;
      RECT 17019.935 187.44 17077.895 8613.565 ;
      RECT 17016.015 187.44 17018.815 8613.565 ;
      RECT 17012.095 187.44 17014.895 8613.565 ;
      RECT 17008.175 187.44 17010.975 8613.565 ;
      RECT 17004.255 187.44 17007.055 8613.565 ;
      RECT 16957.215 187.44 17003.135 8613.565 ;
      RECT 16953.575 187.44 16956.095 8613.565 ;
      RECT 16949.935 187.44 16952.455 8613.565 ;
      RECT 16946.295 187.44 16948.815 8613.565 ;
      RECT 16942.655 187.44 16945.175 8613.565 ;
      RECT 16879.935 187.44 16937.895 8613.565 ;
      RECT 16876.015 187.44 16878.815 8613.565 ;
      RECT 16872.095 187.44 16874.895 8613.565 ;
      RECT 16868.175 187.44 16870.975 8613.565 ;
      RECT 16864.255 187.44 16867.055 8613.565 ;
      RECT 16817.215 187.44 16863.135 8613.565 ;
      RECT 16813.575 187.44 16816.095 8613.565 ;
      RECT 16809.935 187.44 16812.455 8613.565 ;
      RECT 16806.295 187.44 16808.815 8613.565 ;
      RECT 16802.655 187.44 16805.175 8613.565 ;
      RECT 16739.935 187.44 16797.895 8613.565 ;
      RECT 16736.015 187.44 16738.815 8613.565 ;
      RECT 16732.095 187.44 16734.895 8613.565 ;
      RECT 16728.175 187.44 16730.975 8613.565 ;
      RECT 16724.255 187.44 16727.055 8613.565 ;
      RECT 16677.215 187.44 16723.135 8613.565 ;
      RECT 16673.575 187.44 16676.095 8613.565 ;
      RECT 16669.935 187.44 16672.455 8613.565 ;
      RECT 16666.295 187.44 16668.815 8613.565 ;
      RECT 16662.655 187.44 16665.175 8613.565 ;
      RECT 16599.935 187.44 16657.895 8613.565 ;
      RECT 16596.015 187.44 16598.815 8613.565 ;
      RECT 16592.095 187.44 16594.895 8613.565 ;
      RECT 16588.175 187.44 16590.975 8613.565 ;
      RECT 16584.255 187.44 16587.055 8613.565 ;
      RECT 16537.215 187.44 16583.135 8613.565 ;
      RECT 16533.575 187.44 16536.095 8613.565 ;
      RECT 16529.935 187.44 16532.455 8613.565 ;
      RECT 16526.295 187.44 16528.815 8613.565 ;
      RECT 16522.655 187.44 16525.175 8613.565 ;
      RECT 16459.935 187.44 16517.895 8613.565 ;
      RECT 16456.015 187.44 16458.815 8613.565 ;
      RECT 16452.095 187.44 16454.895 8613.565 ;
      RECT 16448.175 187.44 16450.975 8613.565 ;
      RECT 16444.255 187.44 16447.055 8613.565 ;
      RECT 16397.215 187.44 16443.135 8613.565 ;
      RECT 16393.575 187.44 16396.095 8613.565 ;
      RECT 16389.935 187.44 16392.455 8613.565 ;
      RECT 16386.295 187.44 16388.815 8613.565 ;
      RECT 16382.655 187.44 16385.175 8613.565 ;
      RECT 16319.935 187.44 16377.895 8613.565 ;
      RECT 16316.015 187.44 16318.815 8613.565 ;
      RECT 16312.095 187.44 16314.895 8613.565 ;
      RECT 16308.175 187.44 16310.975 8613.565 ;
      RECT 16304.255 187.44 16307.055 8613.565 ;
      RECT 16257.215 187.44 16303.135 8613.565 ;
      RECT 16253.575 187.44 16256.095 8613.565 ;
      RECT 16249.935 187.44 16252.455 8613.565 ;
      RECT 16246.295 187.44 16248.815 8613.565 ;
      RECT 16242.655 187.44 16245.175 8613.565 ;
      RECT 16179.935 187.44 16237.895 8613.565 ;
      RECT 16176.015 187.44 16178.815 8613.565 ;
      RECT 16172.095 187.44 16174.895 8613.565 ;
      RECT 16168.175 187.44 16170.975 8613.565 ;
      RECT 16164.255 187.44 16167.055 8613.565 ;
      RECT 16117.215 187.44 16163.135 8613.565 ;
      RECT 16113.575 187.44 16116.095 8613.565 ;
      RECT 16109.935 187.44 16112.455 8613.565 ;
      RECT 16106.295 187.44 16108.815 8613.565 ;
      RECT 16102.655 187.44 16105.175 8613.565 ;
      RECT 16039.935 187.44 16097.895 8613.565 ;
      RECT 16036.015 187.44 16038.815 8613.565 ;
      RECT 16032.095 187.44 16034.895 8613.565 ;
      RECT 16028.175 187.44 16030.975 8613.565 ;
      RECT 16024.255 187.44 16027.055 8613.565 ;
      RECT 15977.215 187.44 16023.135 8613.565 ;
      RECT 15973.575 187.44 15976.095 8613.565 ;
      RECT 15969.935 187.44 15972.455 8613.565 ;
      RECT 15966.295 187.44 15968.815 8613.565 ;
      RECT 15962.655 187.44 15965.175 8613.565 ;
      RECT 15899.935 187.44 15957.895 8613.565 ;
      RECT 15896.015 187.44 15898.815 8613.565 ;
      RECT 15892.095 187.44 15894.895 8613.565 ;
      RECT 15888.175 187.44 15890.975 8613.565 ;
      RECT 15884.255 187.44 15887.055 8613.565 ;
      RECT 15837.215 187.44 15883.135 8613.565 ;
      RECT 15833.575 187.44 15836.095 8613.565 ;
      RECT 15829.935 187.44 15832.455 8613.565 ;
      RECT 15826.295 187.44 15828.815 8613.565 ;
      RECT 15822.655 187.44 15825.175 8613.565 ;
      RECT 15759.935 187.44 15817.895 8613.565 ;
      RECT 15756.015 187.44 15758.815 8613.565 ;
      RECT 15752.095 187.44 15754.895 8613.565 ;
      RECT 15748.175 187.44 15750.975 8613.565 ;
      RECT 15744.255 187.44 15747.055 8613.565 ;
      RECT 15697.215 187.44 15743.135 8613.565 ;
      RECT 15693.575 187.44 15696.095 8613.565 ;
      RECT 15689.935 187.44 15692.455 8613.565 ;
      RECT 15686.295 187.44 15688.815 8613.565 ;
      RECT 15682.655 187.44 15685.175 8613.565 ;
      RECT 15619.935 187.44 15677.895 8613.565 ;
      RECT 15616.015 187.44 15618.815 8613.565 ;
      RECT 15612.095 187.44 15614.895 8613.565 ;
      RECT 15608.175 187.44 15610.975 8613.565 ;
      RECT 15604.255 187.44 15607.055 8613.565 ;
      RECT 15557.215 187.44 15603.135 8613.565 ;
      RECT 15553.575 187.44 15556.095 8613.565 ;
      RECT 15549.935 187.44 15552.455 8613.565 ;
      RECT 15546.295 187.44 15548.815 8613.565 ;
      RECT 15542.655 187.44 15545.175 8613.565 ;
      RECT 15479.935 187.44 15537.895 8613.565 ;
      RECT 15476.015 187.44 15478.815 8613.565 ;
      RECT 15472.095 187.44 15474.895 8613.565 ;
      RECT 15468.175 187.44 15470.975 8613.565 ;
      RECT 15464.255 187.44 15467.055 8613.565 ;
      RECT 15417.215 187.44 15463.135 8613.565 ;
      RECT 15413.575 187.44 15416.095 8613.565 ;
      RECT 15409.935 187.44 15412.455 8613.565 ;
      RECT 15406.295 187.44 15408.815 8613.565 ;
      RECT 15402.655 187.44 15405.175 8613.565 ;
      RECT 15339.935 187.44 15397.895 8613.565 ;
      RECT 15336.015 187.44 15338.815 8613.565 ;
      RECT 15332.095 187.44 15334.895 8613.565 ;
      RECT 15328.175 187.44 15330.975 8613.565 ;
      RECT 15324.255 187.44 15327.055 8613.565 ;
      RECT 15277.215 187.44 15323.135 8613.565 ;
      RECT 15273.575 187.44 15276.095 8613.565 ;
      RECT 15269.935 187.44 15272.455 8613.565 ;
      RECT 15266.295 187.44 15268.815 8613.565 ;
      RECT 15262.655 187.44 15265.175 8613.565 ;
      RECT 15199.935 187.44 15257.895 8613.565 ;
      RECT 15196.015 187.44 15198.815 8613.565 ;
      RECT 15192.095 187.44 15194.895 8613.565 ;
      RECT 15188.175 187.44 15190.975 8613.565 ;
      RECT 15184.255 187.44 15187.055 8613.565 ;
      RECT 15137.215 187.44 15183.135 8613.565 ;
      RECT 15133.575 187.44 15136.095 8613.565 ;
      RECT 15129.935 187.44 15132.455 8613.565 ;
      RECT 15126.295 187.44 15128.815 8613.565 ;
      RECT 15122.655 187.44 15125.175 8613.565 ;
      RECT 15059.935 187.44 15117.895 8613.565 ;
      RECT 15056.015 187.44 15058.815 8613.565 ;
      RECT 15052.095 187.44 15054.895 8613.565 ;
      RECT 15048.175 187.44 15050.975 8613.565 ;
      RECT 15044.255 187.44 15047.055 8613.565 ;
      RECT 14997.215 187.44 15043.135 8613.565 ;
      RECT 14993.575 187.44 14996.095 8613.565 ;
      RECT 14989.935 187.44 14992.455 8613.565 ;
      RECT 14986.295 187.44 14988.815 8613.565 ;
      RECT 14982.655 187.44 14985.175 8613.565 ;
      RECT 14919.935 187.44 14977.895 8613.565 ;
      RECT 14916.015 187.44 14918.815 8613.565 ;
      RECT 14912.095 187.44 14914.895 8613.565 ;
      RECT 14908.175 187.44 14910.975 8613.565 ;
      RECT 14904.255 187.44 14907.055 8613.565 ;
      RECT 14857.215 187.44 14903.135 8613.565 ;
      RECT 14853.575 187.44 14856.095 8613.565 ;
      RECT 14849.935 187.44 14852.455 8613.565 ;
      RECT 14846.295 187.44 14848.815 8613.565 ;
      RECT 14842.655 187.44 14845.175 8613.565 ;
      RECT 14779.935 187.44 14837.895 8613.565 ;
      RECT 14776.015 187.44 14778.815 8613.565 ;
      RECT 14772.095 187.44 14774.895 8613.565 ;
      RECT 14768.175 187.44 14770.975 8613.565 ;
      RECT 14764.255 187.44 14767.055 8613.565 ;
      RECT 14717.215 187.44 14763.135 8613.565 ;
      RECT 14713.575 187.44 14716.095 8613.565 ;
      RECT 14709.935 187.44 14712.455 8613.565 ;
      RECT 14706.295 187.44 14708.815 8613.565 ;
      RECT 14702.655 187.44 14705.175 8613.565 ;
      RECT 14639.935 187.44 14697.895 8613.565 ;
      RECT 14636.015 187.44 14638.815 8613.565 ;
      RECT 14632.095 187.44 14634.895 8613.565 ;
      RECT 14628.175 187.44 14630.975 8613.565 ;
      RECT 14624.255 187.44 14627.055 8613.565 ;
      RECT 14577.215 187.44 14623.135 8613.565 ;
      RECT 14573.575 187.44 14576.095 8613.565 ;
      RECT 14569.935 187.44 14572.455 8613.565 ;
      RECT 14566.295 187.44 14568.815 8613.565 ;
      RECT 14562.655 187.44 14565.175 8613.565 ;
      RECT 14499.935 187.44 14557.895 8613.565 ;
      RECT 14496.015 187.44 14498.815 8613.565 ;
      RECT 14492.095 187.44 14494.895 8613.565 ;
      RECT 14488.175 187.44 14490.975 8613.565 ;
      RECT 14484.255 187.44 14487.055 8613.565 ;
      RECT 14437.215 187.44 14483.135 8613.565 ;
      RECT 14433.575 187.44 14436.095 8613.565 ;
      RECT 14429.935 187.44 14432.455 8613.565 ;
      RECT 14426.295 187.44 14428.815 8613.565 ;
      RECT 14422.655 187.44 14425.175 8613.565 ;
      RECT 14359.935 187.44 14417.895 8613.565 ;
      RECT 14356.015 187.44 14358.815 8613.565 ;
      RECT 14352.095 187.44 14354.895 8613.565 ;
      RECT 14348.175 187.44 14350.975 8613.565 ;
      RECT 14344.255 187.44 14347.055 8613.565 ;
      RECT 14297.215 187.44 14343.135 8613.565 ;
      RECT 14293.575 187.44 14296.095 8613.565 ;
      RECT 14289.935 187.44 14292.455 8613.565 ;
      RECT 14286.295 187.44 14288.815 8613.565 ;
      RECT 14282.655 187.44 14285.175 8613.565 ;
      RECT 14219.935 187.44 14277.895 8613.565 ;
      RECT 14216.015 187.44 14218.815 8613.565 ;
      RECT 14212.095 187.44 14214.895 8613.565 ;
      RECT 14208.175 187.44 14210.975 8613.565 ;
      RECT 14204.255 187.44 14207.055 8613.565 ;
      RECT 14157.215 187.44 14203.135 8613.565 ;
      RECT 14153.575 187.44 14156.095 8613.565 ;
      RECT 14149.935 187.44 14152.455 8613.565 ;
      RECT 14146.295 187.44 14148.815 8613.565 ;
      RECT 14142.655 187.44 14145.175 8613.565 ;
      RECT 14079.935 187.44 14137.895 8613.565 ;
      RECT 14076.015 187.44 14078.815 8613.565 ;
      RECT 14072.095 187.44 14074.895 8613.565 ;
      RECT 14068.175 187.44 14070.975 8613.565 ;
      RECT 14064.255 187.44 14067.055 8613.565 ;
      RECT 14017.215 187.44 14063.135 8613.565 ;
      RECT 14013.575 187.44 14016.095 8613.565 ;
      RECT 14009.935 187.44 14012.455 8613.565 ;
      RECT 14006.295 187.44 14008.815 8613.565 ;
      RECT 14002.655 187.44 14005.175 8613.565 ;
      RECT 13939.935 187.44 13997.895 8613.565 ;
      RECT 13936.015 187.44 13938.815 8613.565 ;
      RECT 13932.095 187.44 13934.895 8613.565 ;
      RECT 13928.175 187.44 13930.975 8613.565 ;
      RECT 13924.255 187.44 13927.055 8613.565 ;
      RECT 13877.215 187.44 13923.135 8613.565 ;
      RECT 13873.575 187.44 13876.095 8613.565 ;
      RECT 13869.935 187.44 13872.455 8613.565 ;
      RECT 13866.295 187.44 13868.815 8613.565 ;
      RECT 13862.655 187.44 13865.175 8613.565 ;
      RECT 13799.935 187.44 13857.895 8613.565 ;
      RECT 13796.015 187.44 13798.815 8613.565 ;
      RECT 13792.095 187.44 13794.895 8613.565 ;
      RECT 13788.175 187.44 13790.975 8613.565 ;
      RECT 13784.255 187.44 13787.055 8613.565 ;
      RECT 13737.215 187.44 13783.135 8613.565 ;
      RECT 13733.575 187.44 13736.095 8613.565 ;
      RECT 13729.935 187.44 13732.455 8613.565 ;
      RECT 13726.295 187.44 13728.815 8613.565 ;
      RECT 13722.655 187.44 13725.175 8613.565 ;
      RECT 13659.935 187.44 13717.895 8613.565 ;
      RECT 13656.015 187.44 13658.815 8613.565 ;
      RECT 13652.095 187.44 13654.895 8613.565 ;
      RECT 13648.175 187.44 13650.975 8613.565 ;
      RECT 13644.255 187.44 13647.055 8613.565 ;
      RECT 13597.215 187.44 13643.135 8613.565 ;
      RECT 13593.575 187.44 13596.095 8613.565 ;
      RECT 13589.935 187.44 13592.455 8613.565 ;
      RECT 13586.295 187.44 13588.815 8613.565 ;
      RECT 13582.655 187.44 13585.175 8613.565 ;
      RECT 13519.935 187.44 13577.895 8613.565 ;
      RECT 13516.015 187.44 13518.815 8613.565 ;
      RECT 13512.095 187.44 13514.895 8613.565 ;
      RECT 13508.175 187.44 13510.975 8613.565 ;
      RECT 13504.255 187.44 13507.055 8613.565 ;
      RECT 13457.215 187.44 13503.135 8613.565 ;
      RECT 13453.575 187.44 13456.095 8613.565 ;
      RECT 13449.935 187.44 13452.455 8613.565 ;
      RECT 13446.295 187.44 13448.815 8613.565 ;
      RECT 13442.655 187.44 13445.175 8613.565 ;
      RECT 13379.935 187.44 13437.895 8613.565 ;
      RECT 13376.015 187.44 13378.815 8613.565 ;
      RECT 13372.095 187.44 13374.895 8613.565 ;
      RECT 13368.175 187.44 13370.975 8613.565 ;
      RECT 13364.255 187.44 13367.055 8613.565 ;
      RECT 13317.215 187.44 13363.135 8613.565 ;
      RECT 13313.575 187.44 13316.095 8613.565 ;
      RECT 13309.935 187.44 13312.455 8613.565 ;
      RECT 13306.295 187.44 13308.815 8613.565 ;
      RECT 13302.655 187.44 13305.175 8613.565 ;
      RECT 13239.935 187.44 13297.895 8613.565 ;
      RECT 13236.015 187.44 13238.815 8613.565 ;
      RECT 13232.095 187.44 13234.895 8613.565 ;
      RECT 13228.175 187.44 13230.975 8613.565 ;
      RECT 13224.255 187.44 13227.055 8613.565 ;
      RECT 13177.215 187.44 13223.135 8613.565 ;
      RECT 13173.575 187.44 13176.095 8613.565 ;
      RECT 13169.935 187.44 13172.455 8613.565 ;
      RECT 13166.295 187.44 13168.815 8613.565 ;
      RECT 13162.655 187.44 13165.175 8613.565 ;
      RECT 13099.935 187.44 13157.895 8613.565 ;
      RECT 13096.015 187.44 13098.815 8613.565 ;
      RECT 13092.095 187.44 13094.895 8613.565 ;
      RECT 13088.175 187.44 13090.975 8613.565 ;
      RECT 13084.255 187.44 13087.055 8613.565 ;
      RECT 13037.215 187.44 13083.135 8613.565 ;
      RECT 13033.575 187.44 13036.095 8613.565 ;
      RECT 13029.935 187.44 13032.455 8613.565 ;
      RECT 13026.295 187.44 13028.815 8613.565 ;
      RECT 13022.655 187.44 13025.175 8613.565 ;
      RECT 12959.935 187.44 13017.895 8613.565 ;
      RECT 12956.015 187.44 12958.815 8613.565 ;
      RECT 12952.095 187.44 12954.895 8613.565 ;
      RECT 326.66 188.86 12952.095 8613.565 ;
      RECT 12882.655 187.94 12952.095 8613.565 ;
      RECT 12742.655 187.94 12881.535 8613.565 ;
      RECT 12879.015 187.44 12881.535 8613.565 ;
      RECT 12602.655 187.94 12741.535 8613.565 ;
      RECT 12739.015 187.44 12741.535 8613.565 ;
      RECT 12462.655 187.94 12601.535 8613.565 ;
      RECT 12599.015 187.44 12601.535 8613.565 ;
      RECT 12322.655 187.94 12461.535 8613.565 ;
      RECT 12459.015 187.44 12461.535 8613.565 ;
      RECT 12182.655 187.94 12321.535 8613.565 ;
      RECT 12319.015 187.44 12321.535 8613.565 ;
      RECT 12042.655 187.94 12181.535 8613.565 ;
      RECT 12179.015 187.44 12181.535 8613.565 ;
      RECT 11902.655 187.94 12041.535 8613.565 ;
      RECT 12039.015 187.44 12041.535 8613.565 ;
      RECT 11762.655 187.94 11901.535 8613.565 ;
      RECT 11899.015 187.44 11901.535 8613.565 ;
      RECT 11622.655 187.94 11761.535 8613.565 ;
      RECT 11759.015 187.44 11761.535 8613.565 ;
      RECT 11482.655 187.94 11621.535 8613.565 ;
      RECT 11619.015 187.44 11621.535 8613.565 ;
      RECT 11342.655 187.94 11481.535 8613.565 ;
      RECT 11479.015 187.44 11481.535 8613.565 ;
      RECT 11202.655 187.94 11341.535 8613.565 ;
      RECT 11339.015 187.44 11341.535 8613.565 ;
      RECT 11062.655 187.94 11201.535 8613.565 ;
      RECT 11199.015 187.44 11201.535 8613.565 ;
      RECT 10922.655 187.94 11061.535 8613.565 ;
      RECT 11059.015 187.44 11061.535 8613.565 ;
      RECT 10782.655 187.94 10921.535 8613.565 ;
      RECT 10919.015 187.44 10921.535 8613.565 ;
      RECT 10642.655 187.94 10781.535 8613.565 ;
      RECT 10779.015 187.44 10781.535 8613.565 ;
      RECT 10502.655 187.94 10641.535 8613.565 ;
      RECT 10639.015 187.44 10641.535 8613.565 ;
      RECT 10362.655 187.94 10501.535 8613.565 ;
      RECT 10499.015 187.44 10501.535 8613.565 ;
      RECT 10222.655 187.94 10361.535 8613.565 ;
      RECT 10359.015 187.44 10361.535 8613.565 ;
      RECT 10082.655 187.94 10221.535 8613.565 ;
      RECT 10219.015 187.44 10221.535 8613.565 ;
      RECT 9942.655 187.94 10081.535 8613.565 ;
      RECT 10079.015 187.44 10081.535 8613.565 ;
      RECT 9802.655 187.94 9941.535 8613.565 ;
      RECT 9939.015 187.44 9941.535 8613.565 ;
      RECT 9662.655 187.94 9801.535 8613.565 ;
      RECT 9799.015 187.44 9801.535 8613.565 ;
      RECT 9522.655 187.94 9661.535 8613.565 ;
      RECT 9659.015 187.44 9661.535 8613.565 ;
      RECT 9420.305 188.715 9521.535 8613.565 ;
      RECT 9519.015 187.44 9521.535 8613.565 ;
      RECT 9419.175 187.44 9419.455 8613.565 ;
      RECT 9417.495 187.44 9417.775 8613.565 ;
      RECT 9415.815 187.44 9416.095 8613.565 ;
      RECT 9414.135 187.44 9414.415 8613.565 ;
      RECT 9412.455 187.44 9412.735 8613.565 ;
      RECT 9410.775 187.44 9411.055 8613.565 ;
      RECT 9409.095 187.44 9409.375 8613.565 ;
      RECT 9382.655 187.94 9407.915 8613.565 ;
      RECT 9242.655 187.94 9381.535 8613.565 ;
      RECT 9379.015 187.44 9381.535 8613.565 ;
      RECT 9102.655 187.94 9241.535 8613.565 ;
      RECT 9239.015 187.44 9241.535 8613.565 ;
      RECT 8962.655 187.94 9101.535 8613.565 ;
      RECT 9099.015 187.44 9101.535 8613.565 ;
      RECT 8822.655 187.94 8961.535 8613.565 ;
      RECT 8959.015 187.44 8961.535 8613.565 ;
      RECT 8682.655 187.94 8821.535 8613.565 ;
      RECT 8819.015 187.44 8821.535 8613.565 ;
      RECT 8542.655 187.94 8681.535 8613.565 ;
      RECT 8679.015 187.44 8681.535 8613.565 ;
      RECT 8402.655 187.94 8541.535 8613.565 ;
      RECT 8539.015 187.44 8541.535 8613.565 ;
      RECT 8262.655 187.94 8401.535 8613.565 ;
      RECT 8399.015 187.44 8401.535 8613.565 ;
      RECT 8122.655 187.94 8261.535 8613.565 ;
      RECT 8259.015 187.44 8261.535 8613.565 ;
      RECT 7982.655 187.94 8121.535 8613.565 ;
      RECT 8119.015 187.44 8121.535 8613.565 ;
      RECT 7842.655 187.94 7981.535 8613.565 ;
      RECT 7979.015 187.44 7981.535 8613.565 ;
      RECT 7702.655 187.94 7841.535 8613.565 ;
      RECT 7839.015 187.44 7841.535 8613.565 ;
      RECT 7562.655 187.94 7701.535 8613.565 ;
      RECT 7699.015 187.44 7701.535 8613.565 ;
      RECT 7422.655 187.94 7561.535 8613.565 ;
      RECT 7559.015 187.44 7561.535 8613.565 ;
      RECT 7282.655 187.94 7421.535 8613.565 ;
      RECT 7419.015 187.44 7421.535 8613.565 ;
      RECT 7142.655 187.94 7281.535 8613.565 ;
      RECT 7279.015 187.44 7281.535 8613.565 ;
      RECT 7002.655 187.94 7141.535 8613.565 ;
      RECT 7139.015 187.44 7141.535 8613.565 ;
      RECT 6862.655 187.94 7001.535 8613.565 ;
      RECT 6999.015 187.44 7001.535 8613.565 ;
      RECT 6722.655 187.94 6861.535 8613.565 ;
      RECT 6859.015 187.44 6861.535 8613.565 ;
      RECT 6582.655 187.94 6721.535 8613.565 ;
      RECT 6719.015 187.44 6721.535 8613.565 ;
      RECT 6442.655 187.94 6581.535 8613.565 ;
      RECT 6579.015 187.44 6581.535 8613.565 ;
      RECT 6302.655 187.94 6441.535 8613.565 ;
      RECT 6439.015 187.44 6441.535 8613.565 ;
      RECT 6162.655 187.94 6301.535 8613.565 ;
      RECT 6299.015 187.44 6301.535 8613.565 ;
      RECT 6022.655 187.94 6161.535 8613.565 ;
      RECT 6159.015 187.44 6161.535 8613.565 ;
      RECT 5882.655 187.94 6021.535 8613.565 ;
      RECT 6019.015 187.44 6021.535 8613.565 ;
      RECT 5742.655 187.94 5881.535 8613.565 ;
      RECT 5879.015 187.44 5881.535 8613.565 ;
      RECT 5602.655 187.94 5741.535 8613.565 ;
      RECT 5739.015 187.44 5741.535 8613.565 ;
      RECT 5462.655 187.94 5601.535 8613.565 ;
      RECT 5599.015 187.44 5601.535 8613.565 ;
      RECT 5322.655 187.94 5461.535 8613.565 ;
      RECT 5459.015 187.44 5461.535 8613.565 ;
      RECT 5182.655 187.94 5321.535 8613.565 ;
      RECT 5319.015 187.44 5321.535 8613.565 ;
      RECT 5042.655 187.94 5181.535 8613.565 ;
      RECT 5179.015 187.44 5181.535 8613.565 ;
      RECT 4902.655 187.94 5041.535 8613.565 ;
      RECT 5039.015 187.44 5041.535 8613.565 ;
      RECT 4762.655 187.94 4901.535 8613.565 ;
      RECT 4899.015 187.44 4901.535 8613.565 ;
      RECT 4622.655 187.94 4761.535 8613.565 ;
      RECT 4759.015 187.44 4761.535 8613.565 ;
      RECT 4482.655 187.94 4621.535 8613.565 ;
      RECT 4619.015 187.44 4621.535 8613.565 ;
      RECT 4342.655 187.94 4481.535 8613.565 ;
      RECT 4479.015 187.44 4481.535 8613.565 ;
      RECT 4202.655 187.94 4341.535 8613.565 ;
      RECT 4339.015 187.44 4341.535 8613.565 ;
      RECT 4062.655 187.94 4201.535 8613.565 ;
      RECT 4199.015 187.44 4201.535 8613.565 ;
      RECT 3922.655 187.94 4061.535 8613.565 ;
      RECT 4059.015 187.44 4061.535 8613.565 ;
      RECT 3782.655 187.94 3921.535 8613.565 ;
      RECT 3919.015 187.44 3921.535 8613.565 ;
      RECT 3642.655 187.94 3781.535 8613.565 ;
      RECT 3779.015 187.44 3781.535 8613.565 ;
      RECT 3502.655 187.94 3641.535 8613.565 ;
      RECT 3639.015 187.44 3641.535 8613.565 ;
      RECT 3362.655 187.94 3501.535 8613.565 ;
      RECT 3499.015 187.44 3501.535 8613.565 ;
      RECT 3222.655 187.94 3361.535 8613.565 ;
      RECT 3359.015 187.44 3361.535 8613.565 ;
      RECT 3082.655 187.94 3221.535 8613.565 ;
      RECT 3219.015 187.44 3221.535 8613.565 ;
      RECT 2942.655 187.94 3081.535 8613.565 ;
      RECT 3079.015 187.44 3081.535 8613.565 ;
      RECT 2802.655 187.94 2941.535 8613.565 ;
      RECT 2939.015 187.44 2941.535 8613.565 ;
      RECT 2662.655 187.94 2801.535 8613.565 ;
      RECT 2799.015 187.44 2801.535 8613.565 ;
      RECT 2522.655 187.94 2661.535 8613.565 ;
      RECT 2659.015 187.44 2661.535 8613.565 ;
      RECT 2382.655 187.94 2521.535 8613.565 ;
      RECT 2519.015 187.44 2521.535 8613.565 ;
      RECT 2242.655 187.94 2381.535 8613.565 ;
      RECT 2379.015 187.44 2381.535 8613.565 ;
      RECT 2102.655 187.94 2241.535 8613.565 ;
      RECT 2239.015 187.44 2241.535 8613.565 ;
      RECT 1962.655 187.94 2101.535 8613.565 ;
      RECT 2099.015 187.44 2101.535 8613.565 ;
      RECT 1822.655 187.94 1961.535 8613.565 ;
      RECT 1959.015 187.44 1961.535 8613.565 ;
      RECT 1682.655 187.94 1821.535 8613.565 ;
      RECT 1819.015 187.44 1821.535 8613.565 ;
      RECT 1542.655 187.94 1681.535 8613.565 ;
      RECT 1679.015 187.44 1681.535 8613.565 ;
      RECT 1402.655 187.94 1541.535 8613.565 ;
      RECT 1539.015 187.44 1541.535 8613.565 ;
      RECT 1262.655 187.94 1401.535 8613.565 ;
      RECT 1399.015 187.44 1401.535 8613.565 ;
      RECT 1122.655 187.94 1261.535 8613.565 ;
      RECT 1259.015 187.44 1261.535 8613.565 ;
      RECT 982.655 187.94 1121.535 8613.565 ;
      RECT 1119.015 187.44 1121.535 8613.565 ;
      RECT 842.655 187.94 981.535 8613.565 ;
      RECT 979.015 187.44 981.535 8613.565 ;
      RECT 702.655 187.94 841.535 8613.565 ;
      RECT 839.015 187.44 841.535 8613.565 ;
      RECT 562.655 187.94 701.535 8613.565 ;
      RECT 699.015 187.44 701.535 8613.565 ;
      RECT 337.025 187.94 561.535 8613.565 ;
      RECT 559.015 187.44 561.535 8613.565 ;
      RECT 326.66 187.44 331.985 8613.565 ;
      RECT 9432.615 187.94 9521.535 8613.565 ;
      RECT 9420.305 187.94 9431.305 8613.565 ;
      RECT 12948.175 187.44 12950.975 8613.565 ;
      RECT 12944.255 187.44 12947.055 8613.565 ;
      RECT 12897.215 187.44 12943.135 8613.565 ;
      RECT 12893.575 187.44 12896.095 8613.565 ;
      RECT 12889.935 187.44 12892.455 8613.565 ;
      RECT 12886.295 187.44 12888.815 8613.565 ;
      RECT 12882.655 187.44 12885.175 8613.565 ;
      RECT 12819.935 187.44 12877.895 8613.565 ;
      RECT 12816.015 187.44 12818.815 8613.565 ;
      RECT 12812.095 187.44 12814.895 8613.565 ;
      RECT 12808.175 187.44 12810.975 8613.565 ;
      RECT 12804.255 187.44 12807.055 8613.565 ;
      RECT 12757.215 187.44 12803.135 8613.565 ;
      RECT 12753.575 187.44 12756.095 8613.565 ;
      RECT 12749.935 187.44 12752.455 8613.565 ;
      RECT 12746.295 187.44 12748.815 8613.565 ;
      RECT 12742.655 187.44 12745.175 8613.565 ;
      RECT 12679.935 187.44 12737.895 8613.565 ;
      RECT 12676.015 187.44 12678.815 8613.565 ;
      RECT 12672.095 187.44 12674.895 8613.565 ;
      RECT 12668.175 187.44 12670.975 8613.565 ;
      RECT 12664.255 187.44 12667.055 8613.565 ;
      RECT 12617.215 187.44 12663.135 8613.565 ;
      RECT 12613.575 187.44 12616.095 8613.565 ;
      RECT 12609.935 187.44 12612.455 8613.565 ;
      RECT 12606.295 187.44 12608.815 8613.565 ;
      RECT 12602.655 187.44 12605.175 8613.565 ;
      RECT 12539.935 187.44 12597.895 8613.565 ;
      RECT 12536.015 187.44 12538.815 8613.565 ;
      RECT 12532.095 187.44 12534.895 8613.565 ;
      RECT 12528.175 187.44 12530.975 8613.565 ;
      RECT 12524.255 187.44 12527.055 8613.565 ;
      RECT 12477.215 187.44 12523.135 8613.565 ;
      RECT 12473.575 187.44 12476.095 8613.565 ;
      RECT 12469.935 187.44 12472.455 8613.565 ;
      RECT 12466.295 187.44 12468.815 8613.565 ;
      RECT 12462.655 187.44 12465.175 8613.565 ;
      RECT 12399.935 187.44 12457.895 8613.565 ;
      RECT 12396.015 187.44 12398.815 8613.565 ;
      RECT 12392.095 187.44 12394.895 8613.565 ;
      RECT 12388.175 187.44 12390.975 8613.565 ;
      RECT 12384.255 187.44 12387.055 8613.565 ;
      RECT 12337.215 187.44 12383.135 8613.565 ;
      RECT 12333.575 187.44 12336.095 8613.565 ;
      RECT 12329.935 187.44 12332.455 8613.565 ;
      RECT 12326.295 187.44 12328.815 8613.565 ;
      RECT 12322.655 187.44 12325.175 8613.565 ;
      RECT 12259.935 187.44 12317.895 8613.565 ;
      RECT 12256.015 187.44 12258.815 8613.565 ;
      RECT 12252.095 187.44 12254.895 8613.565 ;
      RECT 12248.175 187.44 12250.975 8613.565 ;
      RECT 12244.255 187.44 12247.055 8613.565 ;
      RECT 12197.215 187.44 12243.135 8613.565 ;
      RECT 12193.575 187.44 12196.095 8613.565 ;
      RECT 12189.935 187.44 12192.455 8613.565 ;
      RECT 12186.295 187.44 12188.815 8613.565 ;
      RECT 12182.655 187.44 12185.175 8613.565 ;
      RECT 12119.935 187.44 12177.895 8613.565 ;
      RECT 12116.015 187.44 12118.815 8613.565 ;
      RECT 12112.095 187.44 12114.895 8613.565 ;
      RECT 12108.175 187.44 12110.975 8613.565 ;
      RECT 12104.255 187.44 12107.055 8613.565 ;
      RECT 12057.215 187.44 12103.135 8613.565 ;
      RECT 12053.575 187.44 12056.095 8613.565 ;
      RECT 12049.935 187.44 12052.455 8613.565 ;
      RECT 12046.295 187.44 12048.815 8613.565 ;
      RECT 12042.655 187.44 12045.175 8613.565 ;
      RECT 11979.935 187.44 12037.895 8613.565 ;
      RECT 11976.015 187.44 11978.815 8613.565 ;
      RECT 11972.095 187.44 11974.895 8613.565 ;
      RECT 11968.175 187.44 11970.975 8613.565 ;
      RECT 11964.255 187.44 11967.055 8613.565 ;
      RECT 11917.215 187.44 11963.135 8613.565 ;
      RECT 11913.575 187.44 11916.095 8613.565 ;
      RECT 11909.935 187.44 11912.455 8613.565 ;
      RECT 11906.295 187.44 11908.815 8613.565 ;
      RECT 11902.655 187.44 11905.175 8613.565 ;
      RECT 11839.935 187.44 11897.895 8613.565 ;
      RECT 11836.015 187.44 11838.815 8613.565 ;
      RECT 11832.095 187.44 11834.895 8613.565 ;
      RECT 11828.175 187.44 11830.975 8613.565 ;
      RECT 11824.255 187.44 11827.055 8613.565 ;
      RECT 11777.215 187.44 11823.135 8613.565 ;
      RECT 11773.575 187.44 11776.095 8613.565 ;
      RECT 11769.935 187.44 11772.455 8613.565 ;
      RECT 11766.295 187.44 11768.815 8613.565 ;
      RECT 11762.655 187.44 11765.175 8613.565 ;
      RECT 11699.935 187.44 11757.895 8613.565 ;
      RECT 11696.015 187.44 11698.815 8613.565 ;
      RECT 11692.095 187.44 11694.895 8613.565 ;
      RECT 11688.175 187.44 11690.975 8613.565 ;
      RECT 11684.255 187.44 11687.055 8613.565 ;
      RECT 11637.215 187.44 11683.135 8613.565 ;
      RECT 11633.575 187.44 11636.095 8613.565 ;
      RECT 11629.935 187.44 11632.455 8613.565 ;
      RECT 11626.295 187.44 11628.815 8613.565 ;
      RECT 11622.655 187.44 11625.175 8613.565 ;
      RECT 11559.935 187.44 11617.895 8613.565 ;
      RECT 11556.015 187.44 11558.815 8613.565 ;
      RECT 11552.095 187.44 11554.895 8613.565 ;
      RECT 11548.175 187.44 11550.975 8613.565 ;
      RECT 11544.255 187.44 11547.055 8613.565 ;
      RECT 11497.215 187.44 11543.135 8613.565 ;
      RECT 11493.575 187.44 11496.095 8613.565 ;
      RECT 11489.935 187.44 11492.455 8613.565 ;
      RECT 11486.295 187.44 11488.815 8613.565 ;
      RECT 11482.655 187.44 11485.175 8613.565 ;
      RECT 11419.935 187.44 11477.895 8613.565 ;
      RECT 11416.015 187.44 11418.815 8613.565 ;
      RECT 11412.095 187.44 11414.895 8613.565 ;
      RECT 11408.175 187.44 11410.975 8613.565 ;
      RECT 11404.255 187.44 11407.055 8613.565 ;
      RECT 11357.215 187.44 11403.135 8613.565 ;
      RECT 11353.575 187.44 11356.095 8613.565 ;
      RECT 11349.935 187.44 11352.455 8613.565 ;
      RECT 11346.295 187.44 11348.815 8613.565 ;
      RECT 11342.655 187.44 11345.175 8613.565 ;
      RECT 11279.935 187.44 11337.895 8613.565 ;
      RECT 11276.015 187.44 11278.815 8613.565 ;
      RECT 11272.095 187.44 11274.895 8613.565 ;
      RECT 11268.175 187.44 11270.975 8613.565 ;
      RECT 11264.255 187.44 11267.055 8613.565 ;
      RECT 11217.215 187.44 11263.135 8613.565 ;
      RECT 11213.575 187.44 11216.095 8613.565 ;
      RECT 11209.935 187.44 11212.455 8613.565 ;
      RECT 11206.295 187.44 11208.815 8613.565 ;
      RECT 11202.655 187.44 11205.175 8613.565 ;
      RECT 11139.935 187.44 11197.895 8613.565 ;
      RECT 11136.015 187.44 11138.815 8613.565 ;
      RECT 11132.095 187.44 11134.895 8613.565 ;
      RECT 11128.175 187.44 11130.975 8613.565 ;
      RECT 11124.255 187.44 11127.055 8613.565 ;
      RECT 11077.215 187.44 11123.135 8613.565 ;
      RECT 11073.575 187.44 11076.095 8613.565 ;
      RECT 11069.935 187.44 11072.455 8613.565 ;
      RECT 11066.295 187.44 11068.815 8613.565 ;
      RECT 11062.655 187.44 11065.175 8613.565 ;
      RECT 10999.935 187.44 11057.895 8613.565 ;
      RECT 10996.015 187.44 10998.815 8613.565 ;
      RECT 10992.095 187.44 10994.895 8613.565 ;
      RECT 10988.175 187.44 10990.975 8613.565 ;
      RECT 10984.255 187.44 10987.055 8613.565 ;
      RECT 10937.215 187.44 10983.135 8613.565 ;
      RECT 10933.575 187.44 10936.095 8613.565 ;
      RECT 10929.935 187.44 10932.455 8613.565 ;
      RECT 10926.295 187.44 10928.815 8613.565 ;
      RECT 10922.655 187.44 10925.175 8613.565 ;
      RECT 10859.935 187.44 10917.895 8613.565 ;
      RECT 10856.015 187.44 10858.815 8613.565 ;
      RECT 10852.095 187.44 10854.895 8613.565 ;
      RECT 10848.175 187.44 10850.975 8613.565 ;
      RECT 10844.255 187.44 10847.055 8613.565 ;
      RECT 10797.215 187.44 10843.135 8613.565 ;
      RECT 10793.575 187.44 10796.095 8613.565 ;
      RECT 10789.935 187.44 10792.455 8613.565 ;
      RECT 10786.295 187.44 10788.815 8613.565 ;
      RECT 10782.655 187.44 10785.175 8613.565 ;
      RECT 10719.935 187.44 10777.895 8613.565 ;
      RECT 10716.015 187.44 10718.815 8613.565 ;
      RECT 10712.095 187.44 10714.895 8613.565 ;
      RECT 10708.175 187.44 10710.975 8613.565 ;
      RECT 10704.255 187.44 10707.055 8613.565 ;
      RECT 10657.215 187.44 10703.135 8613.565 ;
      RECT 10653.575 187.44 10656.095 8613.565 ;
      RECT 10649.935 187.44 10652.455 8613.565 ;
      RECT 10646.295 187.44 10648.815 8613.565 ;
      RECT 10642.655 187.44 10645.175 8613.565 ;
      RECT 10579.935 187.44 10637.895 8613.565 ;
      RECT 10576.015 187.44 10578.815 8613.565 ;
      RECT 10572.095 187.44 10574.895 8613.565 ;
      RECT 10568.175 187.44 10570.975 8613.565 ;
      RECT 10564.255 187.44 10567.055 8613.565 ;
      RECT 10517.215 187.44 10563.135 8613.565 ;
      RECT 10513.575 187.44 10516.095 8613.565 ;
      RECT 10509.935 187.44 10512.455 8613.565 ;
      RECT 10506.295 187.44 10508.815 8613.565 ;
      RECT 10502.655 187.44 10505.175 8613.565 ;
      RECT 10439.935 187.44 10497.895 8613.565 ;
      RECT 10436.015 187.44 10438.815 8613.565 ;
      RECT 10432.095 187.44 10434.895 8613.565 ;
      RECT 10428.175 187.44 10430.975 8613.565 ;
      RECT 10424.255 187.44 10427.055 8613.565 ;
      RECT 10377.215 187.44 10423.135 8613.565 ;
      RECT 10373.575 187.44 10376.095 8613.565 ;
      RECT 10369.935 187.44 10372.455 8613.565 ;
      RECT 10366.295 187.44 10368.815 8613.565 ;
      RECT 10362.655 187.44 10365.175 8613.565 ;
      RECT 10299.935 187.44 10357.895 8613.565 ;
      RECT 10296.015 187.44 10298.815 8613.565 ;
      RECT 10292.095 187.44 10294.895 8613.565 ;
      RECT 10288.175 187.44 10290.975 8613.565 ;
      RECT 10284.255 187.44 10287.055 8613.565 ;
      RECT 10237.215 187.44 10283.135 8613.565 ;
      RECT 10233.575 187.44 10236.095 8613.565 ;
      RECT 10229.935 187.44 10232.455 8613.565 ;
      RECT 10226.295 187.44 10228.815 8613.565 ;
      RECT 10222.655 187.44 10225.175 8613.565 ;
      RECT 10159.935 187.44 10217.895 8613.565 ;
      RECT 10156.015 187.44 10158.815 8613.565 ;
      RECT 10152.095 187.44 10154.895 8613.565 ;
      RECT 10148.175 187.44 10150.975 8613.565 ;
      RECT 10144.255 187.44 10147.055 8613.565 ;
      RECT 10097.215 187.44 10143.135 8613.565 ;
      RECT 10093.575 187.44 10096.095 8613.565 ;
      RECT 10089.935 187.44 10092.455 8613.565 ;
      RECT 10086.295 187.44 10088.815 8613.565 ;
      RECT 10082.655 187.44 10085.175 8613.565 ;
      RECT 10019.935 187.44 10077.895 8613.565 ;
      RECT 10016.015 187.44 10018.815 8613.565 ;
      RECT 10012.095 187.44 10014.895 8613.565 ;
      RECT 10008.175 187.44 10010.975 8613.565 ;
      RECT 10004.255 187.44 10007.055 8613.565 ;
      RECT 9957.215 187.44 10003.135 8613.565 ;
      RECT 9953.575 187.44 9956.095 8613.565 ;
      RECT 9949.935 187.44 9952.455 8613.565 ;
      RECT 9946.295 187.44 9948.815 8613.565 ;
      RECT 9942.655 187.44 9945.175 8613.565 ;
      RECT 9879.935 187.44 9937.895 8613.565 ;
      RECT 9876.015 187.44 9878.815 8613.565 ;
      RECT 9872.095 187.44 9874.895 8613.565 ;
      RECT 9868.175 187.44 9870.975 8613.565 ;
      RECT 9864.255 187.44 9867.055 8613.565 ;
      RECT 9817.215 187.44 9863.135 8613.565 ;
      RECT 9813.575 187.44 9816.095 8613.565 ;
      RECT 9809.935 187.44 9812.455 8613.565 ;
      RECT 9806.295 187.44 9808.815 8613.565 ;
      RECT 9802.655 187.44 9805.175 8613.565 ;
      RECT 9739.935 187.44 9797.895 8613.565 ;
      RECT 9736.015 187.44 9738.815 8613.565 ;
      RECT 9732.095 187.44 9734.895 8613.565 ;
      RECT 9728.175 187.44 9730.975 8613.565 ;
      RECT 9724.255 187.44 9727.055 8613.565 ;
      RECT 9677.215 187.44 9723.135 8613.565 ;
      RECT 9673.575 187.44 9676.095 8613.565 ;
      RECT 9669.935 187.44 9672.455 8613.565 ;
      RECT 9666.295 187.44 9668.815 8613.565 ;
      RECT 9662.655 187.44 9665.175 8613.565 ;
      RECT 9599.935 187.44 9657.895 8613.565 ;
      RECT 9596.015 187.44 9598.815 8613.565 ;
      RECT 9592.095 187.44 9594.895 8613.565 ;
      RECT 9588.175 187.44 9590.975 8613.565 ;
      RECT 9584.255 187.44 9587.055 8613.565 ;
      RECT 9537.215 187.44 9583.135 8613.565 ;
      RECT 9533.575 187.44 9536.095 8613.565 ;
      RECT 9529.935 187.44 9532.455 8613.565 ;
      RECT 9526.295 187.44 9528.815 8613.565 ;
      RECT 9522.655 187.44 9525.175 8613.565 ;
      RECT 9459.935 187.44 9517.895 8613.565 ;
      RECT 9456.015 187.44 9458.815 8613.565 ;
      RECT 9452.095 187.44 9454.895 8613.565 ;
      RECT 9448.175 187.44 9450.975 8613.565 ;
      RECT 9444.255 187.44 9447.055 8613.565 ;
      RECT 9432.615 187.44 9443.135 8613.565 ;
      RECT 9430.935 187.44 9431.215 8613.565 ;
      RECT 9429.255 187.44 9429.535 8613.565 ;
      RECT 9427.575 187.44 9427.855 8613.565 ;
      RECT 9425.895 187.44 9426.175 8613.565 ;
      RECT 9424.215 187.44 9424.495 8613.565 ;
      RECT 9422.535 187.44 9422.815 8613.565 ;
      RECT 9420.855 187.44 9421.135 8613.565 ;
      RECT 9397.215 187.44 9407.695 8613.565 ;
      RECT 9393.575 187.44 9396.095 8613.565 ;
      RECT 9389.935 187.44 9392.455 8613.565 ;
      RECT 9386.295 187.44 9388.815 8613.565 ;
      RECT 9382.655 187.44 9385.175 8613.565 ;
      RECT 9319.935 187.44 9377.895 8613.565 ;
      RECT 9316.015 187.44 9318.815 8613.565 ;
      RECT 9312.095 187.44 9314.895 8613.565 ;
      RECT 9308.175 187.44 9310.975 8613.565 ;
      RECT 9304.255 187.44 9307.055 8613.565 ;
      RECT 9257.215 187.44 9303.135 8613.565 ;
      RECT 9253.575 187.44 9256.095 8613.565 ;
      RECT 9249.935 187.44 9252.455 8613.565 ;
      RECT 9246.295 187.44 9248.815 8613.565 ;
      RECT 9242.655 187.44 9245.175 8613.565 ;
      RECT 9179.935 187.44 9237.895 8613.565 ;
      RECT 9176.015 187.44 9178.815 8613.565 ;
      RECT 9172.095 187.44 9174.895 8613.565 ;
      RECT 9168.175 187.44 9170.975 8613.565 ;
      RECT 9164.255 187.44 9167.055 8613.565 ;
      RECT 9117.215 187.44 9163.135 8613.565 ;
      RECT 9113.575 187.44 9116.095 8613.565 ;
      RECT 9109.935 187.44 9112.455 8613.565 ;
      RECT 9106.295 187.44 9108.815 8613.565 ;
      RECT 9102.655 187.44 9105.175 8613.565 ;
      RECT 9039.935 187.44 9097.895 8613.565 ;
      RECT 9036.015 187.44 9038.815 8613.565 ;
      RECT 9032.095 187.44 9034.895 8613.565 ;
      RECT 9028.175 187.44 9030.975 8613.565 ;
      RECT 9024.255 187.44 9027.055 8613.565 ;
      RECT 8977.215 187.44 9023.135 8613.565 ;
      RECT 8973.575 187.44 8976.095 8613.565 ;
      RECT 8969.935 187.44 8972.455 8613.565 ;
      RECT 8966.295 187.44 8968.815 8613.565 ;
      RECT 8962.655 187.44 8965.175 8613.565 ;
      RECT 8899.935 187.44 8957.895 8613.565 ;
      RECT 8896.015 187.44 8898.815 8613.565 ;
      RECT 8892.095 187.44 8894.895 8613.565 ;
      RECT 8888.175 187.44 8890.975 8613.565 ;
      RECT 8884.255 187.44 8887.055 8613.565 ;
      RECT 8837.215 187.44 8883.135 8613.565 ;
      RECT 8833.575 187.44 8836.095 8613.565 ;
      RECT 8829.935 187.44 8832.455 8613.565 ;
      RECT 8826.295 187.44 8828.815 8613.565 ;
      RECT 8822.655 187.44 8825.175 8613.565 ;
      RECT 8759.935 187.44 8817.895 8613.565 ;
      RECT 8756.015 187.44 8758.815 8613.565 ;
      RECT 8752.095 187.44 8754.895 8613.565 ;
      RECT 8748.175 187.44 8750.975 8613.565 ;
      RECT 8744.255 187.44 8747.055 8613.565 ;
      RECT 8697.215 187.44 8743.135 8613.565 ;
      RECT 8693.575 187.44 8696.095 8613.565 ;
      RECT 8689.935 187.44 8692.455 8613.565 ;
      RECT 8686.295 187.44 8688.815 8613.565 ;
      RECT 8682.655 187.44 8685.175 8613.565 ;
      RECT 8619.935 187.44 8677.895 8613.565 ;
      RECT 8616.015 187.44 8618.815 8613.565 ;
      RECT 8612.095 187.44 8614.895 8613.565 ;
      RECT 8608.175 187.44 8610.975 8613.565 ;
      RECT 8604.255 187.44 8607.055 8613.565 ;
      RECT 8557.215 187.44 8603.135 8613.565 ;
      RECT 8553.575 187.44 8556.095 8613.565 ;
      RECT 8549.935 187.44 8552.455 8613.565 ;
      RECT 8546.295 187.44 8548.815 8613.565 ;
      RECT 8542.655 187.44 8545.175 8613.565 ;
      RECT 8479.935 187.44 8537.895 8613.565 ;
      RECT 8476.015 187.44 8478.815 8613.565 ;
      RECT 8472.095 187.44 8474.895 8613.565 ;
      RECT 8468.175 187.44 8470.975 8613.565 ;
      RECT 8464.255 187.44 8467.055 8613.565 ;
      RECT 8417.215 187.44 8463.135 8613.565 ;
      RECT 8413.575 187.44 8416.095 8613.565 ;
      RECT 8409.935 187.44 8412.455 8613.565 ;
      RECT 8406.295 187.44 8408.815 8613.565 ;
      RECT 8402.655 187.44 8405.175 8613.565 ;
      RECT 8339.935 187.44 8397.895 8613.565 ;
      RECT 8336.015 187.44 8338.815 8613.565 ;
      RECT 8332.095 187.44 8334.895 8613.565 ;
      RECT 8328.175 187.44 8330.975 8613.565 ;
      RECT 8324.255 187.44 8327.055 8613.565 ;
      RECT 8277.215 187.44 8323.135 8613.565 ;
      RECT 8273.575 187.44 8276.095 8613.565 ;
      RECT 8269.935 187.44 8272.455 8613.565 ;
      RECT 8266.295 187.44 8268.815 8613.565 ;
      RECT 8262.655 187.44 8265.175 8613.565 ;
      RECT 8199.935 187.44 8257.895 8613.565 ;
      RECT 8196.015 187.44 8198.815 8613.565 ;
      RECT 8192.095 187.44 8194.895 8613.565 ;
      RECT 8188.175 187.44 8190.975 8613.565 ;
      RECT 8184.255 187.44 8187.055 8613.565 ;
      RECT 8137.215 187.44 8183.135 8613.565 ;
      RECT 8133.575 187.44 8136.095 8613.565 ;
      RECT 8129.935 187.44 8132.455 8613.565 ;
      RECT 8126.295 187.44 8128.815 8613.565 ;
      RECT 8122.655 187.44 8125.175 8613.565 ;
      RECT 8059.935 187.44 8117.895 8613.565 ;
      RECT 8056.015 187.44 8058.815 8613.565 ;
      RECT 8052.095 187.44 8054.895 8613.565 ;
      RECT 8048.175 187.44 8050.975 8613.565 ;
      RECT 8044.255 187.44 8047.055 8613.565 ;
      RECT 7997.215 187.44 8043.135 8613.565 ;
      RECT 7993.575 187.44 7996.095 8613.565 ;
      RECT 7989.935 187.44 7992.455 8613.565 ;
      RECT 7986.295 187.44 7988.815 8613.565 ;
      RECT 7982.655 187.44 7985.175 8613.565 ;
      RECT 7919.935 187.44 7977.895 8613.565 ;
      RECT 7916.015 187.44 7918.815 8613.565 ;
      RECT 7912.095 187.44 7914.895 8613.565 ;
      RECT 7908.175 187.44 7910.975 8613.565 ;
      RECT 7904.255 187.44 7907.055 8613.565 ;
      RECT 7857.215 187.44 7903.135 8613.565 ;
      RECT 7853.575 187.44 7856.095 8613.565 ;
      RECT 7849.935 187.44 7852.455 8613.565 ;
      RECT 7846.295 187.44 7848.815 8613.565 ;
      RECT 7842.655 187.44 7845.175 8613.565 ;
      RECT 7779.935 187.44 7837.895 8613.565 ;
      RECT 7776.015 187.44 7778.815 8613.565 ;
      RECT 7772.095 187.44 7774.895 8613.565 ;
      RECT 7768.175 187.44 7770.975 8613.565 ;
      RECT 7764.255 187.44 7767.055 8613.565 ;
      RECT 7717.215 187.44 7763.135 8613.565 ;
      RECT 7713.575 187.44 7716.095 8613.565 ;
      RECT 7709.935 187.44 7712.455 8613.565 ;
      RECT 7706.295 187.44 7708.815 8613.565 ;
      RECT 7702.655 187.44 7705.175 8613.565 ;
      RECT 7639.935 187.44 7697.895 8613.565 ;
      RECT 7636.015 187.44 7638.815 8613.565 ;
      RECT 7632.095 187.44 7634.895 8613.565 ;
      RECT 7628.175 187.44 7630.975 8613.565 ;
      RECT 7624.255 187.44 7627.055 8613.565 ;
      RECT 7577.215 187.44 7623.135 8613.565 ;
      RECT 7573.575 187.44 7576.095 8613.565 ;
      RECT 7569.935 187.44 7572.455 8613.565 ;
      RECT 7566.295 187.44 7568.815 8613.565 ;
      RECT 7562.655 187.44 7565.175 8613.565 ;
      RECT 7499.935 187.44 7557.895 8613.565 ;
      RECT 7496.015 187.44 7498.815 8613.565 ;
      RECT 7492.095 187.44 7494.895 8613.565 ;
      RECT 7488.175 187.44 7490.975 8613.565 ;
      RECT 7484.255 187.44 7487.055 8613.565 ;
      RECT 7437.215 187.44 7483.135 8613.565 ;
      RECT 7433.575 187.44 7436.095 8613.565 ;
      RECT 7429.935 187.44 7432.455 8613.565 ;
      RECT 7426.295 187.44 7428.815 8613.565 ;
      RECT 7422.655 187.44 7425.175 8613.565 ;
      RECT 7359.935 187.44 7417.895 8613.565 ;
      RECT 7356.015 187.44 7358.815 8613.565 ;
      RECT 7352.095 187.44 7354.895 8613.565 ;
      RECT 7348.175 187.44 7350.975 8613.565 ;
      RECT 7344.255 187.44 7347.055 8613.565 ;
      RECT 7297.215 187.44 7343.135 8613.565 ;
      RECT 7293.575 187.44 7296.095 8613.565 ;
      RECT 7289.935 187.44 7292.455 8613.565 ;
      RECT 7286.295 187.44 7288.815 8613.565 ;
      RECT 7282.655 187.44 7285.175 8613.565 ;
      RECT 7219.935 187.44 7277.895 8613.565 ;
      RECT 7216.015 187.44 7218.815 8613.565 ;
      RECT 7212.095 187.44 7214.895 8613.565 ;
      RECT 7208.175 187.44 7210.975 8613.565 ;
      RECT 7204.255 187.44 7207.055 8613.565 ;
      RECT 7157.215 187.44 7203.135 8613.565 ;
      RECT 7153.575 187.44 7156.095 8613.565 ;
      RECT 7149.935 187.44 7152.455 8613.565 ;
      RECT 7146.295 187.44 7148.815 8613.565 ;
      RECT 7142.655 187.44 7145.175 8613.565 ;
      RECT 7079.935 187.44 7137.895 8613.565 ;
      RECT 7076.015 187.44 7078.815 8613.565 ;
      RECT 7072.095 187.44 7074.895 8613.565 ;
      RECT 7068.175 187.44 7070.975 8613.565 ;
      RECT 7064.255 187.44 7067.055 8613.565 ;
      RECT 7017.215 187.44 7063.135 8613.565 ;
      RECT 7013.575 187.44 7016.095 8613.565 ;
      RECT 7009.935 187.44 7012.455 8613.565 ;
      RECT 7006.295 187.44 7008.815 8613.565 ;
      RECT 7002.655 187.44 7005.175 8613.565 ;
      RECT 6939.935 187.44 6997.895 8613.565 ;
      RECT 6936.015 187.44 6938.815 8613.565 ;
      RECT 6932.095 187.44 6934.895 8613.565 ;
      RECT 6928.175 187.44 6930.975 8613.565 ;
      RECT 6924.255 187.44 6927.055 8613.565 ;
      RECT 6877.215 187.44 6923.135 8613.565 ;
      RECT 6873.575 187.44 6876.095 8613.565 ;
      RECT 6869.935 187.44 6872.455 8613.565 ;
      RECT 6866.295 187.44 6868.815 8613.565 ;
      RECT 6862.655 187.44 6865.175 8613.565 ;
      RECT 6799.935 187.44 6857.895 8613.565 ;
      RECT 6796.015 187.44 6798.815 8613.565 ;
      RECT 6792.095 187.44 6794.895 8613.565 ;
      RECT 6788.175 187.44 6790.975 8613.565 ;
      RECT 6784.255 187.44 6787.055 8613.565 ;
      RECT 6737.215 187.44 6783.135 8613.565 ;
      RECT 6733.575 187.44 6736.095 8613.565 ;
      RECT 6729.935 187.44 6732.455 8613.565 ;
      RECT 6726.295 187.44 6728.815 8613.565 ;
      RECT 6722.655 187.44 6725.175 8613.565 ;
      RECT 6659.935 187.44 6717.895 8613.565 ;
      RECT 6656.015 187.44 6658.815 8613.565 ;
      RECT 6652.095 187.44 6654.895 8613.565 ;
      RECT 6648.175 187.44 6650.975 8613.565 ;
      RECT 6644.255 187.44 6647.055 8613.565 ;
      RECT 6597.215 187.44 6643.135 8613.565 ;
      RECT 6593.575 187.44 6596.095 8613.565 ;
      RECT 6589.935 187.44 6592.455 8613.565 ;
      RECT 6586.295 187.44 6588.815 8613.565 ;
      RECT 6582.655 187.44 6585.175 8613.565 ;
      RECT 6519.935 187.44 6577.895 8613.565 ;
      RECT 6516.015 187.44 6518.815 8613.565 ;
      RECT 6512.095 187.44 6514.895 8613.565 ;
      RECT 6508.175 187.44 6510.975 8613.565 ;
      RECT 6504.255 187.44 6507.055 8613.565 ;
      RECT 6457.215 187.44 6503.135 8613.565 ;
      RECT 6453.575 187.44 6456.095 8613.565 ;
      RECT 6449.935 187.44 6452.455 8613.565 ;
      RECT 6446.295 187.44 6448.815 8613.565 ;
      RECT 6442.655 187.44 6445.175 8613.565 ;
      RECT 6379.935 187.44 6437.895 8613.565 ;
      RECT 6376.015 187.44 6378.815 8613.565 ;
      RECT 6372.095 187.44 6374.895 8613.565 ;
      RECT 6368.175 187.44 6370.975 8613.565 ;
      RECT 6364.255 187.44 6367.055 8613.565 ;
      RECT 6317.215 187.44 6363.135 8613.565 ;
      RECT 6313.575 187.44 6316.095 8613.565 ;
      RECT 6309.935 187.44 6312.455 8613.565 ;
      RECT 6306.295 187.44 6308.815 8613.565 ;
      RECT 6302.655 187.44 6305.175 8613.565 ;
      RECT 6239.935 187.44 6297.895 8613.565 ;
      RECT 6236.015 187.44 6238.815 8613.565 ;
      RECT 6232.095 187.44 6234.895 8613.565 ;
      RECT 6228.175 187.44 6230.975 8613.565 ;
      RECT 6224.255 187.44 6227.055 8613.565 ;
      RECT 6177.215 187.44 6223.135 8613.565 ;
      RECT 6173.575 187.44 6176.095 8613.565 ;
      RECT 6169.935 187.44 6172.455 8613.565 ;
      RECT 6166.295 187.44 6168.815 8613.565 ;
      RECT 6162.655 187.44 6165.175 8613.565 ;
      RECT 6099.935 187.44 6157.895 8613.565 ;
      RECT 6096.015 187.44 6098.815 8613.565 ;
      RECT 6092.095 187.44 6094.895 8613.565 ;
      RECT 6088.175 187.44 6090.975 8613.565 ;
      RECT 6084.255 187.44 6087.055 8613.565 ;
      RECT 6037.215 187.44 6083.135 8613.565 ;
      RECT 6033.575 187.44 6036.095 8613.565 ;
      RECT 6029.935 187.44 6032.455 8613.565 ;
      RECT 6026.295 187.44 6028.815 8613.565 ;
      RECT 6022.655 187.44 6025.175 8613.565 ;
      RECT 5959.935 187.44 6017.895 8613.565 ;
      RECT 5956.015 187.44 5958.815 8613.565 ;
      RECT 5952.095 187.44 5954.895 8613.565 ;
      RECT 5948.175 187.44 5950.975 8613.565 ;
      RECT 5944.255 187.44 5947.055 8613.565 ;
      RECT 5897.215 187.44 5943.135 8613.565 ;
      RECT 5893.575 187.44 5896.095 8613.565 ;
      RECT 5889.935 187.44 5892.455 8613.565 ;
      RECT 5886.295 187.44 5888.815 8613.565 ;
      RECT 5882.655 187.44 5885.175 8613.565 ;
      RECT 5819.935 187.44 5877.895 8613.565 ;
      RECT 5816.015 187.44 5818.815 8613.565 ;
      RECT 5812.095 187.44 5814.895 8613.565 ;
      RECT 5808.175 187.44 5810.975 8613.565 ;
      RECT 5804.255 187.44 5807.055 8613.565 ;
      RECT 5757.215 187.44 5803.135 8613.565 ;
      RECT 5753.575 187.44 5756.095 8613.565 ;
      RECT 5749.935 187.44 5752.455 8613.565 ;
      RECT 5746.295 187.44 5748.815 8613.565 ;
      RECT 5742.655 187.44 5745.175 8613.565 ;
      RECT 5679.935 187.44 5737.895 8613.565 ;
      RECT 5676.015 187.44 5678.815 8613.565 ;
      RECT 5672.095 187.44 5674.895 8613.565 ;
      RECT 5668.175 187.44 5670.975 8613.565 ;
      RECT 5664.255 187.44 5667.055 8613.565 ;
      RECT 5617.215 187.44 5663.135 8613.565 ;
      RECT 5613.575 187.44 5616.095 8613.565 ;
      RECT 5609.935 187.44 5612.455 8613.565 ;
      RECT 5606.295 187.44 5608.815 8613.565 ;
      RECT 5602.655 187.44 5605.175 8613.565 ;
      RECT 5539.935 187.44 5597.895 8613.565 ;
      RECT 5536.015 187.44 5538.815 8613.565 ;
      RECT 5532.095 187.44 5534.895 8613.565 ;
      RECT 5528.175 187.44 5530.975 8613.565 ;
      RECT 5524.255 187.44 5527.055 8613.565 ;
      RECT 5477.215 187.44 5523.135 8613.565 ;
      RECT 5473.575 187.44 5476.095 8613.565 ;
      RECT 5469.935 187.44 5472.455 8613.565 ;
      RECT 5466.295 187.44 5468.815 8613.565 ;
      RECT 5462.655 187.44 5465.175 8613.565 ;
      RECT 5399.935 187.44 5457.895 8613.565 ;
      RECT 5396.015 187.44 5398.815 8613.565 ;
      RECT 5392.095 187.44 5394.895 8613.565 ;
      RECT 5388.175 187.44 5390.975 8613.565 ;
      RECT 5384.255 187.44 5387.055 8613.565 ;
      RECT 5337.215 187.44 5383.135 8613.565 ;
      RECT 5333.575 187.44 5336.095 8613.565 ;
      RECT 5329.935 187.44 5332.455 8613.565 ;
      RECT 5326.295 187.44 5328.815 8613.565 ;
      RECT 5322.655 187.44 5325.175 8613.565 ;
      RECT 5259.935 187.44 5317.895 8613.565 ;
      RECT 5256.015 187.44 5258.815 8613.565 ;
      RECT 5252.095 187.44 5254.895 8613.565 ;
      RECT 5248.175 187.44 5250.975 8613.565 ;
      RECT 5244.255 187.44 5247.055 8613.565 ;
      RECT 5197.215 187.44 5243.135 8613.565 ;
      RECT 5193.575 187.44 5196.095 8613.565 ;
      RECT 5189.935 187.44 5192.455 8613.565 ;
      RECT 5186.295 187.44 5188.815 8613.565 ;
      RECT 5182.655 187.44 5185.175 8613.565 ;
      RECT 5119.935 187.44 5177.895 8613.565 ;
      RECT 5116.015 187.44 5118.815 8613.565 ;
      RECT 5112.095 187.44 5114.895 8613.565 ;
      RECT 5108.175 187.44 5110.975 8613.565 ;
      RECT 5104.255 187.44 5107.055 8613.565 ;
      RECT 5057.215 187.44 5103.135 8613.565 ;
      RECT 5053.575 187.44 5056.095 8613.565 ;
      RECT 5049.935 187.44 5052.455 8613.565 ;
      RECT 5046.295 187.44 5048.815 8613.565 ;
      RECT 5042.655 187.44 5045.175 8613.565 ;
      RECT 4979.935 187.44 5037.895 8613.565 ;
      RECT 4976.015 187.44 4978.815 8613.565 ;
      RECT 4972.095 187.44 4974.895 8613.565 ;
      RECT 4968.175 187.44 4970.975 8613.565 ;
      RECT 4964.255 187.44 4967.055 8613.565 ;
      RECT 4917.215 187.44 4963.135 8613.565 ;
      RECT 4913.575 187.44 4916.095 8613.565 ;
      RECT 4909.935 187.44 4912.455 8613.565 ;
      RECT 4906.295 187.44 4908.815 8613.565 ;
      RECT 4902.655 187.44 4905.175 8613.565 ;
      RECT 4839.935 187.44 4897.895 8613.565 ;
      RECT 4836.015 187.44 4838.815 8613.565 ;
      RECT 4832.095 187.44 4834.895 8613.565 ;
      RECT 4828.175 187.44 4830.975 8613.565 ;
      RECT 4824.255 187.44 4827.055 8613.565 ;
      RECT 4777.215 187.44 4823.135 8613.565 ;
      RECT 4773.575 187.44 4776.095 8613.565 ;
      RECT 4769.935 187.44 4772.455 8613.565 ;
      RECT 4766.295 187.44 4768.815 8613.565 ;
      RECT 4762.655 187.44 4765.175 8613.565 ;
      RECT 4699.935 187.44 4757.895 8613.565 ;
      RECT 4696.015 187.44 4698.815 8613.565 ;
      RECT 4692.095 187.44 4694.895 8613.565 ;
      RECT 4688.175 187.44 4690.975 8613.565 ;
      RECT 4684.255 187.44 4687.055 8613.565 ;
      RECT 4637.215 187.44 4683.135 8613.565 ;
      RECT 4633.575 187.44 4636.095 8613.565 ;
      RECT 4629.935 187.44 4632.455 8613.565 ;
      RECT 4626.295 187.44 4628.815 8613.565 ;
      RECT 4622.655 187.44 4625.175 8613.565 ;
      RECT 4559.935 187.44 4617.895 8613.565 ;
      RECT 4556.015 187.44 4558.815 8613.565 ;
      RECT 4552.095 187.44 4554.895 8613.565 ;
      RECT 4548.175 187.44 4550.975 8613.565 ;
      RECT 4544.255 187.44 4547.055 8613.565 ;
      RECT 4497.215 187.44 4543.135 8613.565 ;
      RECT 4493.575 187.44 4496.095 8613.565 ;
      RECT 4489.935 187.44 4492.455 8613.565 ;
      RECT 4486.295 187.44 4488.815 8613.565 ;
      RECT 4482.655 187.44 4485.175 8613.565 ;
      RECT 4419.935 187.44 4477.895 8613.565 ;
      RECT 4416.015 187.44 4418.815 8613.565 ;
      RECT 4412.095 187.44 4414.895 8613.565 ;
      RECT 4408.175 187.44 4410.975 8613.565 ;
      RECT 4404.255 187.44 4407.055 8613.565 ;
      RECT 4357.215 187.44 4403.135 8613.565 ;
      RECT 4353.575 187.44 4356.095 8613.565 ;
      RECT 4349.935 187.44 4352.455 8613.565 ;
      RECT 4346.295 187.44 4348.815 8613.565 ;
      RECT 4342.655 187.44 4345.175 8613.565 ;
      RECT 4279.935 187.44 4337.895 8613.565 ;
      RECT 4276.015 187.44 4278.815 8613.565 ;
      RECT 4272.095 187.44 4274.895 8613.565 ;
      RECT 4268.175 187.44 4270.975 8613.565 ;
      RECT 4264.255 187.44 4267.055 8613.565 ;
      RECT 4217.215 187.44 4263.135 8613.565 ;
      RECT 4213.575 187.44 4216.095 8613.565 ;
      RECT 4209.935 187.44 4212.455 8613.565 ;
      RECT 4206.295 187.44 4208.815 8613.565 ;
      RECT 4202.655 187.44 4205.175 8613.565 ;
      RECT 4139.935 187.44 4197.895 8613.565 ;
      RECT 4136.015 187.44 4138.815 8613.565 ;
      RECT 4132.095 187.44 4134.895 8613.565 ;
      RECT 4128.175 187.44 4130.975 8613.565 ;
      RECT 4124.255 187.44 4127.055 8613.565 ;
      RECT 4077.215 187.44 4123.135 8613.565 ;
      RECT 4073.575 187.44 4076.095 8613.565 ;
      RECT 4069.935 187.44 4072.455 8613.565 ;
      RECT 4066.295 187.44 4068.815 8613.565 ;
      RECT 4062.655 187.44 4065.175 8613.565 ;
      RECT 3999.935 187.44 4057.895 8613.565 ;
      RECT 3996.015 187.44 3998.815 8613.565 ;
      RECT 3992.095 187.44 3994.895 8613.565 ;
      RECT 3988.175 187.44 3990.975 8613.565 ;
      RECT 3984.255 187.44 3987.055 8613.565 ;
      RECT 3937.215 187.44 3983.135 8613.565 ;
      RECT 3933.575 187.44 3936.095 8613.565 ;
      RECT 3929.935 187.44 3932.455 8613.565 ;
      RECT 3926.295 187.44 3928.815 8613.565 ;
      RECT 3922.655 187.44 3925.175 8613.565 ;
      RECT 3859.935 187.44 3917.895 8613.565 ;
      RECT 3856.015 187.44 3858.815 8613.565 ;
      RECT 3852.095 187.44 3854.895 8613.565 ;
      RECT 3848.175 187.44 3850.975 8613.565 ;
      RECT 3844.255 187.44 3847.055 8613.565 ;
      RECT 3797.215 187.44 3843.135 8613.565 ;
      RECT 3793.575 187.44 3796.095 8613.565 ;
      RECT 3789.935 187.44 3792.455 8613.565 ;
      RECT 3786.295 187.44 3788.815 8613.565 ;
      RECT 3782.655 187.44 3785.175 8613.565 ;
      RECT 3719.935 187.44 3777.895 8613.565 ;
      RECT 3716.015 187.44 3718.815 8613.565 ;
      RECT 3712.095 187.44 3714.895 8613.565 ;
      RECT 3708.175 187.44 3710.975 8613.565 ;
      RECT 3704.255 187.44 3707.055 8613.565 ;
      RECT 3657.215 187.44 3703.135 8613.565 ;
      RECT 3653.575 187.44 3656.095 8613.565 ;
      RECT 3649.935 187.44 3652.455 8613.565 ;
      RECT 3646.295 187.44 3648.815 8613.565 ;
      RECT 3642.655 187.44 3645.175 8613.565 ;
      RECT 3579.935 187.44 3637.895 8613.565 ;
      RECT 3576.015 187.44 3578.815 8613.565 ;
      RECT 3572.095 187.44 3574.895 8613.565 ;
      RECT 3568.175 187.44 3570.975 8613.565 ;
      RECT 3564.255 187.44 3567.055 8613.565 ;
      RECT 3517.215 187.44 3563.135 8613.565 ;
      RECT 3513.575 187.44 3516.095 8613.565 ;
      RECT 3509.935 187.44 3512.455 8613.565 ;
      RECT 3506.295 187.44 3508.815 8613.565 ;
      RECT 3502.655 187.44 3505.175 8613.565 ;
      RECT 3439.935 187.44 3497.895 8613.565 ;
      RECT 3436.015 187.44 3438.815 8613.565 ;
      RECT 3432.095 187.44 3434.895 8613.565 ;
      RECT 3428.175 187.44 3430.975 8613.565 ;
      RECT 3424.255 187.44 3427.055 8613.565 ;
      RECT 3377.215 187.44 3423.135 8613.565 ;
      RECT 3373.575 187.44 3376.095 8613.565 ;
      RECT 3369.935 187.44 3372.455 8613.565 ;
      RECT 3366.295 187.44 3368.815 8613.565 ;
      RECT 3362.655 187.44 3365.175 8613.565 ;
      RECT 3299.935 187.44 3357.895 8613.565 ;
      RECT 3296.015 187.44 3298.815 8613.565 ;
      RECT 3292.095 187.44 3294.895 8613.565 ;
      RECT 3288.175 187.44 3290.975 8613.565 ;
      RECT 3284.255 187.44 3287.055 8613.565 ;
      RECT 3237.215 187.44 3283.135 8613.565 ;
      RECT 3233.575 187.44 3236.095 8613.565 ;
      RECT 3229.935 187.44 3232.455 8613.565 ;
      RECT 3226.295 187.44 3228.815 8613.565 ;
      RECT 3222.655 187.44 3225.175 8613.565 ;
      RECT 3159.935 187.44 3217.895 8613.565 ;
      RECT 3156.015 187.44 3158.815 8613.565 ;
      RECT 3152.095 187.44 3154.895 8613.565 ;
      RECT 3148.175 187.44 3150.975 8613.565 ;
      RECT 3144.255 187.44 3147.055 8613.565 ;
      RECT 3097.215 187.44 3143.135 8613.565 ;
      RECT 3093.575 187.44 3096.095 8613.565 ;
      RECT 3089.935 187.44 3092.455 8613.565 ;
      RECT 3086.295 187.44 3088.815 8613.565 ;
      RECT 3082.655 187.44 3085.175 8613.565 ;
      RECT 3019.935 187.44 3077.895 8613.565 ;
      RECT 3016.015 187.44 3018.815 8613.565 ;
      RECT 3012.095 187.44 3014.895 8613.565 ;
      RECT 3008.175 187.44 3010.975 8613.565 ;
      RECT 3004.255 187.44 3007.055 8613.565 ;
      RECT 2957.215 187.44 3003.135 8613.565 ;
      RECT 2953.575 187.44 2956.095 8613.565 ;
      RECT 2949.935 187.44 2952.455 8613.565 ;
      RECT 2946.295 187.44 2948.815 8613.565 ;
      RECT 2942.655 187.44 2945.175 8613.565 ;
      RECT 2879.935 187.44 2937.895 8613.565 ;
      RECT 2876.015 187.44 2878.815 8613.565 ;
      RECT 2872.095 187.44 2874.895 8613.565 ;
      RECT 2868.175 187.44 2870.975 8613.565 ;
      RECT 2864.255 187.44 2867.055 8613.565 ;
      RECT 2817.215 187.44 2863.135 8613.565 ;
      RECT 2813.575 187.44 2816.095 8613.565 ;
      RECT 2809.935 187.44 2812.455 8613.565 ;
      RECT 2806.295 187.44 2808.815 8613.565 ;
      RECT 2802.655 187.44 2805.175 8613.565 ;
      RECT 2739.935 187.44 2797.895 8613.565 ;
      RECT 2736.015 187.44 2738.815 8613.565 ;
      RECT 2732.095 187.44 2734.895 8613.565 ;
      RECT 2728.175 187.44 2730.975 8613.565 ;
      RECT 2724.255 187.44 2727.055 8613.565 ;
      RECT 2677.215 187.44 2723.135 8613.565 ;
      RECT 2673.575 187.44 2676.095 8613.565 ;
      RECT 2669.935 187.44 2672.455 8613.565 ;
      RECT 2666.295 187.44 2668.815 8613.565 ;
      RECT 2662.655 187.44 2665.175 8613.565 ;
      RECT 2599.935 187.44 2657.895 8613.565 ;
      RECT 2596.015 187.44 2598.815 8613.565 ;
      RECT 2592.095 187.44 2594.895 8613.565 ;
      RECT 2588.175 187.44 2590.975 8613.565 ;
      RECT 2584.255 187.44 2587.055 8613.565 ;
      RECT 2537.215 187.44 2583.135 8613.565 ;
      RECT 2533.575 187.44 2536.095 8613.565 ;
      RECT 2529.935 187.44 2532.455 8613.565 ;
      RECT 2526.295 187.44 2528.815 8613.565 ;
      RECT 2522.655 187.44 2525.175 8613.565 ;
      RECT 2459.935 187.44 2517.895 8613.565 ;
      RECT 2456.015 187.44 2458.815 8613.565 ;
      RECT 2452.095 187.44 2454.895 8613.565 ;
      RECT 2448.175 187.44 2450.975 8613.565 ;
      RECT 2444.255 187.44 2447.055 8613.565 ;
      RECT 2397.215 187.44 2443.135 8613.565 ;
      RECT 2393.575 187.44 2396.095 8613.565 ;
      RECT 2389.935 187.44 2392.455 8613.565 ;
      RECT 2386.295 187.44 2388.815 8613.565 ;
      RECT 2382.655 187.44 2385.175 8613.565 ;
      RECT 2319.935 187.44 2377.895 8613.565 ;
      RECT 2316.015 187.44 2318.815 8613.565 ;
      RECT 2312.095 187.44 2314.895 8613.565 ;
      RECT 2308.175 187.44 2310.975 8613.565 ;
      RECT 2304.255 187.44 2307.055 8613.565 ;
      RECT 2257.215 187.44 2303.135 8613.565 ;
      RECT 2253.575 187.44 2256.095 8613.565 ;
      RECT 2249.935 187.44 2252.455 8613.565 ;
      RECT 2246.295 187.44 2248.815 8613.565 ;
      RECT 2242.655 187.44 2245.175 8613.565 ;
      RECT 2179.935 187.44 2237.895 8613.565 ;
      RECT 2176.015 187.44 2178.815 8613.565 ;
      RECT 2172.095 187.44 2174.895 8613.565 ;
      RECT 2168.175 187.44 2170.975 8613.565 ;
      RECT 2164.255 187.44 2167.055 8613.565 ;
      RECT 2117.215 187.44 2163.135 8613.565 ;
      RECT 2113.575 187.44 2116.095 8613.565 ;
      RECT 2109.935 187.44 2112.455 8613.565 ;
      RECT 2106.295 187.44 2108.815 8613.565 ;
      RECT 2102.655 187.44 2105.175 8613.565 ;
      RECT 2039.935 187.44 2097.895 8613.565 ;
      RECT 2036.015 187.44 2038.815 8613.565 ;
      RECT 2032.095 187.44 2034.895 8613.565 ;
      RECT 2028.175 187.44 2030.975 8613.565 ;
      RECT 2024.255 187.44 2027.055 8613.565 ;
      RECT 1977.215 187.44 2023.135 8613.565 ;
      RECT 1973.575 187.44 1976.095 8613.565 ;
      RECT 1969.935 187.44 1972.455 8613.565 ;
      RECT 1966.295 187.44 1968.815 8613.565 ;
      RECT 1962.655 187.44 1965.175 8613.565 ;
      RECT 1899.935 187.44 1957.895 8613.565 ;
      RECT 1896.015 187.44 1898.815 8613.565 ;
      RECT 1892.095 187.44 1894.895 8613.565 ;
      RECT 1888.175 187.44 1890.975 8613.565 ;
      RECT 1884.255 187.44 1887.055 8613.565 ;
      RECT 1837.215 187.44 1883.135 8613.565 ;
      RECT 1833.575 187.44 1836.095 8613.565 ;
      RECT 1829.935 187.44 1832.455 8613.565 ;
      RECT 1826.295 187.44 1828.815 8613.565 ;
      RECT 1822.655 187.44 1825.175 8613.565 ;
      RECT 1759.935 187.44 1817.895 8613.565 ;
      RECT 1756.015 187.44 1758.815 8613.565 ;
      RECT 1752.095 187.44 1754.895 8613.565 ;
      RECT 1748.175 187.44 1750.975 8613.565 ;
      RECT 1744.255 187.44 1747.055 8613.565 ;
      RECT 1697.215 187.44 1743.135 8613.565 ;
      RECT 1693.575 187.44 1696.095 8613.565 ;
      RECT 1689.935 187.44 1692.455 8613.565 ;
      RECT 1686.295 187.44 1688.815 8613.565 ;
      RECT 1682.655 187.44 1685.175 8613.565 ;
      RECT 1619.935 187.44 1677.895 8613.565 ;
      RECT 1616.015 187.44 1618.815 8613.565 ;
      RECT 1612.095 187.44 1614.895 8613.565 ;
      RECT 1608.175 187.44 1610.975 8613.565 ;
      RECT 1604.255 187.44 1607.055 8613.565 ;
      RECT 1557.215 187.44 1603.135 8613.565 ;
      RECT 1553.575 187.44 1556.095 8613.565 ;
      RECT 1549.935 187.44 1552.455 8613.565 ;
      RECT 1546.295 187.44 1548.815 8613.565 ;
      RECT 1542.655 187.44 1545.175 8613.565 ;
      RECT 1479.935 187.44 1537.895 8613.565 ;
      RECT 1476.015 187.44 1478.815 8613.565 ;
      RECT 1472.095 187.44 1474.895 8613.565 ;
      RECT 1468.175 187.44 1470.975 8613.565 ;
      RECT 1464.255 187.44 1467.055 8613.565 ;
      RECT 1417.215 187.44 1463.135 8613.565 ;
      RECT 1413.575 187.44 1416.095 8613.565 ;
      RECT 1409.935 187.44 1412.455 8613.565 ;
      RECT 1406.295 187.44 1408.815 8613.565 ;
      RECT 1402.655 187.44 1405.175 8613.565 ;
      RECT 1339.935 187.44 1397.895 8613.565 ;
      RECT 1336.015 187.44 1338.815 8613.565 ;
      RECT 1332.095 187.44 1334.895 8613.565 ;
      RECT 1328.175 187.44 1330.975 8613.565 ;
      RECT 1324.255 187.44 1327.055 8613.565 ;
      RECT 1277.215 187.44 1323.135 8613.565 ;
      RECT 1273.575 187.44 1276.095 8613.565 ;
      RECT 1269.935 187.44 1272.455 8613.565 ;
      RECT 1266.295 187.44 1268.815 8613.565 ;
      RECT 1262.655 187.44 1265.175 8613.565 ;
      RECT 1199.935 187.44 1257.895 8613.565 ;
      RECT 1196.015 187.44 1198.815 8613.565 ;
      RECT 1192.095 187.44 1194.895 8613.565 ;
      RECT 1188.175 187.44 1190.975 8613.565 ;
      RECT 1184.255 187.44 1187.055 8613.565 ;
      RECT 1137.215 187.44 1183.135 8613.565 ;
      RECT 1133.575 187.44 1136.095 8613.565 ;
      RECT 1129.935 187.44 1132.455 8613.565 ;
      RECT 1126.295 187.44 1128.815 8613.565 ;
      RECT 1122.655 187.44 1125.175 8613.565 ;
      RECT 1059.935 187.44 1117.895 8613.565 ;
      RECT 1056.015 187.44 1058.815 8613.565 ;
      RECT 1052.095 187.44 1054.895 8613.565 ;
      RECT 1048.175 187.44 1050.975 8613.565 ;
      RECT 1044.255 187.44 1047.055 8613.565 ;
      RECT 997.215 187.44 1043.135 8613.565 ;
      RECT 993.575 187.44 996.095 8613.565 ;
      RECT 989.935 187.44 992.455 8613.565 ;
      RECT 986.295 187.44 988.815 8613.565 ;
      RECT 982.655 187.44 985.175 8613.565 ;
      RECT 919.935 187.44 977.895 8613.565 ;
      RECT 916.015 187.44 918.815 8613.565 ;
      RECT 912.095 187.44 914.895 8613.565 ;
      RECT 908.175 187.44 910.975 8613.565 ;
      RECT 904.255 187.44 907.055 8613.565 ;
      RECT 857.215 187.44 903.135 8613.565 ;
      RECT 853.575 187.44 856.095 8613.565 ;
      RECT 849.935 187.44 852.455 8613.565 ;
      RECT 846.295 187.44 848.815 8613.565 ;
      RECT 842.655 187.44 845.175 8613.565 ;
      RECT 779.935 187.44 837.895 8613.565 ;
      RECT 776.015 187.44 778.815 8613.565 ;
      RECT 772.095 187.44 774.895 8613.565 ;
      RECT 768.175 187.44 770.975 8613.565 ;
      RECT 764.255 187.44 767.055 8613.565 ;
      RECT 717.215 187.44 763.135 8613.565 ;
      RECT 713.575 187.44 716.095 8613.565 ;
      RECT 709.935 187.44 712.455 8613.565 ;
      RECT 706.295 187.44 708.815 8613.565 ;
      RECT 702.655 187.44 705.175 8613.565 ;
      RECT 639.935 187.44 697.895 8613.565 ;
      RECT 636.015 187.44 638.815 8613.565 ;
      RECT 632.095 187.44 634.895 8613.565 ;
      RECT 628.175 187.44 630.975 8613.565 ;
      RECT 624.255 187.44 627.055 8613.565 ;
      RECT 577.215 187.44 623.135 8613.565 ;
      RECT 573.575 187.44 576.095 8613.565 ;
      RECT 569.935 187.44 572.455 8613.565 ;
      RECT 566.295 187.44 568.815 8613.565 ;
      RECT 562.655 187.44 565.175 8613.565 ;
      RECT 499.935 187.44 557.895 8613.565 ;
      RECT 496.015 187.44 498.815 8613.565 ;
      RECT 492.095 187.44 494.895 8613.565 ;
      RECT 488.175 187.44 490.975 8613.565 ;
      RECT 484.255 187.44 487.055 8613.565 ;
      RECT 337.025 187.44 483.135 8613.565 ;
    LAYER M4 ;
      RECT 18465.79 8399.58 18488.86 8401 ;
      RECT 18465.79 8438.095 18488.86 8439.515 ;
      RECT 18465.79 8471.58 18488.86 8473 ;
      RECT 18465.79 8510.095 18488.86 8511.515 ;
      RECT 18465.79 8543.58 18488.86 8545 ;
      RECT 18465.79 8582.095 18488.86 8583.515 ;
      RECT 18361.065 189.04 18361.345 318.595 ;
      RECT 18360.505 189.04 18360.785 342.165 ;
      RECT 18359.945 187.94 18360.225 342.405 ;
      RECT 18359.385 189.04 18359.665 342.645 ;
      RECT 18358.825 187.94 18359.105 342.89 ;
      RECT 18358.265 189.04 18358.545 343.13 ;
      RECT 18357.705 187.94 18357.985 343.37 ;
      RECT 18357.145 189.04 18357.425 343.61 ;
      RECT 18356.585 189.04 18356.865 343.85 ;
      RECT 18356.025 189.04 18356.305 329.47 ;
      RECT 18355.465 189.04 18355.745 329.23 ;
      RECT 18354.905 189.04 18355.185 328.99 ;
      RECT 18354.345 189.04 18354.625 328.75 ;
      RECT 18353.785 189.04 18354.065 328.51 ;
      RECT 18353.225 189.04 18353.505 328.27 ;
      RECT 18352.665 189.04 18352.945 328.03 ;
      RECT 18352.105 189.04 18352.385 327.79 ;
      RECT 18351.545 189.04 18351.825 327.55 ;
      RECT 18350.985 189.04 18351.265 327.31 ;
      RECT 18350.425 187.94 18350.705 327.07 ;
      RECT 18349.865 189.04 18350.145 326.83 ;
      RECT 18349.305 187.94 18349.585 326.59 ;
      RECT 18348.745 189.04 18349.025 326.35 ;
      RECT 18334.745 187.94 18335.025 332.47 ;
      RECT 18334.185 189.04 18334.465 332.23 ;
      RECT 18333.625 189.04 18333.905 331.99 ;
      RECT 18333.065 189.04 18333.345 331.75 ;
      RECT 18332.505 189.04 18332.785 331.51 ;
      RECT 18331.945 189.04 18332.225 331.27 ;
      RECT 18331.385 189.04 18331.665 331.03 ;
      RECT 18330.825 189.04 18331.105 330.79 ;
      RECT 18330.265 189.04 18330.545 330.55 ;
      RECT 18329.705 187.94 18329.985 330.31 ;
      RECT 18329.145 189.04 18329.425 330.07 ;
      RECT 18328.585 187.94 18328.865 329.83 ;
      RECT 18328.025 189.04 18328.305 329.59 ;
      RECT 18327.465 189.04 18327.745 329.35 ;
      RECT 18326.905 189.04 18327.185 329.11 ;
      RECT 18326.345 189.04 18326.625 328.87 ;
      RECT 18325.785 189.04 18326.065 328.63 ;
      RECT 18325.225 189.04 18325.505 328.39 ;
      RECT 18324.665 189.04 18324.945 328.15 ;
      RECT 18324.105 189.04 18324.385 327.91 ;
      RECT 18323.545 189.04 18323.825 327.67 ;
      RECT 18322.985 189.04 18323.265 327.43 ;
      RECT 18322.425 189.04 18322.705 327.19 ;
      RECT 18283.225 189.04 18283.505 334.095 ;
      RECT 18282.665 189.04 18282.945 334.335 ;
      RECT 18282.105 189.04 18282.385 334.575 ;
      RECT 18281.545 187.94 18281.825 334.815 ;
      RECT 18280.985 189.04 18281.265 335.055 ;
      RECT 18280.425 187.94 18280.705 335.295 ;
      RECT 18279.865 189.04 18280.145 335.535 ;
      RECT 18279.305 189.04 18279.585 335.775 ;
      RECT 18278.745 189.04 18279.025 336.015 ;
      RECT 18278.185 187.94 18278.465 336.255 ;
      RECT 18277.625 189.04 18277.905 336.495 ;
      RECT 18277.065 187.94 18277.345 336.735 ;
      RECT 18276.505 189.04 18276.785 336.975 ;
      RECT 18275.945 187.94 18276.225 337.215 ;
      RECT 18275.385 189.04 18275.665 337.455 ;
      RECT 18274.825 189.04 18275.105 337.695 ;
      RECT 18274.265 189.04 18274.545 337.695 ;
      RECT 18273.705 189.04 18273.985 337.455 ;
      RECT 18273.145 189.04 18273.425 337.215 ;
      RECT 18272.585 189.04 18272.865 336.975 ;
      RECT 18272.025 189.04 18272.305 336.735 ;
      RECT 18271.465 189.04 18271.745 336.495 ;
      RECT 18270.905 189.04 18271.185 336.255 ;
      RECT 18270.345 189.04 18270.625 336.015 ;
      RECT 18269.785 189.04 18270.065 335.775 ;
      RECT 18260.825 189.04 18261.105 335.29 ;
      RECT 18260.265 187.94 18260.545 335.05 ;
      RECT 18259.705 189.04 18259.985 334.81 ;
      RECT 18259.145 187.94 18259.425 334.57 ;
      RECT 18258.585 189.04 18258.865 334.33 ;
      RECT 18258.025 187.94 18258.305 334.09 ;
      RECT 18257.465 189.04 18257.745 333.85 ;
      RECT 18256.905 189.04 18257.185 333.61 ;
      RECT 18256.345 189.04 18256.625 333.37 ;
      RECT 18255.785 189.04 18256.065 333.13 ;
      RECT 18255.225 189.04 18255.505 332.89 ;
      RECT 18254.665 189.04 18254.945 332.65 ;
      RECT 18254.105 189.04 18254.385 332.41 ;
      RECT 18253.545 189.04 18253.825 332.17 ;
      RECT 18251.025 187.94 18251.305 333.89 ;
      RECT 18250.465 189.04 18250.745 333.65 ;
      RECT 18249.905 187.94 18250.185 333.41 ;
      RECT 18249.345 189.04 18249.625 333.17 ;
      RECT 18248.785 189.04 18249.065 332.93 ;
      RECT 18248.225 189.04 18248.505 332.69 ;
      RECT 18247.665 189.04 18247.945 332.45 ;
      RECT 18247.105 189.04 18247.385 332.21 ;
      RECT 18221.065 189.04 18221.345 329.86 ;
      RECT 18220.505 189.04 18220.785 330.1 ;
      RECT 18219.945 189.04 18220.225 330.34 ;
      RECT 18219.385 189.04 18219.665 330.585 ;
      RECT 18218.825 189.04 18219.105 330.825 ;
      RECT 18218.265 189.04 18218.545 331.065 ;
      RECT 18217.705 189.04 18217.985 331.065 ;
      RECT 18217.145 189.04 18217.425 330.825 ;
      RECT 18216.585 189.04 18216.865 330.585 ;
      RECT 18216.025 187.94 18216.305 330.345 ;
      RECT 18215.465 189.04 18215.745 330.105 ;
      RECT 18214.905 187.94 18215.185 329.865 ;
      RECT 18214.345 189.04 18214.625 329.625 ;
      RECT 18213.785 189.04 18214.065 329.385 ;
      RECT 18213.225 189.04 18213.505 329.145 ;
      RECT 18212.665 187.94 18212.945 328.905 ;
      RECT 18212.105 189.04 18212.385 328.665 ;
      RECT 18211.545 187.94 18211.825 328.425 ;
      RECT 18210.985 189.04 18211.265 328.185 ;
      RECT 18210.425 187.94 18210.705 327.945 ;
      RECT 18209.865 189.04 18210.145 327.705 ;
      RECT 18209.305 189.04 18209.585 327.465 ;
      RECT 18208.745 189.04 18209.025 327.225 ;
      RECT 18208.185 189.04 18208.465 326.985 ;
      RECT 18194.745 189.04 18195.025 332.785 ;
      RECT 18194.185 189.04 18194.465 332.545 ;
      RECT 18193.625 189.04 18193.905 332.305 ;
      RECT 18193.065 189.04 18193.345 332.065 ;
      RECT 18192.505 189.04 18192.785 331.825 ;
      RECT 18191.945 189.04 18192.225 331.585 ;
      RECT 18191.385 189.04 18191.665 331.345 ;
      RECT 18190.825 189.04 18191.105 331.105 ;
      RECT 18190.265 187.94 18190.545 330.865 ;
      RECT 18189.705 189.04 18189.985 330.625 ;
      RECT 18189.145 187.94 18189.425 330.305 ;
      RECT 18188.585 189.04 18188.865 330.145 ;
      RECT 18188.025 187.94 18188.305 329.905 ;
      RECT 18187.465 189.04 18187.745 329.665 ;
      RECT 18186.905 189.04 18187.185 329.425 ;
      RECT 18186.345 189.04 18186.625 329.185 ;
      RECT 18185.785 189.04 18186.065 328.945 ;
      RECT 18185.225 189.04 18185.505 328.705 ;
      RECT 18184.665 189.04 18184.945 328.465 ;
      RECT 18184.105 189.04 18184.385 328.225 ;
      RECT 18183.545 189.04 18183.825 327.985 ;
      RECT 18182.985 187.94 18183.265 327.745 ;
      RECT 18182.425 189.04 18182.705 327.505 ;
      RECT 18181.865 187.94 18182.145 327.265 ;
      RECT 18142.665 189.04 18142.945 332.875 ;
      RECT 18142.105 189.04 18142.385 333.115 ;
      RECT 18141.545 189.04 18141.825 333.355 ;
      RECT 18140.985 189.04 18141.265 333.595 ;
      RECT 18140.425 189.04 18140.705 333.835 ;
      RECT 18139.865 189.04 18140.145 334.075 ;
      RECT 18139.305 189.04 18139.585 334.315 ;
      RECT 18138.745 189.04 18139.025 334.555 ;
      RECT 18138.185 189.04 18138.465 334.795 ;
      RECT 18137.625 189.04 18137.905 335.035 ;
      RECT 18137.065 189.04 18137.345 335.275 ;
      RECT 18136.505 189.04 18136.785 335.515 ;
      RECT 18135.945 189.04 18136.225 335.755 ;
      RECT 18135.385 189.04 18135.665 335.755 ;
      RECT 18134.825 187.94 18135.105 335.515 ;
      RECT 18134.265 189.04 18134.545 335.275 ;
      RECT 18133.705 187.94 18133.985 335.035 ;
      RECT 18133.145 189.04 18133.425 334.795 ;
      RECT 18132.585 189.04 18132.865 334.555 ;
      RECT 18132.025 189.04 18132.305 334.315 ;
      RECT 18131.465 187.94 18131.745 334.05 ;
      RECT 18130.905 189.04 18131.185 333.81 ;
      RECT 18130.345 187.94 18130.625 333.57 ;
      RECT 18129.785 189.04 18130.065 333.33 ;
      RECT 18120.825 187.94 18121.105 327.165 ;
      RECT 18120.265 189.04 18120.545 327.405 ;
      RECT 18119.705 189.04 18119.985 327.645 ;
      RECT 18119.145 189.04 18119.425 327.645 ;
      RECT 18118.585 189.04 18118.865 327.405 ;
      RECT 18118.025 189.04 18118.305 327.165 ;
      RECT 18117.465 189.04 18117.745 326.925 ;
      RECT 18116.905 189.04 18117.185 326.685 ;
      RECT 18116.345 189.04 18116.625 326.445 ;
      RECT 18115.785 189.04 18116.065 326.205 ;
      RECT 18115.225 189.04 18115.505 325.965 ;
      RECT 18114.665 189.04 18114.945 325.725 ;
      RECT 18114.105 189.04 18114.385 325.485 ;
      RECT 18113.545 187.94 18113.825 325.245 ;
      RECT 18111.025 189.04 18111.305 326.965 ;
      RECT 18110.465 187.94 18110.745 326.725 ;
      RECT 18109.905 189.04 18110.185 326.485 ;
      RECT 18109.345 187.94 18109.625 326.245 ;
      RECT 18108.785 189.04 18109.065 326.005 ;
      RECT 18108.225 189.04 18108.505 325.765 ;
      RECT 18107.665 189.04 18107.945 325.525 ;
      RECT 18081.625 189.04 18081.905 328.31 ;
      RECT 18081.065 189.04 18081.345 328.55 ;
      RECT 18080.505 189.04 18080.785 328.79 ;
      RECT 18079.945 189.04 18080.225 329.03 ;
      RECT 18079.385 189.04 18079.665 329.27 ;
      RECT 18078.825 187.94 18079.105 329.51 ;
      RECT 18078.265 189.04 18078.545 329.75 ;
      RECT 18077.705 187.94 18077.985 329.99 ;
      RECT 18077.145 189.04 18077.425 330.23 ;
      RECT 18076.585 189.04 18076.865 330.47 ;
      RECT 18076.025 189.04 18076.305 330.71 ;
      RECT 18075.465 189.04 18075.745 330.95 ;
      RECT 18074.905 189.04 18075.185 331.19 ;
      RECT 18074.345 189.04 18074.625 331.43 ;
      RECT 18073.785 189.04 18074.065 331.67 ;
      RECT 18073.225 189.04 18073.505 331.67 ;
      RECT 18072.665 189.04 18072.945 331.43 ;
      RECT 18072.105 189.04 18072.385 331.19 ;
      RECT 18071.545 189.04 18071.825 330.95 ;
      RECT 18070.985 189.04 18071.265 330.705 ;
      RECT 18070.425 189.04 18070.705 330.465 ;
      RECT 18069.865 189.04 18070.145 330.225 ;
      RECT 18069.305 187.94 18069.585 329.985 ;
      RECT 18068.745 189.04 18069.025 329.745 ;
      RECT 18055.305 187.94 18055.585 327.225 ;
      RECT 18054.745 189.04 18055.025 326.985 ;
      RECT 18054.185 189.04 18054.465 326.745 ;
      RECT 18053.625 189.04 18053.905 326.505 ;
      RECT 18053.065 187.94 18053.345 326.265 ;
      RECT 18052.505 189.04 18052.785 326.025 ;
      RECT 18051.945 187.94 18052.225 325.785 ;
      RECT 18051.385 189.04 18051.665 325.545 ;
      RECT 18050.825 187.94 18051.105 325.305 ;
      RECT 18050.265 189.04 18050.545 325.065 ;
      RECT 18049.705 189.04 18049.985 324.825 ;
      RECT 18049.145 189.04 18049.425 324.585 ;
      RECT 18048.585 189.04 18048.865 324.345 ;
      RECT 18048.025 189.04 18048.305 324.105 ;
      RECT 18047.465 189.04 18047.745 323.865 ;
      RECT 18046.905 189.04 18047.185 323.625 ;
      RECT 18046.345 189.04 18046.625 323.385 ;
      RECT 18045.785 189.04 18046.065 323.145 ;
      RECT 18045.225 189.04 18045.505 322.905 ;
      RECT 18044.665 189.04 18044.945 322.665 ;
      RECT 18044.105 189.04 18044.385 322.425 ;
      RECT 18043.545 187.94 18043.825 322.185 ;
      RECT 18042.985 189.04 18043.265 321.945 ;
      RECT 18042.425 187.94 18042.705 321.705 ;
      RECT 18002.665 189.04 18002.945 332.175 ;
      RECT 18002.105 187.94 18002.385 332.415 ;
      RECT 18001.545 189.04 18001.825 332.655 ;
      RECT 18000.985 189.04 18001.265 332.895 ;
      RECT 18000.425 189.04 18000.705 333.135 ;
      RECT 17999.865 189.04 18000.145 333.375 ;
      RECT 17999.305 189.04 17999.585 333.615 ;
      RECT 17998.745 189.04 17999.025 333.86 ;
      RECT 17998.185 189.04 17998.465 334.1 ;
      RECT 17997.625 189.04 17997.905 334.34 ;
      RECT 17997.065 187.94 17997.345 334.58 ;
      RECT 17996.505 189.04 17996.785 334.82 ;
      RECT 17995.945 187.94 17996.225 335.06 ;
      RECT 17995.385 189.04 17995.665 335.3 ;
      RECT 17994.825 189.04 17995.105 335.54 ;
      RECT 17994.265 189.04 17994.545 335.78 ;
      RECT 17993.705 189.04 17993.985 336.02 ;
      RECT 17993.145 189.04 17993.425 336.26 ;
      RECT 17992.585 189.04 17992.865 336.5 ;
      RECT 17992.025 189.04 17992.305 336.74 ;
      RECT 17991.465 189.04 17991.745 336.98 ;
      RECT 17990.905 189.04 17991.185 337.22 ;
      RECT 17990.345 189.04 17990.625 337.46 ;
      RECT 17989.785 189.04 17990.065 337.7 ;
      RECT 17980.825 189.04 17981.105 333.285 ;
      RECT 17980.265 189.04 17980.545 333.045 ;
      RECT 17979.705 189.04 17979.985 332.805 ;
      RECT 17979.145 187.94 17979.425 332.565 ;
      RECT 17978.585 189.04 17978.865 332.325 ;
      RECT 17978.025 187.94 17978.305 332.085 ;
      RECT 17977.465 189.04 17977.745 331.845 ;
      RECT 17976.905 189.04 17977.185 331.605 ;
      RECT 17976.345 189.04 17976.625 331.365 ;
      RECT 17975.785 187.94 17976.065 331.125 ;
      RECT 17975.225 189.04 17975.505 330.885 ;
      RECT 17974.665 187.94 17974.945 330.645 ;
      RECT 17974.105 189.04 17974.385 330.405 ;
      RECT 17973.545 187.94 17973.825 330.165 ;
      RECT 17971.025 189.04 17971.305 322.565 ;
      RECT 17970.465 189.04 17970.745 322.325 ;
      RECT 17969.905 189.04 17970.185 322.085 ;
      RECT 17969.345 189.04 17969.625 321.845 ;
      RECT 17968.785 189.04 17969.065 321.605 ;
      RECT 17968.225 189.04 17968.505 321.365 ;
      RECT 17967.665 189.04 17967.945 321.125 ;
      RECT 17941.625 189.04 17941.905 335 ;
      RECT 17941.065 189.04 17941.345 335.24 ;
      RECT 17940.505 189.04 17940.785 335.48 ;
      RECT 17939.945 189.04 17940.225 335.72 ;
      RECT 17939.385 189.04 17939.665 335.96 ;
      RECT 17938.825 187.94 17939.105 335.96 ;
      RECT 17938.265 189.04 17938.545 335.72 ;
      RECT 17937.705 187.94 17937.985 335.475 ;
      RECT 17937.145 189.04 17937.425 335.235 ;
      RECT 17936.585 187.94 17936.865 334.995 ;
      RECT 17936.025 189.04 17936.305 334.755 ;
      RECT 17935.465 189.04 17935.745 334.515 ;
      RECT 17934.905 189.04 17935.185 334.275 ;
      RECT 17934.345 189.04 17934.625 334.035 ;
      RECT 17933.785 189.04 17934.065 333.795 ;
      RECT 17933.225 189.04 17933.505 333.555 ;
      RECT 17932.665 189.04 17932.945 333.315 ;
      RECT 17932.105 189.04 17932.385 333.075 ;
      RECT 17931.545 187.94 17931.825 332.835 ;
      RECT 17930.985 189.04 17931.265 332.595 ;
      RECT 17930.425 187.94 17930.705 332.355 ;
      RECT 17929.865 189.04 17930.145 332.115 ;
      RECT 17929.305 189.04 17929.585 331.875 ;
      RECT 17928.745 189.04 17929.025 331.635 ;
      RECT 17915.305 189.04 17915.585 335.035 ;
      RECT 17914.745 189.04 17915.025 335.275 ;
      RECT 17914.185 189.04 17914.465 335.52 ;
      RECT 17913.625 189.04 17913.905 335.76 ;
      RECT 17913.065 189.04 17913.345 336 ;
      RECT 17912.505 189.04 17912.785 336 ;
      RECT 17911.945 189.04 17912.225 335.76 ;
      RECT 17911.385 189.04 17911.665 335.52 ;
      RECT 17910.825 189.04 17911.105 328.505 ;
      RECT 17910.265 189.04 17910.545 328.265 ;
      RECT 17909.705 189.04 17909.985 328.025 ;
      RECT 17909.145 187.94 17909.425 327.785 ;
      RECT 17908.585 189.04 17908.865 327.545 ;
      RECT 17908.025 187.94 17908.305 327.305 ;
      RECT 17907.465 189.04 17907.745 327.065 ;
      RECT 17906.905 189.04 17907.185 326.825 ;
      RECT 17906.345 189.04 17906.625 326.585 ;
      RECT 17905.785 187.94 17906.065 326.345 ;
      RECT 17905.225 189.04 17905.505 326.105 ;
      RECT 17904.665 187.94 17904.945 325.865 ;
      RECT 17904.105 189.04 17904.385 325.625 ;
      RECT 17903.545 187.94 17903.825 325.385 ;
      RECT 17902.985 189.04 17903.265 325.145 ;
      RECT 17902.425 189.04 17902.705 324.905 ;
      RECT 17862.105 189.04 17862.385 333.8 ;
      RECT 17861.545 189.04 17861.825 334.04 ;
      RECT 17860.985 189.04 17861.265 334.285 ;
      RECT 17860.425 189.04 17860.705 334.525 ;
      RECT 17859.865 189.04 17860.145 334.765 ;
      RECT 17859.305 189.04 17859.585 335.005 ;
      RECT 17858.745 189.04 17859.025 335.245 ;
      RECT 17858.185 189.04 17858.465 335.485 ;
      RECT 17857.625 189.04 17857.905 335.725 ;
      RECT 17857.065 189.04 17857.345 335.965 ;
      RECT 17856.505 187.94 17856.785 336.205 ;
      RECT 17855.945 189.04 17856.225 336.445 ;
      RECT 17855.385 187.94 17855.665 336.685 ;
      RECT 17854.825 189.04 17855.105 336.925 ;
      RECT 17854.265 187.94 17854.545 337.165 ;
      RECT 17853.705 189.04 17853.985 337.165 ;
      RECT 17853.145 189.04 17853.425 336.925 ;
      RECT 17852.585 189.04 17852.865 336.685 ;
      RECT 17852.025 189.04 17852.305 336.445 ;
      RECT 17851.465 189.04 17851.745 336.205 ;
      RECT 17850.905 189.04 17851.185 335.965 ;
      RECT 17850.345 189.04 17850.625 335.725 ;
      RECT 17849.785 189.04 17850.065 335.485 ;
      RECT 17840.825 187.94 17841.105 335.515 ;
      RECT 17840.265 189.04 17840.545 335.755 ;
      RECT 17839.705 187.94 17839.985 335.995 ;
      RECT 17839.145 189.04 17839.425 336.21 ;
      RECT 17838.585 189.04 17838.865 335.785 ;
      RECT 17838.025 189.04 17838.305 335.545 ;
      RECT 17837.465 189.04 17837.745 335.305 ;
      RECT 17836.905 189.04 17837.185 335.065 ;
      RECT 17836.345 189.04 17836.625 334.825 ;
      RECT 17835.785 189.04 17836.065 334.585 ;
      RECT 17835.225 189.04 17835.505 334.345 ;
      RECT 17834.665 189.04 17834.945 334.105 ;
      RECT 17834.105 189.04 17834.385 333.865 ;
      RECT 17833.545 189.04 17833.825 333.625 ;
      RECT 17831.025 189.04 17831.305 332.8 ;
      RECT 17830.465 189.04 17830.745 332.56 ;
      RECT 17829.905 189.04 17830.185 332.32 ;
      RECT 17829.345 187.94 17829.625 332.08 ;
      RECT 17828.785 189.04 17829.065 331.84 ;
      RECT 17828.225 187.94 17828.505 331.6 ;
      RECT 17827.665 189.04 17827.945 331.36 ;
      RECT 17827.105 189.04 17827.385 331.12 ;
      RECT 17800.505 189.04 17800.785 342.165 ;
      RECT 17799.945 187.94 17800.225 342.405 ;
      RECT 17799.385 189.04 17799.665 342.645 ;
      RECT 17798.825 187.94 17799.105 342.89 ;
      RECT 17798.265 189.04 17798.545 343.13 ;
      RECT 17797.705 187.94 17797.985 343.37 ;
      RECT 17797.145 189.04 17797.425 343.61 ;
      RECT 17796.585 189.04 17796.865 343.85 ;
      RECT 17796.025 189.04 17796.305 329.47 ;
      RECT 17795.465 189.04 17795.745 329.23 ;
      RECT 17794.905 189.04 17795.185 328.99 ;
      RECT 17794.345 189.04 17794.625 328.75 ;
      RECT 17793.785 189.04 17794.065 328.51 ;
      RECT 17793.225 189.04 17793.505 328.27 ;
      RECT 17792.665 189.04 17792.945 328.03 ;
      RECT 17792.105 189.04 17792.385 327.79 ;
      RECT 17791.545 189.04 17791.825 327.55 ;
      RECT 17790.985 189.04 17791.265 327.31 ;
      RECT 17790.425 187.94 17790.705 327.07 ;
      RECT 17789.865 189.04 17790.145 326.83 ;
      RECT 17789.305 187.94 17789.585 326.59 ;
      RECT 17788.745 189.04 17789.025 326.35 ;
      RECT 17774.745 187.94 17775.025 332.47 ;
      RECT 17774.185 189.04 17774.465 332.23 ;
      RECT 17773.625 189.04 17773.905 331.99 ;
      RECT 17773.065 189.04 17773.345 331.75 ;
      RECT 17772.505 189.04 17772.785 331.51 ;
      RECT 17771.945 189.04 17772.225 331.27 ;
      RECT 17771.385 189.04 17771.665 331.03 ;
      RECT 17770.825 189.04 17771.105 330.79 ;
      RECT 17770.265 189.04 17770.545 330.55 ;
      RECT 17769.705 187.94 17769.985 330.31 ;
      RECT 17769.145 189.04 17769.425 330.07 ;
      RECT 17768.585 187.94 17768.865 329.83 ;
      RECT 17768.025 189.04 17768.305 329.59 ;
      RECT 17767.465 189.04 17767.745 329.35 ;
      RECT 17766.905 189.04 17767.185 329.11 ;
      RECT 17766.345 189.04 17766.625 328.87 ;
      RECT 17765.785 189.04 17766.065 328.63 ;
      RECT 17765.225 189.04 17765.505 328.39 ;
      RECT 17764.665 189.04 17764.945 328.15 ;
      RECT 17764.105 189.04 17764.385 327.91 ;
      RECT 17763.545 189.04 17763.825 327.67 ;
      RECT 17762.985 189.04 17763.265 327.43 ;
      RECT 17762.425 189.04 17762.705 327.19 ;
      RECT 17723.225 189.04 17723.505 334.095 ;
      RECT 17722.665 189.04 17722.945 334.335 ;
      RECT 17722.105 189.04 17722.385 334.575 ;
      RECT 17721.545 187.94 17721.825 334.815 ;
      RECT 17720.985 189.04 17721.265 335.055 ;
      RECT 17720.425 187.94 17720.705 335.295 ;
      RECT 17719.865 189.04 17720.145 335.535 ;
      RECT 17719.305 189.04 17719.585 335.775 ;
      RECT 17718.745 189.04 17719.025 336.015 ;
      RECT 17718.185 187.94 17718.465 336.255 ;
      RECT 17717.625 189.04 17717.905 336.495 ;
      RECT 17717.065 187.94 17717.345 336.735 ;
      RECT 17716.505 189.04 17716.785 336.975 ;
      RECT 17715.945 187.94 17716.225 337.215 ;
      RECT 17715.385 189.04 17715.665 337.455 ;
      RECT 17714.825 189.04 17715.105 337.695 ;
      RECT 17714.265 189.04 17714.545 337.695 ;
      RECT 17713.705 189.04 17713.985 337.455 ;
      RECT 17713.145 189.04 17713.425 337.215 ;
      RECT 17712.585 189.04 17712.865 336.975 ;
      RECT 17712.025 189.04 17712.305 336.735 ;
      RECT 17711.465 189.04 17711.745 336.495 ;
      RECT 17710.905 189.04 17711.185 336.255 ;
      RECT 17710.345 189.04 17710.625 336.015 ;
      RECT 17709.785 189.04 17710.065 335.775 ;
      RECT 17700.825 189.04 17701.105 335.29 ;
      RECT 17700.265 187.94 17700.545 335.05 ;
      RECT 17699.705 189.04 17699.985 334.81 ;
      RECT 17699.145 187.94 17699.425 334.57 ;
      RECT 17698.585 189.04 17698.865 334.33 ;
      RECT 17698.025 187.94 17698.305 334.09 ;
      RECT 17697.465 189.04 17697.745 333.85 ;
      RECT 17696.905 189.04 17697.185 333.61 ;
      RECT 17696.345 189.04 17696.625 333.37 ;
      RECT 17695.785 189.04 17696.065 333.13 ;
      RECT 17695.225 189.04 17695.505 332.89 ;
      RECT 17694.665 189.04 17694.945 332.65 ;
      RECT 17694.105 189.04 17694.385 332.41 ;
      RECT 17693.545 189.04 17693.825 332.17 ;
      RECT 17691.025 187.94 17691.305 333.89 ;
      RECT 17690.465 189.04 17690.745 333.65 ;
      RECT 17689.905 187.94 17690.185 333.41 ;
      RECT 17689.345 189.04 17689.625 333.17 ;
      RECT 17688.785 189.04 17689.065 332.93 ;
      RECT 17688.225 189.04 17688.505 332.69 ;
      RECT 17687.665 189.04 17687.945 332.45 ;
      RECT 17687.105 189.04 17687.385 332.21 ;
      RECT 17661.065 189.04 17661.345 329.86 ;
      RECT 17660.505 189.04 17660.785 330.1 ;
      RECT 17659.945 189.04 17660.225 330.34 ;
      RECT 17659.385 189.04 17659.665 330.585 ;
      RECT 17658.825 189.04 17659.105 330.825 ;
      RECT 17658.265 189.04 17658.545 331.065 ;
      RECT 17657.705 189.04 17657.985 331.065 ;
      RECT 17657.145 189.04 17657.425 330.825 ;
      RECT 17656.585 189.04 17656.865 330.585 ;
      RECT 17656.025 187.94 17656.305 330.345 ;
      RECT 17655.465 189.04 17655.745 330.105 ;
      RECT 17654.905 187.94 17655.185 329.865 ;
      RECT 17654.345 189.04 17654.625 329.625 ;
      RECT 17653.785 189.04 17654.065 329.385 ;
      RECT 17653.225 189.04 17653.505 329.145 ;
      RECT 17652.665 187.94 17652.945 328.905 ;
      RECT 17652.105 189.04 17652.385 328.665 ;
      RECT 17651.545 187.94 17651.825 328.425 ;
      RECT 17650.985 189.04 17651.265 328.185 ;
      RECT 17650.425 187.94 17650.705 327.945 ;
      RECT 17649.865 189.04 17650.145 327.705 ;
      RECT 17649.305 189.04 17649.585 327.465 ;
      RECT 17648.745 189.04 17649.025 327.225 ;
      RECT 17648.185 189.04 17648.465 326.985 ;
      RECT 17634.745 189.04 17635.025 332.785 ;
      RECT 17634.185 189.04 17634.465 332.545 ;
      RECT 17633.625 189.04 17633.905 332.305 ;
      RECT 17633.065 189.04 17633.345 332.065 ;
      RECT 17632.505 189.04 17632.785 331.825 ;
      RECT 17631.945 189.04 17632.225 331.585 ;
      RECT 17631.385 189.04 17631.665 331.345 ;
      RECT 17630.825 189.04 17631.105 331.105 ;
      RECT 17630.265 187.94 17630.545 330.865 ;
      RECT 17629.705 189.04 17629.985 330.625 ;
      RECT 17629.145 187.94 17629.425 330.305 ;
      RECT 17628.585 189.04 17628.865 330.145 ;
      RECT 17628.025 187.94 17628.305 329.905 ;
      RECT 17627.465 189.04 17627.745 329.665 ;
      RECT 17626.905 189.04 17627.185 329.425 ;
      RECT 17626.345 189.04 17626.625 329.185 ;
      RECT 17625.785 189.04 17626.065 328.945 ;
      RECT 17625.225 189.04 17625.505 328.705 ;
      RECT 17624.665 189.04 17624.945 328.465 ;
      RECT 17624.105 189.04 17624.385 328.225 ;
      RECT 17623.545 189.04 17623.825 327.985 ;
      RECT 17622.985 187.94 17623.265 327.745 ;
      RECT 17622.425 189.04 17622.705 327.505 ;
      RECT 17621.865 187.94 17622.145 327.265 ;
      RECT 17582.665 189.04 17582.945 332.875 ;
      RECT 17582.105 189.04 17582.385 333.115 ;
      RECT 17581.545 189.04 17581.825 333.355 ;
      RECT 17580.985 189.04 17581.265 333.595 ;
      RECT 17580.425 189.04 17580.705 333.835 ;
      RECT 17579.865 189.04 17580.145 334.075 ;
      RECT 17579.305 189.04 17579.585 334.315 ;
      RECT 17578.745 189.04 17579.025 334.555 ;
      RECT 17578.185 189.04 17578.465 334.795 ;
      RECT 17577.625 189.04 17577.905 335.035 ;
      RECT 17577.065 189.04 17577.345 335.275 ;
      RECT 17576.505 189.04 17576.785 335.515 ;
      RECT 17575.945 189.04 17576.225 335.755 ;
      RECT 17575.385 189.04 17575.665 335.755 ;
      RECT 17574.825 187.94 17575.105 335.515 ;
      RECT 17574.265 189.04 17574.545 335.275 ;
      RECT 17573.705 187.94 17573.985 335.035 ;
      RECT 17573.145 189.04 17573.425 334.795 ;
      RECT 17572.585 189.04 17572.865 334.555 ;
      RECT 17572.025 189.04 17572.305 334.315 ;
      RECT 17571.465 187.94 17571.745 334.05 ;
      RECT 17570.905 189.04 17571.185 333.81 ;
      RECT 17570.345 187.94 17570.625 333.57 ;
      RECT 17569.785 189.04 17570.065 333.33 ;
      RECT 17560.825 187.94 17561.105 327.165 ;
      RECT 17560.265 189.04 17560.545 327.405 ;
      RECT 17559.705 189.04 17559.985 327.645 ;
      RECT 17559.145 189.04 17559.425 327.645 ;
      RECT 17558.585 189.04 17558.865 327.405 ;
      RECT 17558.025 189.04 17558.305 327.165 ;
      RECT 17557.465 189.04 17557.745 326.925 ;
      RECT 17556.905 189.04 17557.185 326.685 ;
      RECT 17556.345 189.04 17556.625 326.445 ;
      RECT 17555.785 189.04 17556.065 326.205 ;
      RECT 17555.225 189.04 17555.505 325.965 ;
      RECT 17554.665 189.04 17554.945 325.725 ;
      RECT 17554.105 189.04 17554.385 325.485 ;
      RECT 17553.545 187.94 17553.825 325.245 ;
      RECT 17551.025 189.04 17551.305 326.965 ;
      RECT 17550.465 187.94 17550.745 326.725 ;
      RECT 17549.905 189.04 17550.185 326.485 ;
      RECT 17549.345 187.94 17549.625 326.245 ;
      RECT 17548.785 189.04 17549.065 326.005 ;
      RECT 17548.225 189.04 17548.505 325.765 ;
      RECT 17547.665 189.04 17547.945 325.525 ;
      RECT 17521.625 189.04 17521.905 328.31 ;
      RECT 17521.065 189.04 17521.345 328.55 ;
      RECT 17520.505 189.04 17520.785 328.79 ;
      RECT 17519.945 189.04 17520.225 329.03 ;
      RECT 17519.385 189.04 17519.665 329.27 ;
      RECT 17518.825 187.94 17519.105 329.51 ;
      RECT 17518.265 189.04 17518.545 329.75 ;
      RECT 17517.705 187.94 17517.985 329.99 ;
      RECT 17517.145 189.04 17517.425 330.23 ;
      RECT 17516.585 189.04 17516.865 330.47 ;
      RECT 17516.025 189.04 17516.305 330.71 ;
      RECT 17515.465 189.04 17515.745 330.95 ;
      RECT 17514.905 189.04 17515.185 331.19 ;
      RECT 17514.345 189.04 17514.625 331.43 ;
      RECT 17513.785 189.04 17514.065 331.67 ;
      RECT 17513.225 189.04 17513.505 331.67 ;
      RECT 17512.665 189.04 17512.945 331.43 ;
      RECT 17512.105 189.04 17512.385 331.19 ;
      RECT 17511.545 189.04 17511.825 330.95 ;
      RECT 17510.985 189.04 17511.265 330.705 ;
      RECT 17510.425 189.04 17510.705 330.465 ;
      RECT 17509.865 189.04 17510.145 330.225 ;
      RECT 17509.305 187.94 17509.585 329.985 ;
      RECT 17508.745 189.04 17509.025 329.745 ;
      RECT 17495.305 187.94 17495.585 327.225 ;
      RECT 17494.745 189.04 17495.025 326.985 ;
      RECT 17494.185 189.04 17494.465 326.745 ;
      RECT 17493.625 189.04 17493.905 326.505 ;
      RECT 17493.065 187.94 17493.345 326.265 ;
      RECT 17492.505 189.04 17492.785 326.025 ;
      RECT 17491.945 187.94 17492.225 325.785 ;
      RECT 17491.385 189.04 17491.665 325.545 ;
      RECT 17490.825 187.94 17491.105 325.305 ;
      RECT 17490.265 189.04 17490.545 325.065 ;
      RECT 17489.705 189.04 17489.985 324.825 ;
      RECT 17489.145 189.04 17489.425 324.585 ;
      RECT 17488.585 189.04 17488.865 324.345 ;
      RECT 17488.025 189.04 17488.305 324.105 ;
      RECT 17487.465 189.04 17487.745 323.865 ;
      RECT 17486.905 189.04 17487.185 323.625 ;
      RECT 17486.345 189.04 17486.625 323.385 ;
      RECT 17485.785 189.04 17486.065 323.145 ;
      RECT 17485.225 189.04 17485.505 322.905 ;
      RECT 17484.665 189.04 17484.945 322.665 ;
      RECT 17484.105 189.04 17484.385 322.425 ;
      RECT 17483.545 187.94 17483.825 322.185 ;
      RECT 17482.985 189.04 17483.265 321.945 ;
      RECT 17482.425 187.94 17482.705 321.705 ;
      RECT 17442.665 189.04 17442.945 332.175 ;
      RECT 17442.105 187.94 17442.385 332.415 ;
      RECT 17441.545 189.04 17441.825 332.655 ;
      RECT 17440.985 189.04 17441.265 332.895 ;
      RECT 17440.425 189.04 17440.705 333.135 ;
      RECT 17439.865 189.04 17440.145 333.375 ;
      RECT 17439.305 189.04 17439.585 333.615 ;
      RECT 17438.745 189.04 17439.025 333.86 ;
      RECT 17438.185 189.04 17438.465 334.1 ;
      RECT 17437.625 189.04 17437.905 334.34 ;
      RECT 17437.065 187.94 17437.345 334.58 ;
      RECT 17436.505 189.04 17436.785 334.82 ;
      RECT 17435.945 187.94 17436.225 335.06 ;
      RECT 17435.385 189.04 17435.665 335.3 ;
      RECT 17434.825 189.04 17435.105 335.54 ;
      RECT 17434.265 189.04 17434.545 335.78 ;
      RECT 17433.705 189.04 17433.985 336.02 ;
      RECT 17433.145 189.04 17433.425 336.26 ;
      RECT 17432.585 189.04 17432.865 336.5 ;
      RECT 17432.025 189.04 17432.305 336.74 ;
      RECT 17431.465 189.04 17431.745 336.98 ;
      RECT 17430.905 189.04 17431.185 337.22 ;
      RECT 17430.345 189.04 17430.625 337.46 ;
      RECT 17429.785 189.04 17430.065 337.7 ;
      RECT 17420.825 189.04 17421.105 333.285 ;
      RECT 17420.265 189.04 17420.545 333.045 ;
      RECT 17419.705 189.04 17419.985 332.805 ;
      RECT 17419.145 187.94 17419.425 332.565 ;
      RECT 17418.585 189.04 17418.865 332.325 ;
      RECT 17418.025 187.94 17418.305 332.085 ;
      RECT 17417.465 189.04 17417.745 331.845 ;
      RECT 17416.905 189.04 17417.185 331.605 ;
      RECT 17416.345 189.04 17416.625 331.365 ;
      RECT 17415.785 187.94 17416.065 331.125 ;
      RECT 17415.225 189.04 17415.505 330.885 ;
      RECT 17414.665 187.94 17414.945 330.645 ;
      RECT 17414.105 189.04 17414.385 330.405 ;
      RECT 17413.545 187.94 17413.825 330.165 ;
      RECT 17411.025 189.04 17411.305 322.565 ;
      RECT 17410.465 189.04 17410.745 322.325 ;
      RECT 17409.905 189.04 17410.185 322.085 ;
      RECT 17409.345 189.04 17409.625 321.845 ;
      RECT 17408.785 189.04 17409.065 321.605 ;
      RECT 17408.225 189.04 17408.505 321.365 ;
      RECT 17407.665 189.04 17407.945 321.125 ;
      RECT 17381.625 189.04 17381.905 335 ;
      RECT 17381.065 189.04 17381.345 335.24 ;
      RECT 17380.505 189.04 17380.785 335.48 ;
      RECT 17379.945 189.04 17380.225 335.72 ;
      RECT 17379.385 189.04 17379.665 335.96 ;
      RECT 17378.825 187.94 17379.105 335.96 ;
      RECT 17378.265 189.04 17378.545 335.72 ;
      RECT 17377.705 187.94 17377.985 335.475 ;
      RECT 17377.145 189.04 17377.425 335.235 ;
      RECT 17376.585 187.94 17376.865 334.995 ;
      RECT 17376.025 189.04 17376.305 334.755 ;
      RECT 17375.465 189.04 17375.745 334.515 ;
      RECT 17374.905 189.04 17375.185 334.275 ;
      RECT 17374.345 189.04 17374.625 334.035 ;
      RECT 17373.785 189.04 17374.065 333.795 ;
      RECT 17373.225 189.04 17373.505 333.555 ;
      RECT 17372.665 189.04 17372.945 333.315 ;
      RECT 17372.105 189.04 17372.385 333.075 ;
      RECT 17371.545 187.94 17371.825 332.835 ;
      RECT 17370.985 189.04 17371.265 332.595 ;
      RECT 17370.425 187.94 17370.705 332.355 ;
      RECT 17369.865 189.04 17370.145 332.115 ;
      RECT 17369.305 189.04 17369.585 331.875 ;
      RECT 17368.745 189.04 17369.025 331.635 ;
      RECT 17355.305 189.04 17355.585 335.035 ;
      RECT 17354.745 189.04 17355.025 335.275 ;
      RECT 17354.185 189.04 17354.465 335.52 ;
      RECT 17353.625 189.04 17353.905 335.76 ;
      RECT 17353.065 189.04 17353.345 336 ;
      RECT 17352.505 189.04 17352.785 336 ;
      RECT 17351.945 189.04 17352.225 335.76 ;
      RECT 17351.385 189.04 17351.665 335.52 ;
      RECT 17350.825 189.04 17351.105 328.505 ;
      RECT 17350.265 189.04 17350.545 328.265 ;
      RECT 17349.705 189.04 17349.985 328.025 ;
      RECT 17349.145 187.94 17349.425 327.785 ;
      RECT 17348.585 189.04 17348.865 327.545 ;
      RECT 17348.025 187.94 17348.305 327.305 ;
      RECT 17347.465 189.04 17347.745 327.065 ;
      RECT 17346.905 189.04 17347.185 326.825 ;
      RECT 17346.345 189.04 17346.625 326.585 ;
      RECT 17345.785 187.94 17346.065 326.345 ;
      RECT 17345.225 189.04 17345.505 326.105 ;
      RECT 17344.665 187.94 17344.945 325.865 ;
      RECT 17344.105 189.04 17344.385 325.625 ;
      RECT 17343.545 187.94 17343.825 325.385 ;
      RECT 17342.985 189.04 17343.265 325.145 ;
      RECT 17342.425 189.04 17342.705 324.905 ;
      RECT 17302.105 189.04 17302.385 333.8 ;
      RECT 17301.545 189.04 17301.825 334.04 ;
      RECT 17300.985 189.04 17301.265 334.285 ;
      RECT 17300.425 189.04 17300.705 334.525 ;
      RECT 17299.865 189.04 17300.145 334.765 ;
      RECT 17299.305 189.04 17299.585 335.005 ;
      RECT 17298.745 189.04 17299.025 335.245 ;
      RECT 17298.185 189.04 17298.465 335.485 ;
      RECT 17297.625 189.04 17297.905 335.725 ;
      RECT 17297.065 189.04 17297.345 335.965 ;
      RECT 17296.505 187.94 17296.785 336.205 ;
      RECT 17295.945 189.04 17296.225 336.445 ;
      RECT 17295.385 187.94 17295.665 336.685 ;
      RECT 17294.825 189.04 17295.105 336.925 ;
      RECT 17294.265 187.94 17294.545 337.165 ;
      RECT 17293.705 189.04 17293.985 337.165 ;
      RECT 17293.145 189.04 17293.425 336.925 ;
      RECT 17292.585 189.04 17292.865 336.685 ;
      RECT 17292.025 189.04 17292.305 336.445 ;
      RECT 17291.465 189.04 17291.745 336.205 ;
      RECT 17290.905 189.04 17291.185 335.965 ;
      RECT 17290.345 189.04 17290.625 335.725 ;
      RECT 17289.785 189.04 17290.065 335.485 ;
      RECT 17280.825 187.94 17281.105 335.515 ;
      RECT 17280.265 189.04 17280.545 335.755 ;
      RECT 17279.705 187.94 17279.985 335.995 ;
      RECT 17279.145 189.04 17279.425 336.21 ;
      RECT 17278.585 189.04 17278.865 335.785 ;
      RECT 17278.025 189.04 17278.305 335.545 ;
      RECT 17277.465 189.04 17277.745 335.305 ;
      RECT 17276.905 189.04 17277.185 335.065 ;
      RECT 17276.345 189.04 17276.625 334.825 ;
      RECT 17275.785 189.04 17276.065 334.585 ;
      RECT 17275.225 189.04 17275.505 334.345 ;
      RECT 17274.665 189.04 17274.945 334.105 ;
      RECT 17274.105 189.04 17274.385 333.865 ;
      RECT 17273.545 189.04 17273.825 333.625 ;
      RECT 17271.025 189.04 17271.305 332.8 ;
      RECT 17270.465 189.04 17270.745 332.56 ;
      RECT 17269.905 189.04 17270.185 332.32 ;
      RECT 17269.345 187.94 17269.625 332.08 ;
      RECT 17268.785 189.04 17269.065 331.84 ;
      RECT 17268.225 187.94 17268.505 331.6 ;
      RECT 17267.665 189.04 17267.945 331.36 ;
      RECT 17267.105 189.04 17267.385 331.12 ;
      RECT 17240.505 189.04 17240.785 342.165 ;
      RECT 17239.945 187.94 17240.225 342.405 ;
      RECT 17239.385 189.04 17239.665 342.645 ;
      RECT 17238.825 187.94 17239.105 342.89 ;
      RECT 17238.265 189.04 17238.545 343.13 ;
      RECT 17237.705 187.94 17237.985 343.37 ;
      RECT 17237.145 189.04 17237.425 343.61 ;
      RECT 17236.585 189.04 17236.865 343.85 ;
      RECT 17236.025 189.04 17236.305 329.47 ;
      RECT 17235.465 189.04 17235.745 329.23 ;
      RECT 17234.905 189.04 17235.185 328.99 ;
      RECT 17234.345 189.04 17234.625 328.75 ;
      RECT 17233.785 189.04 17234.065 328.51 ;
      RECT 17233.225 189.04 17233.505 328.27 ;
      RECT 17232.665 189.04 17232.945 328.03 ;
      RECT 17232.105 189.04 17232.385 327.79 ;
      RECT 17231.545 189.04 17231.825 327.55 ;
      RECT 17230.985 189.04 17231.265 327.31 ;
      RECT 17230.425 187.94 17230.705 327.07 ;
      RECT 17229.865 189.04 17230.145 326.83 ;
      RECT 17229.305 187.94 17229.585 326.59 ;
      RECT 17228.745 189.04 17229.025 326.35 ;
      RECT 17214.745 187.94 17215.025 332.47 ;
      RECT 17214.185 189.04 17214.465 332.23 ;
      RECT 17213.625 189.04 17213.905 331.99 ;
      RECT 17213.065 189.04 17213.345 331.75 ;
      RECT 17212.505 189.04 17212.785 331.51 ;
      RECT 17211.945 189.04 17212.225 331.27 ;
      RECT 17211.385 189.04 17211.665 331.03 ;
      RECT 17210.825 189.04 17211.105 330.79 ;
      RECT 17210.265 189.04 17210.545 330.55 ;
      RECT 17209.705 187.94 17209.985 330.31 ;
      RECT 17209.145 189.04 17209.425 330.07 ;
      RECT 17208.585 187.94 17208.865 329.83 ;
      RECT 17208.025 189.04 17208.305 329.59 ;
      RECT 17207.465 189.04 17207.745 329.35 ;
      RECT 17206.905 189.04 17207.185 329.11 ;
      RECT 17206.345 189.04 17206.625 328.87 ;
      RECT 17205.785 189.04 17206.065 328.63 ;
      RECT 17205.225 189.04 17205.505 328.39 ;
      RECT 17204.665 189.04 17204.945 328.15 ;
      RECT 17204.105 189.04 17204.385 327.91 ;
      RECT 17203.545 189.04 17203.825 327.67 ;
      RECT 17202.985 189.04 17203.265 327.43 ;
      RECT 17202.425 189.04 17202.705 327.19 ;
      RECT 17163.225 189.04 17163.505 334.095 ;
      RECT 17162.665 189.04 17162.945 334.335 ;
      RECT 17162.105 189.04 17162.385 334.575 ;
      RECT 17161.545 187.94 17161.825 334.815 ;
      RECT 17160.985 189.04 17161.265 335.055 ;
      RECT 17160.425 187.94 17160.705 335.295 ;
      RECT 17159.865 189.04 17160.145 335.535 ;
      RECT 17159.305 189.04 17159.585 335.775 ;
      RECT 17158.745 189.04 17159.025 336.015 ;
      RECT 17158.185 187.94 17158.465 336.255 ;
      RECT 17157.625 189.04 17157.905 336.495 ;
      RECT 17157.065 187.94 17157.345 336.735 ;
      RECT 17156.505 189.04 17156.785 336.975 ;
      RECT 17155.945 187.94 17156.225 337.215 ;
      RECT 17155.385 189.04 17155.665 337.455 ;
      RECT 17154.825 189.04 17155.105 337.695 ;
      RECT 17154.265 189.04 17154.545 337.695 ;
      RECT 17153.705 189.04 17153.985 337.455 ;
      RECT 17153.145 189.04 17153.425 337.215 ;
      RECT 17152.585 189.04 17152.865 336.975 ;
      RECT 17152.025 189.04 17152.305 336.735 ;
      RECT 17151.465 189.04 17151.745 336.495 ;
      RECT 17150.905 189.04 17151.185 336.255 ;
      RECT 17150.345 189.04 17150.625 336.015 ;
      RECT 17149.785 189.04 17150.065 335.775 ;
      RECT 17140.825 189.04 17141.105 335.29 ;
      RECT 17140.265 187.94 17140.545 335.05 ;
      RECT 17139.705 189.04 17139.985 334.81 ;
      RECT 17139.145 187.94 17139.425 334.57 ;
      RECT 17138.585 189.04 17138.865 334.33 ;
      RECT 17138.025 187.94 17138.305 334.09 ;
      RECT 17137.465 189.04 17137.745 333.85 ;
      RECT 17136.905 189.04 17137.185 333.61 ;
      RECT 17136.345 189.04 17136.625 333.37 ;
      RECT 17135.785 189.04 17136.065 333.13 ;
      RECT 17135.225 189.04 17135.505 332.89 ;
      RECT 17134.665 189.04 17134.945 332.65 ;
      RECT 17134.105 189.04 17134.385 332.41 ;
      RECT 17133.545 189.04 17133.825 332.17 ;
      RECT 17131.025 187.94 17131.305 333.89 ;
      RECT 17130.465 189.04 17130.745 333.65 ;
      RECT 17129.905 187.94 17130.185 333.41 ;
      RECT 17129.345 189.04 17129.625 333.17 ;
      RECT 17128.785 189.04 17129.065 332.93 ;
      RECT 17128.225 189.04 17128.505 332.69 ;
      RECT 17127.665 189.04 17127.945 332.45 ;
      RECT 17127.105 189.04 17127.385 332.21 ;
      RECT 17101.065 189.04 17101.345 329.86 ;
      RECT 17100.505 189.04 17100.785 330.1 ;
      RECT 17099.945 189.04 17100.225 330.34 ;
      RECT 17099.385 189.04 17099.665 330.585 ;
      RECT 17098.825 189.04 17099.105 330.825 ;
      RECT 17098.265 189.04 17098.545 331.065 ;
      RECT 17097.705 189.04 17097.985 331.065 ;
      RECT 17097.145 189.04 17097.425 330.825 ;
      RECT 17096.585 189.04 17096.865 330.585 ;
      RECT 17096.025 187.94 17096.305 330.345 ;
      RECT 17095.465 189.04 17095.745 330.105 ;
      RECT 17094.905 187.94 17095.185 329.865 ;
      RECT 17094.345 189.04 17094.625 329.625 ;
      RECT 17093.785 189.04 17094.065 329.385 ;
      RECT 17093.225 189.04 17093.505 329.145 ;
      RECT 17092.665 187.94 17092.945 328.905 ;
      RECT 17092.105 189.04 17092.385 328.665 ;
      RECT 17091.545 187.94 17091.825 328.425 ;
      RECT 17090.985 189.04 17091.265 328.185 ;
      RECT 17090.425 187.94 17090.705 327.945 ;
      RECT 17089.865 189.04 17090.145 327.705 ;
      RECT 17089.305 189.04 17089.585 327.465 ;
      RECT 17088.745 189.04 17089.025 327.225 ;
      RECT 17088.185 189.04 17088.465 326.985 ;
      RECT 17074.745 189.04 17075.025 332.785 ;
      RECT 17074.185 189.04 17074.465 332.545 ;
      RECT 17073.625 189.04 17073.905 332.305 ;
      RECT 17073.065 189.04 17073.345 332.065 ;
      RECT 17072.505 189.04 17072.785 331.825 ;
      RECT 17071.945 189.04 17072.225 331.585 ;
      RECT 17071.385 189.04 17071.665 331.345 ;
      RECT 17070.825 189.04 17071.105 331.105 ;
      RECT 17070.265 187.94 17070.545 330.865 ;
      RECT 17069.705 189.04 17069.985 330.625 ;
      RECT 17069.145 187.94 17069.425 330.305 ;
      RECT 17068.585 189.04 17068.865 330.145 ;
      RECT 17068.025 187.94 17068.305 329.905 ;
      RECT 17067.465 189.04 17067.745 329.665 ;
      RECT 17066.905 189.04 17067.185 329.425 ;
      RECT 17066.345 189.04 17066.625 329.185 ;
      RECT 17065.785 189.04 17066.065 328.945 ;
      RECT 17065.225 189.04 17065.505 328.705 ;
      RECT 17064.665 189.04 17064.945 328.465 ;
      RECT 17064.105 189.04 17064.385 328.225 ;
      RECT 17063.545 189.04 17063.825 327.985 ;
      RECT 17062.985 187.94 17063.265 327.745 ;
      RECT 17062.425 189.04 17062.705 327.505 ;
      RECT 17061.865 187.94 17062.145 327.265 ;
      RECT 17022.665 189.04 17022.945 332.875 ;
      RECT 17022.105 189.04 17022.385 333.115 ;
      RECT 17021.545 189.04 17021.825 333.355 ;
      RECT 17020.985 189.04 17021.265 333.595 ;
      RECT 17020.425 189.04 17020.705 333.835 ;
      RECT 17019.865 189.04 17020.145 334.075 ;
      RECT 17019.305 189.04 17019.585 334.315 ;
      RECT 17018.745 189.04 17019.025 334.555 ;
      RECT 17018.185 189.04 17018.465 334.795 ;
      RECT 17017.625 189.04 17017.905 335.035 ;
      RECT 17017.065 189.04 17017.345 335.275 ;
      RECT 17016.505 189.04 17016.785 335.515 ;
      RECT 17015.945 189.04 17016.225 335.755 ;
      RECT 17015.385 189.04 17015.665 335.755 ;
      RECT 17014.825 187.94 17015.105 335.515 ;
      RECT 17014.265 189.04 17014.545 335.275 ;
      RECT 17013.705 187.94 17013.985 335.035 ;
      RECT 17013.145 189.04 17013.425 334.795 ;
      RECT 17012.585 189.04 17012.865 334.555 ;
      RECT 17012.025 189.04 17012.305 334.315 ;
      RECT 17011.465 187.94 17011.745 334.05 ;
      RECT 17010.905 189.04 17011.185 333.81 ;
      RECT 17010.345 187.94 17010.625 333.57 ;
      RECT 17009.785 189.04 17010.065 333.33 ;
      RECT 17000.825 187.94 17001.105 327.165 ;
      RECT 17000.265 189.04 17000.545 327.405 ;
      RECT 16999.705 189.04 16999.985 327.645 ;
      RECT 16999.145 189.04 16999.425 327.645 ;
      RECT 16998.585 189.04 16998.865 327.405 ;
      RECT 16998.025 189.04 16998.305 327.165 ;
      RECT 16997.465 189.04 16997.745 326.925 ;
      RECT 16996.905 189.04 16997.185 326.685 ;
      RECT 16996.345 189.04 16996.625 326.445 ;
      RECT 16995.785 189.04 16996.065 326.205 ;
      RECT 16995.225 189.04 16995.505 325.965 ;
      RECT 16994.665 189.04 16994.945 325.725 ;
      RECT 16994.105 189.04 16994.385 325.485 ;
      RECT 16993.545 187.94 16993.825 325.245 ;
      RECT 16991.025 189.04 16991.305 326.965 ;
      RECT 16990.465 187.94 16990.745 326.725 ;
      RECT 16989.905 189.04 16990.185 326.485 ;
      RECT 16989.345 187.94 16989.625 326.245 ;
      RECT 16988.785 189.04 16989.065 326.005 ;
      RECT 16988.225 189.04 16988.505 325.765 ;
      RECT 16987.665 189.04 16987.945 325.525 ;
      RECT 16961.625 189.04 16961.905 328.31 ;
      RECT 16961.065 189.04 16961.345 328.55 ;
      RECT 16960.505 189.04 16960.785 328.79 ;
      RECT 16959.945 189.04 16960.225 329.03 ;
      RECT 16959.385 189.04 16959.665 329.27 ;
      RECT 16958.825 187.94 16959.105 329.51 ;
      RECT 16958.265 189.04 16958.545 329.75 ;
      RECT 16957.705 187.94 16957.985 329.99 ;
      RECT 16957.145 189.04 16957.425 330.23 ;
      RECT 16956.585 189.04 16956.865 330.47 ;
      RECT 16956.025 189.04 16956.305 330.71 ;
      RECT 16955.465 189.04 16955.745 330.95 ;
      RECT 16954.905 189.04 16955.185 331.19 ;
      RECT 16954.345 189.04 16954.625 331.43 ;
      RECT 16953.785 189.04 16954.065 331.67 ;
      RECT 16953.225 189.04 16953.505 331.67 ;
      RECT 16952.665 189.04 16952.945 331.43 ;
      RECT 16952.105 189.04 16952.385 331.19 ;
      RECT 16951.545 189.04 16951.825 330.95 ;
      RECT 16950.985 189.04 16951.265 330.705 ;
      RECT 16950.425 189.04 16950.705 330.465 ;
      RECT 16949.865 189.04 16950.145 330.225 ;
      RECT 16949.305 187.94 16949.585 329.985 ;
      RECT 16948.745 189.04 16949.025 329.745 ;
      RECT 16935.305 187.94 16935.585 327.225 ;
      RECT 16934.745 189.04 16935.025 326.985 ;
      RECT 16934.185 189.04 16934.465 326.745 ;
      RECT 16933.625 189.04 16933.905 326.505 ;
      RECT 16933.065 187.94 16933.345 326.265 ;
      RECT 16932.505 189.04 16932.785 326.025 ;
      RECT 16931.945 187.94 16932.225 325.785 ;
      RECT 16931.385 189.04 16931.665 325.545 ;
      RECT 16930.825 187.94 16931.105 325.305 ;
      RECT 16930.265 189.04 16930.545 325.065 ;
      RECT 16929.705 189.04 16929.985 324.825 ;
      RECT 16929.145 189.04 16929.425 324.585 ;
      RECT 16928.585 189.04 16928.865 324.345 ;
      RECT 16928.025 189.04 16928.305 324.105 ;
      RECT 16927.465 189.04 16927.745 323.865 ;
      RECT 16926.905 189.04 16927.185 323.625 ;
      RECT 16926.345 189.04 16926.625 323.385 ;
      RECT 16925.785 189.04 16926.065 323.145 ;
      RECT 16925.225 189.04 16925.505 322.905 ;
      RECT 16924.665 189.04 16924.945 322.665 ;
      RECT 16924.105 189.04 16924.385 322.425 ;
      RECT 16923.545 187.94 16923.825 322.185 ;
      RECT 16922.985 189.04 16923.265 321.945 ;
      RECT 16922.425 187.94 16922.705 321.705 ;
      RECT 16882.665 189.04 16882.945 332.175 ;
      RECT 16882.105 187.94 16882.385 332.415 ;
      RECT 16881.545 189.04 16881.825 332.655 ;
      RECT 16880.985 189.04 16881.265 332.895 ;
      RECT 16880.425 189.04 16880.705 333.135 ;
      RECT 16879.865 189.04 16880.145 333.375 ;
      RECT 16879.305 189.04 16879.585 333.615 ;
      RECT 16878.745 189.04 16879.025 333.86 ;
      RECT 16878.185 189.04 16878.465 334.1 ;
      RECT 16877.625 189.04 16877.905 334.34 ;
      RECT 16877.065 187.94 16877.345 334.58 ;
      RECT 16876.505 189.04 16876.785 334.82 ;
      RECT 16875.945 187.94 16876.225 335.06 ;
      RECT 16875.385 189.04 16875.665 335.3 ;
      RECT 16874.825 189.04 16875.105 335.54 ;
      RECT 16874.265 189.04 16874.545 335.78 ;
      RECT 16873.705 189.04 16873.985 336.02 ;
      RECT 16873.145 189.04 16873.425 336.26 ;
      RECT 16872.585 189.04 16872.865 336.5 ;
      RECT 16872.025 189.04 16872.305 336.74 ;
      RECT 16871.465 189.04 16871.745 336.98 ;
      RECT 16870.905 189.04 16871.185 337.22 ;
      RECT 16870.345 189.04 16870.625 337.46 ;
      RECT 16869.785 189.04 16870.065 337.7 ;
      RECT 16860.825 189.04 16861.105 333.285 ;
      RECT 16860.265 189.04 16860.545 333.045 ;
      RECT 16859.705 189.04 16859.985 332.805 ;
      RECT 16859.145 187.94 16859.425 332.565 ;
      RECT 16858.585 189.04 16858.865 332.325 ;
      RECT 16858.025 187.94 16858.305 332.085 ;
      RECT 16857.465 189.04 16857.745 331.845 ;
      RECT 16856.905 189.04 16857.185 331.605 ;
      RECT 16856.345 189.04 16856.625 331.365 ;
      RECT 16855.785 187.94 16856.065 331.125 ;
      RECT 16855.225 189.04 16855.505 330.885 ;
      RECT 16854.665 187.94 16854.945 330.645 ;
      RECT 16854.105 189.04 16854.385 330.405 ;
      RECT 16853.545 187.94 16853.825 330.165 ;
      RECT 16851.025 189.04 16851.305 322.565 ;
      RECT 16850.465 189.04 16850.745 322.325 ;
      RECT 16849.905 189.04 16850.185 322.085 ;
      RECT 16849.345 189.04 16849.625 321.845 ;
      RECT 16848.785 189.04 16849.065 321.605 ;
      RECT 16848.225 189.04 16848.505 321.365 ;
      RECT 16847.665 189.04 16847.945 321.125 ;
      RECT 16821.625 189.04 16821.905 335 ;
      RECT 16821.065 189.04 16821.345 335.24 ;
      RECT 16820.505 189.04 16820.785 335.48 ;
      RECT 16819.945 189.04 16820.225 335.72 ;
      RECT 16819.385 189.04 16819.665 335.96 ;
      RECT 16818.825 187.94 16819.105 335.96 ;
      RECT 16818.265 189.04 16818.545 335.72 ;
      RECT 16817.705 187.94 16817.985 335.475 ;
      RECT 16817.145 189.04 16817.425 335.235 ;
      RECT 16816.585 187.94 16816.865 334.995 ;
      RECT 16816.025 189.04 16816.305 334.755 ;
      RECT 16815.465 189.04 16815.745 334.515 ;
      RECT 16814.905 189.04 16815.185 334.275 ;
      RECT 16814.345 189.04 16814.625 334.035 ;
      RECT 16813.785 189.04 16814.065 333.795 ;
      RECT 16813.225 189.04 16813.505 333.555 ;
      RECT 16812.665 189.04 16812.945 333.315 ;
      RECT 16812.105 189.04 16812.385 333.075 ;
      RECT 16811.545 187.94 16811.825 332.835 ;
      RECT 16810.985 189.04 16811.265 332.595 ;
      RECT 16810.425 187.94 16810.705 332.355 ;
      RECT 16809.865 189.04 16810.145 332.115 ;
      RECT 16809.305 189.04 16809.585 331.875 ;
      RECT 16808.745 189.04 16809.025 331.635 ;
      RECT 16795.305 189.04 16795.585 335.035 ;
      RECT 16794.745 189.04 16795.025 335.275 ;
      RECT 16794.185 189.04 16794.465 335.52 ;
      RECT 16793.625 189.04 16793.905 335.76 ;
      RECT 16793.065 189.04 16793.345 336 ;
      RECT 16792.505 189.04 16792.785 336 ;
      RECT 16791.945 189.04 16792.225 335.76 ;
      RECT 16791.385 189.04 16791.665 335.52 ;
      RECT 16790.825 189.04 16791.105 328.505 ;
      RECT 16790.265 189.04 16790.545 328.265 ;
      RECT 16789.705 189.04 16789.985 328.025 ;
      RECT 16789.145 187.94 16789.425 327.785 ;
      RECT 16788.585 189.04 16788.865 327.545 ;
      RECT 16788.025 187.94 16788.305 327.305 ;
      RECT 16787.465 189.04 16787.745 327.065 ;
      RECT 16786.905 189.04 16787.185 326.825 ;
      RECT 16786.345 189.04 16786.625 326.585 ;
      RECT 16785.785 187.94 16786.065 326.345 ;
      RECT 16785.225 189.04 16785.505 326.105 ;
      RECT 16784.665 187.94 16784.945 325.865 ;
      RECT 16784.105 189.04 16784.385 325.625 ;
      RECT 16783.545 187.94 16783.825 325.385 ;
      RECT 16782.985 189.04 16783.265 325.145 ;
      RECT 16782.425 189.04 16782.705 324.905 ;
      RECT 16742.105 189.04 16742.385 333.8 ;
      RECT 16741.545 189.04 16741.825 334.04 ;
      RECT 16740.985 189.04 16741.265 334.285 ;
      RECT 16740.425 189.04 16740.705 334.525 ;
      RECT 16739.865 189.04 16740.145 334.765 ;
      RECT 16739.305 189.04 16739.585 335.005 ;
      RECT 16738.745 189.04 16739.025 335.245 ;
      RECT 16738.185 189.04 16738.465 335.485 ;
      RECT 16737.625 189.04 16737.905 335.725 ;
      RECT 16737.065 189.04 16737.345 335.965 ;
      RECT 16736.505 187.94 16736.785 336.205 ;
      RECT 16735.945 189.04 16736.225 336.445 ;
      RECT 16735.385 187.94 16735.665 336.685 ;
      RECT 16734.825 189.04 16735.105 336.925 ;
      RECT 16734.265 187.94 16734.545 337.165 ;
      RECT 16733.705 189.04 16733.985 337.165 ;
      RECT 16733.145 189.04 16733.425 336.925 ;
      RECT 16732.585 189.04 16732.865 336.685 ;
      RECT 16732.025 189.04 16732.305 336.445 ;
      RECT 16731.465 189.04 16731.745 336.205 ;
      RECT 16730.905 189.04 16731.185 335.965 ;
      RECT 16730.345 189.04 16730.625 335.725 ;
      RECT 16729.785 189.04 16730.065 335.485 ;
      RECT 16720.825 187.94 16721.105 335.515 ;
      RECT 16720.265 189.04 16720.545 335.755 ;
      RECT 16719.705 187.94 16719.985 335.995 ;
      RECT 16719.145 189.04 16719.425 336.21 ;
      RECT 16718.585 189.04 16718.865 335.785 ;
      RECT 16718.025 189.04 16718.305 335.545 ;
      RECT 16717.465 189.04 16717.745 335.305 ;
      RECT 16716.905 189.04 16717.185 335.065 ;
      RECT 16716.345 189.04 16716.625 334.825 ;
      RECT 16715.785 189.04 16716.065 334.585 ;
      RECT 16715.225 189.04 16715.505 334.345 ;
      RECT 16714.665 189.04 16714.945 334.105 ;
      RECT 16714.105 189.04 16714.385 333.865 ;
      RECT 16713.545 189.04 16713.825 333.625 ;
      RECT 16711.025 189.04 16711.305 332.8 ;
      RECT 16710.465 189.04 16710.745 332.56 ;
      RECT 16709.905 189.04 16710.185 332.32 ;
      RECT 16709.345 187.94 16709.625 332.08 ;
      RECT 16708.785 189.04 16709.065 331.84 ;
      RECT 16708.225 187.94 16708.505 331.6 ;
      RECT 16707.665 189.04 16707.945 331.36 ;
      RECT 16707.105 189.04 16707.385 331.12 ;
      RECT 16680.505 189.04 16680.785 342.165 ;
      RECT 16679.945 187.94 16680.225 342.405 ;
      RECT 16679.385 189.04 16679.665 342.645 ;
      RECT 16678.825 187.94 16679.105 342.89 ;
      RECT 16678.265 189.04 16678.545 343.13 ;
      RECT 16677.705 187.94 16677.985 343.37 ;
      RECT 16677.145 189.04 16677.425 343.61 ;
      RECT 16676.585 189.04 16676.865 343.85 ;
      RECT 16676.025 189.04 16676.305 329.47 ;
      RECT 16675.465 189.04 16675.745 329.23 ;
      RECT 16674.905 189.04 16675.185 328.99 ;
      RECT 16674.345 189.04 16674.625 328.75 ;
      RECT 16673.785 189.04 16674.065 328.51 ;
      RECT 16673.225 189.04 16673.505 328.27 ;
      RECT 16672.665 189.04 16672.945 328.03 ;
      RECT 16672.105 189.04 16672.385 327.79 ;
      RECT 16671.545 189.04 16671.825 327.55 ;
      RECT 16670.985 189.04 16671.265 327.31 ;
      RECT 16670.425 187.94 16670.705 327.07 ;
      RECT 16669.865 189.04 16670.145 326.83 ;
      RECT 16669.305 187.94 16669.585 326.59 ;
      RECT 16668.745 189.04 16669.025 326.35 ;
      RECT 16654.745 187.94 16655.025 332.47 ;
      RECT 16654.185 189.04 16654.465 332.23 ;
      RECT 16653.625 189.04 16653.905 331.99 ;
      RECT 16653.065 189.04 16653.345 331.75 ;
      RECT 16652.505 189.04 16652.785 331.51 ;
      RECT 16651.945 189.04 16652.225 331.27 ;
      RECT 16651.385 189.04 16651.665 331.03 ;
      RECT 16650.825 189.04 16651.105 330.79 ;
      RECT 16650.265 189.04 16650.545 330.55 ;
      RECT 16649.705 187.94 16649.985 330.31 ;
      RECT 16649.145 189.04 16649.425 330.07 ;
      RECT 16648.585 187.94 16648.865 329.83 ;
      RECT 16648.025 189.04 16648.305 329.59 ;
      RECT 16647.465 189.04 16647.745 329.35 ;
      RECT 16646.905 189.04 16647.185 329.11 ;
      RECT 16646.345 189.04 16646.625 328.87 ;
      RECT 16645.785 189.04 16646.065 328.63 ;
      RECT 16645.225 189.04 16645.505 328.39 ;
      RECT 16644.665 189.04 16644.945 328.15 ;
      RECT 16644.105 189.04 16644.385 327.91 ;
      RECT 16643.545 189.04 16643.825 327.67 ;
      RECT 16642.985 189.04 16643.265 327.43 ;
      RECT 16642.425 189.04 16642.705 327.19 ;
      RECT 16603.225 189.04 16603.505 334.095 ;
      RECT 16602.665 189.04 16602.945 334.335 ;
      RECT 16602.105 189.04 16602.385 334.575 ;
      RECT 16601.545 187.94 16601.825 334.815 ;
      RECT 16600.985 189.04 16601.265 335.055 ;
      RECT 16600.425 187.94 16600.705 335.295 ;
      RECT 16599.865 189.04 16600.145 335.535 ;
      RECT 16599.305 189.04 16599.585 335.775 ;
      RECT 16598.745 189.04 16599.025 336.015 ;
      RECT 16598.185 187.94 16598.465 336.255 ;
      RECT 16597.625 189.04 16597.905 336.495 ;
      RECT 16597.065 187.94 16597.345 336.735 ;
      RECT 16596.505 189.04 16596.785 336.975 ;
      RECT 16595.945 187.94 16596.225 337.215 ;
      RECT 16595.385 189.04 16595.665 337.455 ;
      RECT 16594.825 189.04 16595.105 337.695 ;
      RECT 16594.265 189.04 16594.545 337.695 ;
      RECT 16593.705 189.04 16593.985 337.455 ;
      RECT 16593.145 189.04 16593.425 337.215 ;
      RECT 16592.585 189.04 16592.865 336.975 ;
      RECT 16592.025 189.04 16592.305 336.735 ;
      RECT 16591.465 189.04 16591.745 336.495 ;
      RECT 16590.905 189.04 16591.185 336.255 ;
      RECT 16590.345 189.04 16590.625 336.015 ;
      RECT 16589.785 189.04 16590.065 335.775 ;
      RECT 16580.825 189.04 16581.105 335.29 ;
      RECT 16580.265 187.94 16580.545 335.05 ;
      RECT 16579.705 189.04 16579.985 334.81 ;
      RECT 16579.145 187.94 16579.425 334.57 ;
      RECT 16578.585 189.04 16578.865 334.33 ;
      RECT 16578.025 187.94 16578.305 334.09 ;
      RECT 16577.465 189.04 16577.745 333.85 ;
      RECT 16576.905 189.04 16577.185 333.61 ;
      RECT 16576.345 189.04 16576.625 333.37 ;
      RECT 16575.785 189.04 16576.065 333.13 ;
      RECT 16575.225 189.04 16575.505 332.89 ;
      RECT 16574.665 189.04 16574.945 332.65 ;
      RECT 16574.105 189.04 16574.385 332.41 ;
      RECT 16573.545 189.04 16573.825 332.17 ;
      RECT 16571.025 187.94 16571.305 333.89 ;
      RECT 16570.465 189.04 16570.745 333.65 ;
      RECT 16569.905 187.94 16570.185 333.41 ;
      RECT 16569.345 189.04 16569.625 333.17 ;
      RECT 16568.785 189.04 16569.065 332.93 ;
      RECT 16568.225 189.04 16568.505 332.69 ;
      RECT 16567.665 189.04 16567.945 332.45 ;
      RECT 16567.105 189.04 16567.385 332.21 ;
      RECT 16541.065 189.04 16541.345 329.86 ;
      RECT 16540.505 189.04 16540.785 330.1 ;
      RECT 16539.945 189.04 16540.225 330.34 ;
      RECT 16539.385 189.04 16539.665 330.585 ;
      RECT 16538.825 189.04 16539.105 330.825 ;
      RECT 16538.265 189.04 16538.545 331.065 ;
      RECT 16537.705 189.04 16537.985 331.065 ;
      RECT 16537.145 189.04 16537.425 330.825 ;
      RECT 16536.585 189.04 16536.865 330.585 ;
      RECT 16536.025 187.94 16536.305 330.345 ;
      RECT 16535.465 189.04 16535.745 330.105 ;
      RECT 16534.905 187.94 16535.185 329.865 ;
      RECT 16534.345 189.04 16534.625 329.625 ;
      RECT 16533.785 189.04 16534.065 329.385 ;
      RECT 16533.225 189.04 16533.505 329.145 ;
      RECT 16532.665 187.94 16532.945 328.905 ;
      RECT 16532.105 189.04 16532.385 328.665 ;
      RECT 16531.545 187.94 16531.825 328.425 ;
      RECT 16530.985 189.04 16531.265 328.185 ;
      RECT 16530.425 187.94 16530.705 327.945 ;
      RECT 16529.865 189.04 16530.145 327.705 ;
      RECT 16529.305 189.04 16529.585 327.465 ;
      RECT 16528.745 189.04 16529.025 327.225 ;
      RECT 16528.185 189.04 16528.465 326.985 ;
      RECT 16514.745 189.04 16515.025 332.785 ;
      RECT 16514.185 189.04 16514.465 332.545 ;
      RECT 16513.625 189.04 16513.905 332.305 ;
      RECT 16513.065 189.04 16513.345 332.065 ;
      RECT 16512.505 189.04 16512.785 331.825 ;
      RECT 16511.945 189.04 16512.225 331.585 ;
      RECT 16511.385 189.04 16511.665 331.345 ;
      RECT 16510.825 189.04 16511.105 331.105 ;
      RECT 16510.265 187.94 16510.545 330.865 ;
      RECT 16509.705 189.04 16509.985 330.625 ;
      RECT 16509.145 187.94 16509.425 330.305 ;
      RECT 16508.585 189.04 16508.865 330.145 ;
      RECT 16508.025 187.94 16508.305 329.905 ;
      RECT 16507.465 189.04 16507.745 329.665 ;
      RECT 16506.905 189.04 16507.185 329.425 ;
      RECT 16506.345 189.04 16506.625 329.185 ;
      RECT 16505.785 189.04 16506.065 328.945 ;
      RECT 16505.225 189.04 16505.505 328.705 ;
      RECT 16504.665 189.04 16504.945 328.465 ;
      RECT 16504.105 189.04 16504.385 328.225 ;
      RECT 16503.545 189.04 16503.825 327.985 ;
      RECT 16502.985 187.94 16503.265 327.745 ;
      RECT 16502.425 189.04 16502.705 327.505 ;
      RECT 16501.865 187.94 16502.145 327.265 ;
      RECT 16462.665 189.04 16462.945 332.875 ;
      RECT 16462.105 189.04 16462.385 333.115 ;
      RECT 16461.545 189.04 16461.825 333.355 ;
      RECT 16460.985 189.04 16461.265 333.595 ;
      RECT 16460.425 189.04 16460.705 333.835 ;
      RECT 16459.865 189.04 16460.145 334.075 ;
      RECT 16459.305 189.04 16459.585 334.315 ;
      RECT 16458.745 189.04 16459.025 334.555 ;
      RECT 16458.185 189.04 16458.465 334.795 ;
      RECT 16457.625 189.04 16457.905 335.035 ;
      RECT 16457.065 189.04 16457.345 335.275 ;
      RECT 16456.505 189.04 16456.785 335.515 ;
      RECT 16455.945 189.04 16456.225 335.755 ;
      RECT 16455.385 189.04 16455.665 335.755 ;
      RECT 16454.825 187.94 16455.105 335.515 ;
      RECT 16454.265 189.04 16454.545 335.275 ;
      RECT 16453.705 187.94 16453.985 335.035 ;
      RECT 16453.145 189.04 16453.425 334.795 ;
      RECT 16452.585 189.04 16452.865 334.555 ;
      RECT 16452.025 189.04 16452.305 334.315 ;
      RECT 16451.465 187.94 16451.745 334.05 ;
      RECT 16450.905 189.04 16451.185 333.81 ;
      RECT 16450.345 187.94 16450.625 333.57 ;
      RECT 16449.785 189.04 16450.065 333.33 ;
      RECT 16440.825 187.94 16441.105 327.165 ;
      RECT 16440.265 189.04 16440.545 327.405 ;
      RECT 16439.705 189.04 16439.985 327.645 ;
      RECT 16439.145 189.04 16439.425 327.645 ;
      RECT 16438.585 189.04 16438.865 327.405 ;
      RECT 16438.025 189.04 16438.305 327.165 ;
      RECT 16437.465 189.04 16437.745 326.925 ;
      RECT 16436.905 189.04 16437.185 326.685 ;
      RECT 16436.345 189.04 16436.625 326.445 ;
      RECT 16435.785 189.04 16436.065 326.205 ;
      RECT 16435.225 189.04 16435.505 325.965 ;
      RECT 16434.665 189.04 16434.945 325.725 ;
      RECT 16434.105 189.04 16434.385 325.485 ;
      RECT 16433.545 187.94 16433.825 325.245 ;
      RECT 16431.025 189.04 16431.305 326.965 ;
      RECT 16430.465 187.94 16430.745 326.725 ;
      RECT 16429.905 189.04 16430.185 326.485 ;
      RECT 16429.345 187.94 16429.625 326.245 ;
      RECT 16428.785 189.04 16429.065 326.005 ;
      RECT 16428.225 189.04 16428.505 325.765 ;
      RECT 16427.665 189.04 16427.945 325.525 ;
      RECT 16401.625 189.04 16401.905 328.31 ;
      RECT 16401.065 189.04 16401.345 328.55 ;
      RECT 16400.505 189.04 16400.785 328.79 ;
      RECT 16399.945 189.04 16400.225 329.03 ;
      RECT 16399.385 189.04 16399.665 329.27 ;
      RECT 16398.825 187.94 16399.105 329.51 ;
      RECT 16398.265 189.04 16398.545 329.75 ;
      RECT 16397.705 187.94 16397.985 329.99 ;
      RECT 16397.145 189.04 16397.425 330.23 ;
      RECT 16396.585 189.04 16396.865 330.47 ;
      RECT 16396.025 189.04 16396.305 330.71 ;
      RECT 16395.465 189.04 16395.745 330.95 ;
      RECT 16394.905 189.04 16395.185 331.19 ;
      RECT 16394.345 189.04 16394.625 331.43 ;
      RECT 16393.785 189.04 16394.065 331.67 ;
      RECT 16393.225 189.04 16393.505 331.67 ;
      RECT 16392.665 189.04 16392.945 331.43 ;
      RECT 16392.105 189.04 16392.385 331.19 ;
      RECT 16391.545 189.04 16391.825 330.95 ;
      RECT 16390.985 189.04 16391.265 330.705 ;
      RECT 16390.425 189.04 16390.705 330.465 ;
      RECT 16389.865 189.04 16390.145 330.225 ;
      RECT 16389.305 187.94 16389.585 329.985 ;
      RECT 16388.745 189.04 16389.025 329.745 ;
      RECT 16375.305 187.94 16375.585 327.225 ;
      RECT 16374.745 189.04 16375.025 326.985 ;
      RECT 16374.185 189.04 16374.465 326.745 ;
      RECT 16373.625 189.04 16373.905 326.505 ;
      RECT 16373.065 187.94 16373.345 326.265 ;
      RECT 16372.505 189.04 16372.785 326.025 ;
      RECT 16371.945 187.94 16372.225 325.785 ;
      RECT 16371.385 189.04 16371.665 325.545 ;
      RECT 16370.825 187.94 16371.105 325.305 ;
      RECT 16370.265 189.04 16370.545 325.065 ;
      RECT 16369.705 189.04 16369.985 324.825 ;
      RECT 16369.145 189.04 16369.425 324.585 ;
      RECT 16368.585 189.04 16368.865 324.345 ;
      RECT 16368.025 189.04 16368.305 324.105 ;
      RECT 16367.465 189.04 16367.745 323.865 ;
      RECT 16366.905 189.04 16367.185 323.625 ;
      RECT 16366.345 189.04 16366.625 323.385 ;
      RECT 16365.785 189.04 16366.065 323.145 ;
      RECT 16365.225 189.04 16365.505 322.905 ;
      RECT 16364.665 189.04 16364.945 322.665 ;
      RECT 16364.105 189.04 16364.385 322.425 ;
      RECT 16363.545 187.94 16363.825 322.185 ;
      RECT 16362.985 189.04 16363.265 321.945 ;
      RECT 16362.425 187.94 16362.705 321.705 ;
      RECT 16322.665 189.04 16322.945 332.175 ;
      RECT 16322.105 187.94 16322.385 332.415 ;
      RECT 16321.545 189.04 16321.825 332.655 ;
      RECT 16320.985 189.04 16321.265 332.895 ;
      RECT 16320.425 189.04 16320.705 333.135 ;
      RECT 16319.865 189.04 16320.145 333.375 ;
      RECT 16319.305 189.04 16319.585 333.615 ;
      RECT 16318.745 189.04 16319.025 333.86 ;
      RECT 16318.185 189.04 16318.465 334.1 ;
      RECT 16317.625 189.04 16317.905 334.34 ;
      RECT 16317.065 187.94 16317.345 334.58 ;
      RECT 16316.505 189.04 16316.785 334.82 ;
      RECT 16315.945 187.94 16316.225 335.06 ;
      RECT 16315.385 189.04 16315.665 335.3 ;
      RECT 16314.825 189.04 16315.105 335.54 ;
      RECT 16314.265 189.04 16314.545 335.78 ;
      RECT 16313.705 189.04 16313.985 336.02 ;
      RECT 16313.145 189.04 16313.425 336.26 ;
      RECT 16312.585 189.04 16312.865 336.5 ;
      RECT 16312.025 189.04 16312.305 336.74 ;
      RECT 16311.465 189.04 16311.745 336.98 ;
      RECT 16310.905 189.04 16311.185 337.22 ;
      RECT 16310.345 189.04 16310.625 337.46 ;
      RECT 16309.785 189.04 16310.065 337.7 ;
      RECT 16300.825 189.04 16301.105 333.285 ;
      RECT 16300.265 189.04 16300.545 333.045 ;
      RECT 16299.705 189.04 16299.985 332.805 ;
      RECT 16299.145 187.94 16299.425 332.565 ;
      RECT 16298.585 189.04 16298.865 332.325 ;
      RECT 16298.025 187.94 16298.305 332.085 ;
      RECT 16297.465 189.04 16297.745 331.845 ;
      RECT 16296.905 189.04 16297.185 331.605 ;
      RECT 16296.345 189.04 16296.625 331.365 ;
      RECT 16295.785 187.94 16296.065 331.125 ;
      RECT 16295.225 189.04 16295.505 330.885 ;
      RECT 16294.665 187.94 16294.945 330.645 ;
      RECT 16294.105 189.04 16294.385 330.405 ;
      RECT 16293.545 187.94 16293.825 330.165 ;
      RECT 16291.025 189.04 16291.305 322.565 ;
      RECT 16290.465 189.04 16290.745 322.325 ;
      RECT 16289.905 189.04 16290.185 322.085 ;
      RECT 16289.345 189.04 16289.625 321.845 ;
      RECT 16288.785 189.04 16289.065 321.605 ;
      RECT 16288.225 189.04 16288.505 321.365 ;
      RECT 16287.665 189.04 16287.945 321.125 ;
      RECT 16261.625 189.04 16261.905 335 ;
      RECT 16261.065 189.04 16261.345 335.24 ;
      RECT 16260.505 189.04 16260.785 335.48 ;
      RECT 16259.945 189.04 16260.225 335.72 ;
      RECT 16259.385 189.04 16259.665 335.96 ;
      RECT 16258.825 187.94 16259.105 335.96 ;
      RECT 16258.265 189.04 16258.545 335.72 ;
      RECT 16257.705 187.94 16257.985 335.475 ;
      RECT 16257.145 189.04 16257.425 335.235 ;
      RECT 16256.585 187.94 16256.865 334.995 ;
      RECT 16256.025 189.04 16256.305 334.755 ;
      RECT 16255.465 189.04 16255.745 334.515 ;
      RECT 16254.905 189.04 16255.185 334.275 ;
      RECT 16254.345 189.04 16254.625 334.035 ;
      RECT 16253.785 189.04 16254.065 333.795 ;
      RECT 16253.225 189.04 16253.505 333.555 ;
      RECT 16252.665 189.04 16252.945 333.315 ;
      RECT 16252.105 189.04 16252.385 333.075 ;
      RECT 16251.545 187.94 16251.825 332.835 ;
      RECT 16250.985 189.04 16251.265 332.595 ;
      RECT 16250.425 187.94 16250.705 332.355 ;
      RECT 16249.865 189.04 16250.145 332.115 ;
      RECT 16249.305 189.04 16249.585 331.875 ;
      RECT 16248.745 189.04 16249.025 331.635 ;
      RECT 16235.305 189.04 16235.585 335.035 ;
      RECT 16234.745 189.04 16235.025 335.275 ;
      RECT 16234.185 189.04 16234.465 335.52 ;
      RECT 16233.625 189.04 16233.905 335.76 ;
      RECT 16233.065 189.04 16233.345 336 ;
      RECT 16232.505 189.04 16232.785 336 ;
      RECT 16231.945 189.04 16232.225 335.76 ;
      RECT 16231.385 189.04 16231.665 335.52 ;
      RECT 16230.825 189.04 16231.105 328.505 ;
      RECT 16230.265 189.04 16230.545 328.265 ;
      RECT 16229.705 189.04 16229.985 328.025 ;
      RECT 16229.145 187.94 16229.425 327.785 ;
      RECT 16228.585 189.04 16228.865 327.545 ;
      RECT 16228.025 187.94 16228.305 327.305 ;
      RECT 16227.465 189.04 16227.745 327.065 ;
      RECT 16226.905 189.04 16227.185 326.825 ;
      RECT 16226.345 189.04 16226.625 326.585 ;
      RECT 16225.785 187.94 16226.065 326.345 ;
      RECT 16225.225 189.04 16225.505 326.105 ;
      RECT 16224.665 187.94 16224.945 325.865 ;
      RECT 16224.105 189.04 16224.385 325.625 ;
      RECT 16223.545 187.94 16223.825 325.385 ;
      RECT 16222.985 189.04 16223.265 325.145 ;
      RECT 16222.425 189.04 16222.705 324.905 ;
      RECT 16182.105 189.04 16182.385 333.8 ;
      RECT 16181.545 189.04 16181.825 334.04 ;
      RECT 16180.985 189.04 16181.265 334.285 ;
      RECT 16180.425 189.04 16180.705 334.525 ;
      RECT 16179.865 189.04 16180.145 334.765 ;
      RECT 16179.305 189.04 16179.585 335.005 ;
      RECT 16178.745 189.04 16179.025 335.245 ;
      RECT 16178.185 189.04 16178.465 335.485 ;
      RECT 16177.625 189.04 16177.905 335.725 ;
      RECT 16177.065 189.04 16177.345 335.965 ;
      RECT 16176.505 187.94 16176.785 336.205 ;
      RECT 16175.945 189.04 16176.225 336.445 ;
      RECT 16175.385 187.94 16175.665 336.685 ;
      RECT 16174.825 189.04 16175.105 336.925 ;
      RECT 16174.265 187.94 16174.545 337.165 ;
      RECT 16173.705 189.04 16173.985 337.165 ;
      RECT 16173.145 189.04 16173.425 336.925 ;
      RECT 16172.585 189.04 16172.865 336.685 ;
      RECT 16172.025 189.04 16172.305 336.445 ;
      RECT 16171.465 189.04 16171.745 336.205 ;
      RECT 16170.905 189.04 16171.185 335.965 ;
      RECT 16170.345 189.04 16170.625 335.725 ;
      RECT 16169.785 189.04 16170.065 335.485 ;
      RECT 16160.825 187.94 16161.105 335.515 ;
      RECT 16160.265 189.04 16160.545 335.755 ;
      RECT 16159.705 187.94 16159.985 335.995 ;
      RECT 16159.145 189.04 16159.425 336.21 ;
      RECT 16158.585 189.04 16158.865 335.785 ;
      RECT 16158.025 189.04 16158.305 335.545 ;
      RECT 16157.465 189.04 16157.745 335.305 ;
      RECT 16156.905 189.04 16157.185 335.065 ;
      RECT 16156.345 189.04 16156.625 334.825 ;
      RECT 16155.785 189.04 16156.065 334.585 ;
      RECT 16155.225 189.04 16155.505 334.345 ;
      RECT 16154.665 189.04 16154.945 334.105 ;
      RECT 16154.105 189.04 16154.385 333.865 ;
      RECT 16153.545 189.04 16153.825 333.625 ;
      RECT 16151.025 189.04 16151.305 332.8 ;
      RECT 16150.465 189.04 16150.745 332.56 ;
      RECT 16149.905 189.04 16150.185 332.32 ;
      RECT 16149.345 187.94 16149.625 332.08 ;
      RECT 16148.785 189.04 16149.065 331.84 ;
      RECT 16148.225 187.94 16148.505 331.6 ;
      RECT 16147.665 189.04 16147.945 331.36 ;
      RECT 16147.105 189.04 16147.385 331.12 ;
      RECT 16120.505 189.04 16120.785 342.165 ;
      RECT 16119.945 187.94 16120.225 342.405 ;
      RECT 16119.385 189.04 16119.665 342.645 ;
      RECT 16118.825 187.94 16119.105 342.89 ;
      RECT 16118.265 189.04 16118.545 343.13 ;
      RECT 16117.705 187.94 16117.985 343.37 ;
      RECT 16117.145 189.04 16117.425 343.61 ;
      RECT 16116.585 189.04 16116.865 343.85 ;
      RECT 16116.025 189.04 16116.305 329.47 ;
      RECT 16115.465 189.04 16115.745 329.23 ;
      RECT 16114.905 189.04 16115.185 328.99 ;
      RECT 16114.345 189.04 16114.625 328.75 ;
      RECT 16113.785 189.04 16114.065 328.51 ;
      RECT 16113.225 189.04 16113.505 328.27 ;
      RECT 16112.665 189.04 16112.945 328.03 ;
      RECT 16112.105 189.04 16112.385 327.79 ;
      RECT 16111.545 189.04 16111.825 327.55 ;
      RECT 16110.985 189.04 16111.265 327.31 ;
      RECT 16110.425 187.94 16110.705 327.07 ;
      RECT 16109.865 189.04 16110.145 326.83 ;
      RECT 16109.305 187.94 16109.585 326.59 ;
      RECT 16108.745 189.04 16109.025 326.35 ;
      RECT 16094.745 187.94 16095.025 332.47 ;
      RECT 16094.185 189.04 16094.465 332.23 ;
      RECT 16093.625 189.04 16093.905 331.99 ;
      RECT 16093.065 189.04 16093.345 331.75 ;
      RECT 16092.505 189.04 16092.785 331.51 ;
      RECT 16091.945 189.04 16092.225 331.27 ;
      RECT 16091.385 189.04 16091.665 331.03 ;
      RECT 16090.825 189.04 16091.105 330.79 ;
      RECT 16090.265 189.04 16090.545 330.55 ;
      RECT 16089.705 187.94 16089.985 330.31 ;
      RECT 16089.145 189.04 16089.425 330.07 ;
      RECT 16088.585 187.94 16088.865 329.83 ;
      RECT 16088.025 189.04 16088.305 329.59 ;
      RECT 16087.465 189.04 16087.745 329.35 ;
      RECT 16086.905 189.04 16087.185 329.11 ;
      RECT 16086.345 189.04 16086.625 328.87 ;
      RECT 16085.785 189.04 16086.065 328.63 ;
      RECT 16085.225 189.04 16085.505 328.39 ;
      RECT 16084.665 189.04 16084.945 328.15 ;
      RECT 16084.105 189.04 16084.385 327.91 ;
      RECT 16083.545 189.04 16083.825 327.67 ;
      RECT 16082.985 189.04 16083.265 327.43 ;
      RECT 16082.425 189.04 16082.705 327.19 ;
      RECT 16043.225 189.04 16043.505 334.095 ;
      RECT 16042.665 189.04 16042.945 334.335 ;
      RECT 16042.105 189.04 16042.385 334.575 ;
      RECT 16041.545 187.94 16041.825 334.815 ;
      RECT 16040.985 189.04 16041.265 335.055 ;
      RECT 16040.425 187.94 16040.705 335.295 ;
      RECT 16039.865 189.04 16040.145 335.535 ;
      RECT 16039.305 189.04 16039.585 335.775 ;
      RECT 16038.745 189.04 16039.025 336.015 ;
      RECT 16038.185 187.94 16038.465 336.255 ;
      RECT 16037.625 189.04 16037.905 336.495 ;
      RECT 16037.065 187.94 16037.345 336.735 ;
      RECT 16036.505 189.04 16036.785 336.975 ;
      RECT 16035.945 187.94 16036.225 337.215 ;
      RECT 16035.385 189.04 16035.665 337.455 ;
      RECT 16034.825 189.04 16035.105 337.695 ;
      RECT 16034.265 189.04 16034.545 337.695 ;
      RECT 16033.705 189.04 16033.985 337.455 ;
      RECT 16033.145 189.04 16033.425 337.215 ;
      RECT 16032.585 189.04 16032.865 336.975 ;
      RECT 16032.025 189.04 16032.305 336.735 ;
      RECT 16031.465 189.04 16031.745 336.495 ;
      RECT 16030.905 189.04 16031.185 336.255 ;
      RECT 16030.345 189.04 16030.625 336.015 ;
      RECT 16029.785 189.04 16030.065 335.775 ;
      RECT 16020.825 189.04 16021.105 335.29 ;
      RECT 16020.265 187.94 16020.545 335.05 ;
      RECT 16019.705 189.04 16019.985 334.81 ;
      RECT 16019.145 187.94 16019.425 334.57 ;
      RECT 16018.585 189.04 16018.865 334.33 ;
      RECT 16018.025 187.94 16018.305 334.09 ;
      RECT 16017.465 189.04 16017.745 333.85 ;
      RECT 16016.905 189.04 16017.185 333.61 ;
      RECT 16016.345 189.04 16016.625 333.37 ;
      RECT 16015.785 189.04 16016.065 333.13 ;
      RECT 16015.225 189.04 16015.505 332.89 ;
      RECT 16014.665 189.04 16014.945 332.65 ;
      RECT 16014.105 189.04 16014.385 332.41 ;
      RECT 16013.545 189.04 16013.825 332.17 ;
      RECT 16011.025 187.94 16011.305 333.89 ;
      RECT 16010.465 189.04 16010.745 333.65 ;
      RECT 16009.905 187.94 16010.185 333.41 ;
      RECT 16009.345 189.04 16009.625 333.17 ;
      RECT 16008.785 189.04 16009.065 332.93 ;
      RECT 16008.225 189.04 16008.505 332.69 ;
      RECT 16007.665 189.04 16007.945 332.45 ;
      RECT 16007.105 189.04 16007.385 332.21 ;
      RECT 15981.065 189.04 15981.345 329.86 ;
      RECT 15980.505 189.04 15980.785 330.1 ;
      RECT 15979.945 189.04 15980.225 330.34 ;
      RECT 15979.385 189.04 15979.665 330.585 ;
      RECT 15978.825 189.04 15979.105 330.825 ;
      RECT 15978.265 189.04 15978.545 331.065 ;
      RECT 15977.705 189.04 15977.985 331.065 ;
      RECT 15977.145 189.04 15977.425 330.825 ;
      RECT 15976.585 189.04 15976.865 330.585 ;
      RECT 15976.025 187.94 15976.305 330.345 ;
      RECT 15975.465 189.04 15975.745 330.105 ;
      RECT 15974.905 187.94 15975.185 329.865 ;
      RECT 15974.345 189.04 15974.625 329.625 ;
      RECT 15973.785 189.04 15974.065 329.385 ;
      RECT 15973.225 189.04 15973.505 329.145 ;
      RECT 15972.665 187.94 15972.945 328.905 ;
      RECT 15972.105 189.04 15972.385 328.665 ;
      RECT 15971.545 187.94 15971.825 328.425 ;
      RECT 15970.985 189.04 15971.265 328.185 ;
      RECT 15970.425 187.94 15970.705 327.945 ;
      RECT 15969.865 189.04 15970.145 327.705 ;
      RECT 15969.305 189.04 15969.585 327.465 ;
      RECT 15968.745 189.04 15969.025 327.225 ;
      RECT 15968.185 189.04 15968.465 326.985 ;
      RECT 15954.745 189.04 15955.025 332.785 ;
      RECT 15954.185 189.04 15954.465 332.545 ;
      RECT 15953.625 189.04 15953.905 332.305 ;
      RECT 15953.065 189.04 15953.345 332.065 ;
      RECT 15952.505 189.04 15952.785 331.825 ;
      RECT 15951.945 189.04 15952.225 331.585 ;
      RECT 15951.385 189.04 15951.665 331.345 ;
      RECT 15950.825 189.04 15951.105 331.105 ;
      RECT 15950.265 187.94 15950.545 330.865 ;
      RECT 15949.705 189.04 15949.985 330.625 ;
      RECT 15949.145 187.94 15949.425 330.305 ;
      RECT 15948.585 189.04 15948.865 330.145 ;
      RECT 15948.025 187.94 15948.305 329.905 ;
      RECT 15947.465 189.04 15947.745 329.665 ;
      RECT 15946.905 189.04 15947.185 329.425 ;
      RECT 15946.345 189.04 15946.625 329.185 ;
      RECT 15945.785 189.04 15946.065 328.945 ;
      RECT 15945.225 189.04 15945.505 328.705 ;
      RECT 15944.665 189.04 15944.945 328.465 ;
      RECT 15944.105 189.04 15944.385 328.225 ;
      RECT 15943.545 189.04 15943.825 327.985 ;
      RECT 15942.985 187.94 15943.265 327.745 ;
      RECT 15942.425 189.04 15942.705 327.505 ;
      RECT 15941.865 187.94 15942.145 327.265 ;
      RECT 15902.665 189.04 15902.945 332.875 ;
      RECT 15902.105 189.04 15902.385 333.115 ;
      RECT 15901.545 189.04 15901.825 333.355 ;
      RECT 15900.985 189.04 15901.265 333.595 ;
      RECT 15900.425 189.04 15900.705 333.835 ;
      RECT 15899.865 189.04 15900.145 334.075 ;
      RECT 15899.305 189.04 15899.585 334.315 ;
      RECT 15898.745 189.04 15899.025 334.555 ;
      RECT 15898.185 189.04 15898.465 334.795 ;
      RECT 15897.625 189.04 15897.905 335.035 ;
      RECT 15897.065 189.04 15897.345 335.275 ;
      RECT 15896.505 189.04 15896.785 335.515 ;
      RECT 15895.945 189.04 15896.225 335.755 ;
      RECT 15895.385 189.04 15895.665 335.755 ;
      RECT 15894.825 187.94 15895.105 335.515 ;
      RECT 15894.265 189.04 15894.545 335.275 ;
      RECT 15893.705 187.94 15893.985 335.035 ;
      RECT 15893.145 189.04 15893.425 334.795 ;
      RECT 15892.585 189.04 15892.865 334.555 ;
      RECT 15892.025 189.04 15892.305 334.315 ;
      RECT 15891.465 187.94 15891.745 334.05 ;
      RECT 15890.905 189.04 15891.185 333.81 ;
      RECT 15890.345 187.94 15890.625 333.57 ;
      RECT 15889.785 189.04 15890.065 333.33 ;
      RECT 15880.825 187.94 15881.105 327.165 ;
      RECT 15880.265 189.04 15880.545 327.405 ;
      RECT 15879.705 189.04 15879.985 327.645 ;
      RECT 15879.145 189.04 15879.425 327.645 ;
      RECT 15878.585 189.04 15878.865 327.405 ;
      RECT 15878.025 189.04 15878.305 327.165 ;
      RECT 15877.465 189.04 15877.745 326.925 ;
      RECT 15876.905 189.04 15877.185 326.685 ;
      RECT 15876.345 189.04 15876.625 326.445 ;
      RECT 15875.785 189.04 15876.065 326.205 ;
      RECT 15875.225 189.04 15875.505 325.965 ;
      RECT 15874.665 189.04 15874.945 325.725 ;
      RECT 15874.105 189.04 15874.385 325.485 ;
      RECT 15873.545 187.94 15873.825 325.245 ;
      RECT 15871.025 189.04 15871.305 326.965 ;
      RECT 15870.465 187.94 15870.745 326.725 ;
      RECT 15869.905 189.04 15870.185 326.485 ;
      RECT 15869.345 187.94 15869.625 326.245 ;
      RECT 15868.785 189.04 15869.065 326.005 ;
      RECT 15868.225 189.04 15868.505 325.765 ;
      RECT 15867.665 189.04 15867.945 325.525 ;
      RECT 15841.625 189.04 15841.905 328.31 ;
      RECT 15841.065 189.04 15841.345 328.55 ;
      RECT 15840.505 189.04 15840.785 328.79 ;
      RECT 15839.945 189.04 15840.225 329.03 ;
      RECT 15839.385 189.04 15839.665 329.27 ;
      RECT 15838.825 187.94 15839.105 329.51 ;
      RECT 15838.265 189.04 15838.545 329.75 ;
      RECT 15837.705 187.94 15837.985 329.99 ;
      RECT 15837.145 189.04 15837.425 330.23 ;
      RECT 15836.585 189.04 15836.865 330.47 ;
      RECT 15836.025 189.04 15836.305 330.71 ;
      RECT 15835.465 189.04 15835.745 330.95 ;
      RECT 15834.905 189.04 15835.185 331.19 ;
      RECT 15834.345 189.04 15834.625 331.43 ;
      RECT 15833.785 189.04 15834.065 331.67 ;
      RECT 15833.225 189.04 15833.505 331.67 ;
      RECT 15832.665 189.04 15832.945 331.43 ;
      RECT 15832.105 189.04 15832.385 331.19 ;
      RECT 15831.545 189.04 15831.825 330.95 ;
      RECT 15830.985 189.04 15831.265 330.705 ;
      RECT 15830.425 189.04 15830.705 330.465 ;
      RECT 15829.865 189.04 15830.145 330.225 ;
      RECT 15829.305 187.94 15829.585 329.985 ;
      RECT 15828.745 189.04 15829.025 329.745 ;
      RECT 15815.305 187.94 15815.585 327.225 ;
      RECT 15814.745 189.04 15815.025 326.985 ;
      RECT 15814.185 189.04 15814.465 326.745 ;
      RECT 15813.625 189.04 15813.905 326.505 ;
      RECT 15813.065 187.94 15813.345 326.265 ;
      RECT 15812.505 189.04 15812.785 326.025 ;
      RECT 15811.945 187.94 15812.225 325.785 ;
      RECT 15811.385 189.04 15811.665 325.545 ;
      RECT 15810.825 187.94 15811.105 325.305 ;
      RECT 15810.265 189.04 15810.545 325.065 ;
      RECT 15809.705 189.04 15809.985 324.825 ;
      RECT 15809.145 189.04 15809.425 324.585 ;
      RECT 15808.585 189.04 15808.865 324.345 ;
      RECT 15808.025 189.04 15808.305 324.105 ;
      RECT 15807.465 189.04 15807.745 323.865 ;
      RECT 15806.905 189.04 15807.185 323.625 ;
      RECT 15806.345 189.04 15806.625 323.385 ;
      RECT 15805.785 189.04 15806.065 323.145 ;
      RECT 15805.225 189.04 15805.505 322.905 ;
      RECT 15804.665 189.04 15804.945 322.665 ;
      RECT 15804.105 189.04 15804.385 322.425 ;
      RECT 15803.545 187.94 15803.825 322.185 ;
      RECT 15802.985 189.04 15803.265 321.945 ;
      RECT 15802.425 187.94 15802.705 321.705 ;
      RECT 15762.665 189.04 15762.945 332.175 ;
      RECT 15762.105 187.94 15762.385 332.415 ;
      RECT 15761.545 189.04 15761.825 332.655 ;
      RECT 15760.985 189.04 15761.265 332.895 ;
      RECT 15760.425 189.04 15760.705 333.135 ;
      RECT 15759.865 189.04 15760.145 333.375 ;
      RECT 15759.305 189.04 15759.585 333.615 ;
      RECT 15758.745 189.04 15759.025 333.86 ;
      RECT 15758.185 189.04 15758.465 334.1 ;
      RECT 15757.625 189.04 15757.905 334.34 ;
      RECT 15757.065 187.94 15757.345 334.58 ;
      RECT 15756.505 189.04 15756.785 334.82 ;
      RECT 15755.945 187.94 15756.225 335.06 ;
      RECT 15755.385 189.04 15755.665 335.3 ;
      RECT 15754.825 189.04 15755.105 335.54 ;
      RECT 15754.265 189.04 15754.545 335.78 ;
      RECT 15753.705 189.04 15753.985 336.02 ;
      RECT 15753.145 189.04 15753.425 336.26 ;
      RECT 15752.585 189.04 15752.865 336.5 ;
      RECT 15752.025 189.04 15752.305 336.74 ;
      RECT 15751.465 189.04 15751.745 336.98 ;
      RECT 15750.905 189.04 15751.185 337.22 ;
      RECT 15750.345 189.04 15750.625 337.46 ;
      RECT 15749.785 189.04 15750.065 337.7 ;
      RECT 15740.825 189.04 15741.105 333.285 ;
      RECT 15740.265 189.04 15740.545 333.045 ;
      RECT 15739.705 189.04 15739.985 332.805 ;
      RECT 15739.145 187.94 15739.425 332.565 ;
      RECT 15738.585 189.04 15738.865 332.325 ;
      RECT 15738.025 187.94 15738.305 332.085 ;
      RECT 15737.465 189.04 15737.745 331.845 ;
      RECT 15736.905 189.04 15737.185 331.605 ;
      RECT 15736.345 189.04 15736.625 331.365 ;
      RECT 15735.785 187.94 15736.065 331.125 ;
      RECT 15735.225 189.04 15735.505 330.885 ;
      RECT 15734.665 187.94 15734.945 330.645 ;
      RECT 15734.105 189.04 15734.385 330.405 ;
      RECT 15733.545 187.94 15733.825 330.165 ;
      RECT 15731.025 189.04 15731.305 322.565 ;
      RECT 15730.465 189.04 15730.745 322.325 ;
      RECT 15729.905 189.04 15730.185 322.085 ;
      RECT 15729.345 189.04 15729.625 321.845 ;
      RECT 15728.785 189.04 15729.065 321.605 ;
      RECT 15728.225 189.04 15728.505 321.365 ;
      RECT 15727.665 189.04 15727.945 321.125 ;
      RECT 15701.625 189.04 15701.905 335 ;
      RECT 15701.065 189.04 15701.345 335.24 ;
      RECT 15700.505 189.04 15700.785 335.48 ;
      RECT 15699.945 189.04 15700.225 335.72 ;
      RECT 15699.385 189.04 15699.665 335.96 ;
      RECT 15698.825 187.94 15699.105 335.96 ;
      RECT 15698.265 189.04 15698.545 335.72 ;
      RECT 15697.705 187.94 15697.985 335.475 ;
      RECT 15697.145 189.04 15697.425 335.235 ;
      RECT 15696.585 187.94 15696.865 334.995 ;
      RECT 15696.025 189.04 15696.305 334.755 ;
      RECT 15695.465 189.04 15695.745 334.515 ;
      RECT 15694.905 189.04 15695.185 334.275 ;
      RECT 15694.345 189.04 15694.625 334.035 ;
      RECT 15693.785 189.04 15694.065 333.795 ;
      RECT 15693.225 189.04 15693.505 333.555 ;
      RECT 15692.665 189.04 15692.945 333.315 ;
      RECT 15692.105 189.04 15692.385 333.075 ;
      RECT 15691.545 187.94 15691.825 332.835 ;
      RECT 15690.985 189.04 15691.265 332.595 ;
      RECT 15690.425 187.94 15690.705 332.355 ;
      RECT 15689.865 189.04 15690.145 332.115 ;
      RECT 15689.305 189.04 15689.585 331.875 ;
      RECT 15688.745 189.04 15689.025 331.635 ;
      RECT 15675.305 189.04 15675.585 335.035 ;
      RECT 15674.745 189.04 15675.025 335.275 ;
      RECT 15674.185 189.04 15674.465 335.52 ;
      RECT 15673.625 189.04 15673.905 335.76 ;
      RECT 15673.065 189.04 15673.345 336 ;
      RECT 15672.505 189.04 15672.785 336 ;
      RECT 15671.945 189.04 15672.225 335.76 ;
      RECT 15671.385 189.04 15671.665 335.52 ;
      RECT 15670.825 189.04 15671.105 328.505 ;
      RECT 15670.265 189.04 15670.545 328.265 ;
      RECT 15669.705 189.04 15669.985 328.025 ;
      RECT 15669.145 187.94 15669.425 327.785 ;
      RECT 15668.585 189.04 15668.865 327.545 ;
      RECT 15668.025 187.94 15668.305 327.305 ;
      RECT 15667.465 189.04 15667.745 327.065 ;
      RECT 15666.905 189.04 15667.185 326.825 ;
      RECT 15666.345 189.04 15666.625 326.585 ;
      RECT 15665.785 187.94 15666.065 326.345 ;
      RECT 15665.225 189.04 15665.505 326.105 ;
      RECT 15664.665 187.94 15664.945 325.865 ;
      RECT 15664.105 189.04 15664.385 325.625 ;
      RECT 15663.545 187.94 15663.825 325.385 ;
      RECT 15662.985 189.04 15663.265 325.145 ;
      RECT 15662.425 189.04 15662.705 324.905 ;
      RECT 15622.105 189.04 15622.385 333.8 ;
      RECT 15621.545 189.04 15621.825 334.04 ;
      RECT 15620.985 189.04 15621.265 334.285 ;
      RECT 15620.425 189.04 15620.705 334.525 ;
      RECT 15619.865 189.04 15620.145 334.765 ;
      RECT 15619.305 189.04 15619.585 335.005 ;
      RECT 15618.745 189.04 15619.025 335.245 ;
      RECT 15618.185 189.04 15618.465 335.485 ;
      RECT 15617.625 189.04 15617.905 335.725 ;
      RECT 15617.065 189.04 15617.345 335.965 ;
      RECT 15616.505 187.94 15616.785 336.205 ;
      RECT 15615.945 189.04 15616.225 336.445 ;
      RECT 15615.385 187.94 15615.665 336.685 ;
      RECT 15614.825 189.04 15615.105 336.925 ;
      RECT 15614.265 187.94 15614.545 337.165 ;
      RECT 15613.705 189.04 15613.985 337.165 ;
      RECT 15613.145 189.04 15613.425 336.925 ;
      RECT 15612.585 189.04 15612.865 336.685 ;
      RECT 15612.025 189.04 15612.305 336.445 ;
      RECT 15611.465 189.04 15611.745 336.205 ;
      RECT 15610.905 189.04 15611.185 335.965 ;
      RECT 15610.345 189.04 15610.625 335.725 ;
      RECT 15609.785 189.04 15610.065 335.485 ;
      RECT 15600.825 187.94 15601.105 335.515 ;
      RECT 15600.265 189.04 15600.545 335.755 ;
      RECT 15599.705 187.94 15599.985 335.995 ;
      RECT 15599.145 189.04 15599.425 336.21 ;
      RECT 15598.585 189.04 15598.865 335.785 ;
      RECT 15598.025 189.04 15598.305 335.545 ;
      RECT 15597.465 189.04 15597.745 335.305 ;
      RECT 15596.905 189.04 15597.185 335.065 ;
      RECT 15596.345 189.04 15596.625 334.825 ;
      RECT 15595.785 189.04 15596.065 334.585 ;
      RECT 15595.225 189.04 15595.505 334.345 ;
      RECT 15594.665 189.04 15594.945 334.105 ;
      RECT 15594.105 189.04 15594.385 333.865 ;
      RECT 15593.545 189.04 15593.825 333.625 ;
      RECT 15591.025 189.04 15591.305 332.8 ;
      RECT 15590.465 189.04 15590.745 332.56 ;
      RECT 15589.905 189.04 15590.185 332.32 ;
      RECT 15589.345 187.94 15589.625 332.08 ;
      RECT 15588.785 189.04 15589.065 331.84 ;
      RECT 15588.225 187.94 15588.505 331.6 ;
      RECT 15587.665 189.04 15587.945 331.36 ;
      RECT 15587.105 189.04 15587.385 331.12 ;
      RECT 15560.505 189.04 15560.785 342.165 ;
      RECT 15559.945 187.94 15560.225 342.405 ;
      RECT 15559.385 189.04 15559.665 342.645 ;
      RECT 15558.825 187.94 15559.105 342.89 ;
      RECT 15558.265 189.04 15558.545 343.13 ;
      RECT 15557.705 187.94 15557.985 343.37 ;
      RECT 15557.145 189.04 15557.425 343.61 ;
      RECT 15556.585 189.04 15556.865 343.85 ;
      RECT 15556.025 189.04 15556.305 329.47 ;
      RECT 15555.465 189.04 15555.745 329.23 ;
      RECT 15554.905 189.04 15555.185 328.99 ;
      RECT 15554.345 189.04 15554.625 328.75 ;
      RECT 15553.785 189.04 15554.065 328.51 ;
      RECT 15553.225 189.04 15553.505 328.27 ;
      RECT 15552.665 189.04 15552.945 328.03 ;
      RECT 15552.105 189.04 15552.385 327.79 ;
      RECT 15551.545 189.04 15551.825 327.55 ;
      RECT 15550.985 189.04 15551.265 327.31 ;
      RECT 15550.425 187.94 15550.705 327.07 ;
      RECT 15549.865 189.04 15550.145 326.83 ;
      RECT 15549.305 187.94 15549.585 326.59 ;
      RECT 15548.745 189.04 15549.025 326.35 ;
      RECT 15534.745 187.94 15535.025 332.47 ;
      RECT 15534.185 189.04 15534.465 332.23 ;
      RECT 15533.625 189.04 15533.905 331.99 ;
      RECT 15533.065 189.04 15533.345 331.75 ;
      RECT 15532.505 189.04 15532.785 331.51 ;
      RECT 15531.945 189.04 15532.225 331.27 ;
      RECT 15531.385 189.04 15531.665 331.03 ;
      RECT 15530.825 189.04 15531.105 330.79 ;
      RECT 15530.265 189.04 15530.545 330.55 ;
      RECT 15529.705 187.94 15529.985 330.31 ;
      RECT 15529.145 189.04 15529.425 330.07 ;
      RECT 15528.585 187.94 15528.865 329.83 ;
      RECT 15528.025 189.04 15528.305 329.59 ;
      RECT 15527.465 189.04 15527.745 329.35 ;
      RECT 15526.905 189.04 15527.185 329.11 ;
      RECT 15526.345 189.04 15526.625 328.87 ;
      RECT 15525.785 189.04 15526.065 328.63 ;
      RECT 15525.225 189.04 15525.505 328.39 ;
      RECT 15524.665 189.04 15524.945 328.15 ;
      RECT 15524.105 189.04 15524.385 327.91 ;
      RECT 15523.545 189.04 15523.825 327.67 ;
      RECT 15522.985 189.04 15523.265 327.43 ;
      RECT 15522.425 189.04 15522.705 327.19 ;
      RECT 15483.225 189.04 15483.505 334.095 ;
      RECT 15482.665 189.04 15482.945 334.335 ;
      RECT 15482.105 189.04 15482.385 334.575 ;
      RECT 15481.545 187.94 15481.825 334.815 ;
      RECT 15480.985 189.04 15481.265 335.055 ;
      RECT 15480.425 187.94 15480.705 335.295 ;
      RECT 15479.865 189.04 15480.145 335.535 ;
      RECT 15479.305 189.04 15479.585 335.775 ;
      RECT 15478.745 189.04 15479.025 336.015 ;
      RECT 15478.185 187.94 15478.465 336.255 ;
      RECT 15477.625 189.04 15477.905 336.495 ;
      RECT 15477.065 187.94 15477.345 336.735 ;
      RECT 15476.505 189.04 15476.785 336.975 ;
      RECT 15475.945 187.94 15476.225 337.215 ;
      RECT 15475.385 189.04 15475.665 337.455 ;
      RECT 15474.825 189.04 15475.105 337.695 ;
      RECT 15474.265 189.04 15474.545 337.695 ;
      RECT 15473.705 189.04 15473.985 337.455 ;
      RECT 15473.145 189.04 15473.425 337.215 ;
      RECT 15472.585 189.04 15472.865 336.975 ;
      RECT 15472.025 189.04 15472.305 336.735 ;
      RECT 15471.465 189.04 15471.745 336.495 ;
      RECT 15470.905 189.04 15471.185 336.255 ;
      RECT 15470.345 189.04 15470.625 336.015 ;
      RECT 15469.785 189.04 15470.065 335.775 ;
      RECT 15460.825 189.04 15461.105 335.29 ;
      RECT 15460.265 187.94 15460.545 335.05 ;
      RECT 15459.705 189.04 15459.985 334.81 ;
      RECT 15459.145 187.94 15459.425 334.57 ;
      RECT 15458.585 189.04 15458.865 334.33 ;
      RECT 15458.025 187.94 15458.305 334.09 ;
      RECT 15457.465 189.04 15457.745 333.85 ;
      RECT 15456.905 189.04 15457.185 333.61 ;
      RECT 15456.345 189.04 15456.625 333.37 ;
      RECT 15455.785 189.04 15456.065 333.13 ;
      RECT 15455.225 189.04 15455.505 332.89 ;
      RECT 15454.665 189.04 15454.945 332.65 ;
      RECT 15454.105 189.04 15454.385 332.41 ;
      RECT 15453.545 189.04 15453.825 332.17 ;
      RECT 15451.025 187.94 15451.305 333.89 ;
      RECT 15450.465 189.04 15450.745 333.65 ;
      RECT 15449.905 187.94 15450.185 333.41 ;
      RECT 15449.345 189.04 15449.625 333.17 ;
      RECT 15448.785 189.04 15449.065 332.93 ;
      RECT 15448.225 189.04 15448.505 332.69 ;
      RECT 15447.665 189.04 15447.945 332.45 ;
      RECT 15447.105 189.04 15447.385 332.21 ;
      RECT 15421.065 189.04 15421.345 329.86 ;
      RECT 15420.505 189.04 15420.785 330.1 ;
      RECT 15419.945 189.04 15420.225 330.34 ;
      RECT 15419.385 189.04 15419.665 330.585 ;
      RECT 15418.825 189.04 15419.105 330.825 ;
      RECT 15418.265 189.04 15418.545 331.065 ;
      RECT 15417.705 189.04 15417.985 331.065 ;
      RECT 15417.145 189.04 15417.425 330.825 ;
      RECT 15416.585 189.04 15416.865 330.585 ;
      RECT 15416.025 187.94 15416.305 330.345 ;
      RECT 15415.465 189.04 15415.745 330.105 ;
      RECT 15414.905 187.94 15415.185 329.865 ;
      RECT 15414.345 189.04 15414.625 329.625 ;
      RECT 15413.785 189.04 15414.065 329.385 ;
      RECT 15413.225 189.04 15413.505 329.145 ;
      RECT 15412.665 187.94 15412.945 328.905 ;
      RECT 15412.105 189.04 15412.385 328.665 ;
      RECT 15411.545 187.94 15411.825 328.425 ;
      RECT 15410.985 189.04 15411.265 328.185 ;
      RECT 15410.425 187.94 15410.705 327.945 ;
      RECT 15409.865 189.04 15410.145 327.705 ;
      RECT 15409.305 189.04 15409.585 327.465 ;
      RECT 15408.745 189.04 15409.025 327.225 ;
      RECT 15408.185 189.04 15408.465 326.985 ;
      RECT 15394.745 189.04 15395.025 332.785 ;
      RECT 15394.185 189.04 15394.465 332.545 ;
      RECT 15393.625 189.04 15393.905 332.305 ;
      RECT 15393.065 189.04 15393.345 332.065 ;
      RECT 15392.505 189.04 15392.785 331.825 ;
      RECT 15391.945 189.04 15392.225 331.585 ;
      RECT 15391.385 189.04 15391.665 331.345 ;
      RECT 15390.825 189.04 15391.105 331.105 ;
      RECT 15390.265 187.94 15390.545 330.865 ;
      RECT 15389.705 189.04 15389.985 330.625 ;
      RECT 15389.145 187.94 15389.425 330.305 ;
      RECT 15388.585 189.04 15388.865 330.145 ;
      RECT 15388.025 187.94 15388.305 329.905 ;
      RECT 15387.465 189.04 15387.745 329.665 ;
      RECT 15386.905 189.04 15387.185 329.425 ;
      RECT 15386.345 189.04 15386.625 329.185 ;
      RECT 15385.785 189.04 15386.065 328.945 ;
      RECT 15385.225 189.04 15385.505 328.705 ;
      RECT 15384.665 189.04 15384.945 328.465 ;
      RECT 15384.105 189.04 15384.385 328.225 ;
      RECT 15383.545 189.04 15383.825 327.985 ;
      RECT 15382.985 187.94 15383.265 327.745 ;
      RECT 15382.425 189.04 15382.705 327.505 ;
      RECT 15381.865 187.94 15382.145 327.265 ;
      RECT 15342.665 189.04 15342.945 332.875 ;
      RECT 15342.105 189.04 15342.385 333.115 ;
      RECT 15341.545 189.04 15341.825 333.355 ;
      RECT 15340.985 189.04 15341.265 333.595 ;
      RECT 15340.425 189.04 15340.705 333.835 ;
      RECT 15339.865 189.04 15340.145 334.075 ;
      RECT 15339.305 189.04 15339.585 334.315 ;
      RECT 15338.745 189.04 15339.025 334.555 ;
      RECT 15338.185 189.04 15338.465 334.795 ;
      RECT 15337.625 189.04 15337.905 335.035 ;
      RECT 15337.065 189.04 15337.345 335.275 ;
      RECT 15336.505 189.04 15336.785 335.515 ;
      RECT 15335.945 189.04 15336.225 335.755 ;
      RECT 15335.385 189.04 15335.665 335.755 ;
      RECT 15334.825 187.94 15335.105 335.515 ;
      RECT 15334.265 189.04 15334.545 335.275 ;
      RECT 15333.705 187.94 15333.985 335.035 ;
      RECT 15333.145 189.04 15333.425 334.795 ;
      RECT 15332.585 189.04 15332.865 334.555 ;
      RECT 15332.025 189.04 15332.305 334.315 ;
      RECT 15331.465 187.94 15331.745 334.05 ;
      RECT 15330.905 189.04 15331.185 333.81 ;
      RECT 15330.345 187.94 15330.625 333.57 ;
      RECT 15329.785 189.04 15330.065 333.33 ;
      RECT 15320.825 187.94 15321.105 327.165 ;
      RECT 15320.265 189.04 15320.545 327.405 ;
      RECT 15319.705 189.04 15319.985 327.645 ;
      RECT 15319.145 189.04 15319.425 327.645 ;
      RECT 15318.585 189.04 15318.865 327.405 ;
      RECT 15318.025 189.04 15318.305 327.165 ;
      RECT 15317.465 189.04 15317.745 326.925 ;
      RECT 15316.905 189.04 15317.185 326.685 ;
      RECT 15316.345 189.04 15316.625 326.445 ;
      RECT 15315.785 189.04 15316.065 326.205 ;
      RECT 15315.225 189.04 15315.505 325.965 ;
      RECT 15314.665 189.04 15314.945 325.725 ;
      RECT 15314.105 189.04 15314.385 325.485 ;
      RECT 15313.545 187.94 15313.825 325.245 ;
      RECT 15311.025 189.04 15311.305 326.965 ;
      RECT 15310.465 187.94 15310.745 326.725 ;
      RECT 15309.905 189.04 15310.185 326.485 ;
      RECT 15309.345 187.94 15309.625 326.245 ;
      RECT 15308.785 189.04 15309.065 326.005 ;
      RECT 15308.225 189.04 15308.505 325.765 ;
      RECT 15307.665 189.04 15307.945 325.525 ;
      RECT 15281.625 189.04 15281.905 328.31 ;
      RECT 15281.065 189.04 15281.345 328.55 ;
      RECT 15280.505 189.04 15280.785 328.79 ;
      RECT 15279.945 189.04 15280.225 329.03 ;
      RECT 15279.385 189.04 15279.665 329.27 ;
      RECT 15278.825 187.94 15279.105 329.51 ;
      RECT 15278.265 189.04 15278.545 329.75 ;
      RECT 15277.705 187.94 15277.985 329.99 ;
      RECT 15277.145 189.04 15277.425 330.23 ;
      RECT 15276.585 189.04 15276.865 330.47 ;
      RECT 15276.025 189.04 15276.305 330.71 ;
      RECT 15275.465 189.04 15275.745 330.95 ;
      RECT 15274.905 189.04 15275.185 331.19 ;
      RECT 15274.345 189.04 15274.625 331.43 ;
      RECT 15273.785 189.04 15274.065 331.67 ;
      RECT 15273.225 189.04 15273.505 331.67 ;
      RECT 15272.665 189.04 15272.945 331.43 ;
      RECT 15272.105 189.04 15272.385 331.19 ;
      RECT 15271.545 189.04 15271.825 330.95 ;
      RECT 15270.985 189.04 15271.265 330.705 ;
      RECT 15270.425 189.04 15270.705 330.465 ;
      RECT 15269.865 189.04 15270.145 330.225 ;
      RECT 15269.305 187.94 15269.585 329.985 ;
      RECT 15268.745 189.04 15269.025 329.745 ;
      RECT 15255.305 187.94 15255.585 327.225 ;
      RECT 15254.745 189.04 15255.025 326.985 ;
      RECT 15254.185 189.04 15254.465 326.745 ;
      RECT 15253.625 189.04 15253.905 326.505 ;
      RECT 15253.065 187.94 15253.345 326.265 ;
      RECT 15252.505 189.04 15252.785 326.025 ;
      RECT 15251.945 187.94 15252.225 325.785 ;
      RECT 15251.385 189.04 15251.665 325.545 ;
      RECT 15250.825 187.94 15251.105 325.305 ;
      RECT 15250.265 189.04 15250.545 325.065 ;
      RECT 15249.705 189.04 15249.985 324.825 ;
      RECT 15249.145 189.04 15249.425 324.585 ;
      RECT 15248.585 189.04 15248.865 324.345 ;
      RECT 15248.025 189.04 15248.305 324.105 ;
      RECT 15247.465 189.04 15247.745 323.865 ;
      RECT 15246.905 189.04 15247.185 323.625 ;
      RECT 15246.345 189.04 15246.625 323.385 ;
      RECT 15245.785 189.04 15246.065 323.145 ;
      RECT 15245.225 189.04 15245.505 322.905 ;
      RECT 15244.665 189.04 15244.945 322.665 ;
      RECT 15244.105 189.04 15244.385 322.425 ;
      RECT 15243.545 187.94 15243.825 322.185 ;
      RECT 15242.985 189.04 15243.265 321.945 ;
      RECT 15242.425 187.94 15242.705 321.705 ;
      RECT 15202.665 189.04 15202.945 332.175 ;
      RECT 15202.105 187.94 15202.385 332.415 ;
      RECT 15201.545 189.04 15201.825 332.655 ;
      RECT 15200.985 189.04 15201.265 332.895 ;
      RECT 15200.425 189.04 15200.705 333.135 ;
      RECT 15199.865 189.04 15200.145 333.375 ;
      RECT 15199.305 189.04 15199.585 333.615 ;
      RECT 15198.745 189.04 15199.025 333.86 ;
      RECT 15198.185 189.04 15198.465 334.1 ;
      RECT 15197.625 189.04 15197.905 334.34 ;
      RECT 15197.065 187.94 15197.345 334.58 ;
      RECT 15196.505 189.04 15196.785 334.82 ;
      RECT 15195.945 187.94 15196.225 335.06 ;
      RECT 15195.385 189.04 15195.665 335.3 ;
      RECT 15194.825 189.04 15195.105 335.54 ;
      RECT 15194.265 189.04 15194.545 335.78 ;
      RECT 15193.705 189.04 15193.985 336.02 ;
      RECT 15193.145 189.04 15193.425 336.26 ;
      RECT 15192.585 189.04 15192.865 336.5 ;
      RECT 15192.025 189.04 15192.305 336.74 ;
      RECT 15191.465 189.04 15191.745 336.98 ;
      RECT 15190.905 189.04 15191.185 337.22 ;
      RECT 15190.345 189.04 15190.625 337.46 ;
      RECT 15189.785 189.04 15190.065 337.7 ;
      RECT 15180.825 189.04 15181.105 333.285 ;
      RECT 15180.265 189.04 15180.545 333.045 ;
      RECT 15179.705 189.04 15179.985 332.805 ;
      RECT 15179.145 187.94 15179.425 332.565 ;
      RECT 15178.585 189.04 15178.865 332.325 ;
      RECT 15178.025 187.94 15178.305 332.085 ;
      RECT 15177.465 189.04 15177.745 331.845 ;
      RECT 15176.905 189.04 15177.185 331.605 ;
      RECT 15176.345 189.04 15176.625 331.365 ;
      RECT 15175.785 187.94 15176.065 331.125 ;
      RECT 15175.225 189.04 15175.505 330.885 ;
      RECT 15174.665 187.94 15174.945 330.645 ;
      RECT 15174.105 189.04 15174.385 330.405 ;
      RECT 15173.545 187.94 15173.825 330.165 ;
      RECT 15171.025 189.04 15171.305 322.565 ;
      RECT 15170.465 189.04 15170.745 322.325 ;
      RECT 15169.905 189.04 15170.185 322.085 ;
      RECT 15169.345 189.04 15169.625 321.845 ;
      RECT 15168.785 189.04 15169.065 321.605 ;
      RECT 15168.225 189.04 15168.505 321.365 ;
      RECT 15167.665 189.04 15167.945 321.125 ;
      RECT 15141.625 189.04 15141.905 335 ;
      RECT 15141.065 189.04 15141.345 335.24 ;
      RECT 15140.505 189.04 15140.785 335.48 ;
      RECT 15139.945 189.04 15140.225 335.72 ;
      RECT 15139.385 189.04 15139.665 335.96 ;
      RECT 15138.825 187.94 15139.105 335.96 ;
      RECT 15138.265 189.04 15138.545 335.72 ;
      RECT 15137.705 187.94 15137.985 335.475 ;
      RECT 15137.145 189.04 15137.425 335.235 ;
      RECT 15136.585 187.94 15136.865 334.995 ;
      RECT 15136.025 189.04 15136.305 334.755 ;
      RECT 15135.465 189.04 15135.745 334.515 ;
      RECT 15134.905 189.04 15135.185 334.275 ;
      RECT 15134.345 189.04 15134.625 334.035 ;
      RECT 15133.785 189.04 15134.065 333.795 ;
      RECT 15133.225 189.04 15133.505 333.555 ;
      RECT 15132.665 189.04 15132.945 333.315 ;
      RECT 15132.105 189.04 15132.385 333.075 ;
      RECT 15131.545 187.94 15131.825 332.835 ;
      RECT 15130.985 189.04 15131.265 332.595 ;
      RECT 15130.425 187.94 15130.705 332.355 ;
      RECT 15129.865 189.04 15130.145 332.115 ;
      RECT 15129.305 189.04 15129.585 331.875 ;
      RECT 15128.745 189.04 15129.025 331.635 ;
      RECT 15115.305 189.04 15115.585 335.035 ;
      RECT 15114.745 189.04 15115.025 335.275 ;
      RECT 15114.185 189.04 15114.465 335.52 ;
      RECT 15113.625 189.04 15113.905 335.76 ;
      RECT 15113.065 189.04 15113.345 336 ;
      RECT 15112.505 189.04 15112.785 336 ;
      RECT 15111.945 189.04 15112.225 335.76 ;
      RECT 15111.385 189.04 15111.665 335.52 ;
      RECT 15110.825 189.04 15111.105 328.505 ;
      RECT 15110.265 189.04 15110.545 328.265 ;
      RECT 15109.705 189.04 15109.985 328.025 ;
      RECT 15109.145 187.94 15109.425 327.785 ;
      RECT 15108.585 189.04 15108.865 327.545 ;
      RECT 15108.025 187.94 15108.305 327.305 ;
      RECT 15107.465 189.04 15107.745 327.065 ;
      RECT 15106.905 189.04 15107.185 326.825 ;
      RECT 15106.345 189.04 15106.625 326.585 ;
      RECT 15105.785 187.94 15106.065 326.345 ;
      RECT 15105.225 189.04 15105.505 326.105 ;
      RECT 15104.665 187.94 15104.945 325.865 ;
      RECT 15104.105 189.04 15104.385 325.625 ;
      RECT 15103.545 187.94 15103.825 325.385 ;
      RECT 15102.985 189.04 15103.265 325.145 ;
      RECT 15102.425 189.04 15102.705 324.905 ;
      RECT 15062.105 189.04 15062.385 333.8 ;
      RECT 15061.545 189.04 15061.825 334.04 ;
      RECT 15060.985 189.04 15061.265 334.285 ;
      RECT 15060.425 189.04 15060.705 334.525 ;
      RECT 15059.865 189.04 15060.145 334.765 ;
      RECT 15059.305 189.04 15059.585 335.005 ;
      RECT 15058.745 189.04 15059.025 335.245 ;
      RECT 15058.185 189.04 15058.465 335.485 ;
      RECT 15057.625 189.04 15057.905 335.725 ;
      RECT 15057.065 189.04 15057.345 335.965 ;
      RECT 15056.505 187.94 15056.785 336.205 ;
      RECT 15055.945 189.04 15056.225 336.445 ;
      RECT 15055.385 187.94 15055.665 336.685 ;
      RECT 15054.825 189.04 15055.105 336.925 ;
      RECT 15054.265 187.94 15054.545 337.165 ;
      RECT 15053.705 189.04 15053.985 337.165 ;
      RECT 15053.145 189.04 15053.425 336.925 ;
      RECT 15052.585 189.04 15052.865 336.685 ;
      RECT 15052.025 189.04 15052.305 336.445 ;
      RECT 15051.465 189.04 15051.745 336.205 ;
      RECT 15050.905 189.04 15051.185 335.965 ;
      RECT 15050.345 189.04 15050.625 335.725 ;
      RECT 15049.785 189.04 15050.065 335.485 ;
      RECT 15040.825 187.94 15041.105 335.515 ;
      RECT 15040.265 189.04 15040.545 335.755 ;
      RECT 15039.705 187.94 15039.985 335.995 ;
      RECT 15039.145 189.04 15039.425 336.21 ;
      RECT 15038.585 189.04 15038.865 335.785 ;
      RECT 15038.025 189.04 15038.305 335.545 ;
      RECT 15037.465 189.04 15037.745 335.305 ;
      RECT 15036.905 189.04 15037.185 335.065 ;
      RECT 15036.345 189.04 15036.625 334.825 ;
      RECT 15035.785 189.04 15036.065 334.585 ;
      RECT 15035.225 189.04 15035.505 334.345 ;
      RECT 15034.665 189.04 15034.945 334.105 ;
      RECT 15034.105 189.04 15034.385 333.865 ;
      RECT 15033.545 189.04 15033.825 333.625 ;
      RECT 15031.025 189.04 15031.305 332.8 ;
      RECT 15030.465 189.04 15030.745 332.56 ;
      RECT 15029.905 189.04 15030.185 332.32 ;
      RECT 15029.345 187.94 15029.625 332.08 ;
      RECT 15028.785 189.04 15029.065 331.84 ;
      RECT 15028.225 187.94 15028.505 331.6 ;
      RECT 15027.665 189.04 15027.945 331.36 ;
      RECT 15027.105 189.04 15027.385 331.12 ;
      RECT 15000.505 189.04 15000.785 342.165 ;
      RECT 14999.945 187.94 15000.225 342.405 ;
      RECT 14999.385 189.04 14999.665 342.645 ;
      RECT 14998.825 187.94 14999.105 342.89 ;
      RECT 14998.265 189.04 14998.545 343.13 ;
      RECT 14997.705 187.94 14997.985 343.37 ;
      RECT 14997.145 189.04 14997.425 343.61 ;
      RECT 14996.585 189.04 14996.865 343.85 ;
      RECT 14996.025 189.04 14996.305 329.47 ;
      RECT 14995.465 189.04 14995.745 329.23 ;
      RECT 14994.905 189.04 14995.185 328.99 ;
      RECT 14994.345 189.04 14994.625 328.75 ;
      RECT 14993.785 189.04 14994.065 328.51 ;
      RECT 14993.225 189.04 14993.505 328.27 ;
      RECT 14992.665 189.04 14992.945 328.03 ;
      RECT 14992.105 189.04 14992.385 327.79 ;
      RECT 14991.545 189.04 14991.825 327.55 ;
      RECT 14990.985 189.04 14991.265 327.31 ;
      RECT 14990.425 187.94 14990.705 327.07 ;
      RECT 14989.865 189.04 14990.145 326.83 ;
      RECT 14989.305 187.94 14989.585 326.59 ;
      RECT 14988.745 189.04 14989.025 326.35 ;
      RECT 14974.745 187.94 14975.025 332.47 ;
      RECT 14974.185 189.04 14974.465 332.23 ;
      RECT 14973.625 189.04 14973.905 331.99 ;
      RECT 14973.065 189.04 14973.345 331.75 ;
      RECT 14972.505 189.04 14972.785 331.51 ;
      RECT 14971.945 189.04 14972.225 331.27 ;
      RECT 14971.385 189.04 14971.665 331.03 ;
      RECT 14970.825 189.04 14971.105 330.79 ;
      RECT 14970.265 189.04 14970.545 330.55 ;
      RECT 14969.705 187.94 14969.985 330.31 ;
      RECT 14969.145 189.04 14969.425 330.07 ;
      RECT 14968.585 187.94 14968.865 329.83 ;
      RECT 14968.025 189.04 14968.305 329.59 ;
      RECT 14967.465 189.04 14967.745 329.35 ;
      RECT 14966.905 189.04 14967.185 329.11 ;
      RECT 14966.345 189.04 14966.625 328.87 ;
      RECT 14965.785 189.04 14966.065 328.63 ;
      RECT 14965.225 189.04 14965.505 328.39 ;
      RECT 14964.665 189.04 14964.945 328.15 ;
      RECT 14964.105 189.04 14964.385 327.91 ;
      RECT 14963.545 189.04 14963.825 327.67 ;
      RECT 14962.985 189.04 14963.265 327.43 ;
      RECT 14962.425 189.04 14962.705 327.19 ;
      RECT 14923.225 189.04 14923.505 334.095 ;
      RECT 14922.665 189.04 14922.945 334.335 ;
      RECT 14922.105 189.04 14922.385 334.575 ;
      RECT 14921.545 187.94 14921.825 334.815 ;
      RECT 14920.985 189.04 14921.265 335.055 ;
      RECT 14920.425 187.94 14920.705 335.295 ;
      RECT 14919.865 189.04 14920.145 335.535 ;
      RECT 14919.305 189.04 14919.585 335.775 ;
      RECT 14918.745 189.04 14919.025 336.015 ;
      RECT 14918.185 187.94 14918.465 336.255 ;
      RECT 14917.625 189.04 14917.905 336.495 ;
      RECT 14917.065 187.94 14917.345 336.735 ;
      RECT 14916.505 189.04 14916.785 336.975 ;
      RECT 14915.945 187.94 14916.225 337.215 ;
      RECT 14915.385 189.04 14915.665 337.455 ;
      RECT 14914.825 189.04 14915.105 337.695 ;
      RECT 14914.265 189.04 14914.545 337.695 ;
      RECT 14913.705 189.04 14913.985 337.455 ;
      RECT 14913.145 189.04 14913.425 337.215 ;
      RECT 14912.585 189.04 14912.865 336.975 ;
      RECT 14912.025 189.04 14912.305 336.735 ;
      RECT 14911.465 189.04 14911.745 336.495 ;
      RECT 14910.905 189.04 14911.185 336.255 ;
      RECT 14910.345 189.04 14910.625 336.015 ;
      RECT 14909.785 189.04 14910.065 335.775 ;
      RECT 14900.825 189.04 14901.105 335.29 ;
      RECT 14900.265 187.94 14900.545 335.05 ;
      RECT 14899.705 189.04 14899.985 334.81 ;
      RECT 14899.145 187.94 14899.425 334.57 ;
      RECT 14898.585 189.04 14898.865 334.33 ;
      RECT 14898.025 187.94 14898.305 334.09 ;
      RECT 14897.465 189.04 14897.745 333.85 ;
      RECT 14896.905 189.04 14897.185 333.61 ;
      RECT 14896.345 189.04 14896.625 333.37 ;
      RECT 14895.785 189.04 14896.065 333.13 ;
      RECT 14895.225 189.04 14895.505 332.89 ;
      RECT 14894.665 189.04 14894.945 332.65 ;
      RECT 14894.105 189.04 14894.385 332.41 ;
      RECT 14893.545 189.04 14893.825 332.17 ;
      RECT 14891.025 187.94 14891.305 333.89 ;
      RECT 14890.465 189.04 14890.745 333.65 ;
      RECT 14889.905 187.94 14890.185 333.41 ;
      RECT 14889.345 189.04 14889.625 333.17 ;
      RECT 14888.785 189.04 14889.065 332.93 ;
      RECT 14888.225 189.04 14888.505 332.69 ;
      RECT 14887.665 189.04 14887.945 332.45 ;
      RECT 14887.105 189.04 14887.385 332.21 ;
      RECT 14861.065 189.04 14861.345 329.86 ;
      RECT 14860.505 189.04 14860.785 330.1 ;
      RECT 14859.945 189.04 14860.225 330.34 ;
      RECT 14859.385 189.04 14859.665 330.585 ;
      RECT 14858.825 189.04 14859.105 330.825 ;
      RECT 14858.265 189.04 14858.545 331.065 ;
      RECT 14857.705 189.04 14857.985 331.065 ;
      RECT 14857.145 189.04 14857.425 330.825 ;
      RECT 14856.585 189.04 14856.865 330.585 ;
      RECT 14856.025 187.94 14856.305 330.345 ;
      RECT 14855.465 189.04 14855.745 330.105 ;
      RECT 14854.905 187.94 14855.185 329.865 ;
      RECT 14854.345 189.04 14854.625 329.625 ;
      RECT 14853.785 189.04 14854.065 329.385 ;
      RECT 14853.225 189.04 14853.505 329.145 ;
      RECT 14852.665 187.94 14852.945 328.905 ;
      RECT 14852.105 189.04 14852.385 328.665 ;
      RECT 14851.545 187.94 14851.825 328.425 ;
      RECT 14850.985 189.04 14851.265 328.185 ;
      RECT 14850.425 187.94 14850.705 327.945 ;
      RECT 14849.865 189.04 14850.145 327.705 ;
      RECT 14849.305 189.04 14849.585 327.465 ;
      RECT 14848.745 189.04 14849.025 327.225 ;
      RECT 14848.185 189.04 14848.465 326.985 ;
      RECT 14834.745 189.04 14835.025 332.785 ;
      RECT 14834.185 189.04 14834.465 332.545 ;
      RECT 14833.625 189.04 14833.905 332.305 ;
      RECT 14833.065 189.04 14833.345 332.065 ;
      RECT 14832.505 189.04 14832.785 331.825 ;
      RECT 14831.945 189.04 14832.225 331.585 ;
      RECT 14831.385 189.04 14831.665 331.345 ;
      RECT 14830.825 189.04 14831.105 331.105 ;
      RECT 14830.265 187.94 14830.545 330.865 ;
      RECT 14829.705 189.04 14829.985 330.625 ;
      RECT 14829.145 187.94 14829.425 330.305 ;
      RECT 14828.585 189.04 14828.865 330.145 ;
      RECT 14828.025 187.94 14828.305 329.905 ;
      RECT 14827.465 189.04 14827.745 329.665 ;
      RECT 14826.905 189.04 14827.185 329.425 ;
      RECT 14826.345 189.04 14826.625 329.185 ;
      RECT 14825.785 189.04 14826.065 328.945 ;
      RECT 14825.225 189.04 14825.505 328.705 ;
      RECT 14824.665 189.04 14824.945 328.465 ;
      RECT 14824.105 189.04 14824.385 328.225 ;
      RECT 14823.545 189.04 14823.825 327.985 ;
      RECT 14822.985 187.94 14823.265 327.745 ;
      RECT 14822.425 189.04 14822.705 327.505 ;
      RECT 14821.865 187.94 14822.145 327.265 ;
      RECT 14782.665 189.04 14782.945 332.875 ;
      RECT 14782.105 189.04 14782.385 333.115 ;
      RECT 14781.545 189.04 14781.825 333.355 ;
      RECT 14780.985 189.04 14781.265 333.595 ;
      RECT 14780.425 189.04 14780.705 333.835 ;
      RECT 14779.865 189.04 14780.145 334.075 ;
      RECT 14779.305 189.04 14779.585 334.315 ;
      RECT 14778.745 189.04 14779.025 334.555 ;
      RECT 14778.185 189.04 14778.465 334.795 ;
      RECT 14777.625 189.04 14777.905 335.035 ;
      RECT 14777.065 189.04 14777.345 335.275 ;
      RECT 14776.505 189.04 14776.785 335.515 ;
      RECT 14775.945 189.04 14776.225 335.755 ;
      RECT 14775.385 189.04 14775.665 335.755 ;
      RECT 14774.825 187.94 14775.105 335.515 ;
      RECT 14774.265 189.04 14774.545 335.275 ;
      RECT 14773.705 187.94 14773.985 335.035 ;
      RECT 14773.145 189.04 14773.425 334.795 ;
      RECT 14772.585 189.04 14772.865 334.555 ;
      RECT 14772.025 189.04 14772.305 334.315 ;
      RECT 14771.465 187.94 14771.745 334.05 ;
      RECT 14770.905 189.04 14771.185 333.81 ;
      RECT 14770.345 187.94 14770.625 333.57 ;
      RECT 14769.785 189.04 14770.065 333.33 ;
      RECT 14760.825 187.94 14761.105 327.165 ;
      RECT 14760.265 189.04 14760.545 327.405 ;
      RECT 14759.705 189.04 14759.985 327.645 ;
      RECT 14759.145 189.04 14759.425 327.645 ;
      RECT 14758.585 189.04 14758.865 327.405 ;
      RECT 14758.025 189.04 14758.305 327.165 ;
      RECT 14757.465 189.04 14757.745 326.925 ;
      RECT 14756.905 189.04 14757.185 326.685 ;
      RECT 14756.345 189.04 14756.625 326.445 ;
      RECT 14755.785 189.04 14756.065 326.205 ;
      RECT 14755.225 189.04 14755.505 325.965 ;
      RECT 14754.665 189.04 14754.945 325.725 ;
      RECT 14754.105 189.04 14754.385 325.485 ;
      RECT 14753.545 187.94 14753.825 325.245 ;
      RECT 14751.025 189.04 14751.305 326.965 ;
      RECT 14750.465 187.94 14750.745 326.725 ;
      RECT 14749.905 189.04 14750.185 326.485 ;
      RECT 14749.345 187.94 14749.625 326.245 ;
      RECT 14748.785 189.04 14749.065 326.005 ;
      RECT 14748.225 189.04 14748.505 325.765 ;
      RECT 14747.665 189.04 14747.945 325.525 ;
      RECT 14721.625 189.04 14721.905 328.31 ;
      RECT 14721.065 189.04 14721.345 328.55 ;
      RECT 14720.505 189.04 14720.785 328.79 ;
      RECT 14719.945 189.04 14720.225 329.03 ;
      RECT 14719.385 189.04 14719.665 329.27 ;
      RECT 14718.825 187.94 14719.105 329.51 ;
      RECT 14718.265 189.04 14718.545 329.75 ;
      RECT 14717.705 187.94 14717.985 329.99 ;
      RECT 14717.145 189.04 14717.425 330.23 ;
      RECT 14716.585 189.04 14716.865 330.47 ;
      RECT 14716.025 189.04 14716.305 330.71 ;
      RECT 14715.465 189.04 14715.745 330.95 ;
      RECT 14714.905 189.04 14715.185 331.19 ;
      RECT 14714.345 189.04 14714.625 331.43 ;
      RECT 14713.785 189.04 14714.065 331.67 ;
      RECT 14713.225 189.04 14713.505 331.67 ;
      RECT 14712.665 189.04 14712.945 331.43 ;
      RECT 14712.105 189.04 14712.385 331.19 ;
      RECT 14711.545 189.04 14711.825 330.95 ;
      RECT 14710.985 189.04 14711.265 330.705 ;
      RECT 14710.425 189.04 14710.705 330.465 ;
      RECT 14709.865 189.04 14710.145 330.225 ;
      RECT 14709.305 187.94 14709.585 329.985 ;
      RECT 14708.745 189.04 14709.025 329.745 ;
      RECT 14695.305 187.94 14695.585 327.225 ;
      RECT 14694.745 189.04 14695.025 326.985 ;
      RECT 14694.185 189.04 14694.465 326.745 ;
      RECT 14693.625 189.04 14693.905 326.505 ;
      RECT 14693.065 187.94 14693.345 326.265 ;
      RECT 14692.505 189.04 14692.785 326.025 ;
      RECT 14691.945 187.94 14692.225 325.785 ;
      RECT 14691.385 189.04 14691.665 325.545 ;
      RECT 14690.825 187.94 14691.105 325.305 ;
      RECT 14690.265 189.04 14690.545 325.065 ;
      RECT 14689.705 189.04 14689.985 324.825 ;
      RECT 14689.145 189.04 14689.425 324.585 ;
      RECT 14688.585 189.04 14688.865 324.345 ;
      RECT 14688.025 189.04 14688.305 324.105 ;
      RECT 14687.465 189.04 14687.745 323.865 ;
      RECT 14686.905 189.04 14687.185 323.625 ;
      RECT 14686.345 189.04 14686.625 323.385 ;
      RECT 14685.785 189.04 14686.065 323.145 ;
      RECT 14685.225 189.04 14685.505 322.905 ;
      RECT 14684.665 189.04 14684.945 322.665 ;
      RECT 14684.105 189.04 14684.385 322.425 ;
      RECT 14683.545 187.94 14683.825 322.185 ;
      RECT 14682.985 189.04 14683.265 321.945 ;
      RECT 14682.425 187.94 14682.705 321.705 ;
      RECT 14642.665 189.04 14642.945 332.175 ;
      RECT 14642.105 187.94 14642.385 332.415 ;
      RECT 14641.545 189.04 14641.825 332.655 ;
      RECT 14640.985 189.04 14641.265 332.895 ;
      RECT 14640.425 189.04 14640.705 333.135 ;
      RECT 14639.865 189.04 14640.145 333.375 ;
      RECT 14639.305 189.04 14639.585 333.615 ;
      RECT 14638.745 189.04 14639.025 333.86 ;
      RECT 14638.185 189.04 14638.465 334.1 ;
      RECT 14637.625 189.04 14637.905 334.34 ;
      RECT 14637.065 187.94 14637.345 334.58 ;
      RECT 14636.505 189.04 14636.785 334.82 ;
      RECT 14635.945 187.94 14636.225 335.06 ;
      RECT 14635.385 189.04 14635.665 335.3 ;
      RECT 14634.825 189.04 14635.105 335.54 ;
      RECT 14634.265 189.04 14634.545 335.78 ;
      RECT 14633.705 189.04 14633.985 336.02 ;
      RECT 14633.145 189.04 14633.425 336.26 ;
      RECT 14632.585 189.04 14632.865 336.5 ;
      RECT 14632.025 189.04 14632.305 336.74 ;
      RECT 14631.465 189.04 14631.745 336.98 ;
      RECT 14630.905 189.04 14631.185 337.22 ;
      RECT 14630.345 189.04 14630.625 337.46 ;
      RECT 14629.785 189.04 14630.065 337.7 ;
      RECT 14620.825 189.04 14621.105 333.285 ;
      RECT 14620.265 189.04 14620.545 333.045 ;
      RECT 14619.705 189.04 14619.985 332.805 ;
      RECT 14619.145 187.94 14619.425 332.565 ;
      RECT 14618.585 189.04 14618.865 332.325 ;
      RECT 14618.025 187.94 14618.305 332.085 ;
      RECT 14617.465 189.04 14617.745 331.845 ;
      RECT 14616.905 189.04 14617.185 331.605 ;
      RECT 14616.345 189.04 14616.625 331.365 ;
      RECT 14615.785 187.94 14616.065 331.125 ;
      RECT 14615.225 189.04 14615.505 330.885 ;
      RECT 14614.665 187.94 14614.945 330.645 ;
      RECT 14614.105 189.04 14614.385 330.405 ;
      RECT 14613.545 187.94 14613.825 330.165 ;
      RECT 14611.025 189.04 14611.305 322.565 ;
      RECT 14610.465 189.04 14610.745 322.325 ;
      RECT 14609.905 189.04 14610.185 322.085 ;
      RECT 14609.345 189.04 14609.625 321.845 ;
      RECT 14608.785 189.04 14609.065 321.605 ;
      RECT 14608.225 189.04 14608.505 321.365 ;
      RECT 14607.665 189.04 14607.945 321.125 ;
      RECT 14581.625 189.04 14581.905 335 ;
      RECT 14581.065 189.04 14581.345 335.24 ;
      RECT 14580.505 189.04 14580.785 335.48 ;
      RECT 14579.945 189.04 14580.225 335.72 ;
      RECT 14579.385 189.04 14579.665 335.96 ;
      RECT 14578.825 187.94 14579.105 335.96 ;
      RECT 14578.265 189.04 14578.545 335.72 ;
      RECT 14577.705 187.94 14577.985 335.475 ;
      RECT 14577.145 189.04 14577.425 335.235 ;
      RECT 14576.585 187.94 14576.865 334.995 ;
      RECT 14576.025 189.04 14576.305 334.755 ;
      RECT 14575.465 189.04 14575.745 334.515 ;
      RECT 14574.905 189.04 14575.185 334.275 ;
      RECT 14574.345 189.04 14574.625 334.035 ;
      RECT 14573.785 189.04 14574.065 333.795 ;
      RECT 14573.225 189.04 14573.505 333.555 ;
      RECT 14572.665 189.04 14572.945 333.315 ;
      RECT 14572.105 189.04 14572.385 333.075 ;
      RECT 14571.545 187.94 14571.825 332.835 ;
      RECT 14570.985 189.04 14571.265 332.595 ;
      RECT 14570.425 187.94 14570.705 332.355 ;
      RECT 14569.865 189.04 14570.145 332.115 ;
      RECT 14569.305 189.04 14569.585 331.875 ;
      RECT 14568.745 189.04 14569.025 331.635 ;
      RECT 14555.305 189.04 14555.585 335.035 ;
      RECT 14554.745 189.04 14555.025 335.275 ;
      RECT 14554.185 189.04 14554.465 335.52 ;
      RECT 14553.625 189.04 14553.905 335.76 ;
      RECT 14553.065 189.04 14553.345 336 ;
      RECT 14552.505 189.04 14552.785 336 ;
      RECT 14551.945 189.04 14552.225 335.76 ;
      RECT 14551.385 189.04 14551.665 335.52 ;
      RECT 14550.825 189.04 14551.105 328.505 ;
      RECT 14550.265 189.04 14550.545 328.265 ;
      RECT 14549.705 189.04 14549.985 328.025 ;
      RECT 14549.145 187.94 14549.425 327.785 ;
      RECT 14548.585 189.04 14548.865 327.545 ;
      RECT 14548.025 187.94 14548.305 327.305 ;
      RECT 14547.465 189.04 14547.745 327.065 ;
      RECT 14546.905 189.04 14547.185 326.825 ;
      RECT 14546.345 189.04 14546.625 326.585 ;
      RECT 14545.785 187.94 14546.065 326.345 ;
      RECT 14545.225 189.04 14545.505 326.105 ;
      RECT 14544.665 187.94 14544.945 325.865 ;
      RECT 14544.105 189.04 14544.385 325.625 ;
      RECT 14543.545 187.94 14543.825 325.385 ;
      RECT 14542.985 189.04 14543.265 325.145 ;
      RECT 14542.425 189.04 14542.705 324.905 ;
      RECT 14502.105 189.04 14502.385 333.8 ;
      RECT 14501.545 189.04 14501.825 334.04 ;
      RECT 14500.985 189.04 14501.265 334.285 ;
      RECT 14500.425 189.04 14500.705 334.525 ;
      RECT 14499.865 189.04 14500.145 334.765 ;
      RECT 14499.305 189.04 14499.585 335.005 ;
      RECT 14498.745 189.04 14499.025 335.245 ;
      RECT 14498.185 189.04 14498.465 335.485 ;
      RECT 14497.625 189.04 14497.905 335.725 ;
      RECT 14497.065 189.04 14497.345 335.965 ;
      RECT 14496.505 187.94 14496.785 336.205 ;
      RECT 14495.945 189.04 14496.225 336.445 ;
      RECT 14495.385 187.94 14495.665 336.685 ;
      RECT 14494.825 189.04 14495.105 336.925 ;
      RECT 14494.265 187.94 14494.545 337.165 ;
      RECT 14493.705 189.04 14493.985 337.165 ;
      RECT 14493.145 189.04 14493.425 336.925 ;
      RECT 14492.585 189.04 14492.865 336.685 ;
      RECT 14492.025 189.04 14492.305 336.445 ;
      RECT 14491.465 189.04 14491.745 336.205 ;
      RECT 14490.905 189.04 14491.185 335.965 ;
      RECT 14490.345 189.04 14490.625 335.725 ;
      RECT 14489.785 189.04 14490.065 335.485 ;
      RECT 14480.825 187.94 14481.105 335.515 ;
      RECT 14480.265 189.04 14480.545 335.755 ;
      RECT 14479.705 187.94 14479.985 335.995 ;
      RECT 14479.145 189.04 14479.425 336.21 ;
      RECT 14478.585 189.04 14478.865 335.785 ;
      RECT 14478.025 189.04 14478.305 335.545 ;
      RECT 14477.465 189.04 14477.745 335.305 ;
      RECT 14476.905 189.04 14477.185 335.065 ;
      RECT 14476.345 189.04 14476.625 334.825 ;
      RECT 14475.785 189.04 14476.065 334.585 ;
      RECT 14475.225 189.04 14475.505 334.345 ;
      RECT 14474.665 189.04 14474.945 334.105 ;
      RECT 14474.105 189.04 14474.385 333.865 ;
      RECT 14473.545 189.04 14473.825 333.625 ;
      RECT 14471.025 189.04 14471.305 332.8 ;
      RECT 14470.465 189.04 14470.745 332.56 ;
      RECT 14469.905 189.04 14470.185 332.32 ;
      RECT 14469.345 187.94 14469.625 332.08 ;
      RECT 14468.785 189.04 14469.065 331.84 ;
      RECT 14468.225 187.94 14468.505 331.6 ;
      RECT 14467.665 189.04 14467.945 331.36 ;
      RECT 14467.105 189.04 14467.385 331.12 ;
      RECT 14440.505 189.04 14440.785 342.165 ;
      RECT 14439.945 187.94 14440.225 342.405 ;
      RECT 14439.385 189.04 14439.665 342.645 ;
      RECT 14438.825 187.94 14439.105 342.89 ;
      RECT 14438.265 189.04 14438.545 343.13 ;
      RECT 14437.705 187.94 14437.985 343.37 ;
      RECT 14437.145 189.04 14437.425 343.61 ;
      RECT 14436.585 189.04 14436.865 343.85 ;
      RECT 14436.025 189.04 14436.305 329.47 ;
      RECT 14435.465 189.04 14435.745 329.23 ;
      RECT 14434.905 189.04 14435.185 328.99 ;
      RECT 14434.345 189.04 14434.625 328.75 ;
      RECT 14433.785 189.04 14434.065 328.51 ;
      RECT 14433.225 189.04 14433.505 328.27 ;
      RECT 14432.665 189.04 14432.945 328.03 ;
      RECT 14432.105 189.04 14432.385 327.79 ;
      RECT 14431.545 189.04 14431.825 327.55 ;
      RECT 14430.985 189.04 14431.265 327.31 ;
      RECT 14430.425 187.94 14430.705 327.07 ;
      RECT 14429.865 189.04 14430.145 326.83 ;
      RECT 14429.305 187.94 14429.585 326.59 ;
      RECT 14428.745 189.04 14429.025 326.35 ;
      RECT 14414.745 187.94 14415.025 332.47 ;
      RECT 14414.185 189.04 14414.465 332.23 ;
      RECT 14413.625 189.04 14413.905 331.99 ;
      RECT 14413.065 189.04 14413.345 331.75 ;
      RECT 14412.505 189.04 14412.785 331.51 ;
      RECT 14411.945 189.04 14412.225 331.27 ;
      RECT 14411.385 189.04 14411.665 331.03 ;
      RECT 14410.825 189.04 14411.105 330.79 ;
      RECT 14410.265 189.04 14410.545 330.55 ;
      RECT 14409.705 187.94 14409.985 330.31 ;
      RECT 14409.145 189.04 14409.425 330.07 ;
      RECT 14408.585 187.94 14408.865 329.83 ;
      RECT 14408.025 189.04 14408.305 329.59 ;
      RECT 14407.465 189.04 14407.745 329.35 ;
      RECT 14406.905 189.04 14407.185 329.11 ;
      RECT 14406.345 189.04 14406.625 328.87 ;
      RECT 14405.785 189.04 14406.065 328.63 ;
      RECT 14405.225 189.04 14405.505 328.39 ;
      RECT 14404.665 189.04 14404.945 328.15 ;
      RECT 14404.105 189.04 14404.385 327.91 ;
      RECT 14403.545 189.04 14403.825 327.67 ;
      RECT 14402.985 189.04 14403.265 327.43 ;
      RECT 14402.425 189.04 14402.705 327.19 ;
      RECT 14363.225 189.04 14363.505 334.095 ;
      RECT 14362.665 189.04 14362.945 334.335 ;
      RECT 14362.105 189.04 14362.385 334.575 ;
      RECT 14361.545 187.94 14361.825 334.815 ;
      RECT 14360.985 189.04 14361.265 335.055 ;
      RECT 14360.425 187.94 14360.705 335.295 ;
      RECT 14359.865 189.04 14360.145 335.535 ;
      RECT 14359.305 189.04 14359.585 335.775 ;
      RECT 14358.745 189.04 14359.025 336.015 ;
      RECT 14358.185 187.94 14358.465 336.255 ;
      RECT 14357.625 189.04 14357.905 336.495 ;
      RECT 14357.065 187.94 14357.345 336.735 ;
      RECT 14356.505 189.04 14356.785 336.975 ;
      RECT 14355.945 187.94 14356.225 337.215 ;
      RECT 14355.385 189.04 14355.665 337.455 ;
      RECT 14354.825 189.04 14355.105 337.695 ;
      RECT 14354.265 189.04 14354.545 337.695 ;
      RECT 14353.705 189.04 14353.985 337.455 ;
      RECT 14353.145 189.04 14353.425 337.215 ;
      RECT 14352.585 189.04 14352.865 336.975 ;
      RECT 14352.025 189.04 14352.305 336.735 ;
      RECT 14351.465 189.04 14351.745 336.495 ;
      RECT 14350.905 189.04 14351.185 336.255 ;
      RECT 14350.345 189.04 14350.625 336.015 ;
      RECT 14349.785 189.04 14350.065 335.775 ;
      RECT 14340.825 189.04 14341.105 335.29 ;
      RECT 14340.265 187.94 14340.545 335.05 ;
      RECT 14339.705 189.04 14339.985 334.81 ;
      RECT 14339.145 187.94 14339.425 334.57 ;
      RECT 14338.585 189.04 14338.865 334.33 ;
      RECT 14338.025 187.94 14338.305 334.09 ;
      RECT 14337.465 189.04 14337.745 333.85 ;
      RECT 14336.905 189.04 14337.185 333.61 ;
      RECT 14336.345 189.04 14336.625 333.37 ;
      RECT 14335.785 189.04 14336.065 333.13 ;
      RECT 14335.225 189.04 14335.505 332.89 ;
      RECT 14334.665 189.04 14334.945 332.65 ;
      RECT 14334.105 189.04 14334.385 332.41 ;
      RECT 14333.545 189.04 14333.825 332.17 ;
      RECT 14331.025 187.94 14331.305 333.89 ;
      RECT 14330.465 189.04 14330.745 333.65 ;
      RECT 14329.905 187.94 14330.185 333.41 ;
      RECT 14329.345 189.04 14329.625 333.17 ;
      RECT 14328.785 189.04 14329.065 332.93 ;
      RECT 14328.225 189.04 14328.505 332.69 ;
      RECT 14327.665 189.04 14327.945 332.45 ;
      RECT 14327.105 189.04 14327.385 332.21 ;
      RECT 14301.065 189.04 14301.345 329.86 ;
      RECT 14300.505 189.04 14300.785 330.1 ;
      RECT 14299.945 189.04 14300.225 330.34 ;
      RECT 14299.385 189.04 14299.665 330.585 ;
      RECT 14298.825 189.04 14299.105 330.825 ;
      RECT 14298.265 189.04 14298.545 331.065 ;
      RECT 14297.705 189.04 14297.985 331.065 ;
      RECT 14297.145 189.04 14297.425 330.825 ;
      RECT 14296.585 189.04 14296.865 330.585 ;
      RECT 14296.025 187.94 14296.305 330.345 ;
      RECT 14295.465 189.04 14295.745 330.105 ;
      RECT 14294.905 187.94 14295.185 329.865 ;
      RECT 14294.345 189.04 14294.625 329.625 ;
      RECT 14293.785 189.04 14294.065 329.385 ;
      RECT 14293.225 189.04 14293.505 329.145 ;
      RECT 14292.665 187.94 14292.945 328.905 ;
      RECT 14292.105 189.04 14292.385 328.665 ;
      RECT 14291.545 187.94 14291.825 328.425 ;
      RECT 14290.985 189.04 14291.265 328.185 ;
      RECT 14290.425 187.94 14290.705 327.945 ;
      RECT 14289.865 189.04 14290.145 327.705 ;
      RECT 14289.305 189.04 14289.585 327.465 ;
      RECT 14288.745 189.04 14289.025 327.225 ;
      RECT 14288.185 189.04 14288.465 326.985 ;
      RECT 14274.745 189.04 14275.025 332.785 ;
      RECT 14274.185 189.04 14274.465 332.545 ;
      RECT 14273.625 189.04 14273.905 332.305 ;
      RECT 14273.065 189.04 14273.345 332.065 ;
      RECT 14272.505 189.04 14272.785 331.825 ;
      RECT 14271.945 189.04 14272.225 331.585 ;
      RECT 14271.385 189.04 14271.665 331.345 ;
      RECT 14270.825 189.04 14271.105 331.105 ;
      RECT 14270.265 187.94 14270.545 330.865 ;
      RECT 14269.705 189.04 14269.985 330.625 ;
      RECT 14269.145 187.94 14269.425 330.305 ;
      RECT 14268.585 189.04 14268.865 330.145 ;
      RECT 14268.025 187.94 14268.305 329.905 ;
      RECT 14267.465 189.04 14267.745 329.665 ;
      RECT 14266.905 189.04 14267.185 329.425 ;
      RECT 14266.345 189.04 14266.625 329.185 ;
      RECT 14265.785 189.04 14266.065 328.945 ;
      RECT 14265.225 189.04 14265.505 328.705 ;
      RECT 14264.665 189.04 14264.945 328.465 ;
      RECT 14264.105 189.04 14264.385 328.225 ;
      RECT 14263.545 189.04 14263.825 327.985 ;
      RECT 14262.985 187.94 14263.265 327.745 ;
      RECT 14262.425 189.04 14262.705 327.505 ;
      RECT 14261.865 187.94 14262.145 327.265 ;
      RECT 14222.665 189.04 14222.945 332.875 ;
      RECT 14222.105 189.04 14222.385 333.115 ;
      RECT 14221.545 189.04 14221.825 333.355 ;
      RECT 14220.985 189.04 14221.265 333.595 ;
      RECT 14220.425 189.04 14220.705 333.835 ;
      RECT 14219.865 189.04 14220.145 334.075 ;
      RECT 14219.305 189.04 14219.585 334.315 ;
      RECT 14218.745 189.04 14219.025 334.555 ;
      RECT 14218.185 189.04 14218.465 334.795 ;
      RECT 14217.625 189.04 14217.905 335.035 ;
      RECT 14217.065 189.04 14217.345 335.275 ;
      RECT 14216.505 189.04 14216.785 335.515 ;
      RECT 14215.945 189.04 14216.225 335.755 ;
      RECT 14215.385 189.04 14215.665 335.755 ;
      RECT 14214.825 187.94 14215.105 335.515 ;
      RECT 14214.265 189.04 14214.545 335.275 ;
      RECT 14213.705 187.94 14213.985 335.035 ;
      RECT 14213.145 189.04 14213.425 334.795 ;
      RECT 14212.585 189.04 14212.865 334.555 ;
      RECT 14212.025 189.04 14212.305 334.315 ;
      RECT 14211.465 187.94 14211.745 334.05 ;
      RECT 14210.905 189.04 14211.185 333.81 ;
      RECT 14210.345 187.94 14210.625 333.57 ;
      RECT 14209.785 189.04 14210.065 333.33 ;
      RECT 14200.825 187.94 14201.105 327.165 ;
      RECT 14200.265 189.04 14200.545 327.405 ;
      RECT 14199.705 189.04 14199.985 327.645 ;
      RECT 14199.145 189.04 14199.425 327.645 ;
      RECT 14198.585 189.04 14198.865 327.405 ;
      RECT 14198.025 189.04 14198.305 327.165 ;
      RECT 14197.465 189.04 14197.745 326.925 ;
      RECT 14196.905 189.04 14197.185 326.685 ;
      RECT 14196.345 189.04 14196.625 326.445 ;
      RECT 14195.785 189.04 14196.065 326.205 ;
      RECT 14195.225 189.04 14195.505 325.965 ;
      RECT 14194.665 189.04 14194.945 325.725 ;
      RECT 14194.105 189.04 14194.385 325.485 ;
      RECT 14193.545 187.94 14193.825 325.245 ;
      RECT 14191.025 189.04 14191.305 326.965 ;
      RECT 14190.465 187.94 14190.745 326.725 ;
      RECT 14189.905 189.04 14190.185 326.485 ;
      RECT 14189.345 187.94 14189.625 326.245 ;
      RECT 14188.785 189.04 14189.065 326.005 ;
      RECT 14188.225 189.04 14188.505 325.765 ;
      RECT 14187.665 189.04 14187.945 325.525 ;
      RECT 14161.625 189.04 14161.905 328.31 ;
      RECT 14161.065 189.04 14161.345 328.55 ;
      RECT 14160.505 189.04 14160.785 328.79 ;
      RECT 14159.945 189.04 14160.225 329.03 ;
      RECT 14159.385 189.04 14159.665 329.27 ;
      RECT 14158.825 187.94 14159.105 329.51 ;
      RECT 14158.265 189.04 14158.545 329.75 ;
      RECT 14157.705 187.94 14157.985 329.99 ;
      RECT 14157.145 189.04 14157.425 330.23 ;
      RECT 14156.585 189.04 14156.865 330.47 ;
      RECT 14156.025 189.04 14156.305 330.71 ;
      RECT 14155.465 189.04 14155.745 330.95 ;
      RECT 14154.905 189.04 14155.185 331.19 ;
      RECT 14154.345 189.04 14154.625 331.43 ;
      RECT 14153.785 189.04 14154.065 331.67 ;
      RECT 14153.225 189.04 14153.505 331.67 ;
      RECT 14152.665 189.04 14152.945 331.43 ;
      RECT 14152.105 189.04 14152.385 331.19 ;
      RECT 14151.545 189.04 14151.825 330.95 ;
      RECT 14150.985 189.04 14151.265 330.705 ;
      RECT 14150.425 189.04 14150.705 330.465 ;
      RECT 14149.865 189.04 14150.145 330.225 ;
      RECT 14149.305 187.94 14149.585 329.985 ;
      RECT 14148.745 189.04 14149.025 329.745 ;
      RECT 14135.305 187.94 14135.585 327.225 ;
      RECT 14134.745 189.04 14135.025 326.985 ;
      RECT 14134.185 189.04 14134.465 326.745 ;
      RECT 14133.625 189.04 14133.905 326.505 ;
      RECT 14133.065 187.94 14133.345 326.265 ;
      RECT 14132.505 189.04 14132.785 326.025 ;
      RECT 14131.945 187.94 14132.225 325.785 ;
      RECT 14131.385 189.04 14131.665 325.545 ;
      RECT 14130.825 187.94 14131.105 325.305 ;
      RECT 14130.265 189.04 14130.545 325.065 ;
      RECT 14129.705 189.04 14129.985 324.825 ;
      RECT 14129.145 189.04 14129.425 324.585 ;
      RECT 14128.585 189.04 14128.865 324.345 ;
      RECT 14128.025 189.04 14128.305 324.105 ;
      RECT 14127.465 189.04 14127.745 323.865 ;
      RECT 14126.905 189.04 14127.185 323.625 ;
      RECT 14126.345 189.04 14126.625 323.385 ;
      RECT 14125.785 189.04 14126.065 323.145 ;
      RECT 14125.225 189.04 14125.505 322.905 ;
      RECT 14124.665 189.04 14124.945 322.665 ;
      RECT 14124.105 189.04 14124.385 322.425 ;
      RECT 14123.545 187.94 14123.825 322.185 ;
      RECT 14122.985 189.04 14123.265 321.945 ;
      RECT 14122.425 187.94 14122.705 321.705 ;
      RECT 14082.665 189.04 14082.945 332.175 ;
      RECT 14082.105 187.94 14082.385 332.415 ;
      RECT 14081.545 189.04 14081.825 332.655 ;
      RECT 14080.985 189.04 14081.265 332.895 ;
      RECT 14080.425 189.04 14080.705 333.135 ;
      RECT 14079.865 189.04 14080.145 333.375 ;
      RECT 14079.305 189.04 14079.585 333.615 ;
      RECT 14078.745 189.04 14079.025 333.86 ;
      RECT 14078.185 189.04 14078.465 334.1 ;
      RECT 14077.625 189.04 14077.905 334.34 ;
      RECT 14077.065 187.94 14077.345 334.58 ;
      RECT 14076.505 189.04 14076.785 334.82 ;
      RECT 14075.945 187.94 14076.225 335.06 ;
      RECT 14075.385 189.04 14075.665 335.3 ;
      RECT 14074.825 189.04 14075.105 335.54 ;
      RECT 14074.265 189.04 14074.545 335.78 ;
      RECT 14073.705 189.04 14073.985 336.02 ;
      RECT 14073.145 189.04 14073.425 336.26 ;
      RECT 14072.585 189.04 14072.865 336.5 ;
      RECT 14072.025 189.04 14072.305 336.74 ;
      RECT 14071.465 189.04 14071.745 336.98 ;
      RECT 14070.905 189.04 14071.185 337.22 ;
      RECT 14070.345 189.04 14070.625 337.46 ;
      RECT 14069.785 189.04 14070.065 337.7 ;
      RECT 14060.825 189.04 14061.105 333.285 ;
      RECT 14060.265 189.04 14060.545 333.045 ;
      RECT 14059.705 189.04 14059.985 332.805 ;
      RECT 14059.145 187.94 14059.425 332.565 ;
      RECT 14058.585 189.04 14058.865 332.325 ;
      RECT 14058.025 187.94 14058.305 332.085 ;
      RECT 14057.465 189.04 14057.745 331.845 ;
      RECT 14056.905 189.04 14057.185 331.605 ;
      RECT 14056.345 189.04 14056.625 331.365 ;
      RECT 14055.785 187.94 14056.065 331.125 ;
      RECT 14055.225 189.04 14055.505 330.885 ;
      RECT 14054.665 187.94 14054.945 330.645 ;
      RECT 14054.105 189.04 14054.385 330.405 ;
      RECT 14053.545 187.94 14053.825 330.165 ;
      RECT 14051.025 189.04 14051.305 322.565 ;
      RECT 14050.465 189.04 14050.745 322.325 ;
      RECT 14049.905 189.04 14050.185 322.085 ;
      RECT 14049.345 189.04 14049.625 321.845 ;
      RECT 14048.785 189.04 14049.065 321.605 ;
      RECT 14048.225 189.04 14048.505 321.365 ;
      RECT 14047.665 189.04 14047.945 321.125 ;
      RECT 14021.625 189.04 14021.905 335 ;
      RECT 14021.065 189.04 14021.345 335.24 ;
      RECT 14020.505 189.04 14020.785 335.48 ;
      RECT 14019.945 189.04 14020.225 335.72 ;
      RECT 14019.385 189.04 14019.665 335.96 ;
      RECT 14018.825 187.94 14019.105 335.96 ;
      RECT 14018.265 189.04 14018.545 335.72 ;
      RECT 14017.705 187.94 14017.985 335.475 ;
      RECT 14017.145 189.04 14017.425 335.235 ;
      RECT 14016.585 187.94 14016.865 334.995 ;
      RECT 14016.025 189.04 14016.305 334.755 ;
      RECT 14015.465 189.04 14015.745 334.515 ;
      RECT 14014.905 189.04 14015.185 334.275 ;
      RECT 14014.345 189.04 14014.625 334.035 ;
      RECT 14013.785 189.04 14014.065 333.795 ;
      RECT 14013.225 189.04 14013.505 333.555 ;
      RECT 14012.665 189.04 14012.945 333.315 ;
      RECT 14012.105 189.04 14012.385 333.075 ;
      RECT 14011.545 187.94 14011.825 332.835 ;
      RECT 14010.985 189.04 14011.265 332.595 ;
      RECT 14010.425 187.94 14010.705 332.355 ;
      RECT 14009.865 189.04 14010.145 332.115 ;
      RECT 14009.305 189.04 14009.585 331.875 ;
      RECT 14008.745 189.04 14009.025 331.635 ;
      RECT 13995.305 189.04 13995.585 335.035 ;
      RECT 13994.745 189.04 13995.025 335.275 ;
      RECT 13994.185 189.04 13994.465 335.52 ;
      RECT 13993.625 189.04 13993.905 335.76 ;
      RECT 13993.065 189.04 13993.345 336 ;
      RECT 13992.505 189.04 13992.785 336 ;
      RECT 13991.945 189.04 13992.225 335.76 ;
      RECT 13991.385 189.04 13991.665 335.52 ;
      RECT 13990.825 189.04 13991.105 328.505 ;
      RECT 13990.265 189.04 13990.545 328.265 ;
      RECT 13989.705 189.04 13989.985 328.025 ;
      RECT 13989.145 187.94 13989.425 327.785 ;
      RECT 13988.585 189.04 13988.865 327.545 ;
      RECT 13988.025 187.94 13988.305 327.305 ;
      RECT 13987.465 189.04 13987.745 327.065 ;
      RECT 13986.905 189.04 13987.185 326.825 ;
      RECT 13986.345 189.04 13986.625 326.585 ;
      RECT 13985.785 187.94 13986.065 326.345 ;
      RECT 13985.225 189.04 13985.505 326.105 ;
      RECT 13984.665 187.94 13984.945 325.865 ;
      RECT 13984.105 189.04 13984.385 325.625 ;
      RECT 13983.545 187.94 13983.825 325.385 ;
      RECT 13982.985 189.04 13983.265 325.145 ;
      RECT 13982.425 189.04 13982.705 324.905 ;
      RECT 13942.105 189.04 13942.385 333.8 ;
      RECT 13941.545 189.04 13941.825 334.04 ;
      RECT 13940.985 189.04 13941.265 334.285 ;
      RECT 13940.425 189.04 13940.705 334.525 ;
      RECT 13939.865 189.04 13940.145 334.765 ;
      RECT 13939.305 189.04 13939.585 335.005 ;
      RECT 13938.745 189.04 13939.025 335.245 ;
      RECT 13938.185 189.04 13938.465 335.485 ;
      RECT 13937.625 189.04 13937.905 335.725 ;
      RECT 13937.065 189.04 13937.345 335.965 ;
      RECT 13936.505 187.94 13936.785 336.205 ;
      RECT 13935.945 189.04 13936.225 336.445 ;
      RECT 13935.385 187.94 13935.665 336.685 ;
      RECT 13934.825 189.04 13935.105 336.925 ;
      RECT 13934.265 187.94 13934.545 337.165 ;
      RECT 13933.705 189.04 13933.985 337.165 ;
      RECT 13933.145 189.04 13933.425 336.925 ;
      RECT 13932.585 189.04 13932.865 336.685 ;
      RECT 13932.025 189.04 13932.305 336.445 ;
      RECT 13931.465 189.04 13931.745 336.205 ;
      RECT 13930.905 189.04 13931.185 335.965 ;
      RECT 13930.345 189.04 13930.625 335.725 ;
      RECT 13929.785 189.04 13930.065 335.485 ;
      RECT 13920.825 187.94 13921.105 335.515 ;
      RECT 13920.265 189.04 13920.545 335.755 ;
      RECT 13919.705 187.94 13919.985 335.995 ;
      RECT 13919.145 189.04 13919.425 336.21 ;
      RECT 13918.585 189.04 13918.865 335.785 ;
      RECT 13918.025 189.04 13918.305 335.545 ;
      RECT 13917.465 189.04 13917.745 335.305 ;
      RECT 13916.905 189.04 13917.185 335.065 ;
      RECT 13916.345 189.04 13916.625 334.825 ;
      RECT 13915.785 189.04 13916.065 334.585 ;
      RECT 13915.225 189.04 13915.505 334.345 ;
      RECT 13914.665 189.04 13914.945 334.105 ;
      RECT 13914.105 189.04 13914.385 333.865 ;
      RECT 13913.545 189.04 13913.825 333.625 ;
      RECT 13911.025 189.04 13911.305 332.8 ;
      RECT 13910.465 189.04 13910.745 332.56 ;
      RECT 13909.905 189.04 13910.185 332.32 ;
      RECT 13909.345 187.94 13909.625 332.08 ;
      RECT 13908.785 189.04 13909.065 331.84 ;
      RECT 13908.225 187.94 13908.505 331.6 ;
      RECT 13907.665 189.04 13907.945 331.36 ;
      RECT 13907.105 189.04 13907.385 331.12 ;
      RECT 13880.505 189.04 13880.785 342.165 ;
      RECT 13879.945 187.94 13880.225 342.405 ;
      RECT 13879.385 189.04 13879.665 342.645 ;
      RECT 13878.825 187.94 13879.105 342.89 ;
      RECT 13878.265 189.04 13878.545 343.13 ;
      RECT 13877.705 187.94 13877.985 343.37 ;
      RECT 13877.145 189.04 13877.425 343.61 ;
      RECT 13876.585 189.04 13876.865 343.85 ;
      RECT 13876.025 189.04 13876.305 329.47 ;
      RECT 13875.465 189.04 13875.745 329.23 ;
      RECT 13874.905 189.04 13875.185 328.99 ;
      RECT 13874.345 189.04 13874.625 328.75 ;
      RECT 13873.785 189.04 13874.065 328.51 ;
      RECT 13873.225 189.04 13873.505 328.27 ;
      RECT 13872.665 189.04 13872.945 328.03 ;
      RECT 13872.105 189.04 13872.385 327.79 ;
      RECT 13871.545 189.04 13871.825 327.55 ;
      RECT 13870.985 189.04 13871.265 327.31 ;
      RECT 13870.425 187.94 13870.705 327.07 ;
      RECT 13869.865 189.04 13870.145 326.83 ;
      RECT 13869.305 187.94 13869.585 326.59 ;
      RECT 13868.745 189.04 13869.025 326.35 ;
      RECT 13854.745 187.94 13855.025 332.47 ;
      RECT 13854.185 189.04 13854.465 332.23 ;
      RECT 13853.625 189.04 13853.905 331.99 ;
      RECT 13853.065 189.04 13853.345 331.75 ;
      RECT 13852.505 189.04 13852.785 331.51 ;
      RECT 13851.945 189.04 13852.225 331.27 ;
      RECT 13851.385 189.04 13851.665 331.03 ;
      RECT 13850.825 189.04 13851.105 330.79 ;
      RECT 13850.265 189.04 13850.545 330.55 ;
      RECT 13849.705 187.94 13849.985 330.31 ;
      RECT 13849.145 189.04 13849.425 330.07 ;
      RECT 13848.585 187.94 13848.865 329.83 ;
      RECT 13848.025 189.04 13848.305 329.59 ;
      RECT 13847.465 189.04 13847.745 329.35 ;
      RECT 13846.905 189.04 13847.185 329.11 ;
      RECT 13846.345 189.04 13846.625 328.87 ;
      RECT 13845.785 189.04 13846.065 328.63 ;
      RECT 13845.225 189.04 13845.505 328.39 ;
      RECT 13844.665 189.04 13844.945 328.15 ;
      RECT 13844.105 189.04 13844.385 327.91 ;
      RECT 13843.545 189.04 13843.825 327.67 ;
      RECT 13842.985 189.04 13843.265 327.43 ;
      RECT 13842.425 189.04 13842.705 327.19 ;
      RECT 13803.225 189.04 13803.505 334.095 ;
      RECT 13802.665 189.04 13802.945 334.335 ;
      RECT 13802.105 189.04 13802.385 334.575 ;
      RECT 13801.545 187.94 13801.825 334.815 ;
      RECT 13800.985 189.04 13801.265 335.055 ;
      RECT 13800.425 187.94 13800.705 335.295 ;
      RECT 13799.865 189.04 13800.145 335.535 ;
      RECT 13799.305 189.04 13799.585 335.775 ;
      RECT 13798.745 189.04 13799.025 336.015 ;
      RECT 13798.185 187.94 13798.465 336.255 ;
      RECT 13797.625 189.04 13797.905 336.495 ;
      RECT 13797.065 187.94 13797.345 336.735 ;
      RECT 13796.505 189.04 13796.785 336.975 ;
      RECT 13795.945 187.94 13796.225 337.215 ;
      RECT 13795.385 189.04 13795.665 337.455 ;
      RECT 13794.825 189.04 13795.105 337.695 ;
      RECT 13794.265 189.04 13794.545 337.695 ;
      RECT 13793.705 189.04 13793.985 337.455 ;
      RECT 13793.145 189.04 13793.425 337.215 ;
      RECT 13792.585 189.04 13792.865 336.975 ;
      RECT 13792.025 189.04 13792.305 336.735 ;
      RECT 13791.465 189.04 13791.745 336.495 ;
      RECT 13790.905 189.04 13791.185 336.255 ;
      RECT 13790.345 189.04 13790.625 336.015 ;
      RECT 13789.785 189.04 13790.065 335.775 ;
      RECT 13780.825 189.04 13781.105 335.29 ;
      RECT 13780.265 187.94 13780.545 335.05 ;
      RECT 13779.705 189.04 13779.985 334.81 ;
      RECT 13779.145 187.94 13779.425 334.57 ;
      RECT 13778.585 189.04 13778.865 334.33 ;
      RECT 13778.025 187.94 13778.305 334.09 ;
      RECT 13777.465 189.04 13777.745 333.85 ;
      RECT 13776.905 189.04 13777.185 333.61 ;
      RECT 13776.345 189.04 13776.625 333.37 ;
      RECT 13775.785 189.04 13776.065 333.13 ;
      RECT 13775.225 189.04 13775.505 332.89 ;
      RECT 13774.665 189.04 13774.945 332.65 ;
      RECT 13774.105 189.04 13774.385 332.41 ;
      RECT 13773.545 189.04 13773.825 332.17 ;
      RECT 13771.025 187.94 13771.305 333.89 ;
      RECT 13770.465 189.04 13770.745 333.65 ;
      RECT 13769.905 187.94 13770.185 333.41 ;
      RECT 13769.345 189.04 13769.625 333.17 ;
      RECT 13768.785 189.04 13769.065 332.93 ;
      RECT 13768.225 189.04 13768.505 332.69 ;
      RECT 13767.665 189.04 13767.945 332.45 ;
      RECT 13767.105 189.04 13767.385 332.21 ;
      RECT 13741.065 189.04 13741.345 329.86 ;
      RECT 13740.505 189.04 13740.785 330.1 ;
      RECT 13739.945 189.04 13740.225 330.34 ;
      RECT 13739.385 189.04 13739.665 330.585 ;
      RECT 13738.825 189.04 13739.105 330.825 ;
      RECT 13738.265 189.04 13738.545 331.065 ;
      RECT 13737.705 189.04 13737.985 331.065 ;
      RECT 13737.145 189.04 13737.425 330.825 ;
      RECT 13736.585 189.04 13736.865 330.585 ;
      RECT 13736.025 187.94 13736.305 330.345 ;
      RECT 13735.465 189.04 13735.745 330.105 ;
      RECT 13734.905 187.94 13735.185 329.865 ;
      RECT 13734.345 189.04 13734.625 329.625 ;
      RECT 13733.785 189.04 13734.065 329.385 ;
      RECT 13733.225 189.04 13733.505 329.145 ;
      RECT 13732.665 187.94 13732.945 328.905 ;
      RECT 13732.105 189.04 13732.385 328.665 ;
      RECT 13731.545 187.94 13731.825 328.425 ;
      RECT 13730.985 189.04 13731.265 328.185 ;
      RECT 13730.425 187.94 13730.705 327.945 ;
      RECT 13729.865 189.04 13730.145 327.705 ;
      RECT 13729.305 189.04 13729.585 327.465 ;
      RECT 13728.745 189.04 13729.025 327.225 ;
      RECT 13728.185 189.04 13728.465 326.985 ;
      RECT 13714.745 189.04 13715.025 332.785 ;
      RECT 13714.185 189.04 13714.465 332.545 ;
      RECT 13713.625 189.04 13713.905 332.305 ;
      RECT 13713.065 189.04 13713.345 332.065 ;
      RECT 13712.505 189.04 13712.785 331.825 ;
      RECT 13711.945 189.04 13712.225 331.585 ;
      RECT 13711.385 189.04 13711.665 331.345 ;
      RECT 13710.825 189.04 13711.105 331.105 ;
      RECT 13710.265 187.94 13710.545 330.865 ;
      RECT 13709.705 189.04 13709.985 330.625 ;
      RECT 13709.145 187.94 13709.425 330.305 ;
      RECT 13708.585 189.04 13708.865 330.145 ;
      RECT 13708.025 187.94 13708.305 329.905 ;
      RECT 13707.465 189.04 13707.745 329.665 ;
      RECT 13706.905 189.04 13707.185 329.425 ;
      RECT 13706.345 189.04 13706.625 329.185 ;
      RECT 13705.785 189.04 13706.065 328.945 ;
      RECT 13705.225 189.04 13705.505 328.705 ;
      RECT 13704.665 189.04 13704.945 328.465 ;
      RECT 13704.105 189.04 13704.385 328.225 ;
      RECT 13703.545 189.04 13703.825 327.985 ;
      RECT 13702.985 187.94 13703.265 327.745 ;
      RECT 13702.425 189.04 13702.705 327.505 ;
      RECT 13701.865 187.94 13702.145 327.265 ;
      RECT 13662.665 189.04 13662.945 332.875 ;
      RECT 13662.105 189.04 13662.385 333.115 ;
      RECT 13661.545 189.04 13661.825 333.355 ;
      RECT 13660.985 189.04 13661.265 333.595 ;
      RECT 13660.425 189.04 13660.705 333.835 ;
      RECT 13659.865 189.04 13660.145 334.075 ;
      RECT 13659.305 189.04 13659.585 334.315 ;
      RECT 13658.745 189.04 13659.025 334.555 ;
      RECT 13658.185 189.04 13658.465 334.795 ;
      RECT 13657.625 189.04 13657.905 335.035 ;
      RECT 13657.065 189.04 13657.345 335.275 ;
      RECT 13656.505 189.04 13656.785 335.515 ;
      RECT 13655.945 189.04 13656.225 335.755 ;
      RECT 13655.385 189.04 13655.665 335.755 ;
      RECT 13654.825 187.94 13655.105 335.515 ;
      RECT 13654.265 189.04 13654.545 335.275 ;
      RECT 13653.705 187.94 13653.985 335.035 ;
      RECT 13653.145 189.04 13653.425 334.795 ;
      RECT 13652.585 189.04 13652.865 334.555 ;
      RECT 13652.025 189.04 13652.305 334.315 ;
      RECT 13651.465 187.94 13651.745 334.05 ;
      RECT 13650.905 189.04 13651.185 333.81 ;
      RECT 13650.345 187.94 13650.625 333.57 ;
      RECT 13649.785 189.04 13650.065 333.33 ;
      RECT 13640.825 187.94 13641.105 327.165 ;
      RECT 13640.265 189.04 13640.545 327.405 ;
      RECT 13639.705 189.04 13639.985 327.645 ;
      RECT 13639.145 189.04 13639.425 327.645 ;
      RECT 13638.585 189.04 13638.865 327.405 ;
      RECT 13638.025 189.04 13638.305 327.165 ;
      RECT 13637.465 189.04 13637.745 326.925 ;
      RECT 13636.905 189.04 13637.185 326.685 ;
      RECT 13636.345 189.04 13636.625 326.445 ;
      RECT 13635.785 189.04 13636.065 326.205 ;
      RECT 13635.225 189.04 13635.505 325.965 ;
      RECT 13634.665 189.04 13634.945 325.725 ;
      RECT 13634.105 189.04 13634.385 325.485 ;
      RECT 13633.545 187.94 13633.825 325.245 ;
      RECT 13631.025 189.04 13631.305 326.965 ;
      RECT 13630.465 187.94 13630.745 326.725 ;
      RECT 13629.905 189.04 13630.185 326.485 ;
      RECT 13629.345 187.94 13629.625 326.245 ;
      RECT 13628.785 189.04 13629.065 326.005 ;
      RECT 13628.225 189.04 13628.505 325.765 ;
      RECT 13627.665 189.04 13627.945 325.525 ;
      RECT 13601.625 189.04 13601.905 328.31 ;
      RECT 13601.065 189.04 13601.345 328.55 ;
      RECT 13600.505 189.04 13600.785 328.79 ;
      RECT 13599.945 189.04 13600.225 329.03 ;
      RECT 13599.385 189.04 13599.665 329.27 ;
      RECT 13598.825 187.94 13599.105 329.51 ;
      RECT 13598.265 189.04 13598.545 329.75 ;
      RECT 13597.705 187.94 13597.985 329.99 ;
      RECT 13597.145 189.04 13597.425 330.23 ;
      RECT 13596.585 189.04 13596.865 330.47 ;
      RECT 13596.025 189.04 13596.305 330.71 ;
      RECT 13595.465 189.04 13595.745 330.95 ;
      RECT 13594.905 189.04 13595.185 331.19 ;
      RECT 13594.345 189.04 13594.625 331.43 ;
      RECT 13593.785 189.04 13594.065 331.67 ;
      RECT 13593.225 189.04 13593.505 331.67 ;
      RECT 13592.665 189.04 13592.945 331.43 ;
      RECT 13592.105 189.04 13592.385 331.19 ;
      RECT 13591.545 189.04 13591.825 330.95 ;
      RECT 13590.985 189.04 13591.265 330.705 ;
      RECT 13590.425 189.04 13590.705 330.465 ;
      RECT 13589.865 189.04 13590.145 330.225 ;
      RECT 13589.305 187.94 13589.585 329.985 ;
      RECT 13588.745 189.04 13589.025 329.745 ;
      RECT 13575.305 187.94 13575.585 327.225 ;
      RECT 13574.745 189.04 13575.025 326.985 ;
      RECT 13574.185 189.04 13574.465 326.745 ;
      RECT 13573.625 189.04 13573.905 326.505 ;
      RECT 13573.065 187.94 13573.345 326.265 ;
      RECT 13572.505 189.04 13572.785 326.025 ;
      RECT 13571.945 187.94 13572.225 325.785 ;
      RECT 13571.385 189.04 13571.665 325.545 ;
      RECT 13570.825 187.94 13571.105 325.305 ;
      RECT 13570.265 189.04 13570.545 325.065 ;
      RECT 13569.705 189.04 13569.985 324.825 ;
      RECT 13569.145 189.04 13569.425 324.585 ;
      RECT 13568.585 189.04 13568.865 324.345 ;
      RECT 13568.025 189.04 13568.305 324.105 ;
      RECT 13567.465 189.04 13567.745 323.865 ;
      RECT 13566.905 189.04 13567.185 323.625 ;
      RECT 13566.345 189.04 13566.625 323.385 ;
      RECT 13565.785 189.04 13566.065 323.145 ;
      RECT 13565.225 189.04 13565.505 322.905 ;
      RECT 13564.665 189.04 13564.945 322.665 ;
      RECT 13564.105 189.04 13564.385 322.425 ;
      RECT 13563.545 187.94 13563.825 322.185 ;
      RECT 13562.985 189.04 13563.265 321.945 ;
      RECT 13562.425 187.94 13562.705 321.705 ;
      RECT 13522.665 189.04 13522.945 332.175 ;
      RECT 13522.105 187.94 13522.385 332.415 ;
      RECT 13521.545 189.04 13521.825 332.655 ;
      RECT 13520.985 189.04 13521.265 332.895 ;
      RECT 13520.425 189.04 13520.705 333.135 ;
      RECT 13519.865 189.04 13520.145 333.375 ;
      RECT 13519.305 189.04 13519.585 333.615 ;
      RECT 13518.745 189.04 13519.025 333.86 ;
      RECT 13518.185 189.04 13518.465 334.1 ;
      RECT 13517.625 189.04 13517.905 334.34 ;
      RECT 13517.065 187.94 13517.345 334.58 ;
      RECT 13516.505 189.04 13516.785 334.82 ;
      RECT 13515.945 187.94 13516.225 335.06 ;
      RECT 13515.385 189.04 13515.665 335.3 ;
      RECT 13514.825 189.04 13515.105 335.54 ;
      RECT 13514.265 189.04 13514.545 335.78 ;
      RECT 13513.705 189.04 13513.985 336.02 ;
      RECT 13513.145 189.04 13513.425 336.26 ;
      RECT 13512.585 189.04 13512.865 336.5 ;
      RECT 13512.025 189.04 13512.305 336.74 ;
      RECT 13511.465 189.04 13511.745 336.98 ;
      RECT 13510.905 189.04 13511.185 337.22 ;
      RECT 13510.345 189.04 13510.625 337.46 ;
      RECT 13509.785 189.04 13510.065 337.7 ;
      RECT 13500.825 189.04 13501.105 333.285 ;
      RECT 13500.265 189.04 13500.545 333.045 ;
      RECT 13499.705 189.04 13499.985 332.805 ;
      RECT 13499.145 187.94 13499.425 332.565 ;
      RECT 13498.585 189.04 13498.865 332.325 ;
      RECT 13498.025 187.94 13498.305 332.085 ;
      RECT 13497.465 189.04 13497.745 331.845 ;
      RECT 13496.905 189.04 13497.185 331.605 ;
      RECT 13496.345 189.04 13496.625 331.365 ;
      RECT 13495.785 187.94 13496.065 331.125 ;
      RECT 13495.225 189.04 13495.505 330.885 ;
      RECT 13494.665 187.94 13494.945 330.645 ;
      RECT 13494.105 189.04 13494.385 330.405 ;
      RECT 13493.545 187.94 13493.825 330.165 ;
      RECT 13491.025 189.04 13491.305 322.565 ;
      RECT 13490.465 189.04 13490.745 322.325 ;
      RECT 13489.905 189.04 13490.185 322.085 ;
      RECT 13489.345 189.04 13489.625 321.845 ;
      RECT 13488.785 189.04 13489.065 321.605 ;
      RECT 13488.225 189.04 13488.505 321.365 ;
      RECT 13487.665 189.04 13487.945 321.125 ;
      RECT 13461.625 189.04 13461.905 335 ;
      RECT 13461.065 189.04 13461.345 335.24 ;
      RECT 13460.505 189.04 13460.785 335.48 ;
      RECT 13459.945 189.04 13460.225 335.72 ;
      RECT 13459.385 189.04 13459.665 335.96 ;
      RECT 13458.825 187.94 13459.105 335.96 ;
      RECT 13458.265 189.04 13458.545 335.72 ;
      RECT 13457.705 187.94 13457.985 335.475 ;
      RECT 13457.145 189.04 13457.425 335.235 ;
      RECT 13456.585 187.94 13456.865 334.995 ;
      RECT 13456.025 189.04 13456.305 334.755 ;
      RECT 13455.465 189.04 13455.745 334.515 ;
      RECT 13454.905 189.04 13455.185 334.275 ;
      RECT 13454.345 189.04 13454.625 334.035 ;
      RECT 13453.785 189.04 13454.065 333.795 ;
      RECT 13453.225 189.04 13453.505 333.555 ;
      RECT 13452.665 189.04 13452.945 333.315 ;
      RECT 13452.105 189.04 13452.385 333.075 ;
      RECT 13451.545 187.94 13451.825 332.835 ;
      RECT 13450.985 189.04 13451.265 332.595 ;
      RECT 13450.425 187.94 13450.705 332.355 ;
      RECT 13449.865 189.04 13450.145 332.115 ;
      RECT 13449.305 189.04 13449.585 331.875 ;
      RECT 13448.745 189.04 13449.025 331.635 ;
      RECT 13435.305 189.04 13435.585 335.035 ;
      RECT 13434.745 189.04 13435.025 335.275 ;
      RECT 13434.185 189.04 13434.465 335.52 ;
      RECT 13433.625 189.04 13433.905 335.76 ;
      RECT 13433.065 189.04 13433.345 336 ;
      RECT 13432.505 189.04 13432.785 336 ;
      RECT 13431.945 189.04 13432.225 335.76 ;
      RECT 13431.385 189.04 13431.665 335.52 ;
      RECT 13430.825 189.04 13431.105 328.505 ;
      RECT 13430.265 189.04 13430.545 328.265 ;
      RECT 13429.705 189.04 13429.985 328.025 ;
      RECT 13429.145 187.94 13429.425 327.785 ;
      RECT 13428.585 189.04 13428.865 327.545 ;
      RECT 13428.025 187.94 13428.305 327.305 ;
      RECT 13427.465 189.04 13427.745 327.065 ;
      RECT 13426.905 189.04 13427.185 326.825 ;
      RECT 13426.345 189.04 13426.625 326.585 ;
      RECT 13425.785 187.94 13426.065 326.345 ;
      RECT 13425.225 189.04 13425.505 326.105 ;
      RECT 13424.665 187.94 13424.945 325.865 ;
      RECT 13424.105 189.04 13424.385 325.625 ;
      RECT 13423.545 187.94 13423.825 325.385 ;
      RECT 13422.985 189.04 13423.265 325.145 ;
      RECT 13422.425 189.04 13422.705 324.905 ;
      RECT 13382.105 189.04 13382.385 333.8 ;
      RECT 13381.545 189.04 13381.825 334.04 ;
      RECT 13380.985 189.04 13381.265 334.285 ;
      RECT 13380.425 189.04 13380.705 334.525 ;
      RECT 13379.865 189.04 13380.145 334.765 ;
      RECT 13379.305 189.04 13379.585 335.005 ;
      RECT 13378.745 189.04 13379.025 335.245 ;
      RECT 13378.185 189.04 13378.465 335.485 ;
      RECT 13377.625 189.04 13377.905 335.725 ;
      RECT 13377.065 189.04 13377.345 335.965 ;
      RECT 13376.505 187.94 13376.785 336.205 ;
      RECT 13375.945 189.04 13376.225 336.445 ;
      RECT 13375.385 187.94 13375.665 336.685 ;
      RECT 13374.825 189.04 13375.105 336.925 ;
      RECT 13374.265 187.94 13374.545 337.165 ;
      RECT 13373.705 189.04 13373.985 337.165 ;
      RECT 13373.145 189.04 13373.425 336.925 ;
      RECT 13372.585 189.04 13372.865 336.685 ;
      RECT 13372.025 189.04 13372.305 336.445 ;
      RECT 13371.465 189.04 13371.745 336.205 ;
      RECT 13370.905 189.04 13371.185 335.965 ;
      RECT 13370.345 189.04 13370.625 335.725 ;
      RECT 13369.785 189.04 13370.065 335.485 ;
      RECT 13360.825 187.94 13361.105 335.515 ;
      RECT 13360.265 189.04 13360.545 335.755 ;
      RECT 13359.705 187.94 13359.985 335.995 ;
      RECT 13359.145 189.04 13359.425 336.21 ;
      RECT 13358.585 189.04 13358.865 335.785 ;
      RECT 13358.025 189.04 13358.305 335.545 ;
      RECT 13357.465 189.04 13357.745 335.305 ;
      RECT 13356.905 189.04 13357.185 335.065 ;
      RECT 13356.345 189.04 13356.625 334.825 ;
      RECT 13355.785 189.04 13356.065 334.585 ;
      RECT 13355.225 189.04 13355.505 334.345 ;
      RECT 13354.665 189.04 13354.945 334.105 ;
      RECT 13354.105 189.04 13354.385 333.865 ;
      RECT 13353.545 189.04 13353.825 333.625 ;
      RECT 13351.025 189.04 13351.305 332.8 ;
      RECT 13350.465 189.04 13350.745 332.56 ;
      RECT 13349.905 189.04 13350.185 332.32 ;
      RECT 13349.345 187.94 13349.625 332.08 ;
      RECT 13348.785 189.04 13349.065 331.84 ;
      RECT 13348.225 187.94 13348.505 331.6 ;
      RECT 13347.665 189.04 13347.945 331.36 ;
      RECT 13347.105 189.04 13347.385 331.12 ;
      RECT 13320.505 189.04 13320.785 342.165 ;
      RECT 13319.945 187.94 13320.225 342.405 ;
      RECT 13319.385 189.04 13319.665 342.645 ;
      RECT 13318.825 187.94 13319.105 342.89 ;
      RECT 13318.265 189.04 13318.545 343.13 ;
      RECT 13317.705 187.94 13317.985 343.37 ;
      RECT 13317.145 189.04 13317.425 343.61 ;
      RECT 13316.585 189.04 13316.865 343.85 ;
      RECT 13316.025 189.04 13316.305 329.47 ;
      RECT 13315.465 189.04 13315.745 329.23 ;
      RECT 13314.905 189.04 13315.185 328.99 ;
      RECT 13314.345 189.04 13314.625 328.75 ;
      RECT 13313.785 189.04 13314.065 328.51 ;
      RECT 13313.225 189.04 13313.505 328.27 ;
      RECT 13312.665 189.04 13312.945 328.03 ;
      RECT 13312.105 189.04 13312.385 327.79 ;
      RECT 13311.545 189.04 13311.825 327.55 ;
      RECT 13310.985 189.04 13311.265 327.31 ;
      RECT 13310.425 187.94 13310.705 327.07 ;
      RECT 13309.865 189.04 13310.145 326.83 ;
      RECT 13309.305 187.94 13309.585 326.59 ;
      RECT 13308.745 189.04 13309.025 326.35 ;
      RECT 13294.745 187.94 13295.025 332.47 ;
      RECT 13294.185 189.04 13294.465 332.23 ;
      RECT 13293.625 189.04 13293.905 331.99 ;
      RECT 13293.065 189.04 13293.345 331.75 ;
      RECT 13292.505 189.04 13292.785 331.51 ;
      RECT 13291.945 189.04 13292.225 331.27 ;
      RECT 13291.385 189.04 13291.665 331.03 ;
      RECT 13290.825 189.04 13291.105 330.79 ;
      RECT 13290.265 189.04 13290.545 330.55 ;
      RECT 13289.705 187.94 13289.985 330.31 ;
      RECT 13289.145 189.04 13289.425 330.07 ;
      RECT 13288.585 187.94 13288.865 329.83 ;
      RECT 13288.025 189.04 13288.305 329.59 ;
      RECT 13287.465 189.04 13287.745 329.35 ;
      RECT 13286.905 189.04 13287.185 329.11 ;
      RECT 13286.345 189.04 13286.625 328.87 ;
      RECT 13285.785 189.04 13286.065 328.63 ;
      RECT 13285.225 189.04 13285.505 328.39 ;
      RECT 13284.665 189.04 13284.945 328.15 ;
      RECT 13284.105 189.04 13284.385 327.91 ;
      RECT 13283.545 189.04 13283.825 327.67 ;
      RECT 13282.985 189.04 13283.265 327.43 ;
      RECT 13282.425 189.04 13282.705 327.19 ;
      RECT 13243.225 189.04 13243.505 334.095 ;
      RECT 13242.665 189.04 13242.945 334.335 ;
      RECT 13242.105 189.04 13242.385 334.575 ;
      RECT 13241.545 187.94 13241.825 334.815 ;
      RECT 13240.985 189.04 13241.265 335.055 ;
      RECT 13240.425 187.94 13240.705 335.295 ;
      RECT 13239.865 189.04 13240.145 335.535 ;
      RECT 13239.305 189.04 13239.585 335.775 ;
      RECT 13238.745 189.04 13239.025 336.015 ;
      RECT 13238.185 187.94 13238.465 336.255 ;
      RECT 13237.625 189.04 13237.905 336.495 ;
      RECT 13237.065 187.94 13237.345 336.735 ;
      RECT 13236.505 189.04 13236.785 336.975 ;
      RECT 13235.945 187.94 13236.225 337.215 ;
      RECT 13235.385 189.04 13235.665 337.455 ;
      RECT 13234.825 189.04 13235.105 337.695 ;
      RECT 13234.265 189.04 13234.545 337.695 ;
      RECT 13233.705 189.04 13233.985 337.455 ;
      RECT 13233.145 189.04 13233.425 337.215 ;
      RECT 13232.585 189.04 13232.865 336.975 ;
      RECT 13232.025 189.04 13232.305 336.735 ;
      RECT 13231.465 189.04 13231.745 336.495 ;
      RECT 13230.905 189.04 13231.185 336.255 ;
      RECT 13230.345 189.04 13230.625 336.015 ;
      RECT 13229.785 189.04 13230.065 335.775 ;
      RECT 13220.825 189.04 13221.105 335.29 ;
      RECT 13220.265 187.94 13220.545 335.05 ;
      RECT 13219.705 189.04 13219.985 334.81 ;
      RECT 13219.145 187.94 13219.425 334.57 ;
      RECT 13218.585 189.04 13218.865 334.33 ;
      RECT 13218.025 187.94 13218.305 334.09 ;
      RECT 13217.465 189.04 13217.745 333.85 ;
      RECT 13216.905 189.04 13217.185 333.61 ;
      RECT 13216.345 189.04 13216.625 333.37 ;
      RECT 13215.785 189.04 13216.065 333.13 ;
      RECT 13215.225 189.04 13215.505 332.89 ;
      RECT 13214.665 189.04 13214.945 332.65 ;
      RECT 13214.105 189.04 13214.385 332.41 ;
      RECT 13213.545 189.04 13213.825 332.17 ;
      RECT 13211.025 187.94 13211.305 333.89 ;
      RECT 13210.465 189.04 13210.745 333.65 ;
      RECT 13209.905 187.94 13210.185 333.41 ;
      RECT 13209.345 189.04 13209.625 333.17 ;
      RECT 13208.785 189.04 13209.065 332.93 ;
      RECT 13208.225 189.04 13208.505 332.69 ;
      RECT 13207.665 189.04 13207.945 332.45 ;
      RECT 13207.105 189.04 13207.385 332.21 ;
      RECT 13181.065 189.04 13181.345 329.86 ;
      RECT 13180.505 189.04 13180.785 330.1 ;
      RECT 13179.945 189.04 13180.225 330.34 ;
      RECT 13179.385 189.04 13179.665 330.585 ;
      RECT 13178.825 189.04 13179.105 330.825 ;
      RECT 13178.265 189.04 13178.545 331.065 ;
      RECT 13177.705 189.04 13177.985 331.065 ;
      RECT 13177.145 189.04 13177.425 330.825 ;
      RECT 13176.585 189.04 13176.865 330.585 ;
      RECT 13176.025 187.94 13176.305 330.345 ;
      RECT 13175.465 189.04 13175.745 330.105 ;
      RECT 13174.905 187.94 13175.185 329.865 ;
      RECT 13174.345 189.04 13174.625 329.625 ;
      RECT 13173.785 189.04 13174.065 329.385 ;
      RECT 13173.225 189.04 13173.505 329.145 ;
      RECT 13172.665 187.94 13172.945 328.905 ;
      RECT 13172.105 189.04 13172.385 328.665 ;
      RECT 13171.545 187.94 13171.825 328.425 ;
      RECT 13170.985 189.04 13171.265 328.185 ;
      RECT 13170.425 187.94 13170.705 327.945 ;
      RECT 13169.865 189.04 13170.145 327.705 ;
      RECT 13169.305 189.04 13169.585 327.465 ;
      RECT 13168.745 189.04 13169.025 327.225 ;
      RECT 13168.185 189.04 13168.465 326.985 ;
      RECT 13154.745 189.04 13155.025 332.785 ;
      RECT 13154.185 189.04 13154.465 332.545 ;
      RECT 13153.625 189.04 13153.905 332.305 ;
      RECT 13153.065 189.04 13153.345 332.065 ;
      RECT 13152.505 189.04 13152.785 331.825 ;
      RECT 13151.945 189.04 13152.225 331.585 ;
      RECT 13151.385 189.04 13151.665 331.345 ;
      RECT 13150.825 189.04 13151.105 331.105 ;
      RECT 13150.265 187.94 13150.545 330.865 ;
      RECT 13149.705 189.04 13149.985 330.625 ;
      RECT 13149.145 187.94 13149.425 330.305 ;
      RECT 13148.585 189.04 13148.865 330.145 ;
      RECT 13148.025 187.94 13148.305 329.905 ;
      RECT 13147.465 189.04 13147.745 329.665 ;
      RECT 13146.905 189.04 13147.185 329.425 ;
      RECT 13146.345 189.04 13146.625 329.185 ;
      RECT 13145.785 189.04 13146.065 328.945 ;
      RECT 13145.225 189.04 13145.505 328.705 ;
      RECT 13144.665 189.04 13144.945 328.465 ;
      RECT 13144.105 189.04 13144.385 328.225 ;
      RECT 13143.545 189.04 13143.825 327.985 ;
      RECT 13142.985 187.94 13143.265 327.745 ;
      RECT 13142.425 189.04 13142.705 327.505 ;
      RECT 13141.865 187.94 13142.145 327.265 ;
      RECT 13102.665 189.04 13102.945 332.875 ;
      RECT 13102.105 189.04 13102.385 333.115 ;
      RECT 13101.545 189.04 13101.825 333.355 ;
      RECT 13100.985 189.04 13101.265 333.595 ;
      RECT 13100.425 189.04 13100.705 333.835 ;
      RECT 13099.865 189.04 13100.145 334.075 ;
      RECT 13099.305 189.04 13099.585 334.315 ;
      RECT 13098.745 189.04 13099.025 334.555 ;
      RECT 13098.185 189.04 13098.465 334.795 ;
      RECT 13097.625 189.04 13097.905 335.035 ;
      RECT 13097.065 189.04 13097.345 335.275 ;
      RECT 13096.505 189.04 13096.785 335.515 ;
      RECT 13095.945 189.04 13096.225 335.755 ;
      RECT 13095.385 189.04 13095.665 335.755 ;
      RECT 13094.825 187.94 13095.105 335.515 ;
      RECT 13094.265 189.04 13094.545 335.275 ;
      RECT 13093.705 187.94 13093.985 335.035 ;
      RECT 13093.145 189.04 13093.425 334.795 ;
      RECT 13092.585 189.04 13092.865 334.555 ;
      RECT 13092.025 189.04 13092.305 334.315 ;
      RECT 13091.465 187.94 13091.745 334.05 ;
      RECT 13090.905 189.04 13091.185 333.81 ;
      RECT 13090.345 187.94 13090.625 333.57 ;
      RECT 13089.785 189.04 13090.065 333.33 ;
      RECT 13080.825 187.94 13081.105 327.165 ;
      RECT 13080.265 189.04 13080.545 327.405 ;
      RECT 13079.705 189.04 13079.985 327.645 ;
      RECT 13079.145 189.04 13079.425 327.645 ;
      RECT 13078.585 189.04 13078.865 327.405 ;
      RECT 13078.025 189.04 13078.305 327.165 ;
      RECT 13077.465 189.04 13077.745 326.925 ;
      RECT 13076.905 189.04 13077.185 326.685 ;
      RECT 13076.345 189.04 13076.625 326.445 ;
      RECT 13075.785 189.04 13076.065 326.205 ;
      RECT 13075.225 189.04 13075.505 325.965 ;
      RECT 13074.665 189.04 13074.945 325.725 ;
      RECT 13074.105 189.04 13074.385 325.485 ;
      RECT 13073.545 187.94 13073.825 325.245 ;
      RECT 13071.025 189.04 13071.305 326.965 ;
      RECT 13070.465 187.94 13070.745 326.725 ;
      RECT 13069.905 189.04 13070.185 326.485 ;
      RECT 13069.345 187.94 13069.625 326.245 ;
      RECT 13068.785 189.04 13069.065 326.005 ;
      RECT 13068.225 189.04 13068.505 325.765 ;
      RECT 13067.665 189.04 13067.945 325.525 ;
      RECT 13041.625 189.04 13041.905 328.31 ;
      RECT 13041.065 189.04 13041.345 328.55 ;
      RECT 13040.505 189.04 13040.785 328.79 ;
      RECT 13039.945 189.04 13040.225 329.03 ;
      RECT 13039.385 189.04 13039.665 329.27 ;
      RECT 13038.825 187.94 13039.105 329.51 ;
      RECT 13038.265 189.04 13038.545 329.75 ;
      RECT 13037.705 187.94 13037.985 329.99 ;
      RECT 13037.145 189.04 13037.425 330.23 ;
      RECT 13036.585 189.04 13036.865 330.47 ;
      RECT 13036.025 189.04 13036.305 330.71 ;
      RECT 13035.465 189.04 13035.745 330.95 ;
      RECT 13034.905 189.04 13035.185 331.19 ;
      RECT 13034.345 189.04 13034.625 331.43 ;
      RECT 13033.785 189.04 13034.065 331.67 ;
      RECT 13033.225 189.04 13033.505 331.67 ;
      RECT 13032.665 189.04 13032.945 331.43 ;
      RECT 13032.105 189.04 13032.385 331.19 ;
      RECT 13031.545 189.04 13031.825 330.95 ;
      RECT 13030.985 189.04 13031.265 330.705 ;
      RECT 13030.425 189.04 13030.705 330.465 ;
      RECT 13029.865 189.04 13030.145 330.225 ;
      RECT 13029.305 187.94 13029.585 329.985 ;
      RECT 13028.745 189.04 13029.025 329.745 ;
      RECT 13015.305 187.94 13015.585 327.225 ;
      RECT 13014.745 189.04 13015.025 326.985 ;
      RECT 13014.185 189.04 13014.465 326.745 ;
      RECT 13013.625 189.04 13013.905 326.505 ;
      RECT 13013.065 187.94 13013.345 326.265 ;
      RECT 13012.505 189.04 13012.785 326.025 ;
      RECT 13011.945 187.94 13012.225 325.785 ;
      RECT 13011.385 189.04 13011.665 325.545 ;
      RECT 13010.825 187.94 13011.105 325.305 ;
      RECT 13010.265 189.04 13010.545 325.065 ;
      RECT 13009.705 189.04 13009.985 324.825 ;
      RECT 13009.145 189.04 13009.425 324.585 ;
      RECT 13008.585 189.04 13008.865 324.345 ;
      RECT 13008.025 189.04 13008.305 324.105 ;
      RECT 13007.465 189.04 13007.745 323.865 ;
      RECT 13006.905 189.04 13007.185 323.625 ;
      RECT 13006.345 189.04 13006.625 323.385 ;
      RECT 13005.785 189.04 13006.065 323.145 ;
      RECT 13005.225 189.04 13005.505 322.905 ;
      RECT 13004.665 189.04 13004.945 322.665 ;
      RECT 13004.105 189.04 13004.385 322.425 ;
      RECT 13003.545 187.94 13003.825 322.185 ;
      RECT 13002.985 189.04 13003.265 321.945 ;
      RECT 13002.425 187.94 13002.705 321.705 ;
      RECT 12962.665 189.04 12962.945 332.175 ;
      RECT 12962.105 187.94 12962.385 332.415 ;
      RECT 12961.545 189.04 12961.825 332.655 ;
      RECT 12960.985 189.04 12961.265 332.895 ;
      RECT 12960.425 189.04 12960.705 333.135 ;
      RECT 12959.865 189.04 12960.145 333.375 ;
      RECT 12959.305 189.04 12959.585 333.615 ;
      RECT 12958.745 189.04 12959.025 333.86 ;
      RECT 12958.185 189.04 12958.465 334.1 ;
      RECT 12957.625 189.04 12957.905 334.34 ;
      RECT 12957.065 187.94 12957.345 334.58 ;
      RECT 12956.505 189.04 12956.785 334.82 ;
      RECT 12955.945 187.94 12956.225 335.06 ;
      RECT 12955.385 189.04 12955.665 335.3 ;
      RECT 12954.825 189.04 12955.105 335.54 ;
      RECT 12954.265 189.04 12954.545 335.78 ;
      RECT 12953.705 189.04 12953.985 336.02 ;
      RECT 12953.145 189.04 12953.425 336.26 ;
      RECT 12952.585 189.04 12952.865 336.5 ;
      RECT 12952.025 189.04 12952.305 336.74 ;
      RECT 12951.465 189.04 12951.745 336.98 ;
      RECT 12950.905 189.04 12951.185 337.22 ;
      RECT 12950.345 189.04 12950.625 337.46 ;
      RECT 12949.785 189.04 12950.065 337.7 ;
      RECT 12940.825 189.04 12941.105 333.285 ;
      RECT 12940.265 189.04 12940.545 333.045 ;
      RECT 12939.705 189.04 12939.985 332.805 ;
      RECT 12939.145 187.94 12939.425 332.565 ;
      RECT 12938.585 189.04 12938.865 332.325 ;
      RECT 12938.025 187.94 12938.305 332.085 ;
      RECT 12937.465 189.04 12937.745 331.845 ;
      RECT 12936.905 189.04 12937.185 331.605 ;
      RECT 12936.345 189.04 12936.625 331.365 ;
      RECT 12935.785 187.94 12936.065 331.125 ;
      RECT 12935.225 189.04 12935.505 330.885 ;
      RECT 12934.665 187.94 12934.945 330.645 ;
      RECT 12934.105 189.04 12934.385 330.405 ;
      RECT 12933.545 187.94 12933.825 330.165 ;
      RECT 12931.025 189.04 12931.305 322.565 ;
      RECT 12930.465 189.04 12930.745 322.325 ;
      RECT 12929.905 189.04 12930.185 322.085 ;
      RECT 12929.345 189.04 12929.625 321.845 ;
      RECT 12928.785 189.04 12929.065 321.605 ;
      RECT 12928.225 189.04 12928.505 321.365 ;
      RECT 12927.665 189.04 12927.945 321.125 ;
      RECT 12901.625 189.04 12901.905 335 ;
      RECT 12901.065 189.04 12901.345 335.24 ;
      RECT 12900.505 189.04 12900.785 335.48 ;
      RECT 12899.945 189.04 12900.225 335.72 ;
      RECT 12899.385 189.04 12899.665 335.96 ;
      RECT 12898.825 187.94 12899.105 335.96 ;
      RECT 12898.265 189.04 12898.545 335.72 ;
      RECT 12897.705 187.94 12897.985 335.475 ;
      RECT 12897.145 189.04 12897.425 335.235 ;
      RECT 12896.585 187.94 12896.865 334.995 ;
      RECT 12896.025 189.04 12896.305 334.755 ;
      RECT 12895.465 189.04 12895.745 334.515 ;
      RECT 12894.905 189.04 12895.185 334.275 ;
      RECT 12894.345 189.04 12894.625 334.035 ;
      RECT 12893.785 189.04 12894.065 333.795 ;
      RECT 12893.225 189.04 12893.505 333.555 ;
      RECT 12892.665 189.04 12892.945 333.315 ;
      RECT 12892.105 189.04 12892.385 333.075 ;
      RECT 12891.545 187.94 12891.825 332.835 ;
      RECT 12890.985 189.04 12891.265 332.595 ;
      RECT 12890.425 187.94 12890.705 332.355 ;
      RECT 12889.865 189.04 12890.145 332.115 ;
      RECT 12889.305 189.04 12889.585 331.875 ;
      RECT 12888.745 189.04 12889.025 331.635 ;
      RECT 12875.305 189.04 12875.585 335.035 ;
      RECT 12874.745 189.04 12875.025 335.275 ;
      RECT 12874.185 189.04 12874.465 335.52 ;
      RECT 12873.625 189.04 12873.905 335.76 ;
      RECT 12873.065 189.04 12873.345 336 ;
      RECT 12872.505 189.04 12872.785 336 ;
      RECT 12871.945 189.04 12872.225 335.76 ;
      RECT 12871.385 189.04 12871.665 335.52 ;
      RECT 12870.825 189.04 12871.105 328.505 ;
      RECT 12870.265 189.04 12870.545 328.265 ;
      RECT 12869.705 189.04 12869.985 328.025 ;
      RECT 12869.145 187.94 12869.425 327.785 ;
      RECT 12868.585 189.04 12868.865 327.545 ;
      RECT 12868.025 187.94 12868.305 327.305 ;
      RECT 12867.465 189.04 12867.745 327.065 ;
      RECT 12866.905 189.04 12867.185 326.825 ;
      RECT 12866.345 189.04 12866.625 326.585 ;
      RECT 12865.785 187.94 12866.065 326.345 ;
      RECT 12865.225 189.04 12865.505 326.105 ;
      RECT 12864.665 187.94 12864.945 325.865 ;
      RECT 12864.105 189.04 12864.385 325.625 ;
      RECT 12863.545 187.94 12863.825 325.385 ;
      RECT 12862.985 189.04 12863.265 325.145 ;
      RECT 12862.425 189.04 12862.705 324.905 ;
      RECT 12822.105 189.04 12822.385 333.8 ;
      RECT 12821.545 189.04 12821.825 334.04 ;
      RECT 12820.985 189.04 12821.265 334.285 ;
      RECT 12820.425 189.04 12820.705 334.525 ;
      RECT 12819.865 189.04 12820.145 334.765 ;
      RECT 12819.305 189.04 12819.585 335.005 ;
      RECT 12818.745 189.04 12819.025 335.245 ;
      RECT 12818.185 189.04 12818.465 335.485 ;
      RECT 12817.625 189.04 12817.905 335.725 ;
      RECT 12817.065 189.04 12817.345 335.965 ;
      RECT 12816.505 187.94 12816.785 336.205 ;
      RECT 12815.945 189.04 12816.225 336.445 ;
      RECT 12815.385 187.94 12815.665 336.685 ;
      RECT 12814.825 189.04 12815.105 336.925 ;
      RECT 12814.265 187.94 12814.545 337.165 ;
      RECT 12813.705 189.04 12813.985 337.165 ;
      RECT 12813.145 189.04 12813.425 336.925 ;
      RECT 12812.585 189.04 12812.865 336.685 ;
      RECT 12812.025 189.04 12812.305 336.445 ;
      RECT 12811.465 189.04 12811.745 336.205 ;
      RECT 12810.905 189.04 12811.185 335.965 ;
      RECT 12810.345 189.04 12810.625 335.725 ;
      RECT 12809.785 189.04 12810.065 335.485 ;
      RECT 12800.825 187.94 12801.105 335.515 ;
      RECT 12800.265 189.04 12800.545 335.755 ;
      RECT 12799.705 187.94 12799.985 335.995 ;
      RECT 12799.145 189.04 12799.425 336.21 ;
      RECT 12798.585 189.04 12798.865 335.785 ;
      RECT 12798.025 189.04 12798.305 335.545 ;
      RECT 12797.465 189.04 12797.745 335.305 ;
      RECT 12796.905 189.04 12797.185 335.065 ;
      RECT 12796.345 189.04 12796.625 334.825 ;
      RECT 12795.785 189.04 12796.065 334.585 ;
      RECT 12795.225 189.04 12795.505 334.345 ;
      RECT 12794.665 189.04 12794.945 334.105 ;
      RECT 12794.105 189.04 12794.385 333.865 ;
      RECT 12793.545 189.04 12793.825 333.625 ;
      RECT 12791.025 189.04 12791.305 332.8 ;
      RECT 12790.465 189.04 12790.745 332.56 ;
      RECT 12789.905 189.04 12790.185 332.32 ;
      RECT 12789.345 187.94 12789.625 332.08 ;
      RECT 12788.785 189.04 12789.065 331.84 ;
      RECT 12788.225 187.94 12788.505 331.6 ;
      RECT 12787.665 189.04 12787.945 331.36 ;
      RECT 12787.105 189.04 12787.385 331.12 ;
      RECT 12760.505 189.04 12760.785 342.165 ;
      RECT 12759.945 187.94 12760.225 342.405 ;
      RECT 12759.385 189.04 12759.665 342.645 ;
      RECT 12758.825 187.94 12759.105 342.89 ;
      RECT 12758.265 189.04 12758.545 343.13 ;
      RECT 12757.705 187.94 12757.985 343.37 ;
      RECT 12757.145 189.04 12757.425 343.61 ;
      RECT 12756.585 189.04 12756.865 343.85 ;
      RECT 12756.025 189.04 12756.305 329.47 ;
      RECT 12755.465 189.04 12755.745 329.23 ;
      RECT 12754.905 189.04 12755.185 328.99 ;
      RECT 12754.345 189.04 12754.625 328.75 ;
      RECT 12753.785 189.04 12754.065 328.51 ;
      RECT 12753.225 189.04 12753.505 328.27 ;
      RECT 12752.665 189.04 12752.945 328.03 ;
      RECT 12752.105 189.04 12752.385 327.79 ;
      RECT 12751.545 189.04 12751.825 327.55 ;
      RECT 12750.985 189.04 12751.265 327.31 ;
      RECT 12750.425 187.94 12750.705 327.07 ;
      RECT 12749.865 189.04 12750.145 326.83 ;
      RECT 12749.305 187.94 12749.585 326.59 ;
      RECT 12748.745 189.04 12749.025 326.35 ;
      RECT 12734.745 187.94 12735.025 332.47 ;
      RECT 12734.185 189.04 12734.465 332.23 ;
      RECT 12733.625 189.04 12733.905 331.99 ;
      RECT 12733.065 189.04 12733.345 331.75 ;
      RECT 12732.505 189.04 12732.785 331.51 ;
      RECT 12731.945 189.04 12732.225 331.27 ;
      RECT 12731.385 189.04 12731.665 331.03 ;
      RECT 12730.825 189.04 12731.105 330.79 ;
      RECT 12730.265 189.04 12730.545 330.55 ;
      RECT 12729.705 187.94 12729.985 330.31 ;
      RECT 12729.145 189.04 12729.425 330.07 ;
      RECT 12728.585 187.94 12728.865 329.83 ;
      RECT 12728.025 189.04 12728.305 329.59 ;
      RECT 12727.465 189.04 12727.745 329.35 ;
      RECT 12726.905 189.04 12727.185 329.11 ;
      RECT 12726.345 189.04 12726.625 328.87 ;
      RECT 12725.785 189.04 12726.065 328.63 ;
      RECT 12725.225 189.04 12725.505 328.39 ;
      RECT 12724.665 189.04 12724.945 328.15 ;
      RECT 12724.105 189.04 12724.385 327.91 ;
      RECT 12723.545 189.04 12723.825 327.67 ;
      RECT 12722.985 189.04 12723.265 327.43 ;
      RECT 12722.425 189.04 12722.705 327.19 ;
      RECT 12683.225 189.04 12683.505 334.095 ;
      RECT 12682.665 189.04 12682.945 334.335 ;
      RECT 12682.105 189.04 12682.385 334.575 ;
      RECT 12681.545 187.94 12681.825 334.815 ;
      RECT 12680.985 189.04 12681.265 335.055 ;
      RECT 12680.425 187.94 12680.705 335.295 ;
      RECT 12679.865 189.04 12680.145 335.535 ;
      RECT 12679.305 189.04 12679.585 335.775 ;
      RECT 12678.745 189.04 12679.025 336.015 ;
      RECT 12678.185 187.94 12678.465 336.255 ;
      RECT 12677.625 189.04 12677.905 336.495 ;
      RECT 12677.065 187.94 12677.345 336.735 ;
      RECT 12676.505 189.04 12676.785 336.975 ;
      RECT 12675.945 187.94 12676.225 337.215 ;
      RECT 12675.385 189.04 12675.665 337.455 ;
      RECT 12674.825 189.04 12675.105 337.695 ;
      RECT 12674.265 189.04 12674.545 337.695 ;
      RECT 12673.705 189.04 12673.985 337.455 ;
      RECT 12673.145 189.04 12673.425 337.215 ;
      RECT 12672.585 189.04 12672.865 336.975 ;
      RECT 12672.025 189.04 12672.305 336.735 ;
      RECT 12671.465 189.04 12671.745 336.495 ;
      RECT 12670.905 189.04 12671.185 336.255 ;
      RECT 12670.345 189.04 12670.625 336.015 ;
      RECT 12669.785 189.04 12670.065 335.775 ;
      RECT 12660.825 189.04 12661.105 335.29 ;
      RECT 12660.265 187.94 12660.545 335.05 ;
      RECT 12659.705 189.04 12659.985 334.81 ;
      RECT 12659.145 187.94 12659.425 334.57 ;
      RECT 12658.585 189.04 12658.865 334.33 ;
      RECT 12658.025 187.94 12658.305 334.09 ;
      RECT 12657.465 189.04 12657.745 333.85 ;
      RECT 12656.905 189.04 12657.185 333.61 ;
      RECT 12656.345 189.04 12656.625 333.37 ;
      RECT 12655.785 189.04 12656.065 333.13 ;
      RECT 12655.225 189.04 12655.505 332.89 ;
      RECT 12654.665 189.04 12654.945 332.65 ;
      RECT 12654.105 189.04 12654.385 332.41 ;
      RECT 12653.545 189.04 12653.825 332.17 ;
      RECT 12651.025 187.94 12651.305 333.89 ;
      RECT 12650.465 189.04 12650.745 333.65 ;
      RECT 12649.905 187.94 12650.185 333.41 ;
      RECT 12649.345 189.04 12649.625 333.17 ;
      RECT 12648.785 189.04 12649.065 332.93 ;
      RECT 12648.225 189.04 12648.505 332.69 ;
      RECT 12647.665 189.04 12647.945 332.45 ;
      RECT 12647.105 189.04 12647.385 332.21 ;
      RECT 12621.065 189.04 12621.345 329.86 ;
      RECT 12620.505 189.04 12620.785 330.1 ;
      RECT 12619.945 189.04 12620.225 330.34 ;
      RECT 12619.385 189.04 12619.665 330.585 ;
      RECT 12618.825 189.04 12619.105 330.825 ;
      RECT 12618.265 189.04 12618.545 331.065 ;
      RECT 12617.705 189.04 12617.985 331.065 ;
      RECT 12617.145 189.04 12617.425 330.825 ;
      RECT 12616.585 189.04 12616.865 330.585 ;
      RECT 12616.025 187.94 12616.305 330.345 ;
      RECT 12615.465 189.04 12615.745 330.105 ;
      RECT 12614.905 187.94 12615.185 329.865 ;
      RECT 12614.345 189.04 12614.625 329.625 ;
      RECT 12613.785 189.04 12614.065 329.385 ;
      RECT 12613.225 189.04 12613.505 329.145 ;
      RECT 12612.665 187.94 12612.945 328.905 ;
      RECT 12612.105 189.04 12612.385 328.665 ;
      RECT 12611.545 187.94 12611.825 328.425 ;
      RECT 12610.985 189.04 12611.265 328.185 ;
      RECT 12610.425 187.94 12610.705 327.945 ;
      RECT 12609.865 189.04 12610.145 327.705 ;
      RECT 12609.305 189.04 12609.585 327.465 ;
      RECT 12608.745 189.04 12609.025 327.225 ;
      RECT 12608.185 189.04 12608.465 326.985 ;
      RECT 12594.745 189.04 12595.025 332.785 ;
      RECT 12594.185 189.04 12594.465 332.545 ;
      RECT 12593.625 189.04 12593.905 332.305 ;
      RECT 12593.065 189.04 12593.345 332.065 ;
      RECT 12592.505 189.04 12592.785 331.825 ;
      RECT 12591.945 189.04 12592.225 331.585 ;
      RECT 12591.385 189.04 12591.665 331.345 ;
      RECT 12590.825 189.04 12591.105 331.105 ;
      RECT 12590.265 187.94 12590.545 330.865 ;
      RECT 12589.705 189.04 12589.985 330.625 ;
      RECT 12589.145 187.94 12589.425 330.305 ;
      RECT 12588.585 189.04 12588.865 330.145 ;
      RECT 12588.025 187.94 12588.305 329.905 ;
      RECT 12587.465 189.04 12587.745 329.665 ;
      RECT 12586.905 189.04 12587.185 329.425 ;
      RECT 12586.345 189.04 12586.625 329.185 ;
      RECT 12585.785 189.04 12586.065 328.945 ;
      RECT 12585.225 189.04 12585.505 328.705 ;
      RECT 12584.665 189.04 12584.945 328.465 ;
      RECT 12584.105 189.04 12584.385 328.225 ;
      RECT 12583.545 189.04 12583.825 327.985 ;
      RECT 12582.985 187.94 12583.265 327.745 ;
      RECT 12582.425 189.04 12582.705 327.505 ;
      RECT 12581.865 187.94 12582.145 327.265 ;
      RECT 12542.665 189.04 12542.945 332.875 ;
      RECT 12542.105 189.04 12542.385 333.115 ;
      RECT 12541.545 189.04 12541.825 333.355 ;
      RECT 12540.985 189.04 12541.265 333.595 ;
      RECT 12540.425 189.04 12540.705 333.835 ;
      RECT 12539.865 189.04 12540.145 334.075 ;
      RECT 12539.305 189.04 12539.585 334.315 ;
      RECT 12538.745 189.04 12539.025 334.555 ;
      RECT 12538.185 189.04 12538.465 334.795 ;
      RECT 12537.625 189.04 12537.905 335.035 ;
      RECT 12537.065 189.04 12537.345 335.275 ;
      RECT 12536.505 189.04 12536.785 335.515 ;
      RECT 12535.945 189.04 12536.225 335.755 ;
      RECT 12535.385 189.04 12535.665 335.755 ;
      RECT 12534.825 187.94 12535.105 335.515 ;
      RECT 12534.265 189.04 12534.545 335.275 ;
      RECT 12533.705 187.94 12533.985 335.035 ;
      RECT 12533.145 189.04 12533.425 334.795 ;
      RECT 12532.585 189.04 12532.865 334.555 ;
      RECT 12532.025 189.04 12532.305 334.315 ;
      RECT 12531.465 187.94 12531.745 334.05 ;
      RECT 12530.905 189.04 12531.185 333.81 ;
      RECT 12530.345 187.94 12530.625 333.57 ;
      RECT 12529.785 189.04 12530.065 333.33 ;
      RECT 12520.825 187.94 12521.105 327.165 ;
      RECT 12520.265 189.04 12520.545 327.405 ;
      RECT 12519.705 189.04 12519.985 327.645 ;
      RECT 12519.145 189.04 12519.425 327.645 ;
      RECT 12518.585 189.04 12518.865 327.405 ;
      RECT 12518.025 189.04 12518.305 327.165 ;
      RECT 12517.465 189.04 12517.745 326.925 ;
      RECT 12516.905 189.04 12517.185 326.685 ;
      RECT 12516.345 189.04 12516.625 326.445 ;
      RECT 12515.785 189.04 12516.065 326.205 ;
      RECT 12515.225 189.04 12515.505 325.965 ;
      RECT 12514.665 189.04 12514.945 325.725 ;
      RECT 12514.105 189.04 12514.385 325.485 ;
      RECT 12513.545 187.94 12513.825 325.245 ;
      RECT 12511.025 189.04 12511.305 326.965 ;
      RECT 12510.465 187.94 12510.745 326.725 ;
      RECT 12509.905 189.04 12510.185 326.485 ;
      RECT 12509.345 187.94 12509.625 326.245 ;
      RECT 12508.785 189.04 12509.065 326.005 ;
      RECT 12508.225 189.04 12508.505 325.765 ;
      RECT 12507.665 189.04 12507.945 325.525 ;
      RECT 12481.625 189.04 12481.905 328.31 ;
      RECT 12481.065 189.04 12481.345 328.55 ;
      RECT 12480.505 189.04 12480.785 328.79 ;
      RECT 12479.945 189.04 12480.225 329.03 ;
      RECT 12479.385 189.04 12479.665 329.27 ;
      RECT 12478.825 187.94 12479.105 329.51 ;
      RECT 12478.265 189.04 12478.545 329.75 ;
      RECT 12477.705 187.94 12477.985 329.99 ;
      RECT 12477.145 189.04 12477.425 330.23 ;
      RECT 12476.585 189.04 12476.865 330.47 ;
      RECT 12476.025 189.04 12476.305 330.71 ;
      RECT 12475.465 189.04 12475.745 330.95 ;
      RECT 12474.905 189.04 12475.185 331.19 ;
      RECT 12474.345 189.04 12474.625 331.43 ;
      RECT 12473.785 189.04 12474.065 331.67 ;
      RECT 12473.225 189.04 12473.505 331.67 ;
      RECT 12472.665 189.04 12472.945 331.43 ;
      RECT 12472.105 189.04 12472.385 331.19 ;
      RECT 12471.545 189.04 12471.825 330.95 ;
      RECT 12470.985 189.04 12471.265 330.705 ;
      RECT 12470.425 189.04 12470.705 330.465 ;
      RECT 12469.865 189.04 12470.145 330.225 ;
      RECT 12469.305 187.94 12469.585 329.985 ;
      RECT 12468.745 189.04 12469.025 329.745 ;
      RECT 12455.305 187.94 12455.585 327.225 ;
      RECT 12454.745 189.04 12455.025 326.985 ;
      RECT 12454.185 189.04 12454.465 326.745 ;
      RECT 12453.625 189.04 12453.905 326.505 ;
      RECT 12453.065 187.94 12453.345 326.265 ;
      RECT 12452.505 189.04 12452.785 326.025 ;
      RECT 12451.945 187.94 12452.225 325.785 ;
      RECT 12451.385 189.04 12451.665 325.545 ;
      RECT 12450.825 187.94 12451.105 325.305 ;
      RECT 12450.265 189.04 12450.545 325.065 ;
      RECT 12449.705 189.04 12449.985 324.825 ;
      RECT 12449.145 189.04 12449.425 324.585 ;
      RECT 12448.585 189.04 12448.865 324.345 ;
      RECT 12448.025 189.04 12448.305 324.105 ;
      RECT 12447.465 189.04 12447.745 323.865 ;
      RECT 12446.905 189.04 12447.185 323.625 ;
      RECT 12446.345 189.04 12446.625 323.385 ;
      RECT 12445.785 189.04 12446.065 323.145 ;
      RECT 12445.225 189.04 12445.505 322.905 ;
      RECT 12444.665 189.04 12444.945 322.665 ;
      RECT 12444.105 189.04 12444.385 322.425 ;
      RECT 12443.545 187.94 12443.825 322.185 ;
      RECT 12442.985 189.04 12443.265 321.945 ;
      RECT 12442.425 187.94 12442.705 321.705 ;
      RECT 12402.665 189.04 12402.945 332.175 ;
      RECT 12402.105 187.94 12402.385 332.415 ;
      RECT 12401.545 189.04 12401.825 332.655 ;
      RECT 12400.985 189.04 12401.265 332.895 ;
      RECT 12400.425 189.04 12400.705 333.135 ;
      RECT 12399.865 189.04 12400.145 333.375 ;
      RECT 12399.305 189.04 12399.585 333.615 ;
      RECT 12398.745 189.04 12399.025 333.86 ;
      RECT 12398.185 189.04 12398.465 334.1 ;
      RECT 12397.625 189.04 12397.905 334.34 ;
      RECT 12397.065 187.94 12397.345 334.58 ;
      RECT 12396.505 189.04 12396.785 334.82 ;
      RECT 12395.945 187.94 12396.225 335.06 ;
      RECT 12395.385 189.04 12395.665 335.3 ;
      RECT 12394.825 189.04 12395.105 335.54 ;
      RECT 12394.265 189.04 12394.545 335.78 ;
      RECT 12393.705 189.04 12393.985 336.02 ;
      RECT 12393.145 189.04 12393.425 336.26 ;
      RECT 12392.585 189.04 12392.865 336.5 ;
      RECT 12392.025 189.04 12392.305 336.74 ;
      RECT 12391.465 189.04 12391.745 336.98 ;
      RECT 12390.905 189.04 12391.185 337.22 ;
      RECT 12390.345 189.04 12390.625 337.46 ;
      RECT 12389.785 189.04 12390.065 337.7 ;
      RECT 12380.825 189.04 12381.105 333.285 ;
      RECT 12380.265 189.04 12380.545 333.045 ;
      RECT 12379.705 189.04 12379.985 332.805 ;
      RECT 12379.145 187.94 12379.425 332.565 ;
      RECT 12378.585 189.04 12378.865 332.325 ;
      RECT 12378.025 187.94 12378.305 332.085 ;
      RECT 12377.465 189.04 12377.745 331.845 ;
      RECT 12376.905 189.04 12377.185 331.605 ;
      RECT 12376.345 189.04 12376.625 331.365 ;
      RECT 12375.785 187.94 12376.065 331.125 ;
      RECT 12375.225 189.04 12375.505 330.885 ;
      RECT 12374.665 187.94 12374.945 330.645 ;
      RECT 12374.105 189.04 12374.385 330.405 ;
      RECT 12373.545 187.94 12373.825 330.165 ;
      RECT 12371.025 189.04 12371.305 322.565 ;
      RECT 12370.465 189.04 12370.745 322.325 ;
      RECT 12369.905 189.04 12370.185 322.085 ;
      RECT 12369.345 189.04 12369.625 321.845 ;
      RECT 12368.785 189.04 12369.065 321.605 ;
      RECT 12368.225 189.04 12368.505 321.365 ;
      RECT 12367.665 189.04 12367.945 321.125 ;
      RECT 12341.625 189.04 12341.905 335 ;
      RECT 12341.065 189.04 12341.345 335.24 ;
      RECT 12340.505 189.04 12340.785 335.48 ;
      RECT 12339.945 189.04 12340.225 335.72 ;
      RECT 12339.385 189.04 12339.665 335.96 ;
      RECT 12338.825 187.94 12339.105 335.96 ;
      RECT 12338.265 189.04 12338.545 335.72 ;
      RECT 12337.705 187.94 12337.985 335.475 ;
      RECT 12337.145 189.04 12337.425 335.235 ;
      RECT 12336.585 187.94 12336.865 334.995 ;
      RECT 12336.025 189.04 12336.305 334.755 ;
      RECT 12335.465 189.04 12335.745 334.515 ;
      RECT 12334.905 189.04 12335.185 334.275 ;
      RECT 12334.345 189.04 12334.625 334.035 ;
      RECT 12333.785 189.04 12334.065 333.795 ;
      RECT 12333.225 189.04 12333.505 333.555 ;
      RECT 12332.665 189.04 12332.945 333.315 ;
      RECT 12332.105 189.04 12332.385 333.075 ;
      RECT 12331.545 187.94 12331.825 332.835 ;
      RECT 12330.985 189.04 12331.265 332.595 ;
      RECT 12330.425 187.94 12330.705 332.355 ;
      RECT 12329.865 189.04 12330.145 332.115 ;
      RECT 12329.305 189.04 12329.585 331.875 ;
      RECT 12328.745 189.04 12329.025 331.635 ;
      RECT 12315.305 189.04 12315.585 335.035 ;
      RECT 12314.745 189.04 12315.025 335.275 ;
      RECT 12314.185 189.04 12314.465 335.52 ;
      RECT 12313.625 189.04 12313.905 335.76 ;
      RECT 12313.065 189.04 12313.345 336 ;
      RECT 12312.505 189.04 12312.785 336 ;
      RECT 12311.945 189.04 12312.225 335.76 ;
      RECT 12311.385 189.04 12311.665 335.52 ;
      RECT 12310.825 189.04 12311.105 328.505 ;
      RECT 12310.265 189.04 12310.545 328.265 ;
      RECT 12309.705 189.04 12309.985 328.025 ;
      RECT 12309.145 187.94 12309.425 327.785 ;
      RECT 12308.585 189.04 12308.865 327.545 ;
      RECT 12308.025 187.94 12308.305 327.305 ;
      RECT 12307.465 189.04 12307.745 327.065 ;
      RECT 12306.905 189.04 12307.185 326.825 ;
      RECT 12306.345 189.04 12306.625 326.585 ;
      RECT 12305.785 187.94 12306.065 326.345 ;
      RECT 12305.225 189.04 12305.505 326.105 ;
      RECT 12304.665 187.94 12304.945 325.865 ;
      RECT 12304.105 189.04 12304.385 325.625 ;
      RECT 12303.545 187.94 12303.825 325.385 ;
      RECT 12302.985 189.04 12303.265 325.145 ;
      RECT 12302.425 189.04 12302.705 324.905 ;
      RECT 12262.105 189.04 12262.385 333.8 ;
      RECT 12261.545 189.04 12261.825 334.04 ;
      RECT 12260.985 189.04 12261.265 334.285 ;
      RECT 12260.425 189.04 12260.705 334.525 ;
      RECT 12259.865 189.04 12260.145 334.765 ;
      RECT 12259.305 189.04 12259.585 335.005 ;
      RECT 12258.745 189.04 12259.025 335.245 ;
      RECT 12258.185 189.04 12258.465 335.485 ;
      RECT 12257.625 189.04 12257.905 335.725 ;
      RECT 12257.065 189.04 12257.345 335.965 ;
      RECT 12256.505 187.94 12256.785 336.205 ;
      RECT 12255.945 189.04 12256.225 336.445 ;
      RECT 12255.385 187.94 12255.665 336.685 ;
      RECT 12254.825 189.04 12255.105 336.925 ;
      RECT 12254.265 187.94 12254.545 337.165 ;
      RECT 12253.705 189.04 12253.985 337.165 ;
      RECT 12253.145 189.04 12253.425 336.925 ;
      RECT 12252.585 189.04 12252.865 336.685 ;
      RECT 12252.025 189.04 12252.305 336.445 ;
      RECT 12251.465 189.04 12251.745 336.205 ;
      RECT 12250.905 189.04 12251.185 335.965 ;
      RECT 12250.345 189.04 12250.625 335.725 ;
      RECT 12249.785 189.04 12250.065 335.485 ;
      RECT 12240.825 187.94 12241.105 335.515 ;
      RECT 12240.265 189.04 12240.545 335.755 ;
      RECT 12239.705 187.94 12239.985 335.995 ;
      RECT 12239.145 189.04 12239.425 336.21 ;
      RECT 12238.585 189.04 12238.865 335.785 ;
      RECT 12238.025 189.04 12238.305 335.545 ;
      RECT 12237.465 189.04 12237.745 335.305 ;
      RECT 12236.905 189.04 12237.185 335.065 ;
      RECT 12236.345 189.04 12236.625 334.825 ;
      RECT 12235.785 189.04 12236.065 334.585 ;
      RECT 12235.225 189.04 12235.505 334.345 ;
      RECT 12234.665 189.04 12234.945 334.105 ;
      RECT 12234.105 189.04 12234.385 333.865 ;
      RECT 12233.545 189.04 12233.825 333.625 ;
      RECT 12231.025 189.04 12231.305 332.8 ;
      RECT 12230.465 189.04 12230.745 332.56 ;
      RECT 12229.905 189.04 12230.185 332.32 ;
      RECT 12229.345 187.94 12229.625 332.08 ;
      RECT 12228.785 189.04 12229.065 331.84 ;
      RECT 12228.225 187.94 12228.505 331.6 ;
      RECT 12227.665 189.04 12227.945 331.36 ;
      RECT 12227.105 189.04 12227.385 331.12 ;
      RECT 12200.505 189.04 12200.785 342.165 ;
      RECT 12199.945 187.94 12200.225 342.405 ;
      RECT 12199.385 189.04 12199.665 342.645 ;
      RECT 12198.825 187.94 12199.105 342.89 ;
      RECT 12198.265 189.04 12198.545 343.13 ;
      RECT 12197.705 187.94 12197.985 343.37 ;
      RECT 12197.145 189.04 12197.425 343.61 ;
      RECT 12196.585 189.04 12196.865 343.85 ;
      RECT 12196.025 189.04 12196.305 329.47 ;
      RECT 12195.465 189.04 12195.745 329.23 ;
      RECT 12194.905 189.04 12195.185 328.99 ;
      RECT 12194.345 189.04 12194.625 328.75 ;
      RECT 12193.785 189.04 12194.065 328.51 ;
      RECT 12193.225 189.04 12193.505 328.27 ;
      RECT 12192.665 189.04 12192.945 328.03 ;
      RECT 12192.105 189.04 12192.385 327.79 ;
      RECT 12191.545 189.04 12191.825 327.55 ;
      RECT 12190.985 189.04 12191.265 327.31 ;
      RECT 12190.425 187.94 12190.705 327.07 ;
      RECT 12189.865 189.04 12190.145 326.83 ;
      RECT 12189.305 187.94 12189.585 326.59 ;
      RECT 12188.745 189.04 12189.025 326.35 ;
      RECT 12174.745 187.94 12175.025 332.47 ;
      RECT 12174.185 189.04 12174.465 332.23 ;
      RECT 12173.625 189.04 12173.905 331.99 ;
      RECT 12173.065 189.04 12173.345 331.75 ;
      RECT 12172.505 189.04 12172.785 331.51 ;
      RECT 12171.945 189.04 12172.225 331.27 ;
      RECT 12171.385 189.04 12171.665 331.03 ;
      RECT 12170.825 189.04 12171.105 330.79 ;
      RECT 12170.265 189.04 12170.545 330.55 ;
      RECT 12169.705 187.94 12169.985 330.31 ;
      RECT 12169.145 189.04 12169.425 330.07 ;
      RECT 12168.585 187.94 12168.865 329.83 ;
      RECT 12168.025 189.04 12168.305 329.59 ;
      RECT 12167.465 189.04 12167.745 329.35 ;
      RECT 12166.905 189.04 12167.185 329.11 ;
      RECT 12166.345 189.04 12166.625 328.87 ;
      RECT 12165.785 189.04 12166.065 328.63 ;
      RECT 12165.225 189.04 12165.505 328.39 ;
      RECT 12164.665 189.04 12164.945 328.15 ;
      RECT 12164.105 189.04 12164.385 327.91 ;
      RECT 12163.545 189.04 12163.825 327.67 ;
      RECT 12162.985 189.04 12163.265 327.43 ;
      RECT 12162.425 189.04 12162.705 327.19 ;
      RECT 12123.225 189.04 12123.505 334.095 ;
      RECT 12122.665 189.04 12122.945 334.335 ;
      RECT 12122.105 189.04 12122.385 334.575 ;
      RECT 12121.545 187.94 12121.825 334.815 ;
      RECT 12120.985 189.04 12121.265 335.055 ;
      RECT 12120.425 187.94 12120.705 335.295 ;
      RECT 12119.865 189.04 12120.145 335.535 ;
      RECT 12119.305 189.04 12119.585 335.775 ;
      RECT 12118.745 189.04 12119.025 336.015 ;
      RECT 12118.185 187.94 12118.465 336.255 ;
      RECT 12117.625 189.04 12117.905 336.495 ;
      RECT 12117.065 187.94 12117.345 336.735 ;
      RECT 12116.505 189.04 12116.785 336.975 ;
      RECT 12115.945 187.94 12116.225 337.215 ;
      RECT 12115.385 189.04 12115.665 337.455 ;
      RECT 12114.825 189.04 12115.105 337.695 ;
      RECT 12114.265 189.04 12114.545 337.695 ;
      RECT 12113.705 189.04 12113.985 337.455 ;
      RECT 12113.145 189.04 12113.425 337.215 ;
      RECT 12112.585 189.04 12112.865 336.975 ;
      RECT 12112.025 189.04 12112.305 336.735 ;
      RECT 12111.465 189.04 12111.745 336.495 ;
      RECT 12110.905 189.04 12111.185 336.255 ;
      RECT 12110.345 189.04 12110.625 336.015 ;
      RECT 12109.785 189.04 12110.065 335.775 ;
      RECT 12100.825 189.04 12101.105 335.29 ;
      RECT 12100.265 187.94 12100.545 335.05 ;
      RECT 12099.705 189.04 12099.985 334.81 ;
      RECT 12099.145 187.94 12099.425 334.57 ;
      RECT 12098.585 189.04 12098.865 334.33 ;
      RECT 12098.025 187.94 12098.305 334.09 ;
      RECT 12097.465 189.04 12097.745 333.85 ;
      RECT 12096.905 189.04 12097.185 333.61 ;
      RECT 12096.345 189.04 12096.625 333.37 ;
      RECT 12095.785 189.04 12096.065 333.13 ;
      RECT 12095.225 189.04 12095.505 332.89 ;
      RECT 12094.665 189.04 12094.945 332.65 ;
      RECT 12094.105 189.04 12094.385 332.41 ;
      RECT 12093.545 189.04 12093.825 332.17 ;
      RECT 12091.025 187.94 12091.305 333.89 ;
      RECT 12090.465 189.04 12090.745 333.65 ;
      RECT 12089.905 187.94 12090.185 333.41 ;
      RECT 12089.345 189.04 12089.625 333.17 ;
      RECT 12088.785 189.04 12089.065 332.93 ;
      RECT 12088.225 189.04 12088.505 332.69 ;
      RECT 12087.665 189.04 12087.945 332.45 ;
      RECT 12087.105 189.04 12087.385 332.21 ;
      RECT 12061.065 189.04 12061.345 329.86 ;
      RECT 12060.505 189.04 12060.785 330.1 ;
      RECT 12059.945 189.04 12060.225 330.34 ;
      RECT 12059.385 189.04 12059.665 330.585 ;
      RECT 12058.825 189.04 12059.105 330.825 ;
      RECT 12058.265 189.04 12058.545 331.065 ;
      RECT 12057.705 189.04 12057.985 331.065 ;
      RECT 12057.145 189.04 12057.425 330.825 ;
      RECT 12056.585 189.04 12056.865 330.585 ;
      RECT 12056.025 187.94 12056.305 330.345 ;
      RECT 12055.465 189.04 12055.745 330.105 ;
      RECT 12054.905 187.94 12055.185 329.865 ;
      RECT 12054.345 189.04 12054.625 329.625 ;
      RECT 12053.785 189.04 12054.065 329.385 ;
      RECT 12053.225 189.04 12053.505 329.145 ;
      RECT 12052.665 187.94 12052.945 328.905 ;
      RECT 12052.105 189.04 12052.385 328.665 ;
      RECT 12051.545 187.94 12051.825 328.425 ;
      RECT 12050.985 189.04 12051.265 328.185 ;
      RECT 12050.425 187.94 12050.705 327.945 ;
      RECT 12049.865 189.04 12050.145 327.705 ;
      RECT 12049.305 189.04 12049.585 327.465 ;
      RECT 12048.745 189.04 12049.025 327.225 ;
      RECT 12048.185 189.04 12048.465 326.985 ;
      RECT 12034.745 189.04 12035.025 332.785 ;
      RECT 12034.185 189.04 12034.465 332.545 ;
      RECT 12033.625 189.04 12033.905 332.305 ;
      RECT 12033.065 189.04 12033.345 332.065 ;
      RECT 12032.505 189.04 12032.785 331.825 ;
      RECT 12031.945 189.04 12032.225 331.585 ;
      RECT 12031.385 189.04 12031.665 331.345 ;
      RECT 12030.825 189.04 12031.105 331.105 ;
      RECT 12030.265 187.94 12030.545 330.865 ;
      RECT 12029.705 189.04 12029.985 330.625 ;
      RECT 12029.145 187.94 12029.425 330.305 ;
      RECT 12028.585 189.04 12028.865 330.145 ;
      RECT 12028.025 187.94 12028.305 329.905 ;
      RECT 12027.465 189.04 12027.745 329.665 ;
      RECT 12026.905 189.04 12027.185 329.425 ;
      RECT 12026.345 189.04 12026.625 329.185 ;
      RECT 12025.785 189.04 12026.065 328.945 ;
      RECT 12025.225 189.04 12025.505 328.705 ;
      RECT 12024.665 189.04 12024.945 328.465 ;
      RECT 12024.105 189.04 12024.385 328.225 ;
      RECT 12023.545 189.04 12023.825 327.985 ;
      RECT 12022.985 187.94 12023.265 327.745 ;
      RECT 12022.425 189.04 12022.705 327.505 ;
      RECT 12021.865 187.94 12022.145 327.265 ;
      RECT 11982.665 189.04 11982.945 332.875 ;
      RECT 11982.105 189.04 11982.385 333.115 ;
      RECT 11981.545 189.04 11981.825 333.355 ;
      RECT 11980.985 189.04 11981.265 333.595 ;
      RECT 11980.425 189.04 11980.705 333.835 ;
      RECT 11979.865 189.04 11980.145 334.075 ;
      RECT 11979.305 189.04 11979.585 334.315 ;
      RECT 11978.745 189.04 11979.025 334.555 ;
      RECT 11978.185 189.04 11978.465 334.795 ;
      RECT 11977.625 189.04 11977.905 335.035 ;
      RECT 11977.065 189.04 11977.345 335.275 ;
      RECT 11976.505 189.04 11976.785 335.515 ;
      RECT 11975.945 189.04 11976.225 335.755 ;
      RECT 11975.385 189.04 11975.665 335.755 ;
      RECT 11974.825 187.94 11975.105 335.515 ;
      RECT 11974.265 189.04 11974.545 335.275 ;
      RECT 11973.705 187.94 11973.985 335.035 ;
      RECT 11973.145 189.04 11973.425 334.795 ;
      RECT 11972.585 189.04 11972.865 334.555 ;
      RECT 11972.025 189.04 11972.305 334.315 ;
      RECT 11971.465 187.94 11971.745 334.05 ;
      RECT 11970.905 189.04 11971.185 333.81 ;
      RECT 11970.345 187.94 11970.625 333.57 ;
      RECT 11969.785 189.04 11970.065 333.33 ;
      RECT 11960.825 187.94 11961.105 327.165 ;
      RECT 11960.265 189.04 11960.545 327.405 ;
      RECT 11959.705 189.04 11959.985 327.645 ;
      RECT 11959.145 189.04 11959.425 327.645 ;
      RECT 11958.585 189.04 11958.865 327.405 ;
      RECT 11958.025 189.04 11958.305 327.165 ;
      RECT 11957.465 189.04 11957.745 326.925 ;
      RECT 11956.905 189.04 11957.185 326.685 ;
      RECT 11956.345 189.04 11956.625 326.445 ;
      RECT 11955.785 189.04 11956.065 326.205 ;
      RECT 11955.225 189.04 11955.505 325.965 ;
      RECT 11954.665 189.04 11954.945 325.725 ;
      RECT 11954.105 189.04 11954.385 325.485 ;
      RECT 11953.545 187.94 11953.825 325.245 ;
      RECT 11951.025 189.04 11951.305 326.965 ;
      RECT 11950.465 187.94 11950.745 326.725 ;
      RECT 11949.905 189.04 11950.185 326.485 ;
      RECT 11949.345 187.94 11949.625 326.245 ;
      RECT 11948.785 189.04 11949.065 326.005 ;
      RECT 11948.225 189.04 11948.505 325.765 ;
      RECT 11947.665 189.04 11947.945 325.525 ;
      RECT 11921.625 189.04 11921.905 328.31 ;
      RECT 11921.065 189.04 11921.345 328.55 ;
      RECT 11920.505 189.04 11920.785 328.79 ;
      RECT 11919.945 189.04 11920.225 329.03 ;
      RECT 11919.385 189.04 11919.665 329.27 ;
      RECT 11918.825 187.94 11919.105 329.51 ;
      RECT 11918.265 189.04 11918.545 329.75 ;
      RECT 11917.705 187.94 11917.985 329.99 ;
      RECT 11917.145 189.04 11917.425 330.23 ;
      RECT 11916.585 189.04 11916.865 330.47 ;
      RECT 11916.025 189.04 11916.305 330.71 ;
      RECT 11915.465 189.04 11915.745 330.95 ;
      RECT 11914.905 189.04 11915.185 331.19 ;
      RECT 11914.345 189.04 11914.625 331.43 ;
      RECT 11913.785 189.04 11914.065 331.67 ;
      RECT 11913.225 189.04 11913.505 331.67 ;
      RECT 11912.665 189.04 11912.945 331.43 ;
      RECT 11912.105 189.04 11912.385 331.19 ;
      RECT 11911.545 189.04 11911.825 330.95 ;
      RECT 11910.985 189.04 11911.265 330.705 ;
      RECT 11910.425 189.04 11910.705 330.465 ;
      RECT 11909.865 189.04 11910.145 330.225 ;
      RECT 11909.305 187.94 11909.585 329.985 ;
      RECT 11908.745 189.04 11909.025 329.745 ;
      RECT 11895.305 187.94 11895.585 327.225 ;
      RECT 11894.745 189.04 11895.025 326.985 ;
      RECT 11894.185 189.04 11894.465 326.745 ;
      RECT 11893.625 189.04 11893.905 326.505 ;
      RECT 11893.065 187.94 11893.345 326.265 ;
      RECT 11892.505 189.04 11892.785 326.025 ;
      RECT 11891.945 187.94 11892.225 325.785 ;
      RECT 11891.385 189.04 11891.665 325.545 ;
      RECT 11890.825 187.94 11891.105 325.305 ;
      RECT 11890.265 189.04 11890.545 325.065 ;
      RECT 11889.705 189.04 11889.985 324.825 ;
      RECT 11889.145 189.04 11889.425 324.585 ;
      RECT 11888.585 189.04 11888.865 324.345 ;
      RECT 11888.025 189.04 11888.305 324.105 ;
      RECT 11887.465 189.04 11887.745 323.865 ;
      RECT 11886.905 189.04 11887.185 323.625 ;
      RECT 11886.345 189.04 11886.625 323.385 ;
      RECT 11885.785 189.04 11886.065 323.145 ;
      RECT 11885.225 189.04 11885.505 322.905 ;
      RECT 11884.665 189.04 11884.945 322.665 ;
      RECT 11884.105 189.04 11884.385 322.425 ;
      RECT 11883.545 187.94 11883.825 322.185 ;
      RECT 11882.985 189.04 11883.265 321.945 ;
      RECT 11882.425 187.94 11882.705 321.705 ;
      RECT 11842.665 189.04 11842.945 332.175 ;
      RECT 11842.105 187.94 11842.385 332.415 ;
      RECT 11841.545 189.04 11841.825 332.655 ;
      RECT 11840.985 189.04 11841.265 332.895 ;
      RECT 11840.425 189.04 11840.705 333.135 ;
      RECT 11839.865 189.04 11840.145 333.375 ;
      RECT 11839.305 189.04 11839.585 333.615 ;
      RECT 11838.745 189.04 11839.025 333.86 ;
      RECT 11838.185 189.04 11838.465 334.1 ;
      RECT 11837.625 189.04 11837.905 334.34 ;
      RECT 11837.065 187.94 11837.345 334.58 ;
      RECT 11836.505 189.04 11836.785 334.82 ;
      RECT 11835.945 187.94 11836.225 335.06 ;
      RECT 11835.385 189.04 11835.665 335.3 ;
      RECT 11834.825 189.04 11835.105 335.54 ;
      RECT 11834.265 189.04 11834.545 335.78 ;
      RECT 11833.705 189.04 11833.985 336.02 ;
      RECT 11833.145 189.04 11833.425 336.26 ;
      RECT 11832.585 189.04 11832.865 336.5 ;
      RECT 11832.025 189.04 11832.305 336.74 ;
      RECT 11831.465 189.04 11831.745 336.98 ;
      RECT 11830.905 189.04 11831.185 337.22 ;
      RECT 11830.345 189.04 11830.625 337.46 ;
      RECT 11829.785 189.04 11830.065 337.7 ;
      RECT 11820.825 189.04 11821.105 333.285 ;
      RECT 11820.265 189.04 11820.545 333.045 ;
      RECT 11819.705 189.04 11819.985 332.805 ;
      RECT 11819.145 187.94 11819.425 332.565 ;
      RECT 11818.585 189.04 11818.865 332.325 ;
      RECT 11818.025 187.94 11818.305 332.085 ;
      RECT 11817.465 189.04 11817.745 331.845 ;
      RECT 11816.905 189.04 11817.185 331.605 ;
      RECT 11816.345 189.04 11816.625 331.365 ;
      RECT 11815.785 187.94 11816.065 331.125 ;
      RECT 11815.225 189.04 11815.505 330.885 ;
      RECT 11814.665 187.94 11814.945 330.645 ;
      RECT 11814.105 189.04 11814.385 330.405 ;
      RECT 11813.545 187.94 11813.825 330.165 ;
      RECT 11811.025 189.04 11811.305 322.565 ;
      RECT 11810.465 189.04 11810.745 322.325 ;
      RECT 11809.905 189.04 11810.185 322.085 ;
      RECT 11809.345 189.04 11809.625 321.845 ;
      RECT 11808.785 189.04 11809.065 321.605 ;
      RECT 11808.225 189.04 11808.505 321.365 ;
      RECT 11807.665 189.04 11807.945 321.125 ;
      RECT 11781.625 189.04 11781.905 335 ;
      RECT 11781.065 189.04 11781.345 335.24 ;
      RECT 11780.505 189.04 11780.785 335.48 ;
      RECT 11779.945 189.04 11780.225 335.72 ;
      RECT 11779.385 189.04 11779.665 335.96 ;
      RECT 11778.825 187.94 11779.105 335.96 ;
      RECT 11778.265 189.04 11778.545 335.72 ;
      RECT 11777.705 187.94 11777.985 335.475 ;
      RECT 11777.145 189.04 11777.425 335.235 ;
      RECT 11776.585 187.94 11776.865 334.995 ;
      RECT 11776.025 189.04 11776.305 334.755 ;
      RECT 11775.465 189.04 11775.745 334.515 ;
      RECT 11774.905 189.04 11775.185 334.275 ;
      RECT 11774.345 189.04 11774.625 334.035 ;
      RECT 11773.785 189.04 11774.065 333.795 ;
      RECT 11773.225 189.04 11773.505 333.555 ;
      RECT 11772.665 189.04 11772.945 333.315 ;
      RECT 11772.105 189.04 11772.385 333.075 ;
      RECT 11771.545 187.94 11771.825 332.835 ;
      RECT 11770.985 189.04 11771.265 332.595 ;
      RECT 11770.425 187.94 11770.705 332.355 ;
      RECT 11769.865 189.04 11770.145 332.115 ;
      RECT 11769.305 189.04 11769.585 331.875 ;
      RECT 11768.745 189.04 11769.025 331.635 ;
      RECT 11755.305 189.04 11755.585 335.035 ;
      RECT 11754.745 189.04 11755.025 335.275 ;
      RECT 11754.185 189.04 11754.465 335.52 ;
      RECT 11753.625 189.04 11753.905 335.76 ;
      RECT 11753.065 189.04 11753.345 336 ;
      RECT 11752.505 189.04 11752.785 336 ;
      RECT 11751.945 189.04 11752.225 335.76 ;
      RECT 11751.385 189.04 11751.665 335.52 ;
      RECT 11750.825 189.04 11751.105 328.505 ;
      RECT 11750.265 189.04 11750.545 328.265 ;
      RECT 11749.705 189.04 11749.985 328.025 ;
      RECT 11749.145 187.94 11749.425 327.785 ;
      RECT 11748.585 189.04 11748.865 327.545 ;
      RECT 11748.025 187.94 11748.305 327.305 ;
      RECT 11747.465 189.04 11747.745 327.065 ;
      RECT 11746.905 189.04 11747.185 326.825 ;
      RECT 11746.345 189.04 11746.625 326.585 ;
      RECT 11745.785 187.94 11746.065 326.345 ;
      RECT 11745.225 189.04 11745.505 326.105 ;
      RECT 11744.665 187.94 11744.945 325.865 ;
      RECT 11744.105 189.04 11744.385 325.625 ;
      RECT 11743.545 187.94 11743.825 325.385 ;
      RECT 11742.985 189.04 11743.265 325.145 ;
      RECT 11742.425 189.04 11742.705 324.905 ;
      RECT 11702.105 189.04 11702.385 333.8 ;
      RECT 11701.545 189.04 11701.825 334.04 ;
      RECT 11700.985 189.04 11701.265 334.285 ;
      RECT 11700.425 189.04 11700.705 334.525 ;
      RECT 11699.865 189.04 11700.145 334.765 ;
      RECT 11699.305 189.04 11699.585 335.005 ;
      RECT 11698.745 189.04 11699.025 335.245 ;
      RECT 11698.185 189.04 11698.465 335.485 ;
      RECT 11697.625 189.04 11697.905 335.725 ;
      RECT 11697.065 189.04 11697.345 335.965 ;
      RECT 11696.505 187.94 11696.785 336.205 ;
      RECT 11695.945 189.04 11696.225 336.445 ;
      RECT 11695.385 187.94 11695.665 336.685 ;
      RECT 11694.825 189.04 11695.105 336.925 ;
      RECT 11694.265 187.94 11694.545 337.165 ;
      RECT 11693.705 189.04 11693.985 337.165 ;
      RECT 11693.145 189.04 11693.425 336.925 ;
      RECT 11692.585 189.04 11692.865 336.685 ;
      RECT 11692.025 189.04 11692.305 336.445 ;
      RECT 11691.465 189.04 11691.745 336.205 ;
      RECT 11690.905 189.04 11691.185 335.965 ;
      RECT 11690.345 189.04 11690.625 335.725 ;
      RECT 11689.785 189.04 11690.065 335.485 ;
      RECT 11680.825 187.94 11681.105 335.515 ;
      RECT 11680.265 189.04 11680.545 335.755 ;
      RECT 11679.705 187.94 11679.985 335.995 ;
      RECT 11679.145 189.04 11679.425 336.21 ;
      RECT 11678.585 189.04 11678.865 335.785 ;
      RECT 11678.025 189.04 11678.305 335.545 ;
      RECT 11677.465 189.04 11677.745 335.305 ;
      RECT 11676.905 189.04 11677.185 335.065 ;
      RECT 11676.345 189.04 11676.625 334.825 ;
      RECT 11675.785 189.04 11676.065 334.585 ;
      RECT 11675.225 189.04 11675.505 334.345 ;
      RECT 11674.665 189.04 11674.945 334.105 ;
      RECT 11674.105 189.04 11674.385 333.865 ;
      RECT 11673.545 189.04 11673.825 333.625 ;
      RECT 11671.025 189.04 11671.305 332.8 ;
      RECT 11670.465 189.04 11670.745 332.56 ;
      RECT 11669.905 189.04 11670.185 332.32 ;
      RECT 11669.345 187.94 11669.625 332.08 ;
      RECT 11668.785 189.04 11669.065 331.84 ;
      RECT 11668.225 187.94 11668.505 331.6 ;
      RECT 11667.665 189.04 11667.945 331.36 ;
      RECT 11667.105 189.04 11667.385 331.12 ;
      RECT 11640.505 189.04 11640.785 342.165 ;
      RECT 11639.945 187.94 11640.225 342.405 ;
      RECT 11639.385 189.04 11639.665 342.645 ;
      RECT 11638.825 187.94 11639.105 342.89 ;
      RECT 11638.265 189.04 11638.545 343.13 ;
      RECT 11637.705 187.94 11637.985 343.37 ;
      RECT 11637.145 189.04 11637.425 343.61 ;
      RECT 11636.585 189.04 11636.865 343.85 ;
      RECT 11636.025 189.04 11636.305 329.47 ;
      RECT 11635.465 189.04 11635.745 329.23 ;
      RECT 11634.905 189.04 11635.185 328.99 ;
      RECT 11634.345 189.04 11634.625 328.75 ;
      RECT 11633.785 189.04 11634.065 328.51 ;
      RECT 11633.225 189.04 11633.505 328.27 ;
      RECT 11632.665 189.04 11632.945 328.03 ;
      RECT 11632.105 189.04 11632.385 327.79 ;
      RECT 11631.545 189.04 11631.825 327.55 ;
      RECT 11630.985 189.04 11631.265 327.31 ;
      RECT 11630.425 187.94 11630.705 327.07 ;
      RECT 11629.865 189.04 11630.145 326.83 ;
      RECT 11629.305 187.94 11629.585 326.59 ;
      RECT 11628.745 189.04 11629.025 326.35 ;
      RECT 11614.745 187.94 11615.025 332.47 ;
      RECT 11614.185 189.04 11614.465 332.23 ;
      RECT 11613.625 189.04 11613.905 331.99 ;
      RECT 11613.065 189.04 11613.345 331.75 ;
      RECT 11612.505 189.04 11612.785 331.51 ;
      RECT 11611.945 189.04 11612.225 331.27 ;
      RECT 11611.385 189.04 11611.665 331.03 ;
      RECT 11610.825 189.04 11611.105 330.79 ;
      RECT 11610.265 189.04 11610.545 330.55 ;
      RECT 11609.705 187.94 11609.985 330.31 ;
      RECT 11609.145 189.04 11609.425 330.07 ;
      RECT 11608.585 187.94 11608.865 329.83 ;
      RECT 11608.025 189.04 11608.305 329.59 ;
      RECT 11607.465 189.04 11607.745 329.35 ;
      RECT 11606.905 189.04 11607.185 329.11 ;
      RECT 11606.345 189.04 11606.625 328.87 ;
      RECT 11605.785 189.04 11606.065 328.63 ;
      RECT 11605.225 189.04 11605.505 328.39 ;
      RECT 11604.665 189.04 11604.945 328.15 ;
      RECT 11604.105 189.04 11604.385 327.91 ;
      RECT 11603.545 189.04 11603.825 327.67 ;
      RECT 11602.985 189.04 11603.265 327.43 ;
      RECT 11602.425 189.04 11602.705 327.19 ;
      RECT 11563.225 189.04 11563.505 334.095 ;
      RECT 11562.665 189.04 11562.945 334.335 ;
      RECT 11562.105 189.04 11562.385 334.575 ;
      RECT 11561.545 187.94 11561.825 334.815 ;
      RECT 11560.985 189.04 11561.265 335.055 ;
      RECT 11560.425 187.94 11560.705 335.295 ;
      RECT 11559.865 189.04 11560.145 335.535 ;
      RECT 11559.305 189.04 11559.585 335.775 ;
      RECT 11558.745 189.04 11559.025 336.015 ;
      RECT 11558.185 187.94 11558.465 336.255 ;
      RECT 11557.625 189.04 11557.905 336.495 ;
      RECT 11557.065 187.94 11557.345 336.735 ;
      RECT 11556.505 189.04 11556.785 336.975 ;
      RECT 11555.945 187.94 11556.225 337.215 ;
      RECT 11555.385 189.04 11555.665 337.455 ;
      RECT 11554.825 189.04 11555.105 337.695 ;
      RECT 11554.265 189.04 11554.545 337.695 ;
      RECT 11553.705 189.04 11553.985 337.455 ;
      RECT 11553.145 189.04 11553.425 337.215 ;
      RECT 11552.585 189.04 11552.865 336.975 ;
      RECT 11552.025 189.04 11552.305 336.735 ;
      RECT 11551.465 189.04 11551.745 336.495 ;
      RECT 11550.905 189.04 11551.185 336.255 ;
      RECT 11550.345 189.04 11550.625 336.015 ;
      RECT 11549.785 189.04 11550.065 335.775 ;
      RECT 11540.825 189.04 11541.105 335.29 ;
      RECT 11540.265 187.94 11540.545 335.05 ;
      RECT 11539.705 189.04 11539.985 334.81 ;
      RECT 11539.145 187.94 11539.425 334.57 ;
      RECT 11538.585 189.04 11538.865 334.33 ;
      RECT 11538.025 187.94 11538.305 334.09 ;
      RECT 11537.465 189.04 11537.745 333.85 ;
      RECT 11536.905 189.04 11537.185 333.61 ;
      RECT 11536.345 189.04 11536.625 333.37 ;
      RECT 11535.785 189.04 11536.065 333.13 ;
      RECT 11535.225 189.04 11535.505 332.89 ;
      RECT 11534.665 189.04 11534.945 332.65 ;
      RECT 11534.105 189.04 11534.385 332.41 ;
      RECT 11533.545 189.04 11533.825 332.17 ;
      RECT 11531.025 187.94 11531.305 333.89 ;
      RECT 11530.465 189.04 11530.745 333.65 ;
      RECT 11529.905 187.94 11530.185 333.41 ;
      RECT 11529.345 189.04 11529.625 333.17 ;
      RECT 11528.785 189.04 11529.065 332.93 ;
      RECT 11528.225 189.04 11528.505 332.69 ;
      RECT 11527.665 189.04 11527.945 332.45 ;
      RECT 11527.105 189.04 11527.385 332.21 ;
      RECT 11501.065 189.04 11501.345 329.86 ;
      RECT 11500.505 189.04 11500.785 330.1 ;
      RECT 11499.945 189.04 11500.225 330.34 ;
      RECT 11499.385 189.04 11499.665 330.585 ;
      RECT 11498.825 189.04 11499.105 330.825 ;
      RECT 11498.265 189.04 11498.545 331.065 ;
      RECT 11497.705 189.04 11497.985 331.065 ;
      RECT 11497.145 189.04 11497.425 330.825 ;
      RECT 11496.585 189.04 11496.865 330.585 ;
      RECT 11496.025 187.94 11496.305 330.345 ;
      RECT 11495.465 189.04 11495.745 330.105 ;
      RECT 11494.905 187.94 11495.185 329.865 ;
      RECT 11494.345 189.04 11494.625 329.625 ;
      RECT 11493.785 189.04 11494.065 329.385 ;
      RECT 11493.225 189.04 11493.505 329.145 ;
      RECT 11492.665 187.94 11492.945 328.905 ;
      RECT 11492.105 189.04 11492.385 328.665 ;
      RECT 11491.545 187.94 11491.825 328.425 ;
      RECT 11490.985 189.04 11491.265 328.185 ;
      RECT 11490.425 187.94 11490.705 327.945 ;
      RECT 11489.865 189.04 11490.145 327.705 ;
      RECT 11489.305 189.04 11489.585 327.465 ;
      RECT 11488.745 189.04 11489.025 327.225 ;
      RECT 11488.185 189.04 11488.465 326.985 ;
      RECT 11474.745 189.04 11475.025 332.785 ;
      RECT 11474.185 189.04 11474.465 332.545 ;
      RECT 11473.625 189.04 11473.905 332.305 ;
      RECT 11473.065 189.04 11473.345 332.065 ;
      RECT 11472.505 189.04 11472.785 331.825 ;
      RECT 11471.945 189.04 11472.225 331.585 ;
      RECT 11471.385 189.04 11471.665 331.345 ;
      RECT 11470.825 189.04 11471.105 331.105 ;
      RECT 11470.265 187.94 11470.545 330.865 ;
      RECT 11469.705 189.04 11469.985 330.625 ;
      RECT 11469.145 187.94 11469.425 330.305 ;
      RECT 11468.585 189.04 11468.865 330.145 ;
      RECT 11468.025 187.94 11468.305 329.905 ;
      RECT 11467.465 189.04 11467.745 329.665 ;
      RECT 11466.905 189.04 11467.185 329.425 ;
      RECT 11466.345 189.04 11466.625 329.185 ;
      RECT 11465.785 189.04 11466.065 328.945 ;
      RECT 11465.225 189.04 11465.505 328.705 ;
      RECT 11464.665 189.04 11464.945 328.465 ;
      RECT 11464.105 189.04 11464.385 328.225 ;
      RECT 11463.545 189.04 11463.825 327.985 ;
      RECT 11462.985 187.94 11463.265 327.745 ;
      RECT 11462.425 189.04 11462.705 327.505 ;
      RECT 11461.865 187.94 11462.145 327.265 ;
      RECT 11422.665 189.04 11422.945 332.875 ;
      RECT 11422.105 189.04 11422.385 333.115 ;
      RECT 11421.545 189.04 11421.825 333.355 ;
      RECT 11420.985 189.04 11421.265 333.595 ;
      RECT 11420.425 189.04 11420.705 333.835 ;
      RECT 11419.865 189.04 11420.145 334.075 ;
      RECT 11419.305 189.04 11419.585 334.315 ;
      RECT 11418.745 189.04 11419.025 334.555 ;
      RECT 11418.185 189.04 11418.465 334.795 ;
      RECT 11417.625 189.04 11417.905 335.035 ;
      RECT 11417.065 189.04 11417.345 335.275 ;
      RECT 11416.505 189.04 11416.785 335.515 ;
      RECT 11415.945 189.04 11416.225 335.755 ;
      RECT 11415.385 189.04 11415.665 335.755 ;
      RECT 11414.825 187.94 11415.105 335.515 ;
      RECT 11414.265 189.04 11414.545 335.275 ;
      RECT 11413.705 187.94 11413.985 335.035 ;
      RECT 11413.145 189.04 11413.425 334.795 ;
      RECT 11412.585 189.04 11412.865 334.555 ;
      RECT 11412.025 189.04 11412.305 334.315 ;
      RECT 11411.465 187.94 11411.745 334.05 ;
      RECT 11410.905 189.04 11411.185 333.81 ;
      RECT 11410.345 187.94 11410.625 333.57 ;
      RECT 11409.785 189.04 11410.065 333.33 ;
      RECT 11400.825 187.94 11401.105 327.165 ;
      RECT 11400.265 189.04 11400.545 327.405 ;
      RECT 11399.705 189.04 11399.985 327.645 ;
      RECT 11399.145 189.04 11399.425 327.645 ;
      RECT 11398.585 189.04 11398.865 327.405 ;
      RECT 11398.025 189.04 11398.305 327.165 ;
      RECT 11397.465 189.04 11397.745 326.925 ;
      RECT 11396.905 189.04 11397.185 326.685 ;
      RECT 11396.345 189.04 11396.625 326.445 ;
      RECT 11395.785 189.04 11396.065 326.205 ;
      RECT 11395.225 189.04 11395.505 325.965 ;
      RECT 11394.665 189.04 11394.945 325.725 ;
      RECT 11394.105 189.04 11394.385 325.485 ;
      RECT 11393.545 187.94 11393.825 325.245 ;
      RECT 11391.025 189.04 11391.305 326.965 ;
      RECT 11390.465 187.94 11390.745 326.725 ;
      RECT 11389.905 189.04 11390.185 326.485 ;
      RECT 11389.345 187.94 11389.625 326.245 ;
      RECT 11388.785 189.04 11389.065 326.005 ;
      RECT 11388.225 189.04 11388.505 325.765 ;
      RECT 11387.665 189.04 11387.945 325.525 ;
      RECT 11361.625 189.04 11361.905 328.31 ;
      RECT 11361.065 189.04 11361.345 328.55 ;
      RECT 11360.505 189.04 11360.785 328.79 ;
      RECT 11359.945 189.04 11360.225 329.03 ;
      RECT 11359.385 189.04 11359.665 329.27 ;
      RECT 11358.825 187.94 11359.105 329.51 ;
      RECT 11358.265 189.04 11358.545 329.75 ;
      RECT 11357.705 187.94 11357.985 329.99 ;
      RECT 11357.145 189.04 11357.425 330.23 ;
      RECT 11356.585 189.04 11356.865 330.47 ;
      RECT 11356.025 189.04 11356.305 330.71 ;
      RECT 11355.465 189.04 11355.745 330.95 ;
      RECT 11354.905 189.04 11355.185 331.19 ;
      RECT 11354.345 189.04 11354.625 331.43 ;
      RECT 11353.785 189.04 11354.065 331.67 ;
      RECT 11353.225 189.04 11353.505 331.67 ;
      RECT 11352.665 189.04 11352.945 331.43 ;
      RECT 11352.105 189.04 11352.385 331.19 ;
      RECT 11351.545 189.04 11351.825 330.95 ;
      RECT 11350.985 189.04 11351.265 330.705 ;
      RECT 11350.425 189.04 11350.705 330.465 ;
      RECT 11349.865 189.04 11350.145 330.225 ;
      RECT 11349.305 187.94 11349.585 329.985 ;
      RECT 11348.745 189.04 11349.025 329.745 ;
      RECT 11335.305 187.94 11335.585 327.225 ;
      RECT 11334.745 189.04 11335.025 326.985 ;
      RECT 11334.185 189.04 11334.465 326.745 ;
      RECT 11333.625 189.04 11333.905 326.505 ;
      RECT 11333.065 187.94 11333.345 326.265 ;
      RECT 11332.505 189.04 11332.785 326.025 ;
      RECT 11331.945 187.94 11332.225 325.785 ;
      RECT 11331.385 189.04 11331.665 325.545 ;
      RECT 11330.825 187.94 11331.105 325.305 ;
      RECT 11330.265 189.04 11330.545 325.065 ;
      RECT 11329.705 189.04 11329.985 324.825 ;
      RECT 11329.145 189.04 11329.425 324.585 ;
      RECT 11328.585 189.04 11328.865 324.345 ;
      RECT 11328.025 189.04 11328.305 324.105 ;
      RECT 11327.465 189.04 11327.745 323.865 ;
      RECT 11326.905 189.04 11327.185 323.625 ;
      RECT 11326.345 189.04 11326.625 323.385 ;
      RECT 11325.785 189.04 11326.065 323.145 ;
      RECT 11325.225 189.04 11325.505 322.905 ;
      RECT 11324.665 189.04 11324.945 322.665 ;
      RECT 11324.105 189.04 11324.385 322.425 ;
      RECT 11323.545 187.94 11323.825 322.185 ;
      RECT 11322.985 189.04 11323.265 321.945 ;
      RECT 11322.425 187.94 11322.705 321.705 ;
      RECT 11282.665 189.04 11282.945 332.175 ;
      RECT 11282.105 187.94 11282.385 332.415 ;
      RECT 11281.545 189.04 11281.825 332.655 ;
      RECT 11280.985 189.04 11281.265 332.895 ;
      RECT 11280.425 189.04 11280.705 333.135 ;
      RECT 11279.865 189.04 11280.145 333.375 ;
      RECT 11279.305 189.04 11279.585 333.615 ;
      RECT 11278.745 189.04 11279.025 333.86 ;
      RECT 11278.185 189.04 11278.465 334.1 ;
      RECT 11277.625 189.04 11277.905 334.34 ;
      RECT 11277.065 187.94 11277.345 334.58 ;
      RECT 11276.505 189.04 11276.785 334.82 ;
      RECT 11275.945 187.94 11276.225 335.06 ;
      RECT 11275.385 189.04 11275.665 335.3 ;
      RECT 11274.825 189.04 11275.105 335.54 ;
      RECT 11274.265 189.04 11274.545 335.78 ;
      RECT 11273.705 189.04 11273.985 336.02 ;
      RECT 11273.145 189.04 11273.425 336.26 ;
      RECT 11272.585 189.04 11272.865 336.5 ;
      RECT 11272.025 189.04 11272.305 336.74 ;
      RECT 11271.465 189.04 11271.745 336.98 ;
      RECT 11270.905 189.04 11271.185 337.22 ;
      RECT 11270.345 189.04 11270.625 337.46 ;
      RECT 11269.785 189.04 11270.065 337.7 ;
      RECT 11260.825 189.04 11261.105 333.285 ;
      RECT 11260.265 189.04 11260.545 333.045 ;
      RECT 11259.705 189.04 11259.985 332.805 ;
      RECT 11259.145 187.94 11259.425 332.565 ;
      RECT 11258.585 189.04 11258.865 332.325 ;
      RECT 11258.025 187.94 11258.305 332.085 ;
      RECT 11257.465 189.04 11257.745 331.845 ;
      RECT 11256.905 189.04 11257.185 331.605 ;
      RECT 11256.345 189.04 11256.625 331.365 ;
      RECT 11255.785 187.94 11256.065 331.125 ;
      RECT 11255.225 189.04 11255.505 330.885 ;
      RECT 11254.665 187.94 11254.945 330.645 ;
      RECT 11254.105 189.04 11254.385 330.405 ;
      RECT 11253.545 187.94 11253.825 330.165 ;
      RECT 11251.025 189.04 11251.305 322.565 ;
      RECT 11250.465 189.04 11250.745 322.325 ;
      RECT 11249.905 189.04 11250.185 322.085 ;
      RECT 11249.345 189.04 11249.625 321.845 ;
      RECT 11248.785 189.04 11249.065 321.605 ;
      RECT 11248.225 189.04 11248.505 321.365 ;
      RECT 11247.665 189.04 11247.945 321.125 ;
      RECT 11221.625 189.04 11221.905 335 ;
      RECT 11221.065 189.04 11221.345 335.24 ;
      RECT 11220.505 189.04 11220.785 335.48 ;
      RECT 11219.945 189.04 11220.225 335.72 ;
      RECT 11219.385 189.04 11219.665 335.96 ;
      RECT 11218.825 187.94 11219.105 335.96 ;
      RECT 11218.265 189.04 11218.545 335.72 ;
      RECT 11217.705 187.94 11217.985 335.475 ;
      RECT 11217.145 189.04 11217.425 335.235 ;
      RECT 11216.585 187.94 11216.865 334.995 ;
      RECT 11216.025 189.04 11216.305 334.755 ;
      RECT 11215.465 189.04 11215.745 334.515 ;
      RECT 11214.905 189.04 11215.185 334.275 ;
      RECT 11214.345 189.04 11214.625 334.035 ;
      RECT 11213.785 189.04 11214.065 333.795 ;
      RECT 11213.225 189.04 11213.505 333.555 ;
      RECT 11212.665 189.04 11212.945 333.315 ;
      RECT 11212.105 189.04 11212.385 333.075 ;
      RECT 11211.545 187.94 11211.825 332.835 ;
      RECT 11210.985 189.04 11211.265 332.595 ;
      RECT 11210.425 187.94 11210.705 332.355 ;
      RECT 11209.865 189.04 11210.145 332.115 ;
      RECT 11209.305 189.04 11209.585 331.875 ;
      RECT 11208.745 189.04 11209.025 331.635 ;
      RECT 11195.305 189.04 11195.585 335.035 ;
      RECT 11194.745 189.04 11195.025 335.275 ;
      RECT 11194.185 189.04 11194.465 335.52 ;
      RECT 11193.625 189.04 11193.905 335.76 ;
      RECT 11193.065 189.04 11193.345 336 ;
      RECT 11192.505 189.04 11192.785 336 ;
      RECT 11191.945 189.04 11192.225 335.76 ;
      RECT 11191.385 189.04 11191.665 335.52 ;
      RECT 11190.825 189.04 11191.105 328.505 ;
      RECT 11190.265 189.04 11190.545 328.265 ;
      RECT 11189.705 189.04 11189.985 328.025 ;
      RECT 11189.145 187.94 11189.425 327.785 ;
      RECT 11188.585 189.04 11188.865 327.545 ;
      RECT 11188.025 187.94 11188.305 327.305 ;
      RECT 11187.465 189.04 11187.745 327.065 ;
      RECT 11186.905 189.04 11187.185 326.825 ;
      RECT 11186.345 189.04 11186.625 326.585 ;
      RECT 11185.785 187.94 11186.065 326.345 ;
      RECT 11185.225 189.04 11185.505 326.105 ;
      RECT 11184.665 187.94 11184.945 325.865 ;
      RECT 11184.105 189.04 11184.385 325.625 ;
      RECT 11183.545 187.94 11183.825 325.385 ;
      RECT 11182.985 189.04 11183.265 325.145 ;
      RECT 11182.425 189.04 11182.705 324.905 ;
      RECT 11142.105 189.04 11142.385 333.8 ;
      RECT 11141.545 189.04 11141.825 334.04 ;
      RECT 11140.985 189.04 11141.265 334.285 ;
      RECT 11140.425 189.04 11140.705 334.525 ;
      RECT 11139.865 189.04 11140.145 334.765 ;
      RECT 11139.305 189.04 11139.585 335.005 ;
      RECT 11138.745 189.04 11139.025 335.245 ;
      RECT 11138.185 189.04 11138.465 335.485 ;
      RECT 11137.625 189.04 11137.905 335.725 ;
      RECT 11137.065 189.04 11137.345 335.965 ;
      RECT 11136.505 187.94 11136.785 336.205 ;
      RECT 11135.945 189.04 11136.225 336.445 ;
      RECT 11135.385 187.94 11135.665 336.685 ;
      RECT 11134.825 189.04 11135.105 336.925 ;
      RECT 11134.265 187.94 11134.545 337.165 ;
      RECT 11133.705 189.04 11133.985 337.165 ;
      RECT 11133.145 189.04 11133.425 336.925 ;
      RECT 11132.585 189.04 11132.865 336.685 ;
      RECT 11132.025 189.04 11132.305 336.445 ;
      RECT 11131.465 189.04 11131.745 336.205 ;
      RECT 11130.905 189.04 11131.185 335.965 ;
      RECT 11130.345 189.04 11130.625 335.725 ;
      RECT 11129.785 189.04 11130.065 335.485 ;
      RECT 11120.825 187.94 11121.105 335.515 ;
      RECT 11120.265 189.04 11120.545 335.755 ;
      RECT 11119.705 187.94 11119.985 335.995 ;
      RECT 11119.145 189.04 11119.425 336.21 ;
      RECT 11118.585 189.04 11118.865 335.785 ;
      RECT 11118.025 189.04 11118.305 335.545 ;
      RECT 11117.465 189.04 11117.745 335.305 ;
      RECT 11116.905 189.04 11117.185 335.065 ;
      RECT 11116.345 189.04 11116.625 334.825 ;
      RECT 11115.785 189.04 11116.065 334.585 ;
      RECT 11115.225 189.04 11115.505 334.345 ;
      RECT 11114.665 189.04 11114.945 334.105 ;
      RECT 11114.105 189.04 11114.385 333.865 ;
      RECT 11113.545 189.04 11113.825 333.625 ;
      RECT 11111.025 189.04 11111.305 332.8 ;
      RECT 11110.465 189.04 11110.745 332.56 ;
      RECT 11109.905 189.04 11110.185 332.32 ;
      RECT 11109.345 187.94 11109.625 332.08 ;
      RECT 11108.785 189.04 11109.065 331.84 ;
      RECT 11108.225 187.94 11108.505 331.6 ;
      RECT 11107.665 189.04 11107.945 331.36 ;
      RECT 11107.105 189.04 11107.385 331.12 ;
      RECT 11080.505 189.04 11080.785 342.165 ;
      RECT 11079.945 187.94 11080.225 342.405 ;
      RECT 11079.385 189.04 11079.665 342.645 ;
      RECT 11078.825 187.94 11079.105 342.89 ;
      RECT 11078.265 189.04 11078.545 343.13 ;
      RECT 11077.705 187.94 11077.985 343.37 ;
      RECT 11077.145 189.04 11077.425 343.61 ;
      RECT 11076.585 189.04 11076.865 343.85 ;
      RECT 11076.025 189.04 11076.305 329.47 ;
      RECT 11075.465 189.04 11075.745 329.23 ;
      RECT 11074.905 189.04 11075.185 328.99 ;
      RECT 11074.345 189.04 11074.625 328.75 ;
      RECT 11073.785 189.04 11074.065 328.51 ;
      RECT 11073.225 189.04 11073.505 328.27 ;
      RECT 11072.665 189.04 11072.945 328.03 ;
      RECT 11072.105 189.04 11072.385 327.79 ;
      RECT 11071.545 189.04 11071.825 327.55 ;
      RECT 11070.985 189.04 11071.265 327.31 ;
      RECT 11070.425 187.94 11070.705 327.07 ;
      RECT 11069.865 189.04 11070.145 326.83 ;
      RECT 11069.305 187.94 11069.585 326.59 ;
      RECT 11068.745 189.04 11069.025 326.35 ;
      RECT 11054.745 187.94 11055.025 332.47 ;
      RECT 11054.185 189.04 11054.465 332.23 ;
      RECT 11053.625 189.04 11053.905 331.99 ;
      RECT 11053.065 189.04 11053.345 331.75 ;
      RECT 11052.505 189.04 11052.785 331.51 ;
      RECT 11051.945 189.04 11052.225 331.27 ;
      RECT 11051.385 189.04 11051.665 331.03 ;
      RECT 11050.825 189.04 11051.105 330.79 ;
      RECT 11050.265 189.04 11050.545 330.55 ;
      RECT 11049.705 187.94 11049.985 330.31 ;
      RECT 11049.145 189.04 11049.425 330.07 ;
      RECT 11048.585 187.94 11048.865 329.83 ;
      RECT 11048.025 189.04 11048.305 329.59 ;
      RECT 11047.465 189.04 11047.745 329.35 ;
      RECT 11046.905 189.04 11047.185 329.11 ;
      RECT 11046.345 189.04 11046.625 328.87 ;
      RECT 11045.785 189.04 11046.065 328.63 ;
      RECT 11045.225 189.04 11045.505 328.39 ;
      RECT 11044.665 189.04 11044.945 328.15 ;
      RECT 11044.105 189.04 11044.385 327.91 ;
      RECT 11043.545 189.04 11043.825 327.67 ;
      RECT 11042.985 189.04 11043.265 327.43 ;
      RECT 11042.425 189.04 11042.705 327.19 ;
      RECT 11003.225 189.04 11003.505 334.095 ;
      RECT 11002.665 189.04 11002.945 334.335 ;
      RECT 11002.105 189.04 11002.385 334.575 ;
      RECT 11001.545 187.94 11001.825 334.815 ;
      RECT 11000.985 189.04 11001.265 335.055 ;
      RECT 11000.425 187.94 11000.705 335.295 ;
      RECT 10999.865 189.04 11000.145 335.535 ;
      RECT 10999.305 189.04 10999.585 335.775 ;
      RECT 10998.745 189.04 10999.025 336.015 ;
      RECT 10998.185 187.94 10998.465 336.255 ;
      RECT 10997.625 189.04 10997.905 336.495 ;
      RECT 10997.065 187.94 10997.345 336.735 ;
      RECT 10996.505 189.04 10996.785 336.975 ;
      RECT 10995.945 187.94 10996.225 337.215 ;
      RECT 10995.385 189.04 10995.665 337.455 ;
      RECT 10994.825 189.04 10995.105 337.695 ;
      RECT 10994.265 189.04 10994.545 337.695 ;
      RECT 10993.705 189.04 10993.985 337.455 ;
      RECT 10993.145 189.04 10993.425 337.215 ;
      RECT 10992.585 189.04 10992.865 336.975 ;
      RECT 10992.025 189.04 10992.305 336.735 ;
      RECT 10991.465 189.04 10991.745 336.495 ;
      RECT 10990.905 189.04 10991.185 336.255 ;
      RECT 10990.345 189.04 10990.625 336.015 ;
      RECT 10989.785 189.04 10990.065 335.775 ;
      RECT 10980.825 189.04 10981.105 335.29 ;
      RECT 10980.265 187.94 10980.545 335.05 ;
      RECT 10979.705 189.04 10979.985 334.81 ;
      RECT 10979.145 187.94 10979.425 334.57 ;
      RECT 10978.585 189.04 10978.865 334.33 ;
      RECT 10978.025 187.94 10978.305 334.09 ;
      RECT 10977.465 189.04 10977.745 333.85 ;
      RECT 10976.905 189.04 10977.185 333.61 ;
      RECT 10976.345 189.04 10976.625 333.37 ;
      RECT 10975.785 189.04 10976.065 333.13 ;
      RECT 10975.225 189.04 10975.505 332.89 ;
      RECT 10974.665 189.04 10974.945 332.65 ;
      RECT 10974.105 189.04 10974.385 332.41 ;
      RECT 10973.545 189.04 10973.825 332.17 ;
      RECT 10971.025 187.94 10971.305 333.89 ;
      RECT 10970.465 189.04 10970.745 333.65 ;
      RECT 10969.905 187.94 10970.185 333.41 ;
      RECT 10969.345 189.04 10969.625 333.17 ;
      RECT 10968.785 189.04 10969.065 332.93 ;
      RECT 10968.225 189.04 10968.505 332.69 ;
      RECT 10967.665 189.04 10967.945 332.45 ;
      RECT 10967.105 189.04 10967.385 332.21 ;
      RECT 10941.065 189.04 10941.345 329.86 ;
      RECT 10940.505 189.04 10940.785 330.1 ;
      RECT 10939.945 189.04 10940.225 330.34 ;
      RECT 10939.385 189.04 10939.665 330.585 ;
      RECT 10938.825 189.04 10939.105 330.825 ;
      RECT 10938.265 189.04 10938.545 331.065 ;
      RECT 10937.705 189.04 10937.985 331.065 ;
      RECT 10937.145 189.04 10937.425 330.825 ;
      RECT 10936.585 189.04 10936.865 330.585 ;
      RECT 10936.025 187.94 10936.305 330.345 ;
      RECT 10935.465 189.04 10935.745 330.105 ;
      RECT 10934.905 187.94 10935.185 329.865 ;
      RECT 10934.345 189.04 10934.625 329.625 ;
      RECT 10933.785 189.04 10934.065 329.385 ;
      RECT 10933.225 189.04 10933.505 329.145 ;
      RECT 10932.665 187.94 10932.945 328.905 ;
      RECT 10932.105 189.04 10932.385 328.665 ;
      RECT 10931.545 187.94 10931.825 328.425 ;
      RECT 10930.985 189.04 10931.265 328.185 ;
      RECT 10930.425 187.94 10930.705 327.945 ;
      RECT 10929.865 189.04 10930.145 327.705 ;
      RECT 10929.305 189.04 10929.585 327.465 ;
      RECT 10928.745 189.04 10929.025 327.225 ;
      RECT 10928.185 189.04 10928.465 326.985 ;
      RECT 10914.745 189.04 10915.025 332.785 ;
      RECT 10914.185 189.04 10914.465 332.545 ;
      RECT 10913.625 189.04 10913.905 332.305 ;
      RECT 10913.065 189.04 10913.345 332.065 ;
      RECT 10912.505 189.04 10912.785 331.825 ;
      RECT 10911.945 189.04 10912.225 331.585 ;
      RECT 10911.385 189.04 10911.665 331.345 ;
      RECT 10910.825 189.04 10911.105 331.105 ;
      RECT 10910.265 187.94 10910.545 330.865 ;
      RECT 10909.705 189.04 10909.985 330.625 ;
      RECT 10909.145 187.94 10909.425 330.305 ;
      RECT 10908.585 189.04 10908.865 330.145 ;
      RECT 10908.025 187.94 10908.305 329.905 ;
      RECT 10907.465 189.04 10907.745 329.665 ;
      RECT 10906.905 189.04 10907.185 329.425 ;
      RECT 10906.345 189.04 10906.625 329.185 ;
      RECT 10905.785 189.04 10906.065 328.945 ;
      RECT 10905.225 189.04 10905.505 328.705 ;
      RECT 10904.665 189.04 10904.945 328.465 ;
      RECT 10904.105 189.04 10904.385 328.225 ;
      RECT 10903.545 189.04 10903.825 327.985 ;
      RECT 10902.985 187.94 10903.265 327.745 ;
      RECT 10902.425 189.04 10902.705 327.505 ;
      RECT 10901.865 187.94 10902.145 327.265 ;
      RECT 10862.665 189.04 10862.945 332.875 ;
      RECT 10862.105 189.04 10862.385 333.115 ;
      RECT 10861.545 189.04 10861.825 333.355 ;
      RECT 10860.985 189.04 10861.265 333.595 ;
      RECT 10860.425 189.04 10860.705 333.835 ;
      RECT 10859.865 189.04 10860.145 334.075 ;
      RECT 10859.305 189.04 10859.585 334.315 ;
      RECT 10858.745 189.04 10859.025 334.555 ;
      RECT 10858.185 189.04 10858.465 334.795 ;
      RECT 10857.625 189.04 10857.905 335.035 ;
      RECT 10857.065 189.04 10857.345 335.275 ;
      RECT 10856.505 189.04 10856.785 335.515 ;
      RECT 10855.945 189.04 10856.225 335.755 ;
      RECT 10855.385 189.04 10855.665 335.755 ;
      RECT 10854.825 187.94 10855.105 335.515 ;
      RECT 10854.265 189.04 10854.545 335.275 ;
      RECT 10853.705 187.94 10853.985 335.035 ;
      RECT 10853.145 189.04 10853.425 334.795 ;
      RECT 10852.585 189.04 10852.865 334.555 ;
      RECT 10852.025 189.04 10852.305 334.315 ;
      RECT 10851.465 187.94 10851.745 334.05 ;
      RECT 10850.905 189.04 10851.185 333.81 ;
      RECT 10850.345 187.94 10850.625 333.57 ;
      RECT 10849.785 189.04 10850.065 333.33 ;
      RECT 10840.825 187.94 10841.105 327.165 ;
      RECT 10840.265 189.04 10840.545 327.405 ;
      RECT 10839.705 189.04 10839.985 327.645 ;
      RECT 10839.145 189.04 10839.425 327.645 ;
      RECT 10838.585 189.04 10838.865 327.405 ;
      RECT 10838.025 189.04 10838.305 327.165 ;
      RECT 10837.465 189.04 10837.745 326.925 ;
      RECT 10836.905 189.04 10837.185 326.685 ;
      RECT 10836.345 189.04 10836.625 326.445 ;
      RECT 10835.785 189.04 10836.065 326.205 ;
      RECT 10835.225 189.04 10835.505 325.965 ;
      RECT 10834.665 189.04 10834.945 325.725 ;
      RECT 10834.105 189.04 10834.385 325.485 ;
      RECT 10833.545 187.94 10833.825 325.245 ;
      RECT 10831.025 189.04 10831.305 326.965 ;
      RECT 10830.465 187.94 10830.745 326.725 ;
      RECT 10829.905 189.04 10830.185 326.485 ;
      RECT 10829.345 187.94 10829.625 326.245 ;
      RECT 10828.785 189.04 10829.065 326.005 ;
      RECT 10828.225 189.04 10828.505 325.765 ;
      RECT 10827.665 189.04 10827.945 325.525 ;
      RECT 10801.625 189.04 10801.905 328.31 ;
      RECT 10801.065 189.04 10801.345 328.55 ;
      RECT 10800.505 189.04 10800.785 328.79 ;
      RECT 10799.945 189.04 10800.225 329.03 ;
      RECT 10799.385 189.04 10799.665 329.27 ;
      RECT 10798.825 187.94 10799.105 329.51 ;
      RECT 10798.265 189.04 10798.545 329.75 ;
      RECT 10797.705 187.94 10797.985 329.99 ;
      RECT 10797.145 189.04 10797.425 330.23 ;
      RECT 10796.585 189.04 10796.865 330.47 ;
      RECT 10796.025 189.04 10796.305 330.71 ;
      RECT 10795.465 189.04 10795.745 330.95 ;
      RECT 10794.905 189.04 10795.185 331.19 ;
      RECT 10794.345 189.04 10794.625 331.43 ;
      RECT 10793.785 189.04 10794.065 331.67 ;
      RECT 10793.225 189.04 10793.505 331.67 ;
      RECT 10792.665 189.04 10792.945 331.43 ;
      RECT 10792.105 189.04 10792.385 331.19 ;
      RECT 10791.545 189.04 10791.825 330.95 ;
      RECT 10790.985 189.04 10791.265 330.705 ;
      RECT 10790.425 189.04 10790.705 330.465 ;
      RECT 10789.865 189.04 10790.145 330.225 ;
      RECT 10789.305 187.94 10789.585 329.985 ;
      RECT 10788.745 189.04 10789.025 329.745 ;
      RECT 10775.305 187.94 10775.585 327.225 ;
      RECT 10774.745 189.04 10775.025 326.985 ;
      RECT 10774.185 189.04 10774.465 326.745 ;
      RECT 10773.625 189.04 10773.905 326.505 ;
      RECT 10773.065 187.94 10773.345 326.265 ;
      RECT 10772.505 189.04 10772.785 326.025 ;
      RECT 10771.945 187.94 10772.225 325.785 ;
      RECT 10771.385 189.04 10771.665 325.545 ;
      RECT 10770.825 187.94 10771.105 325.305 ;
      RECT 10770.265 189.04 10770.545 325.065 ;
      RECT 10769.705 189.04 10769.985 324.825 ;
      RECT 10769.145 189.04 10769.425 324.585 ;
      RECT 10768.585 189.04 10768.865 324.345 ;
      RECT 10768.025 189.04 10768.305 324.105 ;
      RECT 10767.465 189.04 10767.745 323.865 ;
      RECT 10766.905 189.04 10767.185 323.625 ;
      RECT 10766.345 189.04 10766.625 323.385 ;
      RECT 10765.785 189.04 10766.065 323.145 ;
      RECT 10765.225 189.04 10765.505 322.905 ;
      RECT 10764.665 189.04 10764.945 322.665 ;
      RECT 10764.105 189.04 10764.385 322.425 ;
      RECT 10763.545 187.94 10763.825 322.185 ;
      RECT 10762.985 189.04 10763.265 321.945 ;
      RECT 10762.425 187.94 10762.705 321.705 ;
      RECT 10722.665 189.04 10722.945 332.175 ;
      RECT 10722.105 187.94 10722.385 332.415 ;
      RECT 10721.545 189.04 10721.825 332.655 ;
      RECT 10720.985 189.04 10721.265 332.895 ;
      RECT 10720.425 189.04 10720.705 333.135 ;
      RECT 10719.865 189.04 10720.145 333.375 ;
      RECT 10719.305 189.04 10719.585 333.615 ;
      RECT 10718.745 189.04 10719.025 333.86 ;
      RECT 10718.185 189.04 10718.465 334.1 ;
      RECT 10717.625 189.04 10717.905 334.34 ;
      RECT 10717.065 187.94 10717.345 334.58 ;
      RECT 10716.505 189.04 10716.785 334.82 ;
      RECT 10715.945 187.94 10716.225 335.06 ;
      RECT 10715.385 189.04 10715.665 335.3 ;
      RECT 10714.825 189.04 10715.105 335.54 ;
      RECT 10714.265 189.04 10714.545 335.78 ;
      RECT 10713.705 189.04 10713.985 336.02 ;
      RECT 10713.145 189.04 10713.425 336.26 ;
      RECT 10712.585 189.04 10712.865 336.5 ;
      RECT 10712.025 189.04 10712.305 336.74 ;
      RECT 10711.465 189.04 10711.745 336.98 ;
      RECT 10710.905 189.04 10711.185 337.22 ;
      RECT 10710.345 189.04 10710.625 337.46 ;
      RECT 10709.785 189.04 10710.065 337.7 ;
      RECT 10700.825 189.04 10701.105 333.285 ;
      RECT 10700.265 189.04 10700.545 333.045 ;
      RECT 10699.705 189.04 10699.985 332.805 ;
      RECT 10699.145 187.94 10699.425 332.565 ;
      RECT 10698.585 189.04 10698.865 332.325 ;
      RECT 10698.025 187.94 10698.305 332.085 ;
      RECT 10697.465 189.04 10697.745 331.845 ;
      RECT 10696.905 189.04 10697.185 331.605 ;
      RECT 10696.345 189.04 10696.625 331.365 ;
      RECT 10695.785 187.94 10696.065 331.125 ;
      RECT 10695.225 189.04 10695.505 330.885 ;
      RECT 10694.665 187.94 10694.945 330.645 ;
      RECT 10694.105 189.04 10694.385 330.405 ;
      RECT 10693.545 187.94 10693.825 330.165 ;
      RECT 10691.025 189.04 10691.305 322.565 ;
      RECT 10690.465 189.04 10690.745 322.325 ;
      RECT 10689.905 189.04 10690.185 322.085 ;
      RECT 10689.345 189.04 10689.625 321.845 ;
      RECT 10688.785 189.04 10689.065 321.605 ;
      RECT 10688.225 189.04 10688.505 321.365 ;
      RECT 10687.665 189.04 10687.945 321.125 ;
      RECT 10661.625 189.04 10661.905 335 ;
      RECT 10661.065 189.04 10661.345 335.24 ;
      RECT 10660.505 189.04 10660.785 335.48 ;
      RECT 10659.945 189.04 10660.225 335.72 ;
      RECT 10659.385 189.04 10659.665 335.96 ;
      RECT 10658.825 187.94 10659.105 335.96 ;
      RECT 10658.265 189.04 10658.545 335.72 ;
      RECT 10657.705 187.94 10657.985 335.475 ;
      RECT 10657.145 189.04 10657.425 335.235 ;
      RECT 10656.585 187.94 10656.865 334.995 ;
      RECT 10656.025 189.04 10656.305 334.755 ;
      RECT 10655.465 189.04 10655.745 334.515 ;
      RECT 10654.905 189.04 10655.185 334.275 ;
      RECT 10654.345 189.04 10654.625 334.035 ;
      RECT 10653.785 189.04 10654.065 333.795 ;
      RECT 10653.225 189.04 10653.505 333.555 ;
      RECT 10652.665 189.04 10652.945 333.315 ;
      RECT 10652.105 189.04 10652.385 333.075 ;
      RECT 10651.545 187.94 10651.825 332.835 ;
      RECT 10650.985 189.04 10651.265 332.595 ;
      RECT 10650.425 187.94 10650.705 332.355 ;
      RECT 10649.865 189.04 10650.145 332.115 ;
      RECT 10649.305 189.04 10649.585 331.875 ;
      RECT 10648.745 189.04 10649.025 331.635 ;
      RECT 10635.305 189.04 10635.585 335.035 ;
      RECT 10634.745 189.04 10635.025 335.275 ;
      RECT 10634.185 189.04 10634.465 335.52 ;
      RECT 10633.625 189.04 10633.905 335.76 ;
      RECT 10633.065 189.04 10633.345 336 ;
      RECT 10632.505 189.04 10632.785 336 ;
      RECT 10631.945 189.04 10632.225 335.76 ;
      RECT 10631.385 189.04 10631.665 335.52 ;
      RECT 10630.825 189.04 10631.105 328.505 ;
      RECT 10630.265 189.04 10630.545 328.265 ;
      RECT 10629.705 189.04 10629.985 328.025 ;
      RECT 10629.145 187.94 10629.425 327.785 ;
      RECT 10628.585 189.04 10628.865 327.545 ;
      RECT 10628.025 187.94 10628.305 327.305 ;
      RECT 10627.465 189.04 10627.745 327.065 ;
      RECT 10626.905 189.04 10627.185 326.825 ;
      RECT 10626.345 189.04 10626.625 326.585 ;
      RECT 10625.785 187.94 10626.065 326.345 ;
      RECT 10625.225 189.04 10625.505 326.105 ;
      RECT 10624.665 187.94 10624.945 325.865 ;
      RECT 10624.105 189.04 10624.385 325.625 ;
      RECT 10623.545 187.94 10623.825 325.385 ;
      RECT 10622.985 189.04 10623.265 325.145 ;
      RECT 10622.425 189.04 10622.705 324.905 ;
      RECT 10582.105 189.04 10582.385 333.8 ;
      RECT 10581.545 189.04 10581.825 334.04 ;
      RECT 10580.985 189.04 10581.265 334.285 ;
      RECT 10580.425 189.04 10580.705 334.525 ;
      RECT 10579.865 189.04 10580.145 334.765 ;
      RECT 10579.305 189.04 10579.585 335.005 ;
      RECT 10578.745 189.04 10579.025 335.245 ;
      RECT 10578.185 189.04 10578.465 335.485 ;
      RECT 10577.625 189.04 10577.905 335.725 ;
      RECT 10577.065 189.04 10577.345 335.965 ;
      RECT 10576.505 187.94 10576.785 336.205 ;
      RECT 10575.945 189.04 10576.225 336.445 ;
      RECT 10575.385 187.94 10575.665 336.685 ;
      RECT 10574.825 189.04 10575.105 336.925 ;
      RECT 10574.265 187.94 10574.545 337.165 ;
      RECT 10573.705 189.04 10573.985 337.165 ;
      RECT 10573.145 189.04 10573.425 336.925 ;
      RECT 10572.585 189.04 10572.865 336.685 ;
      RECT 10572.025 189.04 10572.305 336.445 ;
      RECT 10571.465 189.04 10571.745 336.205 ;
      RECT 10570.905 189.04 10571.185 335.965 ;
      RECT 10570.345 189.04 10570.625 335.725 ;
      RECT 10569.785 189.04 10570.065 335.485 ;
      RECT 10560.825 187.94 10561.105 335.515 ;
      RECT 10560.265 189.04 10560.545 335.755 ;
      RECT 10559.705 187.94 10559.985 335.995 ;
      RECT 10559.145 189.04 10559.425 336.21 ;
      RECT 10558.585 189.04 10558.865 335.785 ;
      RECT 10558.025 189.04 10558.305 335.545 ;
      RECT 10557.465 189.04 10557.745 335.305 ;
      RECT 10556.905 189.04 10557.185 335.065 ;
      RECT 10556.345 189.04 10556.625 334.825 ;
      RECT 10555.785 189.04 10556.065 334.585 ;
      RECT 10555.225 189.04 10555.505 334.345 ;
      RECT 10554.665 189.04 10554.945 334.105 ;
      RECT 10554.105 189.04 10554.385 333.865 ;
      RECT 10553.545 189.04 10553.825 333.625 ;
      RECT 10551.025 189.04 10551.305 332.8 ;
      RECT 10550.465 189.04 10550.745 332.56 ;
      RECT 10549.905 189.04 10550.185 332.32 ;
      RECT 10549.345 187.94 10549.625 332.08 ;
      RECT 10548.785 189.04 10549.065 331.84 ;
      RECT 10548.225 187.94 10548.505 331.6 ;
      RECT 10547.665 189.04 10547.945 331.36 ;
      RECT 10547.105 189.04 10547.385 331.12 ;
      RECT 10520.505 189.04 10520.785 342.165 ;
      RECT 10519.945 187.94 10520.225 342.405 ;
      RECT 10519.385 189.04 10519.665 342.645 ;
      RECT 10518.825 187.94 10519.105 342.89 ;
      RECT 10518.265 189.04 10518.545 343.13 ;
      RECT 10517.705 187.94 10517.985 343.37 ;
      RECT 10517.145 189.04 10517.425 343.61 ;
      RECT 10516.585 189.04 10516.865 343.85 ;
      RECT 10516.025 189.04 10516.305 329.47 ;
      RECT 10515.465 189.04 10515.745 329.23 ;
      RECT 10514.905 189.04 10515.185 328.99 ;
      RECT 10514.345 189.04 10514.625 328.75 ;
      RECT 10513.785 189.04 10514.065 328.51 ;
      RECT 10513.225 189.04 10513.505 328.27 ;
      RECT 10512.665 189.04 10512.945 328.03 ;
      RECT 10512.105 189.04 10512.385 327.79 ;
      RECT 10511.545 189.04 10511.825 327.55 ;
      RECT 10510.985 189.04 10511.265 327.31 ;
      RECT 10510.425 187.94 10510.705 327.07 ;
      RECT 10509.865 189.04 10510.145 326.83 ;
      RECT 10509.305 187.94 10509.585 326.59 ;
      RECT 10508.745 189.04 10509.025 326.35 ;
      RECT 10494.745 187.94 10495.025 332.47 ;
      RECT 10494.185 189.04 10494.465 332.23 ;
      RECT 10493.625 189.04 10493.905 331.99 ;
      RECT 10493.065 189.04 10493.345 331.75 ;
      RECT 10492.505 189.04 10492.785 331.51 ;
      RECT 10491.945 189.04 10492.225 331.27 ;
      RECT 10491.385 189.04 10491.665 331.03 ;
      RECT 10490.825 189.04 10491.105 330.79 ;
      RECT 10490.265 189.04 10490.545 330.55 ;
      RECT 10489.705 187.94 10489.985 330.31 ;
      RECT 10489.145 189.04 10489.425 330.07 ;
      RECT 10488.585 187.94 10488.865 329.83 ;
      RECT 10488.025 189.04 10488.305 329.59 ;
      RECT 10487.465 189.04 10487.745 329.35 ;
      RECT 10486.905 189.04 10487.185 329.11 ;
      RECT 10486.345 189.04 10486.625 328.87 ;
      RECT 10485.785 189.04 10486.065 328.63 ;
      RECT 10485.225 189.04 10485.505 328.39 ;
      RECT 10484.665 189.04 10484.945 328.15 ;
      RECT 10484.105 189.04 10484.385 327.91 ;
      RECT 10483.545 189.04 10483.825 327.67 ;
      RECT 10482.985 189.04 10483.265 327.43 ;
      RECT 10482.425 189.04 10482.705 327.19 ;
      RECT 10443.225 189.04 10443.505 334.095 ;
      RECT 10442.665 189.04 10442.945 334.335 ;
      RECT 10442.105 189.04 10442.385 334.575 ;
      RECT 10441.545 187.94 10441.825 334.815 ;
      RECT 10440.985 189.04 10441.265 335.055 ;
      RECT 10440.425 187.94 10440.705 335.295 ;
      RECT 10439.865 189.04 10440.145 335.535 ;
      RECT 10439.305 189.04 10439.585 335.775 ;
      RECT 10438.745 189.04 10439.025 336.015 ;
      RECT 10438.185 187.94 10438.465 336.255 ;
      RECT 10437.625 189.04 10437.905 336.495 ;
      RECT 10437.065 187.94 10437.345 336.735 ;
      RECT 10436.505 189.04 10436.785 336.975 ;
      RECT 10435.945 187.94 10436.225 337.215 ;
      RECT 10435.385 189.04 10435.665 337.455 ;
      RECT 10434.825 189.04 10435.105 337.695 ;
      RECT 10434.265 189.04 10434.545 337.695 ;
      RECT 10433.705 189.04 10433.985 337.455 ;
      RECT 10433.145 189.04 10433.425 337.215 ;
      RECT 10432.585 189.04 10432.865 336.975 ;
      RECT 10432.025 189.04 10432.305 336.735 ;
      RECT 10431.465 189.04 10431.745 336.495 ;
      RECT 10430.905 189.04 10431.185 336.255 ;
      RECT 10430.345 189.04 10430.625 336.015 ;
      RECT 10429.785 189.04 10430.065 335.775 ;
      RECT 10420.825 189.04 10421.105 335.29 ;
      RECT 10420.265 187.94 10420.545 335.05 ;
      RECT 10419.705 189.04 10419.985 334.81 ;
      RECT 10419.145 187.94 10419.425 334.57 ;
      RECT 10418.585 189.04 10418.865 334.33 ;
      RECT 10418.025 187.94 10418.305 334.09 ;
      RECT 10417.465 189.04 10417.745 333.85 ;
      RECT 10416.905 189.04 10417.185 333.61 ;
      RECT 10416.345 189.04 10416.625 333.37 ;
      RECT 10415.785 189.04 10416.065 333.13 ;
      RECT 10415.225 189.04 10415.505 332.89 ;
      RECT 10414.665 189.04 10414.945 332.65 ;
      RECT 10414.105 189.04 10414.385 332.41 ;
      RECT 10413.545 189.04 10413.825 332.17 ;
      RECT 10411.025 187.94 10411.305 333.89 ;
      RECT 10410.465 189.04 10410.745 333.65 ;
      RECT 10409.905 187.94 10410.185 333.41 ;
      RECT 10409.345 189.04 10409.625 333.17 ;
      RECT 10408.785 189.04 10409.065 332.93 ;
      RECT 10408.225 189.04 10408.505 332.69 ;
      RECT 10407.665 189.04 10407.945 332.45 ;
      RECT 10407.105 189.04 10407.385 332.21 ;
      RECT 10381.065 189.04 10381.345 329.86 ;
      RECT 10380.505 189.04 10380.785 330.1 ;
      RECT 10379.945 189.04 10380.225 330.34 ;
      RECT 10379.385 189.04 10379.665 330.585 ;
      RECT 10378.825 189.04 10379.105 330.825 ;
      RECT 10378.265 189.04 10378.545 331.065 ;
      RECT 10377.705 189.04 10377.985 331.065 ;
      RECT 10377.145 189.04 10377.425 330.825 ;
      RECT 10376.585 189.04 10376.865 330.585 ;
      RECT 10376.025 187.94 10376.305 330.345 ;
      RECT 10375.465 189.04 10375.745 330.105 ;
      RECT 10374.905 187.94 10375.185 329.865 ;
      RECT 10374.345 189.04 10374.625 329.625 ;
      RECT 10373.785 189.04 10374.065 329.385 ;
      RECT 10373.225 189.04 10373.505 329.145 ;
      RECT 10372.665 187.94 10372.945 328.905 ;
      RECT 10372.105 189.04 10372.385 328.665 ;
      RECT 10371.545 187.94 10371.825 328.425 ;
      RECT 10370.985 189.04 10371.265 328.185 ;
      RECT 10370.425 187.94 10370.705 327.945 ;
      RECT 10369.865 189.04 10370.145 327.705 ;
      RECT 10369.305 189.04 10369.585 327.465 ;
      RECT 10368.745 189.04 10369.025 327.225 ;
      RECT 10368.185 189.04 10368.465 326.985 ;
      RECT 10354.745 189.04 10355.025 332.785 ;
      RECT 10354.185 189.04 10354.465 332.545 ;
      RECT 10353.625 189.04 10353.905 332.305 ;
      RECT 10353.065 189.04 10353.345 332.065 ;
      RECT 10352.505 189.04 10352.785 331.825 ;
      RECT 10351.945 189.04 10352.225 331.585 ;
      RECT 10351.385 189.04 10351.665 331.345 ;
      RECT 10350.825 189.04 10351.105 331.105 ;
      RECT 10350.265 187.94 10350.545 330.865 ;
      RECT 10349.705 189.04 10349.985 330.625 ;
      RECT 10349.145 187.94 10349.425 330.305 ;
      RECT 10348.585 189.04 10348.865 330.145 ;
      RECT 10348.025 187.94 10348.305 329.905 ;
      RECT 10347.465 189.04 10347.745 329.665 ;
      RECT 10346.905 189.04 10347.185 329.425 ;
      RECT 10346.345 189.04 10346.625 329.185 ;
      RECT 10345.785 189.04 10346.065 328.945 ;
      RECT 10345.225 189.04 10345.505 328.705 ;
      RECT 10344.665 189.04 10344.945 328.465 ;
      RECT 10344.105 189.04 10344.385 328.225 ;
      RECT 10343.545 189.04 10343.825 327.985 ;
      RECT 10342.985 187.94 10343.265 327.745 ;
      RECT 10342.425 189.04 10342.705 327.505 ;
      RECT 10341.865 187.94 10342.145 327.265 ;
      RECT 10302.665 189.04 10302.945 332.875 ;
      RECT 10302.105 189.04 10302.385 333.115 ;
      RECT 10301.545 189.04 10301.825 333.355 ;
      RECT 10300.985 189.04 10301.265 333.595 ;
      RECT 10300.425 189.04 10300.705 333.835 ;
      RECT 10299.865 189.04 10300.145 334.075 ;
      RECT 10299.305 189.04 10299.585 334.315 ;
      RECT 10298.745 189.04 10299.025 334.555 ;
      RECT 10298.185 189.04 10298.465 334.795 ;
      RECT 10297.625 189.04 10297.905 335.035 ;
      RECT 10297.065 189.04 10297.345 335.275 ;
      RECT 10296.505 189.04 10296.785 335.515 ;
      RECT 10295.945 189.04 10296.225 335.755 ;
      RECT 10295.385 189.04 10295.665 335.755 ;
      RECT 10294.825 187.94 10295.105 335.515 ;
      RECT 10294.265 189.04 10294.545 335.275 ;
      RECT 10293.705 187.94 10293.985 335.035 ;
      RECT 10293.145 189.04 10293.425 334.795 ;
      RECT 10292.585 189.04 10292.865 334.555 ;
      RECT 10292.025 189.04 10292.305 334.315 ;
      RECT 10291.465 187.94 10291.745 334.05 ;
      RECT 10290.905 189.04 10291.185 333.81 ;
      RECT 10290.345 187.94 10290.625 333.57 ;
      RECT 10289.785 189.04 10290.065 333.33 ;
      RECT 10280.825 187.94 10281.105 327.165 ;
      RECT 10280.265 189.04 10280.545 327.405 ;
      RECT 10279.705 189.04 10279.985 327.645 ;
      RECT 10279.145 189.04 10279.425 327.645 ;
      RECT 10278.585 189.04 10278.865 327.405 ;
      RECT 10278.025 189.04 10278.305 327.165 ;
      RECT 10277.465 189.04 10277.745 326.925 ;
      RECT 10276.905 189.04 10277.185 326.685 ;
      RECT 10276.345 189.04 10276.625 326.445 ;
      RECT 10275.785 189.04 10276.065 326.205 ;
      RECT 10275.225 189.04 10275.505 325.965 ;
      RECT 10274.665 189.04 10274.945 325.725 ;
      RECT 10274.105 189.04 10274.385 325.485 ;
      RECT 10273.545 187.94 10273.825 325.245 ;
      RECT 10271.025 189.04 10271.305 326.965 ;
      RECT 10270.465 187.94 10270.745 326.725 ;
      RECT 10269.905 189.04 10270.185 326.485 ;
      RECT 10269.345 187.94 10269.625 326.245 ;
      RECT 10268.785 189.04 10269.065 326.005 ;
      RECT 10268.225 189.04 10268.505 325.765 ;
      RECT 10267.665 189.04 10267.945 325.525 ;
      RECT 10241.625 189.04 10241.905 328.31 ;
      RECT 10241.065 189.04 10241.345 328.55 ;
      RECT 10240.505 189.04 10240.785 328.79 ;
      RECT 10239.945 189.04 10240.225 329.03 ;
      RECT 10239.385 189.04 10239.665 329.27 ;
      RECT 10238.825 187.94 10239.105 329.51 ;
      RECT 10238.265 189.04 10238.545 329.75 ;
      RECT 10237.705 187.94 10237.985 329.99 ;
      RECT 10237.145 189.04 10237.425 330.23 ;
      RECT 10236.585 189.04 10236.865 330.47 ;
      RECT 10236.025 189.04 10236.305 330.71 ;
      RECT 10235.465 189.04 10235.745 330.95 ;
      RECT 10234.905 189.04 10235.185 331.19 ;
      RECT 10234.345 189.04 10234.625 331.43 ;
      RECT 10233.785 189.04 10234.065 331.67 ;
      RECT 10233.225 189.04 10233.505 331.67 ;
      RECT 10232.665 189.04 10232.945 331.43 ;
      RECT 10232.105 189.04 10232.385 331.19 ;
      RECT 10231.545 189.04 10231.825 330.95 ;
      RECT 10230.985 189.04 10231.265 330.705 ;
      RECT 10230.425 189.04 10230.705 330.465 ;
      RECT 10229.865 189.04 10230.145 330.225 ;
      RECT 10229.305 187.94 10229.585 329.985 ;
      RECT 10228.745 189.04 10229.025 329.745 ;
      RECT 10215.305 187.94 10215.585 327.225 ;
      RECT 10214.745 189.04 10215.025 326.985 ;
      RECT 10214.185 189.04 10214.465 326.745 ;
      RECT 10213.625 189.04 10213.905 326.505 ;
      RECT 10213.065 187.94 10213.345 326.265 ;
      RECT 10212.505 189.04 10212.785 326.025 ;
      RECT 10211.945 187.94 10212.225 325.785 ;
      RECT 10211.385 189.04 10211.665 325.545 ;
      RECT 10210.825 187.94 10211.105 325.305 ;
      RECT 10210.265 189.04 10210.545 325.065 ;
      RECT 10209.705 189.04 10209.985 324.825 ;
      RECT 10209.145 189.04 10209.425 324.585 ;
      RECT 10208.585 189.04 10208.865 324.345 ;
      RECT 10208.025 189.04 10208.305 324.105 ;
      RECT 10207.465 189.04 10207.745 323.865 ;
      RECT 10206.905 189.04 10207.185 323.625 ;
      RECT 10206.345 189.04 10206.625 323.385 ;
      RECT 10205.785 189.04 10206.065 323.145 ;
      RECT 10205.225 189.04 10205.505 322.905 ;
      RECT 10204.665 189.04 10204.945 322.665 ;
      RECT 10204.105 189.04 10204.385 322.425 ;
      RECT 10203.545 187.94 10203.825 322.185 ;
      RECT 10202.985 189.04 10203.265 321.945 ;
      RECT 10202.425 187.94 10202.705 321.705 ;
      RECT 10162.665 189.04 10162.945 332.175 ;
      RECT 10162.105 187.94 10162.385 332.415 ;
      RECT 10161.545 189.04 10161.825 332.655 ;
      RECT 10160.985 189.04 10161.265 332.895 ;
      RECT 10160.425 189.04 10160.705 333.135 ;
      RECT 10159.865 189.04 10160.145 333.375 ;
      RECT 10159.305 189.04 10159.585 333.615 ;
      RECT 10158.745 189.04 10159.025 333.86 ;
      RECT 10158.185 189.04 10158.465 334.1 ;
      RECT 10157.625 189.04 10157.905 334.34 ;
      RECT 10157.065 187.94 10157.345 334.58 ;
      RECT 10156.505 189.04 10156.785 334.82 ;
      RECT 10155.945 187.94 10156.225 335.06 ;
      RECT 10155.385 189.04 10155.665 335.3 ;
      RECT 10154.825 189.04 10155.105 335.54 ;
      RECT 10154.265 189.04 10154.545 335.78 ;
      RECT 10153.705 189.04 10153.985 336.02 ;
      RECT 10153.145 189.04 10153.425 336.26 ;
      RECT 10152.585 189.04 10152.865 336.5 ;
      RECT 10152.025 189.04 10152.305 336.74 ;
      RECT 10151.465 189.04 10151.745 336.98 ;
      RECT 10150.905 189.04 10151.185 337.22 ;
      RECT 10150.345 189.04 10150.625 337.46 ;
      RECT 10149.785 189.04 10150.065 337.7 ;
      RECT 10140.825 189.04 10141.105 333.285 ;
      RECT 10140.265 189.04 10140.545 333.045 ;
      RECT 10139.705 189.04 10139.985 332.805 ;
      RECT 10139.145 187.94 10139.425 332.565 ;
      RECT 10138.585 189.04 10138.865 332.325 ;
      RECT 10138.025 187.94 10138.305 332.085 ;
      RECT 10137.465 189.04 10137.745 331.845 ;
      RECT 10136.905 189.04 10137.185 331.605 ;
      RECT 10136.345 189.04 10136.625 331.365 ;
      RECT 10135.785 187.94 10136.065 331.125 ;
      RECT 10135.225 189.04 10135.505 330.885 ;
      RECT 10134.665 187.94 10134.945 330.645 ;
      RECT 10134.105 189.04 10134.385 330.405 ;
      RECT 10133.545 187.94 10133.825 330.165 ;
      RECT 10131.025 189.04 10131.305 322.565 ;
      RECT 10130.465 189.04 10130.745 322.325 ;
      RECT 10129.905 189.04 10130.185 322.085 ;
      RECT 10129.345 189.04 10129.625 321.845 ;
      RECT 10128.785 189.04 10129.065 321.605 ;
      RECT 10128.225 189.04 10128.505 321.365 ;
      RECT 10127.665 189.04 10127.945 321.125 ;
      RECT 10101.625 189.04 10101.905 335 ;
      RECT 10101.065 189.04 10101.345 335.24 ;
      RECT 10100.505 189.04 10100.785 335.48 ;
      RECT 10099.945 189.04 10100.225 335.72 ;
      RECT 10099.385 189.04 10099.665 335.96 ;
      RECT 10098.825 187.94 10099.105 335.96 ;
      RECT 10098.265 189.04 10098.545 335.72 ;
      RECT 10097.705 187.94 10097.985 335.475 ;
      RECT 10097.145 189.04 10097.425 335.235 ;
      RECT 10096.585 187.94 10096.865 334.995 ;
      RECT 10096.025 189.04 10096.305 334.755 ;
      RECT 10095.465 189.04 10095.745 334.515 ;
      RECT 10094.905 189.04 10095.185 334.275 ;
      RECT 10094.345 189.04 10094.625 334.035 ;
      RECT 10093.785 189.04 10094.065 333.795 ;
      RECT 10093.225 189.04 10093.505 333.555 ;
      RECT 10092.665 189.04 10092.945 333.315 ;
      RECT 10092.105 189.04 10092.385 333.075 ;
      RECT 10091.545 187.94 10091.825 332.835 ;
      RECT 10090.985 189.04 10091.265 332.595 ;
      RECT 10090.425 187.94 10090.705 332.355 ;
      RECT 10089.865 189.04 10090.145 332.115 ;
      RECT 10089.305 189.04 10089.585 331.875 ;
      RECT 10088.745 189.04 10089.025 331.635 ;
      RECT 10075.305 189.04 10075.585 335.035 ;
      RECT 10074.745 189.04 10075.025 335.275 ;
      RECT 10074.185 189.04 10074.465 335.52 ;
      RECT 10073.625 189.04 10073.905 335.76 ;
      RECT 10073.065 189.04 10073.345 336 ;
      RECT 10072.505 189.04 10072.785 336 ;
      RECT 10071.945 189.04 10072.225 335.76 ;
      RECT 10071.385 189.04 10071.665 335.52 ;
      RECT 10070.825 189.04 10071.105 328.505 ;
      RECT 10070.265 189.04 10070.545 328.265 ;
      RECT 10069.705 189.04 10069.985 328.025 ;
      RECT 10069.145 187.94 10069.425 327.785 ;
      RECT 10068.585 189.04 10068.865 327.545 ;
      RECT 10068.025 187.94 10068.305 327.305 ;
      RECT 10067.465 189.04 10067.745 327.065 ;
      RECT 10066.905 189.04 10067.185 326.825 ;
      RECT 10066.345 189.04 10066.625 326.585 ;
      RECT 10065.785 187.94 10066.065 326.345 ;
      RECT 10065.225 189.04 10065.505 326.105 ;
      RECT 10064.665 187.94 10064.945 325.865 ;
      RECT 10064.105 189.04 10064.385 325.625 ;
      RECT 10063.545 187.94 10063.825 325.385 ;
      RECT 10062.985 189.04 10063.265 325.145 ;
      RECT 10062.425 189.04 10062.705 324.905 ;
      RECT 10022.105 189.04 10022.385 333.8 ;
      RECT 10021.545 189.04 10021.825 334.04 ;
      RECT 10020.985 189.04 10021.265 334.285 ;
      RECT 10020.425 189.04 10020.705 334.525 ;
      RECT 10019.865 189.04 10020.145 334.765 ;
      RECT 10019.305 189.04 10019.585 335.005 ;
      RECT 10018.745 189.04 10019.025 335.245 ;
      RECT 10018.185 189.04 10018.465 335.485 ;
      RECT 10017.625 189.04 10017.905 335.725 ;
      RECT 10017.065 189.04 10017.345 335.965 ;
      RECT 10016.505 187.94 10016.785 336.205 ;
      RECT 10015.945 189.04 10016.225 336.445 ;
      RECT 10015.385 187.94 10015.665 336.685 ;
      RECT 10014.825 189.04 10015.105 336.925 ;
      RECT 10014.265 187.94 10014.545 337.165 ;
      RECT 10013.705 189.04 10013.985 337.165 ;
      RECT 10013.145 189.04 10013.425 336.925 ;
      RECT 10012.585 189.04 10012.865 336.685 ;
      RECT 10012.025 189.04 10012.305 336.445 ;
      RECT 10011.465 189.04 10011.745 336.205 ;
      RECT 10010.905 189.04 10011.185 335.965 ;
      RECT 10010.345 189.04 10010.625 335.725 ;
      RECT 10009.785 189.04 10010.065 335.485 ;
      RECT 10000.825 187.94 10001.105 335.515 ;
      RECT 10000.265 189.04 10000.545 335.755 ;
      RECT 9999.705 187.94 9999.985 335.995 ;
      RECT 9999.145 189.04 9999.425 336.21 ;
      RECT 9998.585 189.04 9998.865 335.785 ;
      RECT 9998.025 189.04 9998.305 335.545 ;
      RECT 9997.465 189.04 9997.745 335.305 ;
      RECT 9996.905 189.04 9997.185 335.065 ;
      RECT 9996.345 189.04 9996.625 334.825 ;
      RECT 9995.785 189.04 9996.065 334.585 ;
      RECT 9995.225 189.04 9995.505 334.345 ;
      RECT 9994.665 189.04 9994.945 334.105 ;
      RECT 9994.105 189.04 9994.385 333.865 ;
      RECT 9993.545 189.04 9993.825 333.625 ;
      RECT 9991.025 189.04 9991.305 332.8 ;
      RECT 9990.465 189.04 9990.745 332.56 ;
      RECT 9989.905 189.04 9990.185 332.32 ;
      RECT 9989.345 187.94 9989.625 332.08 ;
      RECT 9988.785 189.04 9989.065 331.84 ;
      RECT 9988.225 187.94 9988.505 331.6 ;
      RECT 9987.665 189.04 9987.945 331.36 ;
      RECT 9987.105 189.04 9987.385 331.12 ;
      RECT 9960.505 189.04 9960.785 342.165 ;
      RECT 9959.945 187.94 9960.225 342.405 ;
      RECT 9959.385 189.04 9959.665 342.645 ;
      RECT 9958.825 187.94 9959.105 342.89 ;
      RECT 9958.265 189.04 9958.545 343.13 ;
      RECT 9957.705 187.94 9957.985 343.37 ;
      RECT 9957.145 189.04 9957.425 343.61 ;
      RECT 9956.585 189.04 9956.865 343.85 ;
      RECT 9956.025 189.04 9956.305 329.47 ;
      RECT 9955.465 189.04 9955.745 329.23 ;
      RECT 9954.905 189.04 9955.185 328.99 ;
      RECT 9954.345 189.04 9954.625 328.75 ;
      RECT 9953.785 189.04 9954.065 328.51 ;
      RECT 9953.225 189.04 9953.505 328.27 ;
      RECT 9952.665 189.04 9952.945 328.03 ;
      RECT 9952.105 189.04 9952.385 327.79 ;
      RECT 9951.545 189.04 9951.825 327.55 ;
      RECT 9950.985 189.04 9951.265 327.31 ;
      RECT 9950.425 187.94 9950.705 327.07 ;
      RECT 9949.865 189.04 9950.145 326.83 ;
      RECT 9949.305 187.94 9949.585 326.59 ;
      RECT 9948.745 189.04 9949.025 326.35 ;
      RECT 9934.745 187.94 9935.025 332.47 ;
      RECT 9934.185 189.04 9934.465 332.23 ;
      RECT 9933.625 189.04 9933.905 331.99 ;
      RECT 9933.065 189.04 9933.345 331.75 ;
      RECT 9932.505 189.04 9932.785 331.51 ;
      RECT 9931.945 189.04 9932.225 331.27 ;
      RECT 9931.385 189.04 9931.665 331.03 ;
      RECT 9930.825 189.04 9931.105 330.79 ;
      RECT 9930.265 189.04 9930.545 330.55 ;
      RECT 9929.705 187.94 9929.985 330.31 ;
      RECT 9929.145 189.04 9929.425 330.07 ;
      RECT 9928.585 187.94 9928.865 329.83 ;
      RECT 9928.025 189.04 9928.305 329.59 ;
      RECT 9927.465 189.04 9927.745 329.35 ;
      RECT 9926.905 189.04 9927.185 329.11 ;
      RECT 9926.345 189.04 9926.625 328.87 ;
      RECT 9925.785 189.04 9926.065 328.63 ;
      RECT 9925.225 189.04 9925.505 328.39 ;
      RECT 9924.665 189.04 9924.945 328.15 ;
      RECT 9924.105 189.04 9924.385 327.91 ;
      RECT 9923.545 189.04 9923.825 327.67 ;
      RECT 9922.985 189.04 9923.265 327.43 ;
      RECT 9922.425 189.04 9922.705 327.19 ;
      RECT 9883.225 189.04 9883.505 334.095 ;
      RECT 9882.665 189.04 9882.945 334.335 ;
      RECT 9882.105 189.04 9882.385 334.575 ;
      RECT 9881.545 187.94 9881.825 334.815 ;
      RECT 9880.985 189.04 9881.265 335.055 ;
      RECT 9880.425 187.94 9880.705 335.295 ;
      RECT 9879.865 189.04 9880.145 335.535 ;
      RECT 9879.305 189.04 9879.585 335.775 ;
      RECT 9878.745 189.04 9879.025 336.015 ;
      RECT 9878.185 187.94 9878.465 336.255 ;
      RECT 9877.625 189.04 9877.905 336.495 ;
      RECT 9877.065 187.94 9877.345 336.735 ;
      RECT 9876.505 189.04 9876.785 336.975 ;
      RECT 9875.945 187.94 9876.225 337.215 ;
      RECT 9875.385 189.04 9875.665 337.455 ;
      RECT 9874.825 189.04 9875.105 337.695 ;
      RECT 9874.265 189.04 9874.545 337.695 ;
      RECT 9873.705 189.04 9873.985 337.455 ;
      RECT 9873.145 189.04 9873.425 337.215 ;
      RECT 9872.585 189.04 9872.865 336.975 ;
      RECT 9872.025 189.04 9872.305 336.735 ;
      RECT 9871.465 189.04 9871.745 336.495 ;
      RECT 9870.905 189.04 9871.185 336.255 ;
      RECT 9870.345 189.04 9870.625 336.015 ;
      RECT 9869.785 189.04 9870.065 335.775 ;
      RECT 9860.825 189.04 9861.105 335.29 ;
      RECT 9860.265 187.94 9860.545 335.05 ;
      RECT 9859.705 189.04 9859.985 334.81 ;
      RECT 9859.145 187.94 9859.425 334.57 ;
      RECT 9858.585 189.04 9858.865 334.33 ;
      RECT 9858.025 187.94 9858.305 334.09 ;
      RECT 9857.465 189.04 9857.745 333.85 ;
      RECT 9856.905 189.04 9857.185 333.61 ;
      RECT 9856.345 189.04 9856.625 333.37 ;
      RECT 9855.785 189.04 9856.065 333.13 ;
      RECT 9855.225 189.04 9855.505 332.89 ;
      RECT 9854.665 189.04 9854.945 332.65 ;
      RECT 9854.105 189.04 9854.385 332.41 ;
      RECT 9853.545 189.04 9853.825 332.17 ;
      RECT 9851.025 187.94 9851.305 333.89 ;
      RECT 9850.465 189.04 9850.745 333.65 ;
      RECT 9849.905 187.94 9850.185 333.41 ;
      RECT 9849.345 189.04 9849.625 333.17 ;
      RECT 9848.785 189.04 9849.065 332.93 ;
      RECT 9848.225 189.04 9848.505 332.69 ;
      RECT 9847.665 189.04 9847.945 332.45 ;
      RECT 9847.105 189.04 9847.385 332.21 ;
      RECT 9821.065 189.04 9821.345 329.86 ;
      RECT 9820.505 189.04 9820.785 330.1 ;
      RECT 9819.945 189.04 9820.225 330.34 ;
      RECT 9819.385 189.04 9819.665 330.585 ;
      RECT 9818.825 189.04 9819.105 330.825 ;
      RECT 9818.265 189.04 9818.545 331.065 ;
      RECT 9817.705 189.04 9817.985 331.065 ;
      RECT 9817.145 189.04 9817.425 330.825 ;
      RECT 9816.585 189.04 9816.865 330.585 ;
      RECT 9816.025 187.94 9816.305 330.345 ;
      RECT 9815.465 189.04 9815.745 330.105 ;
      RECT 9814.905 187.94 9815.185 329.865 ;
      RECT 9814.345 189.04 9814.625 329.625 ;
      RECT 9813.785 189.04 9814.065 329.385 ;
      RECT 9813.225 189.04 9813.505 329.145 ;
      RECT 9812.665 187.94 9812.945 328.905 ;
      RECT 9812.105 189.04 9812.385 328.665 ;
      RECT 9811.545 187.94 9811.825 328.425 ;
      RECT 9810.985 189.04 9811.265 328.185 ;
      RECT 9810.425 187.94 9810.705 327.945 ;
      RECT 9809.865 189.04 9810.145 327.705 ;
      RECT 9809.305 189.04 9809.585 327.465 ;
      RECT 9808.745 189.04 9809.025 327.225 ;
      RECT 9808.185 189.04 9808.465 326.985 ;
      RECT 9794.745 189.04 9795.025 332.785 ;
      RECT 9794.185 189.04 9794.465 332.545 ;
      RECT 9793.625 189.04 9793.905 332.305 ;
      RECT 9793.065 189.04 9793.345 332.065 ;
      RECT 9792.505 189.04 9792.785 331.825 ;
      RECT 9791.945 189.04 9792.225 331.585 ;
      RECT 9791.385 189.04 9791.665 331.345 ;
      RECT 9790.825 189.04 9791.105 331.105 ;
      RECT 9790.265 187.94 9790.545 330.865 ;
      RECT 9789.705 189.04 9789.985 330.625 ;
      RECT 9789.145 187.94 9789.425 330.305 ;
      RECT 9788.585 189.04 9788.865 330.145 ;
      RECT 9788.025 187.94 9788.305 329.905 ;
      RECT 9787.465 189.04 9787.745 329.665 ;
      RECT 9786.905 189.04 9787.185 329.425 ;
      RECT 9786.345 189.04 9786.625 329.185 ;
      RECT 9785.785 189.04 9786.065 328.945 ;
      RECT 9785.225 189.04 9785.505 328.705 ;
      RECT 9784.665 189.04 9784.945 328.465 ;
      RECT 9784.105 189.04 9784.385 328.225 ;
      RECT 9783.545 189.04 9783.825 327.985 ;
      RECT 9782.985 187.94 9783.265 327.745 ;
      RECT 9782.425 189.04 9782.705 327.505 ;
      RECT 9781.865 187.94 9782.145 327.265 ;
      RECT 9742.665 189.04 9742.945 332.875 ;
      RECT 9742.105 189.04 9742.385 333.115 ;
      RECT 9741.545 189.04 9741.825 333.355 ;
      RECT 9740.985 189.04 9741.265 333.595 ;
      RECT 9740.425 189.04 9740.705 333.835 ;
      RECT 9739.865 189.04 9740.145 334.075 ;
      RECT 9739.305 189.04 9739.585 334.315 ;
      RECT 9738.745 189.04 9739.025 334.555 ;
      RECT 9738.185 189.04 9738.465 334.795 ;
      RECT 9737.625 189.04 9737.905 335.035 ;
      RECT 9737.065 189.04 9737.345 335.275 ;
      RECT 9736.505 189.04 9736.785 335.515 ;
      RECT 9735.945 189.04 9736.225 335.755 ;
      RECT 9735.385 189.04 9735.665 335.755 ;
      RECT 9734.825 187.94 9735.105 335.515 ;
      RECT 9734.265 189.04 9734.545 335.275 ;
      RECT 9733.705 187.94 9733.985 335.035 ;
      RECT 9733.145 189.04 9733.425 334.795 ;
      RECT 9732.585 189.04 9732.865 334.555 ;
      RECT 9732.025 189.04 9732.305 334.315 ;
      RECT 9731.465 187.94 9731.745 334.05 ;
      RECT 9730.905 189.04 9731.185 333.81 ;
      RECT 9730.345 187.94 9730.625 333.57 ;
      RECT 9729.785 189.04 9730.065 333.33 ;
      RECT 9720.825 187.94 9721.105 327.165 ;
      RECT 9720.265 189.04 9720.545 327.405 ;
      RECT 9719.705 189.04 9719.985 327.645 ;
      RECT 9719.145 189.04 9719.425 327.645 ;
      RECT 9718.585 189.04 9718.865 327.405 ;
      RECT 9718.025 189.04 9718.305 327.165 ;
      RECT 9717.465 189.04 9717.745 326.925 ;
      RECT 9716.905 189.04 9717.185 326.685 ;
      RECT 9716.345 189.04 9716.625 326.445 ;
      RECT 9715.785 189.04 9716.065 326.205 ;
      RECT 9715.225 189.04 9715.505 325.965 ;
      RECT 9714.665 189.04 9714.945 325.725 ;
      RECT 9714.105 189.04 9714.385 325.485 ;
      RECT 9713.545 187.94 9713.825 325.245 ;
      RECT 9711.025 189.04 9711.305 326.965 ;
      RECT 9710.465 187.94 9710.745 326.725 ;
      RECT 9709.905 189.04 9710.185 326.485 ;
      RECT 9709.345 187.94 9709.625 326.245 ;
      RECT 9708.785 189.04 9709.065 326.005 ;
      RECT 9708.225 189.04 9708.505 325.765 ;
      RECT 9707.665 189.04 9707.945 325.525 ;
      RECT 9681.625 189.04 9681.905 328.31 ;
      RECT 9681.065 189.04 9681.345 328.55 ;
      RECT 9680.505 189.04 9680.785 328.79 ;
      RECT 9679.945 189.04 9680.225 329.03 ;
      RECT 9679.385 189.04 9679.665 329.27 ;
      RECT 9678.825 187.94 9679.105 329.51 ;
      RECT 9678.265 189.04 9678.545 329.75 ;
      RECT 9677.705 187.94 9677.985 329.99 ;
      RECT 9677.145 189.04 9677.425 330.23 ;
      RECT 9676.585 189.04 9676.865 330.47 ;
      RECT 9676.025 189.04 9676.305 330.71 ;
      RECT 9675.465 189.04 9675.745 330.95 ;
      RECT 9674.905 189.04 9675.185 331.19 ;
      RECT 9674.345 189.04 9674.625 331.43 ;
      RECT 9673.785 189.04 9674.065 331.67 ;
      RECT 9673.225 189.04 9673.505 331.67 ;
      RECT 9672.665 189.04 9672.945 331.43 ;
      RECT 9672.105 189.04 9672.385 331.19 ;
      RECT 9671.545 189.04 9671.825 330.95 ;
      RECT 9670.985 189.04 9671.265 330.705 ;
      RECT 9670.425 189.04 9670.705 330.465 ;
      RECT 9669.865 189.04 9670.145 330.225 ;
      RECT 9669.305 187.94 9669.585 329.985 ;
      RECT 9668.745 189.04 9669.025 329.745 ;
      RECT 9655.305 187.94 9655.585 327.225 ;
      RECT 9654.745 189.04 9655.025 326.985 ;
      RECT 9654.185 189.04 9654.465 326.745 ;
      RECT 9653.625 189.04 9653.905 326.505 ;
      RECT 9653.065 187.94 9653.345 326.265 ;
      RECT 9652.505 189.04 9652.785 326.025 ;
      RECT 9651.945 187.94 9652.225 325.785 ;
      RECT 9651.385 189.04 9651.665 325.545 ;
      RECT 9650.825 187.94 9651.105 325.305 ;
      RECT 9650.265 189.04 9650.545 325.065 ;
      RECT 9649.705 189.04 9649.985 324.825 ;
      RECT 9649.145 189.04 9649.425 324.585 ;
      RECT 9648.585 189.04 9648.865 324.345 ;
      RECT 9648.025 189.04 9648.305 324.105 ;
      RECT 9647.465 189.04 9647.745 323.865 ;
      RECT 9646.905 189.04 9647.185 323.625 ;
      RECT 9646.345 189.04 9646.625 323.385 ;
      RECT 9645.785 189.04 9646.065 323.145 ;
      RECT 9645.225 189.04 9645.505 322.905 ;
      RECT 9644.665 189.04 9644.945 322.665 ;
      RECT 9644.105 189.04 9644.385 322.425 ;
      RECT 9643.545 187.94 9643.825 322.185 ;
      RECT 9642.985 189.04 9643.265 321.945 ;
      RECT 9642.425 187.94 9642.705 321.705 ;
      RECT 9602.665 189.04 9602.945 332.175 ;
      RECT 9602.105 187.94 9602.385 332.415 ;
      RECT 9601.545 189.04 9601.825 332.655 ;
      RECT 9600.985 189.04 9601.265 332.895 ;
      RECT 9600.425 189.04 9600.705 333.135 ;
      RECT 9599.865 189.04 9600.145 333.375 ;
      RECT 9599.305 189.04 9599.585 333.615 ;
      RECT 9598.745 189.04 9599.025 333.86 ;
      RECT 9598.185 189.04 9598.465 334.1 ;
      RECT 9597.625 189.04 9597.905 334.34 ;
      RECT 9597.065 187.94 9597.345 334.58 ;
      RECT 9596.505 189.04 9596.785 334.82 ;
      RECT 9595.945 187.94 9596.225 335.06 ;
      RECT 9595.385 189.04 9595.665 335.3 ;
      RECT 9594.825 189.04 9595.105 335.54 ;
      RECT 9594.265 189.04 9594.545 335.78 ;
      RECT 9593.705 189.04 9593.985 336.02 ;
      RECT 9593.145 189.04 9593.425 336.26 ;
      RECT 9592.585 189.04 9592.865 336.5 ;
      RECT 9592.025 189.04 9592.305 336.74 ;
      RECT 9591.465 189.04 9591.745 336.98 ;
      RECT 9590.905 189.04 9591.185 337.22 ;
      RECT 9590.345 189.04 9590.625 337.46 ;
      RECT 9589.785 189.04 9590.065 337.7 ;
      RECT 9580.825 189.04 9581.105 333.285 ;
      RECT 9580.265 189.04 9580.545 333.045 ;
      RECT 9579.705 189.04 9579.985 332.805 ;
      RECT 9579.145 187.94 9579.425 332.565 ;
      RECT 9578.585 189.04 9578.865 332.325 ;
      RECT 9578.025 187.94 9578.305 332.085 ;
      RECT 9577.465 189.04 9577.745 331.845 ;
      RECT 9576.905 189.04 9577.185 331.605 ;
      RECT 9576.345 189.04 9576.625 331.365 ;
      RECT 9575.785 187.94 9576.065 331.125 ;
      RECT 9575.225 189.04 9575.505 330.885 ;
      RECT 9574.665 187.94 9574.945 330.645 ;
      RECT 9574.105 189.04 9574.385 330.405 ;
      RECT 9573.545 187.94 9573.825 330.165 ;
      RECT 9571.025 189.04 9571.305 322.565 ;
      RECT 9570.465 189.04 9570.745 322.325 ;
      RECT 9569.905 189.04 9570.185 322.085 ;
      RECT 9569.345 189.04 9569.625 321.845 ;
      RECT 9568.785 189.04 9569.065 321.605 ;
      RECT 9568.225 189.04 9568.505 321.365 ;
      RECT 9567.665 189.04 9567.945 321.125 ;
      RECT 9541.625 189.04 9541.905 335 ;
      RECT 9541.065 189.04 9541.345 335.24 ;
      RECT 9540.505 189.04 9540.785 335.48 ;
      RECT 9539.945 189.04 9540.225 335.72 ;
      RECT 9539.385 189.04 9539.665 335.96 ;
      RECT 9538.825 187.94 9539.105 335.96 ;
      RECT 9538.265 189.04 9538.545 335.72 ;
      RECT 9537.705 187.94 9537.985 335.475 ;
      RECT 9537.145 189.04 9537.425 335.235 ;
      RECT 9536.585 187.94 9536.865 334.995 ;
      RECT 9536.025 189.04 9536.305 334.755 ;
      RECT 9535.465 189.04 9535.745 334.515 ;
      RECT 9534.905 189.04 9535.185 334.275 ;
      RECT 9534.345 189.04 9534.625 334.035 ;
      RECT 9533.785 189.04 9534.065 333.795 ;
      RECT 9533.225 189.04 9533.505 333.555 ;
      RECT 9532.665 189.04 9532.945 333.315 ;
      RECT 9532.105 189.04 9532.385 333.075 ;
      RECT 9531.545 187.94 9531.825 332.835 ;
      RECT 9530.985 189.04 9531.265 332.595 ;
      RECT 9530.425 187.94 9530.705 332.355 ;
      RECT 9529.865 189.04 9530.145 332.115 ;
      RECT 9529.305 189.04 9529.585 331.875 ;
      RECT 9528.745 189.04 9529.025 331.635 ;
      RECT 9515.305 189.04 9515.585 335.035 ;
      RECT 9514.745 189.04 9515.025 335.275 ;
      RECT 9514.185 189.04 9514.465 335.52 ;
      RECT 9513.625 189.04 9513.905 335.76 ;
      RECT 9513.065 189.04 9513.345 336 ;
      RECT 9512.505 189.04 9512.785 336 ;
      RECT 9511.945 189.04 9512.225 335.76 ;
      RECT 9511.385 189.04 9511.665 335.52 ;
      RECT 9510.825 189.04 9511.105 328.505 ;
      RECT 9510.265 189.04 9510.545 328.265 ;
      RECT 9509.705 189.04 9509.985 328.025 ;
      RECT 9509.145 187.94 9509.425 327.785 ;
      RECT 9508.585 189.04 9508.865 327.545 ;
      RECT 9508.025 187.94 9508.305 327.305 ;
      RECT 9507.465 189.04 9507.745 327.065 ;
      RECT 9506.905 189.04 9507.185 326.825 ;
      RECT 9506.345 189.04 9506.625 326.585 ;
      RECT 9505.785 187.94 9506.065 326.345 ;
      RECT 9505.225 189.04 9505.505 326.105 ;
      RECT 9504.665 187.94 9504.945 325.865 ;
      RECT 9504.105 189.04 9504.385 325.625 ;
      RECT 9503.545 187.94 9503.825 325.385 ;
      RECT 9502.985 189.04 9503.265 325.145 ;
      RECT 9502.425 189.04 9502.705 324.905 ;
      RECT 9462.105 189.04 9462.385 333.8 ;
      RECT 9461.545 189.04 9461.825 334.04 ;
      RECT 9460.985 189.04 9461.265 334.285 ;
      RECT 9460.425 189.04 9460.705 334.525 ;
      RECT 9459.865 189.04 9460.145 334.765 ;
      RECT 9459.305 189.04 9459.585 335.005 ;
      RECT 9458.745 189.04 9459.025 335.245 ;
      RECT 9458.185 189.04 9458.465 335.485 ;
      RECT 9457.625 189.04 9457.905 335.725 ;
      RECT 9457.065 189.04 9457.345 335.965 ;
      RECT 9456.505 187.94 9456.785 336.205 ;
      RECT 9455.945 189.04 9456.225 336.445 ;
      RECT 9455.385 187.94 9455.665 336.685 ;
      RECT 9454.825 189.04 9455.105 336.925 ;
      RECT 9454.265 187.94 9454.545 337.165 ;
      RECT 9453.705 189.04 9453.985 337.165 ;
      RECT 9453.145 189.04 9453.425 336.925 ;
      RECT 9452.585 189.04 9452.865 336.685 ;
      RECT 9452.025 189.04 9452.305 336.445 ;
      RECT 9451.465 189.04 9451.745 336.205 ;
      RECT 9450.905 189.04 9451.185 335.965 ;
      RECT 9450.345 189.04 9450.625 335.725 ;
      RECT 9449.785 189.04 9450.065 335.485 ;
      RECT 9440.825 187.94 9441.105 335.515 ;
      RECT 9440.265 189.04 9440.545 335.755 ;
      RECT 9439.705 187.94 9439.985 335.995 ;
      RECT 9439.145 189.04 9439.425 336.21 ;
      RECT 9438.585 189.04 9438.865 335.785 ;
      RECT 9438.025 189.04 9438.305 335.545 ;
      RECT 9437.465 189.04 9437.745 335.305 ;
      RECT 9436.905 189.04 9437.185 335.065 ;
      RECT 9436.345 189.04 9436.625 334.825 ;
      RECT 9435.785 189.04 9436.065 334.585 ;
      RECT 9435.225 189.04 9435.505 334.345 ;
      RECT 9434.665 189.04 9434.945 334.105 ;
      RECT 9434.105 189.04 9434.385 333.865 ;
      RECT 9433.545 189.04 9433.825 333.625 ;
      RECT 9431.025 189.04 9431.305 332.8 ;
      RECT 9430.465 189.04 9430.745 332.56 ;
      RECT 9429.905 189.04 9430.185 332.32 ;
      RECT 9429.345 187.94 9429.625 332.08 ;
      RECT 9428.785 189.04 9429.065 331.84 ;
      RECT 9428.225 187.94 9428.505 331.6 ;
      RECT 9427.665 189.04 9427.945 331.36 ;
      RECT 9427.105 189.04 9427.385 331.12 ;
      RECT 9400.505 189.04 9400.785 342.165 ;
      RECT 9399.945 187.94 9400.225 342.405 ;
      RECT 9399.385 189.04 9399.665 342.645 ;
      RECT 9398.825 187.94 9399.105 342.89 ;
      RECT 9398.265 189.04 9398.545 343.13 ;
      RECT 9397.705 187.94 9397.985 343.37 ;
      RECT 9397.145 189.04 9397.425 343.61 ;
      RECT 9396.585 189.04 9396.865 343.85 ;
      RECT 9396.025 189.04 9396.305 329.47 ;
      RECT 9395.465 189.04 9395.745 329.23 ;
      RECT 9394.905 189.04 9395.185 328.99 ;
      RECT 9394.345 189.04 9394.625 328.75 ;
      RECT 9393.785 189.04 9394.065 328.51 ;
      RECT 9393.225 189.04 9393.505 328.27 ;
      RECT 9392.665 189.04 9392.945 328.03 ;
      RECT 9392.105 189.04 9392.385 327.79 ;
      RECT 9391.545 189.04 9391.825 327.55 ;
      RECT 9390.985 189.04 9391.265 327.31 ;
      RECT 9390.425 187.94 9390.705 327.07 ;
      RECT 9389.865 189.04 9390.145 326.83 ;
      RECT 9389.305 187.94 9389.585 326.59 ;
      RECT 9388.745 189.04 9389.025 326.35 ;
      RECT 9374.745 187.94 9375.025 332.47 ;
      RECT 9374.185 189.04 9374.465 332.23 ;
      RECT 9373.625 189.04 9373.905 331.99 ;
      RECT 9373.065 189.04 9373.345 331.75 ;
      RECT 9372.505 189.04 9372.785 331.51 ;
      RECT 9371.945 189.04 9372.225 331.27 ;
      RECT 9371.385 189.04 9371.665 331.03 ;
      RECT 9370.825 189.04 9371.105 330.79 ;
      RECT 9370.265 189.04 9370.545 330.55 ;
      RECT 9369.705 187.94 9369.985 330.31 ;
      RECT 9369.145 189.04 9369.425 330.07 ;
      RECT 9368.585 187.94 9368.865 329.83 ;
      RECT 9368.025 189.04 9368.305 329.59 ;
      RECT 9367.465 189.04 9367.745 329.35 ;
      RECT 9366.905 189.04 9367.185 329.11 ;
      RECT 9366.345 189.04 9366.625 328.87 ;
      RECT 9365.785 189.04 9366.065 328.63 ;
      RECT 9365.225 189.04 9365.505 328.39 ;
      RECT 9364.665 189.04 9364.945 328.15 ;
      RECT 9364.105 189.04 9364.385 327.91 ;
      RECT 9363.545 189.04 9363.825 327.67 ;
      RECT 9362.985 189.04 9363.265 327.43 ;
      RECT 9362.425 189.04 9362.705 327.19 ;
      RECT 9323.225 189.04 9323.505 334.095 ;
      RECT 9322.665 189.04 9322.945 334.335 ;
      RECT 9322.105 189.04 9322.385 334.575 ;
      RECT 9321.545 187.94 9321.825 334.815 ;
      RECT 9320.985 189.04 9321.265 335.055 ;
      RECT 9320.425 187.94 9320.705 335.295 ;
      RECT 9319.865 189.04 9320.145 335.535 ;
      RECT 9319.305 189.04 9319.585 335.775 ;
      RECT 9318.745 189.04 9319.025 336.015 ;
      RECT 9318.185 187.94 9318.465 336.255 ;
      RECT 9317.625 189.04 9317.905 336.495 ;
      RECT 9317.065 187.94 9317.345 336.735 ;
      RECT 9316.505 189.04 9316.785 336.975 ;
      RECT 9315.945 187.94 9316.225 337.215 ;
      RECT 9315.385 189.04 9315.665 337.455 ;
      RECT 9314.825 189.04 9315.105 337.695 ;
      RECT 9314.265 189.04 9314.545 337.695 ;
      RECT 9313.705 189.04 9313.985 337.455 ;
      RECT 9313.145 189.04 9313.425 337.215 ;
      RECT 9312.585 189.04 9312.865 336.975 ;
      RECT 9312.025 189.04 9312.305 336.735 ;
      RECT 9311.465 189.04 9311.745 336.495 ;
      RECT 9310.905 189.04 9311.185 336.255 ;
      RECT 9310.345 189.04 9310.625 336.015 ;
      RECT 9309.785 189.04 9310.065 335.775 ;
      RECT 9300.825 189.04 9301.105 335.29 ;
      RECT 9300.265 187.94 9300.545 335.05 ;
      RECT 9299.705 189.04 9299.985 334.81 ;
      RECT 9299.145 187.94 9299.425 334.57 ;
      RECT 9298.585 189.04 9298.865 334.33 ;
      RECT 9298.025 187.94 9298.305 334.09 ;
      RECT 9297.465 189.04 9297.745 333.85 ;
      RECT 9296.905 189.04 9297.185 333.61 ;
      RECT 9296.345 189.04 9296.625 333.37 ;
      RECT 9295.785 189.04 9296.065 333.13 ;
      RECT 9295.225 189.04 9295.505 332.89 ;
      RECT 9294.665 189.04 9294.945 332.65 ;
      RECT 9294.105 189.04 9294.385 332.41 ;
      RECT 9293.545 189.04 9293.825 332.17 ;
      RECT 9291.025 187.94 9291.305 333.89 ;
      RECT 9290.465 189.04 9290.745 333.65 ;
      RECT 9289.905 187.94 9290.185 333.41 ;
      RECT 9289.345 189.04 9289.625 333.17 ;
      RECT 9288.785 189.04 9289.065 332.93 ;
      RECT 9288.225 189.04 9288.505 332.69 ;
      RECT 9287.665 189.04 9287.945 332.45 ;
      RECT 9287.105 189.04 9287.385 332.21 ;
      RECT 9261.065 189.04 9261.345 329.86 ;
      RECT 9260.505 189.04 9260.785 330.1 ;
      RECT 9259.945 189.04 9260.225 330.34 ;
      RECT 9259.385 189.04 9259.665 330.585 ;
      RECT 9258.825 189.04 9259.105 330.825 ;
      RECT 9258.265 189.04 9258.545 331.065 ;
      RECT 9257.705 189.04 9257.985 331.065 ;
      RECT 9257.145 189.04 9257.425 330.825 ;
      RECT 9256.585 189.04 9256.865 330.585 ;
      RECT 9256.025 187.94 9256.305 330.345 ;
      RECT 9255.465 189.04 9255.745 330.105 ;
      RECT 9254.905 187.94 9255.185 329.865 ;
      RECT 9254.345 189.04 9254.625 329.625 ;
      RECT 9253.785 189.04 9254.065 329.385 ;
      RECT 9253.225 189.04 9253.505 329.145 ;
      RECT 9252.665 187.94 9252.945 328.905 ;
      RECT 9252.105 189.04 9252.385 328.665 ;
      RECT 9251.545 187.94 9251.825 328.425 ;
      RECT 9250.985 189.04 9251.265 328.185 ;
      RECT 9250.425 187.94 9250.705 327.945 ;
      RECT 9249.865 189.04 9250.145 327.705 ;
      RECT 9249.305 189.04 9249.585 327.465 ;
      RECT 9248.745 189.04 9249.025 327.225 ;
      RECT 9248.185 189.04 9248.465 326.985 ;
      RECT 9234.745 189.04 9235.025 332.785 ;
      RECT 9234.185 189.04 9234.465 332.545 ;
      RECT 9233.625 189.04 9233.905 332.305 ;
      RECT 9233.065 189.04 9233.345 332.065 ;
      RECT 9232.505 189.04 9232.785 331.825 ;
      RECT 9231.945 189.04 9232.225 331.585 ;
      RECT 9231.385 189.04 9231.665 331.345 ;
      RECT 9230.825 189.04 9231.105 331.105 ;
      RECT 9230.265 187.94 9230.545 330.865 ;
      RECT 9229.705 189.04 9229.985 330.625 ;
      RECT 9229.145 187.94 9229.425 330.305 ;
      RECT 9228.585 189.04 9228.865 330.145 ;
      RECT 9228.025 187.94 9228.305 329.905 ;
      RECT 9227.465 189.04 9227.745 329.665 ;
      RECT 9226.905 189.04 9227.185 329.425 ;
      RECT 9226.345 189.04 9226.625 329.185 ;
      RECT 9225.785 189.04 9226.065 328.945 ;
      RECT 9225.225 189.04 9225.505 328.705 ;
      RECT 9224.665 189.04 9224.945 328.465 ;
      RECT 9224.105 189.04 9224.385 328.225 ;
      RECT 9223.545 189.04 9223.825 327.985 ;
      RECT 9222.985 187.94 9223.265 327.745 ;
      RECT 9222.425 189.04 9222.705 327.505 ;
      RECT 9221.865 187.94 9222.145 327.265 ;
      RECT 9182.665 189.04 9182.945 332.875 ;
      RECT 9182.105 189.04 9182.385 333.115 ;
      RECT 9181.545 189.04 9181.825 333.355 ;
      RECT 9180.985 189.04 9181.265 333.595 ;
      RECT 9180.425 189.04 9180.705 333.835 ;
      RECT 9179.865 189.04 9180.145 334.075 ;
      RECT 9179.305 189.04 9179.585 334.315 ;
      RECT 9178.745 189.04 9179.025 334.555 ;
      RECT 9178.185 189.04 9178.465 334.795 ;
      RECT 9177.625 189.04 9177.905 335.035 ;
      RECT 9177.065 189.04 9177.345 335.275 ;
      RECT 9176.505 189.04 9176.785 335.515 ;
      RECT 9175.945 189.04 9176.225 335.755 ;
      RECT 9175.385 189.04 9175.665 335.755 ;
      RECT 9174.825 187.94 9175.105 335.515 ;
      RECT 9174.265 189.04 9174.545 335.275 ;
      RECT 9173.705 187.94 9173.985 335.035 ;
      RECT 9173.145 189.04 9173.425 334.795 ;
      RECT 9172.585 189.04 9172.865 334.555 ;
      RECT 9172.025 189.04 9172.305 334.315 ;
      RECT 9171.465 187.94 9171.745 334.05 ;
      RECT 9170.905 189.04 9171.185 333.81 ;
      RECT 9170.345 187.94 9170.625 333.57 ;
      RECT 9169.785 189.04 9170.065 333.33 ;
      RECT 9160.825 187.94 9161.105 327.165 ;
      RECT 9160.265 189.04 9160.545 327.405 ;
      RECT 9159.705 189.04 9159.985 327.645 ;
      RECT 9159.145 189.04 9159.425 327.645 ;
      RECT 9158.585 189.04 9158.865 327.405 ;
      RECT 9158.025 189.04 9158.305 327.165 ;
      RECT 9157.465 189.04 9157.745 326.925 ;
      RECT 9156.905 189.04 9157.185 326.685 ;
      RECT 9156.345 189.04 9156.625 326.445 ;
      RECT 9155.785 189.04 9156.065 326.205 ;
      RECT 9155.225 189.04 9155.505 325.965 ;
      RECT 9154.665 189.04 9154.945 325.725 ;
      RECT 9154.105 189.04 9154.385 325.485 ;
      RECT 9153.545 187.94 9153.825 325.245 ;
      RECT 9151.025 189.04 9151.305 326.965 ;
      RECT 9150.465 187.94 9150.745 326.725 ;
      RECT 9149.905 189.04 9150.185 326.485 ;
      RECT 9149.345 187.94 9149.625 326.245 ;
      RECT 9148.785 189.04 9149.065 326.005 ;
      RECT 9148.225 189.04 9148.505 325.765 ;
      RECT 9147.665 189.04 9147.945 325.525 ;
      RECT 9121.625 189.04 9121.905 328.31 ;
      RECT 9121.065 189.04 9121.345 328.55 ;
      RECT 9120.505 189.04 9120.785 328.79 ;
      RECT 9119.945 189.04 9120.225 329.03 ;
      RECT 9119.385 189.04 9119.665 329.27 ;
      RECT 9118.825 187.94 9119.105 329.51 ;
      RECT 9118.265 189.04 9118.545 329.75 ;
      RECT 9117.705 187.94 9117.985 329.99 ;
      RECT 9117.145 189.04 9117.425 330.23 ;
      RECT 9116.585 189.04 9116.865 330.47 ;
      RECT 9116.025 189.04 9116.305 330.71 ;
      RECT 9115.465 189.04 9115.745 330.95 ;
      RECT 9114.905 189.04 9115.185 331.19 ;
      RECT 9114.345 189.04 9114.625 331.43 ;
      RECT 9113.785 189.04 9114.065 331.67 ;
      RECT 9113.225 189.04 9113.505 331.67 ;
      RECT 9112.665 189.04 9112.945 331.43 ;
      RECT 9112.105 189.04 9112.385 331.19 ;
      RECT 9111.545 189.04 9111.825 330.95 ;
      RECT 9110.985 189.04 9111.265 330.705 ;
      RECT 9110.425 189.04 9110.705 330.465 ;
      RECT 9109.865 189.04 9110.145 330.225 ;
      RECT 9109.305 187.94 9109.585 329.985 ;
      RECT 9108.745 189.04 9109.025 329.745 ;
      RECT 9095.305 187.94 9095.585 327.225 ;
      RECT 9094.745 189.04 9095.025 326.985 ;
      RECT 9094.185 189.04 9094.465 326.745 ;
      RECT 9093.625 189.04 9093.905 326.505 ;
      RECT 9093.065 187.94 9093.345 326.265 ;
      RECT 9092.505 189.04 9092.785 326.025 ;
      RECT 9091.945 187.94 9092.225 325.785 ;
      RECT 9091.385 189.04 9091.665 325.545 ;
      RECT 9090.825 187.94 9091.105 325.305 ;
      RECT 9090.265 189.04 9090.545 325.065 ;
      RECT 9089.705 189.04 9089.985 324.825 ;
      RECT 9089.145 189.04 9089.425 324.585 ;
      RECT 9088.585 189.04 9088.865 324.345 ;
      RECT 9088.025 189.04 9088.305 324.105 ;
      RECT 9087.465 189.04 9087.745 323.865 ;
      RECT 9086.905 189.04 9087.185 323.625 ;
      RECT 9086.345 189.04 9086.625 323.385 ;
      RECT 9085.785 189.04 9086.065 323.145 ;
      RECT 9085.225 189.04 9085.505 322.905 ;
      RECT 9084.665 189.04 9084.945 322.665 ;
      RECT 9084.105 189.04 9084.385 322.425 ;
      RECT 9083.545 187.94 9083.825 322.185 ;
      RECT 9082.985 189.04 9083.265 321.945 ;
      RECT 9082.425 187.94 9082.705 321.705 ;
      RECT 9042.665 189.04 9042.945 332.175 ;
      RECT 9042.105 187.94 9042.385 332.415 ;
      RECT 9041.545 189.04 9041.825 332.655 ;
      RECT 9040.985 189.04 9041.265 332.895 ;
      RECT 9040.425 189.04 9040.705 333.135 ;
      RECT 9039.865 189.04 9040.145 333.375 ;
      RECT 9039.305 189.04 9039.585 333.615 ;
      RECT 9038.745 189.04 9039.025 333.86 ;
      RECT 9038.185 189.04 9038.465 334.1 ;
      RECT 9037.625 189.04 9037.905 334.34 ;
      RECT 9037.065 187.94 9037.345 334.58 ;
      RECT 9036.505 189.04 9036.785 334.82 ;
      RECT 9035.945 187.94 9036.225 335.06 ;
      RECT 9035.385 189.04 9035.665 335.3 ;
      RECT 9034.825 189.04 9035.105 335.54 ;
      RECT 9034.265 189.04 9034.545 335.78 ;
      RECT 9033.705 189.04 9033.985 336.02 ;
      RECT 9033.145 189.04 9033.425 336.26 ;
      RECT 9032.585 189.04 9032.865 336.5 ;
      RECT 9032.025 189.04 9032.305 336.74 ;
      RECT 9031.465 189.04 9031.745 336.98 ;
      RECT 9030.905 189.04 9031.185 337.22 ;
      RECT 9030.345 189.04 9030.625 337.46 ;
      RECT 9029.785 189.04 9030.065 337.7 ;
      RECT 9020.825 189.04 9021.105 333.285 ;
      RECT 9020.265 189.04 9020.545 333.045 ;
      RECT 9019.705 189.04 9019.985 332.805 ;
      RECT 9019.145 187.94 9019.425 332.565 ;
      RECT 9018.585 189.04 9018.865 332.325 ;
      RECT 9018.025 187.94 9018.305 332.085 ;
      RECT 9017.465 189.04 9017.745 331.845 ;
      RECT 9016.905 189.04 9017.185 331.605 ;
      RECT 9016.345 189.04 9016.625 331.365 ;
      RECT 9015.785 187.94 9016.065 331.125 ;
      RECT 9015.225 189.04 9015.505 330.885 ;
      RECT 9014.665 187.94 9014.945 330.645 ;
      RECT 9014.105 189.04 9014.385 330.405 ;
      RECT 9013.545 187.94 9013.825 330.165 ;
      RECT 9011.025 189.04 9011.305 322.565 ;
      RECT 9010.465 189.04 9010.745 322.325 ;
      RECT 9009.905 189.04 9010.185 322.085 ;
      RECT 9009.345 189.04 9009.625 321.845 ;
      RECT 9008.785 189.04 9009.065 321.605 ;
      RECT 9008.225 189.04 9008.505 321.365 ;
      RECT 9007.665 189.04 9007.945 321.125 ;
      RECT 8981.625 189.04 8981.905 335 ;
      RECT 8981.065 189.04 8981.345 335.24 ;
      RECT 8980.505 189.04 8980.785 335.48 ;
      RECT 8979.945 189.04 8980.225 335.72 ;
      RECT 8979.385 189.04 8979.665 335.96 ;
      RECT 8978.825 187.94 8979.105 335.96 ;
      RECT 8978.265 189.04 8978.545 335.72 ;
      RECT 8977.705 187.94 8977.985 335.475 ;
      RECT 8977.145 189.04 8977.425 335.235 ;
      RECT 8976.585 187.94 8976.865 334.995 ;
      RECT 8976.025 189.04 8976.305 334.755 ;
      RECT 8975.465 189.04 8975.745 334.515 ;
      RECT 8974.905 189.04 8975.185 334.275 ;
      RECT 8974.345 189.04 8974.625 334.035 ;
      RECT 8973.785 189.04 8974.065 333.795 ;
      RECT 8973.225 189.04 8973.505 333.555 ;
      RECT 8972.665 189.04 8972.945 333.315 ;
      RECT 8972.105 189.04 8972.385 333.075 ;
      RECT 8971.545 187.94 8971.825 332.835 ;
      RECT 8970.985 189.04 8971.265 332.595 ;
      RECT 8970.425 187.94 8970.705 332.355 ;
      RECT 8969.865 189.04 8970.145 332.115 ;
      RECT 8969.305 189.04 8969.585 331.875 ;
      RECT 8968.745 189.04 8969.025 331.635 ;
      RECT 8955.305 189.04 8955.585 335.035 ;
      RECT 8954.745 189.04 8955.025 335.275 ;
      RECT 8954.185 189.04 8954.465 335.52 ;
      RECT 8953.625 189.04 8953.905 335.76 ;
      RECT 8953.065 189.04 8953.345 336 ;
      RECT 8952.505 189.04 8952.785 336 ;
      RECT 8951.945 189.04 8952.225 335.76 ;
      RECT 8951.385 189.04 8951.665 335.52 ;
      RECT 8950.825 189.04 8951.105 328.505 ;
      RECT 8950.265 189.04 8950.545 328.265 ;
      RECT 8949.705 189.04 8949.985 328.025 ;
      RECT 8949.145 187.94 8949.425 327.785 ;
      RECT 8948.585 189.04 8948.865 327.545 ;
      RECT 8948.025 187.94 8948.305 327.305 ;
      RECT 8947.465 189.04 8947.745 327.065 ;
      RECT 8946.905 189.04 8947.185 326.825 ;
      RECT 8946.345 189.04 8946.625 326.585 ;
      RECT 8945.785 187.94 8946.065 326.345 ;
      RECT 8945.225 189.04 8945.505 326.105 ;
      RECT 8944.665 187.94 8944.945 325.865 ;
      RECT 8944.105 189.04 8944.385 325.625 ;
      RECT 8943.545 187.94 8943.825 325.385 ;
      RECT 8942.985 189.04 8943.265 325.145 ;
      RECT 8942.425 189.04 8942.705 324.905 ;
      RECT 8902.105 189.04 8902.385 333.8 ;
      RECT 8901.545 189.04 8901.825 334.04 ;
      RECT 8900.985 189.04 8901.265 334.285 ;
      RECT 8900.425 189.04 8900.705 334.525 ;
      RECT 8899.865 189.04 8900.145 334.765 ;
      RECT 8899.305 189.04 8899.585 335.005 ;
      RECT 8898.745 189.04 8899.025 335.245 ;
      RECT 8898.185 189.04 8898.465 335.485 ;
      RECT 8897.625 189.04 8897.905 335.725 ;
      RECT 8897.065 189.04 8897.345 335.965 ;
      RECT 8896.505 187.94 8896.785 336.205 ;
      RECT 8895.945 189.04 8896.225 336.445 ;
      RECT 8895.385 187.94 8895.665 336.685 ;
      RECT 8894.825 189.04 8895.105 336.925 ;
      RECT 8894.265 187.94 8894.545 337.165 ;
      RECT 8893.705 189.04 8893.985 337.165 ;
      RECT 8893.145 189.04 8893.425 336.925 ;
      RECT 8892.585 189.04 8892.865 336.685 ;
      RECT 8892.025 189.04 8892.305 336.445 ;
      RECT 8891.465 189.04 8891.745 336.205 ;
      RECT 8890.905 189.04 8891.185 335.965 ;
      RECT 8890.345 189.04 8890.625 335.725 ;
      RECT 8889.785 189.04 8890.065 335.485 ;
      RECT 8880.825 187.94 8881.105 335.515 ;
      RECT 8880.265 189.04 8880.545 335.755 ;
      RECT 8879.705 187.94 8879.985 335.995 ;
      RECT 8879.145 189.04 8879.425 336.21 ;
      RECT 8878.585 189.04 8878.865 335.785 ;
      RECT 8878.025 189.04 8878.305 335.545 ;
      RECT 8877.465 189.04 8877.745 335.305 ;
      RECT 8876.905 189.04 8877.185 335.065 ;
      RECT 8876.345 189.04 8876.625 334.825 ;
      RECT 8875.785 189.04 8876.065 334.585 ;
      RECT 8875.225 189.04 8875.505 334.345 ;
      RECT 8874.665 189.04 8874.945 334.105 ;
      RECT 8874.105 189.04 8874.385 333.865 ;
      RECT 8873.545 189.04 8873.825 333.625 ;
      RECT 8871.025 189.04 8871.305 332.8 ;
      RECT 8870.465 189.04 8870.745 332.56 ;
      RECT 8869.905 189.04 8870.185 332.32 ;
      RECT 8869.345 187.94 8869.625 332.08 ;
      RECT 8868.785 189.04 8869.065 331.84 ;
      RECT 8868.225 187.94 8868.505 331.6 ;
      RECT 8867.665 189.04 8867.945 331.36 ;
      RECT 8867.105 189.04 8867.385 331.12 ;
      RECT 8840.505 189.04 8840.785 342.165 ;
      RECT 8839.945 187.94 8840.225 342.405 ;
      RECT 8839.385 189.04 8839.665 342.645 ;
      RECT 8838.825 187.94 8839.105 342.89 ;
      RECT 8838.265 189.04 8838.545 343.13 ;
      RECT 8837.705 187.94 8837.985 343.37 ;
      RECT 8837.145 189.04 8837.425 343.61 ;
      RECT 8836.585 189.04 8836.865 343.85 ;
      RECT 8836.025 189.04 8836.305 329.47 ;
      RECT 8835.465 189.04 8835.745 329.23 ;
      RECT 8834.905 189.04 8835.185 328.99 ;
      RECT 8834.345 189.04 8834.625 328.75 ;
      RECT 8833.785 189.04 8834.065 328.51 ;
      RECT 8833.225 189.04 8833.505 328.27 ;
      RECT 8832.665 189.04 8832.945 328.03 ;
      RECT 8832.105 189.04 8832.385 327.79 ;
      RECT 8831.545 189.04 8831.825 327.55 ;
      RECT 8830.985 189.04 8831.265 327.31 ;
      RECT 8830.425 187.94 8830.705 327.07 ;
      RECT 8829.865 189.04 8830.145 326.83 ;
      RECT 8829.305 187.94 8829.585 326.59 ;
      RECT 8828.745 189.04 8829.025 326.35 ;
      RECT 8814.745 187.94 8815.025 332.47 ;
      RECT 8814.185 189.04 8814.465 332.23 ;
      RECT 8813.625 189.04 8813.905 331.99 ;
      RECT 8813.065 189.04 8813.345 331.75 ;
      RECT 8812.505 189.04 8812.785 331.51 ;
      RECT 8811.945 189.04 8812.225 331.27 ;
      RECT 8811.385 189.04 8811.665 331.03 ;
      RECT 8810.825 189.04 8811.105 330.79 ;
      RECT 8810.265 189.04 8810.545 330.55 ;
      RECT 8809.705 187.94 8809.985 330.31 ;
      RECT 8809.145 189.04 8809.425 330.07 ;
      RECT 8808.585 187.94 8808.865 329.83 ;
      RECT 8808.025 189.04 8808.305 329.59 ;
      RECT 8807.465 189.04 8807.745 329.35 ;
      RECT 8806.905 189.04 8807.185 329.11 ;
      RECT 8806.345 189.04 8806.625 328.87 ;
      RECT 8805.785 189.04 8806.065 328.63 ;
      RECT 8805.225 189.04 8805.505 328.39 ;
      RECT 8804.665 189.04 8804.945 328.15 ;
      RECT 8804.105 189.04 8804.385 327.91 ;
      RECT 8803.545 189.04 8803.825 327.67 ;
      RECT 8802.985 189.04 8803.265 327.43 ;
      RECT 8802.425 189.04 8802.705 327.19 ;
      RECT 8763.225 189.04 8763.505 334.095 ;
      RECT 8762.665 189.04 8762.945 334.335 ;
      RECT 8762.105 189.04 8762.385 334.575 ;
      RECT 8761.545 187.94 8761.825 334.815 ;
      RECT 8760.985 189.04 8761.265 335.055 ;
      RECT 8760.425 187.94 8760.705 335.295 ;
      RECT 8759.865 189.04 8760.145 335.535 ;
      RECT 8759.305 189.04 8759.585 335.775 ;
      RECT 8758.745 189.04 8759.025 336.015 ;
      RECT 8758.185 187.94 8758.465 336.255 ;
      RECT 8757.625 189.04 8757.905 336.495 ;
      RECT 8757.065 187.94 8757.345 336.735 ;
      RECT 8756.505 189.04 8756.785 336.975 ;
      RECT 8755.945 187.94 8756.225 337.215 ;
      RECT 8755.385 189.04 8755.665 337.455 ;
      RECT 8754.825 189.04 8755.105 337.695 ;
      RECT 8754.265 189.04 8754.545 337.695 ;
      RECT 8753.705 189.04 8753.985 337.455 ;
      RECT 8753.145 189.04 8753.425 337.215 ;
      RECT 8752.585 189.04 8752.865 336.975 ;
      RECT 8752.025 189.04 8752.305 336.735 ;
      RECT 8751.465 189.04 8751.745 336.495 ;
      RECT 8750.905 189.04 8751.185 336.255 ;
      RECT 8750.345 189.04 8750.625 336.015 ;
      RECT 8749.785 189.04 8750.065 335.775 ;
      RECT 8740.825 189.04 8741.105 335.29 ;
      RECT 8740.265 187.94 8740.545 335.05 ;
      RECT 8739.705 189.04 8739.985 334.81 ;
      RECT 8739.145 187.94 8739.425 334.57 ;
      RECT 8738.585 189.04 8738.865 334.33 ;
      RECT 8738.025 187.94 8738.305 334.09 ;
      RECT 8737.465 189.04 8737.745 333.85 ;
      RECT 8736.905 189.04 8737.185 333.61 ;
      RECT 8736.345 189.04 8736.625 333.37 ;
      RECT 8735.785 189.04 8736.065 333.13 ;
      RECT 8735.225 189.04 8735.505 332.89 ;
      RECT 8734.665 189.04 8734.945 332.65 ;
      RECT 8734.105 189.04 8734.385 332.41 ;
      RECT 8733.545 189.04 8733.825 332.17 ;
      RECT 8731.025 187.94 8731.305 333.89 ;
      RECT 8730.465 189.04 8730.745 333.65 ;
      RECT 8729.905 187.94 8730.185 333.41 ;
      RECT 8729.345 189.04 8729.625 333.17 ;
      RECT 8728.785 189.04 8729.065 332.93 ;
      RECT 8728.225 189.04 8728.505 332.69 ;
      RECT 8727.665 189.04 8727.945 332.45 ;
      RECT 8727.105 189.04 8727.385 332.21 ;
      RECT 8701.065 189.04 8701.345 329.86 ;
      RECT 8700.505 189.04 8700.785 330.1 ;
      RECT 8699.945 189.04 8700.225 330.34 ;
      RECT 8699.385 189.04 8699.665 330.585 ;
      RECT 8698.825 189.04 8699.105 330.825 ;
      RECT 8698.265 189.04 8698.545 331.065 ;
      RECT 8697.705 189.04 8697.985 331.065 ;
      RECT 8697.145 189.04 8697.425 330.825 ;
      RECT 8696.585 189.04 8696.865 330.585 ;
      RECT 8696.025 187.94 8696.305 330.345 ;
      RECT 8695.465 189.04 8695.745 330.105 ;
      RECT 8694.905 187.94 8695.185 329.865 ;
      RECT 8694.345 189.04 8694.625 329.625 ;
      RECT 8693.785 189.04 8694.065 329.385 ;
      RECT 8693.225 189.04 8693.505 329.145 ;
      RECT 8692.665 187.94 8692.945 328.905 ;
      RECT 8692.105 189.04 8692.385 328.665 ;
      RECT 8691.545 187.94 8691.825 328.425 ;
      RECT 8690.985 189.04 8691.265 328.185 ;
      RECT 8690.425 187.94 8690.705 327.945 ;
      RECT 8689.865 189.04 8690.145 327.705 ;
      RECT 8689.305 189.04 8689.585 327.465 ;
      RECT 8688.745 189.04 8689.025 327.225 ;
      RECT 8688.185 189.04 8688.465 326.985 ;
      RECT 8674.745 189.04 8675.025 332.785 ;
      RECT 8674.185 189.04 8674.465 332.545 ;
      RECT 8673.625 189.04 8673.905 332.305 ;
      RECT 8673.065 189.04 8673.345 332.065 ;
      RECT 8672.505 189.04 8672.785 331.825 ;
      RECT 8671.945 189.04 8672.225 331.585 ;
      RECT 8671.385 189.04 8671.665 331.345 ;
      RECT 8670.825 189.04 8671.105 331.105 ;
      RECT 8670.265 187.94 8670.545 330.865 ;
      RECT 8669.705 189.04 8669.985 330.625 ;
      RECT 8669.145 187.94 8669.425 330.305 ;
      RECT 8668.585 189.04 8668.865 330.145 ;
      RECT 8668.025 187.94 8668.305 329.905 ;
      RECT 8667.465 189.04 8667.745 329.665 ;
      RECT 8666.905 189.04 8667.185 329.425 ;
      RECT 8666.345 189.04 8666.625 329.185 ;
      RECT 8665.785 189.04 8666.065 328.945 ;
      RECT 8665.225 189.04 8665.505 328.705 ;
      RECT 8664.665 189.04 8664.945 328.465 ;
      RECT 8664.105 189.04 8664.385 328.225 ;
      RECT 8663.545 189.04 8663.825 327.985 ;
      RECT 8662.985 187.94 8663.265 327.745 ;
      RECT 8662.425 189.04 8662.705 327.505 ;
      RECT 8661.865 187.94 8662.145 327.265 ;
      RECT 8622.665 189.04 8622.945 332.875 ;
      RECT 8622.105 189.04 8622.385 333.115 ;
      RECT 8621.545 189.04 8621.825 333.355 ;
      RECT 8620.985 189.04 8621.265 333.595 ;
      RECT 8620.425 189.04 8620.705 333.835 ;
      RECT 8619.865 189.04 8620.145 334.075 ;
      RECT 8619.305 189.04 8619.585 334.315 ;
      RECT 8618.745 189.04 8619.025 334.555 ;
      RECT 8618.185 189.04 8618.465 334.795 ;
      RECT 8617.625 189.04 8617.905 335.035 ;
      RECT 8617.065 189.04 8617.345 335.275 ;
      RECT 8616.505 189.04 8616.785 335.515 ;
      RECT 8615.945 189.04 8616.225 335.755 ;
      RECT 8615.385 189.04 8615.665 335.755 ;
      RECT 8614.825 187.94 8615.105 335.515 ;
      RECT 8614.265 189.04 8614.545 335.275 ;
      RECT 8613.705 187.94 8613.985 335.035 ;
      RECT 8613.145 189.04 8613.425 334.795 ;
      RECT 8612.585 189.04 8612.865 334.555 ;
      RECT 8612.025 189.04 8612.305 334.315 ;
      RECT 8611.465 187.94 8611.745 334.05 ;
      RECT 8610.905 189.04 8611.185 333.81 ;
      RECT 8610.345 187.94 8610.625 333.57 ;
      RECT 8609.785 189.04 8610.065 333.33 ;
      RECT 8600.825 187.94 8601.105 327.165 ;
      RECT 8600.265 189.04 8600.545 327.405 ;
      RECT 8599.705 189.04 8599.985 327.645 ;
      RECT 8599.145 189.04 8599.425 327.645 ;
      RECT 8598.585 189.04 8598.865 327.405 ;
      RECT 8598.025 189.04 8598.305 327.165 ;
      RECT 8597.465 189.04 8597.745 326.925 ;
      RECT 8596.905 189.04 8597.185 326.685 ;
      RECT 8596.345 189.04 8596.625 326.445 ;
      RECT 8595.785 189.04 8596.065 326.205 ;
      RECT 8595.225 189.04 8595.505 325.965 ;
      RECT 8594.665 189.04 8594.945 325.725 ;
      RECT 8594.105 189.04 8594.385 325.485 ;
      RECT 8593.545 187.94 8593.825 325.245 ;
      RECT 8591.025 189.04 8591.305 326.965 ;
      RECT 8590.465 187.94 8590.745 326.725 ;
      RECT 8589.905 189.04 8590.185 326.485 ;
      RECT 8589.345 187.94 8589.625 326.245 ;
      RECT 8588.785 189.04 8589.065 326.005 ;
      RECT 8588.225 189.04 8588.505 325.765 ;
      RECT 8587.665 189.04 8587.945 325.525 ;
      RECT 8561.625 189.04 8561.905 328.31 ;
      RECT 8561.065 189.04 8561.345 328.55 ;
      RECT 8560.505 189.04 8560.785 328.79 ;
      RECT 8559.945 189.04 8560.225 329.03 ;
      RECT 8559.385 189.04 8559.665 329.27 ;
      RECT 8558.825 187.94 8559.105 329.51 ;
      RECT 8558.265 189.04 8558.545 329.75 ;
      RECT 8557.705 187.94 8557.985 329.99 ;
      RECT 8557.145 189.04 8557.425 330.23 ;
      RECT 8556.585 189.04 8556.865 330.47 ;
      RECT 8556.025 189.04 8556.305 330.71 ;
      RECT 8555.465 189.04 8555.745 330.95 ;
      RECT 8554.905 189.04 8555.185 331.19 ;
      RECT 8554.345 189.04 8554.625 331.43 ;
      RECT 8553.785 189.04 8554.065 331.67 ;
      RECT 8553.225 189.04 8553.505 331.67 ;
      RECT 8552.665 189.04 8552.945 331.43 ;
      RECT 8552.105 189.04 8552.385 331.19 ;
      RECT 8551.545 189.04 8551.825 330.95 ;
      RECT 8550.985 189.04 8551.265 330.705 ;
      RECT 8550.425 189.04 8550.705 330.465 ;
      RECT 8549.865 189.04 8550.145 330.225 ;
      RECT 8549.305 187.94 8549.585 329.985 ;
      RECT 8548.745 189.04 8549.025 329.745 ;
      RECT 8535.305 187.94 8535.585 327.225 ;
      RECT 8534.745 189.04 8535.025 326.985 ;
      RECT 8534.185 189.04 8534.465 326.745 ;
      RECT 8533.625 189.04 8533.905 326.505 ;
      RECT 8533.065 187.94 8533.345 326.265 ;
      RECT 8532.505 189.04 8532.785 326.025 ;
      RECT 8531.945 187.94 8532.225 325.785 ;
      RECT 8531.385 189.04 8531.665 325.545 ;
      RECT 8530.825 187.94 8531.105 325.305 ;
      RECT 8530.265 189.04 8530.545 325.065 ;
      RECT 8529.705 189.04 8529.985 324.825 ;
      RECT 8529.145 189.04 8529.425 324.585 ;
      RECT 8528.585 189.04 8528.865 324.345 ;
      RECT 8528.025 189.04 8528.305 324.105 ;
      RECT 8527.465 189.04 8527.745 323.865 ;
      RECT 8526.905 189.04 8527.185 323.625 ;
      RECT 8526.345 189.04 8526.625 323.385 ;
      RECT 8525.785 189.04 8526.065 323.145 ;
      RECT 8525.225 189.04 8525.505 322.905 ;
      RECT 8524.665 189.04 8524.945 322.665 ;
      RECT 8524.105 189.04 8524.385 322.425 ;
      RECT 8523.545 187.94 8523.825 322.185 ;
      RECT 8522.985 189.04 8523.265 321.945 ;
      RECT 8522.425 187.94 8522.705 321.705 ;
      RECT 8482.665 189.04 8482.945 332.175 ;
      RECT 8482.105 187.94 8482.385 332.415 ;
      RECT 8481.545 189.04 8481.825 332.655 ;
      RECT 8480.985 189.04 8481.265 332.895 ;
      RECT 8480.425 189.04 8480.705 333.135 ;
      RECT 8479.865 189.04 8480.145 333.375 ;
      RECT 8479.305 189.04 8479.585 333.615 ;
      RECT 8478.745 189.04 8479.025 333.86 ;
      RECT 8478.185 189.04 8478.465 334.1 ;
      RECT 8477.625 189.04 8477.905 334.34 ;
      RECT 8477.065 187.94 8477.345 334.58 ;
      RECT 8476.505 189.04 8476.785 334.82 ;
      RECT 8475.945 187.94 8476.225 335.06 ;
      RECT 8475.385 189.04 8475.665 335.3 ;
      RECT 8474.825 189.04 8475.105 335.54 ;
      RECT 8474.265 189.04 8474.545 335.78 ;
      RECT 8473.705 189.04 8473.985 336.02 ;
      RECT 8473.145 189.04 8473.425 336.26 ;
      RECT 8472.585 189.04 8472.865 336.5 ;
      RECT 8472.025 189.04 8472.305 336.74 ;
      RECT 8471.465 189.04 8471.745 336.98 ;
      RECT 8470.905 189.04 8471.185 337.22 ;
      RECT 8470.345 189.04 8470.625 337.46 ;
      RECT 8469.785 189.04 8470.065 337.7 ;
      RECT 8460.825 189.04 8461.105 333.285 ;
      RECT 8460.265 189.04 8460.545 333.045 ;
      RECT 8459.705 189.04 8459.985 332.805 ;
      RECT 8459.145 187.94 8459.425 332.565 ;
      RECT 8458.585 189.04 8458.865 332.325 ;
      RECT 8458.025 187.94 8458.305 332.085 ;
      RECT 8457.465 189.04 8457.745 331.845 ;
      RECT 8456.905 189.04 8457.185 331.605 ;
      RECT 8456.345 189.04 8456.625 331.365 ;
      RECT 8455.785 187.94 8456.065 331.125 ;
      RECT 8455.225 189.04 8455.505 330.885 ;
      RECT 8454.665 187.94 8454.945 330.645 ;
      RECT 8454.105 189.04 8454.385 330.405 ;
      RECT 8453.545 187.94 8453.825 330.165 ;
      RECT 8451.025 189.04 8451.305 322.565 ;
      RECT 8450.465 189.04 8450.745 322.325 ;
      RECT 8449.905 189.04 8450.185 322.085 ;
      RECT 8449.345 189.04 8449.625 321.845 ;
      RECT 8448.785 189.04 8449.065 321.605 ;
      RECT 8448.225 189.04 8448.505 321.365 ;
      RECT 8447.665 189.04 8447.945 321.125 ;
      RECT 8421.625 189.04 8421.905 335 ;
      RECT 8421.065 189.04 8421.345 335.24 ;
      RECT 8420.505 189.04 8420.785 335.48 ;
      RECT 8419.945 189.04 8420.225 335.72 ;
      RECT 8419.385 189.04 8419.665 335.96 ;
      RECT 8418.825 187.94 8419.105 335.96 ;
      RECT 8418.265 189.04 8418.545 335.72 ;
      RECT 8417.705 187.94 8417.985 335.475 ;
      RECT 8417.145 189.04 8417.425 335.235 ;
      RECT 8416.585 187.94 8416.865 334.995 ;
      RECT 8416.025 189.04 8416.305 334.755 ;
      RECT 8415.465 189.04 8415.745 334.515 ;
      RECT 8414.905 189.04 8415.185 334.275 ;
      RECT 8414.345 189.04 8414.625 334.035 ;
      RECT 8413.785 189.04 8414.065 333.795 ;
      RECT 8413.225 189.04 8413.505 333.555 ;
      RECT 8412.665 189.04 8412.945 333.315 ;
      RECT 8412.105 189.04 8412.385 333.075 ;
      RECT 8411.545 187.94 8411.825 332.835 ;
      RECT 8410.985 189.04 8411.265 332.595 ;
      RECT 8410.425 187.94 8410.705 332.355 ;
      RECT 8409.865 189.04 8410.145 332.115 ;
      RECT 8409.305 189.04 8409.585 331.875 ;
      RECT 8408.745 189.04 8409.025 331.635 ;
      RECT 8395.305 189.04 8395.585 335.035 ;
      RECT 8394.745 189.04 8395.025 335.275 ;
      RECT 8394.185 189.04 8394.465 335.52 ;
      RECT 8393.625 189.04 8393.905 335.76 ;
      RECT 8393.065 189.04 8393.345 336 ;
      RECT 8392.505 189.04 8392.785 336 ;
      RECT 8391.945 189.04 8392.225 335.76 ;
      RECT 8391.385 189.04 8391.665 335.52 ;
      RECT 8390.825 189.04 8391.105 328.505 ;
      RECT 8390.265 189.04 8390.545 328.265 ;
      RECT 8389.705 189.04 8389.985 328.025 ;
      RECT 8389.145 187.94 8389.425 327.785 ;
      RECT 8388.585 189.04 8388.865 327.545 ;
      RECT 8388.025 187.94 8388.305 327.305 ;
      RECT 8387.465 189.04 8387.745 327.065 ;
      RECT 8386.905 189.04 8387.185 326.825 ;
      RECT 8386.345 189.04 8386.625 326.585 ;
      RECT 8385.785 187.94 8386.065 326.345 ;
      RECT 8385.225 189.04 8385.505 326.105 ;
      RECT 8384.665 187.94 8384.945 325.865 ;
      RECT 8384.105 189.04 8384.385 325.625 ;
      RECT 8383.545 187.94 8383.825 325.385 ;
      RECT 8382.985 189.04 8383.265 325.145 ;
      RECT 8382.425 189.04 8382.705 324.905 ;
      RECT 8342.105 189.04 8342.385 333.8 ;
      RECT 8341.545 189.04 8341.825 334.04 ;
      RECT 8340.985 189.04 8341.265 334.285 ;
      RECT 8340.425 189.04 8340.705 334.525 ;
      RECT 8339.865 189.04 8340.145 334.765 ;
      RECT 8339.305 189.04 8339.585 335.005 ;
      RECT 8338.745 189.04 8339.025 335.245 ;
      RECT 8338.185 189.04 8338.465 335.485 ;
      RECT 8337.625 189.04 8337.905 335.725 ;
      RECT 8337.065 189.04 8337.345 335.965 ;
      RECT 8336.505 187.94 8336.785 336.205 ;
      RECT 8335.945 189.04 8336.225 336.445 ;
      RECT 8335.385 187.94 8335.665 336.685 ;
      RECT 8334.825 189.04 8335.105 336.925 ;
      RECT 8334.265 187.94 8334.545 337.165 ;
      RECT 8333.705 189.04 8333.985 337.165 ;
      RECT 8333.145 189.04 8333.425 336.925 ;
      RECT 8332.585 189.04 8332.865 336.685 ;
      RECT 8332.025 189.04 8332.305 336.445 ;
      RECT 8331.465 189.04 8331.745 336.205 ;
      RECT 8330.905 189.04 8331.185 335.965 ;
      RECT 8330.345 189.04 8330.625 335.725 ;
      RECT 8329.785 189.04 8330.065 335.485 ;
      RECT 8320.825 187.94 8321.105 335.515 ;
      RECT 8320.265 189.04 8320.545 335.755 ;
      RECT 8319.705 187.94 8319.985 335.995 ;
      RECT 8319.145 189.04 8319.425 336.21 ;
      RECT 8318.585 189.04 8318.865 335.785 ;
      RECT 8318.025 189.04 8318.305 335.545 ;
      RECT 8317.465 189.04 8317.745 335.305 ;
      RECT 8316.905 189.04 8317.185 335.065 ;
      RECT 8316.345 189.04 8316.625 334.825 ;
      RECT 8315.785 189.04 8316.065 334.585 ;
      RECT 8315.225 189.04 8315.505 334.345 ;
      RECT 8314.665 189.04 8314.945 334.105 ;
      RECT 8314.105 189.04 8314.385 333.865 ;
      RECT 8313.545 189.04 8313.825 333.625 ;
      RECT 8311.025 189.04 8311.305 332.8 ;
      RECT 8310.465 189.04 8310.745 332.56 ;
      RECT 8309.905 189.04 8310.185 332.32 ;
      RECT 8309.345 187.94 8309.625 332.08 ;
      RECT 8308.785 189.04 8309.065 331.84 ;
      RECT 8308.225 187.94 8308.505 331.6 ;
      RECT 8307.665 189.04 8307.945 331.36 ;
      RECT 8307.105 189.04 8307.385 331.12 ;
      RECT 8280.505 189.04 8280.785 342.165 ;
      RECT 8279.945 187.94 8280.225 342.405 ;
      RECT 8279.385 189.04 8279.665 342.645 ;
      RECT 8278.825 187.94 8279.105 342.89 ;
      RECT 8278.265 189.04 8278.545 343.13 ;
      RECT 8277.705 187.94 8277.985 343.37 ;
      RECT 8277.145 189.04 8277.425 343.61 ;
      RECT 8276.585 189.04 8276.865 343.85 ;
      RECT 8276.025 189.04 8276.305 329.47 ;
      RECT 8275.465 189.04 8275.745 329.23 ;
      RECT 8274.905 189.04 8275.185 328.99 ;
      RECT 8274.345 189.04 8274.625 328.75 ;
      RECT 8273.785 189.04 8274.065 328.51 ;
      RECT 8273.225 189.04 8273.505 328.27 ;
      RECT 8272.665 189.04 8272.945 328.03 ;
      RECT 8272.105 189.04 8272.385 327.79 ;
      RECT 8271.545 189.04 8271.825 327.55 ;
      RECT 8270.985 189.04 8271.265 327.31 ;
      RECT 8270.425 187.94 8270.705 327.07 ;
      RECT 8269.865 189.04 8270.145 326.83 ;
      RECT 8269.305 187.94 8269.585 326.59 ;
      RECT 8268.745 189.04 8269.025 326.35 ;
      RECT 8254.745 187.94 8255.025 332.47 ;
      RECT 8254.185 189.04 8254.465 332.23 ;
      RECT 8253.625 189.04 8253.905 331.99 ;
      RECT 8253.065 189.04 8253.345 331.75 ;
      RECT 8252.505 189.04 8252.785 331.51 ;
      RECT 8251.945 189.04 8252.225 331.27 ;
      RECT 8251.385 189.04 8251.665 331.03 ;
      RECT 8250.825 189.04 8251.105 330.79 ;
      RECT 8250.265 189.04 8250.545 330.55 ;
      RECT 8249.705 187.94 8249.985 330.31 ;
      RECT 8249.145 189.04 8249.425 330.07 ;
      RECT 8248.585 187.94 8248.865 329.83 ;
      RECT 8248.025 189.04 8248.305 329.59 ;
      RECT 8247.465 189.04 8247.745 329.35 ;
      RECT 8246.905 189.04 8247.185 329.11 ;
      RECT 8246.345 189.04 8246.625 328.87 ;
      RECT 8245.785 189.04 8246.065 328.63 ;
      RECT 8245.225 189.04 8245.505 328.39 ;
      RECT 8244.665 189.04 8244.945 328.15 ;
      RECT 8244.105 189.04 8244.385 327.91 ;
      RECT 8243.545 189.04 8243.825 327.67 ;
      RECT 8242.985 189.04 8243.265 327.43 ;
      RECT 8242.425 189.04 8242.705 327.19 ;
      RECT 8203.225 189.04 8203.505 334.095 ;
      RECT 8202.665 189.04 8202.945 334.335 ;
      RECT 8202.105 189.04 8202.385 334.575 ;
      RECT 8201.545 187.94 8201.825 334.815 ;
      RECT 8200.985 189.04 8201.265 335.055 ;
      RECT 8200.425 187.94 8200.705 335.295 ;
      RECT 8199.865 189.04 8200.145 335.535 ;
      RECT 8199.305 189.04 8199.585 335.775 ;
      RECT 8198.745 189.04 8199.025 336.015 ;
      RECT 8198.185 187.94 8198.465 336.255 ;
      RECT 8197.625 189.04 8197.905 336.495 ;
      RECT 8197.065 187.94 8197.345 336.735 ;
      RECT 8196.505 189.04 8196.785 336.975 ;
      RECT 8195.945 187.94 8196.225 337.215 ;
      RECT 8195.385 189.04 8195.665 337.455 ;
      RECT 8194.825 189.04 8195.105 337.695 ;
      RECT 8194.265 189.04 8194.545 337.695 ;
      RECT 8193.705 189.04 8193.985 337.455 ;
      RECT 8193.145 189.04 8193.425 337.215 ;
      RECT 8192.585 189.04 8192.865 336.975 ;
      RECT 8192.025 189.04 8192.305 336.735 ;
      RECT 8191.465 189.04 8191.745 336.495 ;
      RECT 8190.905 189.04 8191.185 336.255 ;
      RECT 8190.345 189.04 8190.625 336.015 ;
      RECT 8189.785 189.04 8190.065 335.775 ;
      RECT 8180.825 189.04 8181.105 335.29 ;
      RECT 8180.265 187.94 8180.545 335.05 ;
      RECT 8179.705 189.04 8179.985 334.81 ;
      RECT 8179.145 187.94 8179.425 334.57 ;
      RECT 8178.585 189.04 8178.865 334.33 ;
      RECT 8178.025 187.94 8178.305 334.09 ;
      RECT 8177.465 189.04 8177.745 333.85 ;
      RECT 8176.905 189.04 8177.185 333.61 ;
      RECT 8176.345 189.04 8176.625 333.37 ;
      RECT 8175.785 189.04 8176.065 333.13 ;
      RECT 8175.225 189.04 8175.505 332.89 ;
      RECT 8174.665 189.04 8174.945 332.65 ;
      RECT 8174.105 189.04 8174.385 332.41 ;
      RECT 8173.545 189.04 8173.825 332.17 ;
      RECT 8171.025 187.94 8171.305 333.89 ;
      RECT 8170.465 189.04 8170.745 333.65 ;
      RECT 8169.905 187.94 8170.185 333.41 ;
      RECT 8169.345 189.04 8169.625 333.17 ;
      RECT 8168.785 189.04 8169.065 332.93 ;
      RECT 8168.225 189.04 8168.505 332.69 ;
      RECT 8167.665 189.04 8167.945 332.45 ;
      RECT 8167.105 189.04 8167.385 332.21 ;
      RECT 8141.065 189.04 8141.345 329.86 ;
      RECT 8140.505 189.04 8140.785 330.1 ;
      RECT 8139.945 189.04 8140.225 330.34 ;
      RECT 8139.385 189.04 8139.665 330.585 ;
      RECT 8138.825 189.04 8139.105 330.825 ;
      RECT 8138.265 189.04 8138.545 331.065 ;
      RECT 8137.705 189.04 8137.985 331.065 ;
      RECT 8137.145 189.04 8137.425 330.825 ;
      RECT 8136.585 189.04 8136.865 330.585 ;
      RECT 8136.025 187.94 8136.305 330.345 ;
      RECT 8135.465 189.04 8135.745 330.105 ;
      RECT 8134.905 187.94 8135.185 329.865 ;
      RECT 8134.345 189.04 8134.625 329.625 ;
      RECT 8133.785 189.04 8134.065 329.385 ;
      RECT 8133.225 189.04 8133.505 329.145 ;
      RECT 8132.665 187.94 8132.945 328.905 ;
      RECT 8132.105 189.04 8132.385 328.665 ;
      RECT 8131.545 187.94 8131.825 328.425 ;
      RECT 8130.985 189.04 8131.265 328.185 ;
      RECT 8130.425 187.94 8130.705 327.945 ;
      RECT 8129.865 189.04 8130.145 327.705 ;
      RECT 8129.305 189.04 8129.585 327.465 ;
      RECT 8128.745 189.04 8129.025 327.225 ;
      RECT 8128.185 189.04 8128.465 326.985 ;
      RECT 8114.745 189.04 8115.025 332.785 ;
      RECT 8114.185 189.04 8114.465 332.545 ;
      RECT 8113.625 189.04 8113.905 332.305 ;
      RECT 8113.065 189.04 8113.345 332.065 ;
      RECT 8112.505 189.04 8112.785 331.825 ;
      RECT 8111.945 189.04 8112.225 331.585 ;
      RECT 8111.385 189.04 8111.665 331.345 ;
      RECT 8110.825 189.04 8111.105 331.105 ;
      RECT 8110.265 187.94 8110.545 330.865 ;
      RECT 8109.705 189.04 8109.985 330.625 ;
      RECT 8109.145 187.94 8109.425 330.305 ;
      RECT 8108.585 189.04 8108.865 330.145 ;
      RECT 8108.025 187.94 8108.305 329.905 ;
      RECT 8107.465 189.04 8107.745 329.665 ;
      RECT 8106.905 189.04 8107.185 329.425 ;
      RECT 8106.345 189.04 8106.625 329.185 ;
      RECT 8105.785 189.04 8106.065 328.945 ;
      RECT 8105.225 189.04 8105.505 328.705 ;
      RECT 8104.665 189.04 8104.945 328.465 ;
      RECT 8104.105 189.04 8104.385 328.225 ;
      RECT 8103.545 189.04 8103.825 327.985 ;
      RECT 8102.985 187.94 8103.265 327.745 ;
      RECT 8102.425 189.04 8102.705 327.505 ;
      RECT 8101.865 187.94 8102.145 327.265 ;
      RECT 8062.665 189.04 8062.945 332.875 ;
      RECT 8062.105 189.04 8062.385 333.115 ;
      RECT 8061.545 189.04 8061.825 333.355 ;
      RECT 8060.985 189.04 8061.265 333.595 ;
      RECT 8060.425 189.04 8060.705 333.835 ;
      RECT 8059.865 189.04 8060.145 334.075 ;
      RECT 8059.305 189.04 8059.585 334.315 ;
      RECT 8058.745 189.04 8059.025 334.555 ;
      RECT 8058.185 189.04 8058.465 334.795 ;
      RECT 8057.625 189.04 8057.905 335.035 ;
      RECT 8057.065 189.04 8057.345 335.275 ;
      RECT 8056.505 189.04 8056.785 335.515 ;
      RECT 8055.945 189.04 8056.225 335.755 ;
      RECT 8055.385 189.04 8055.665 335.755 ;
      RECT 8054.825 187.94 8055.105 335.515 ;
      RECT 8054.265 189.04 8054.545 335.275 ;
      RECT 8053.705 187.94 8053.985 335.035 ;
      RECT 8053.145 189.04 8053.425 334.795 ;
      RECT 8052.585 189.04 8052.865 334.555 ;
      RECT 8052.025 189.04 8052.305 334.315 ;
      RECT 8051.465 187.94 8051.745 334.05 ;
      RECT 8050.905 189.04 8051.185 333.81 ;
      RECT 8050.345 187.94 8050.625 333.57 ;
      RECT 8049.785 189.04 8050.065 333.33 ;
      RECT 8040.825 187.94 8041.105 327.165 ;
      RECT 8040.265 189.04 8040.545 327.405 ;
      RECT 8039.705 189.04 8039.985 327.645 ;
      RECT 8039.145 189.04 8039.425 327.645 ;
      RECT 8038.585 189.04 8038.865 327.405 ;
      RECT 8038.025 189.04 8038.305 327.165 ;
      RECT 8037.465 189.04 8037.745 326.925 ;
      RECT 8036.905 189.04 8037.185 326.685 ;
      RECT 8036.345 189.04 8036.625 326.445 ;
      RECT 8035.785 189.04 8036.065 326.205 ;
      RECT 8035.225 189.04 8035.505 325.965 ;
      RECT 8034.665 189.04 8034.945 325.725 ;
      RECT 8034.105 189.04 8034.385 325.485 ;
      RECT 8033.545 187.94 8033.825 325.245 ;
      RECT 8031.025 189.04 8031.305 326.965 ;
      RECT 8030.465 187.94 8030.745 326.725 ;
      RECT 8029.905 189.04 8030.185 326.485 ;
      RECT 8029.345 187.94 8029.625 326.245 ;
      RECT 8028.785 189.04 8029.065 326.005 ;
      RECT 8028.225 189.04 8028.505 325.765 ;
      RECT 8027.665 189.04 8027.945 325.525 ;
      RECT 8001.625 189.04 8001.905 328.31 ;
      RECT 8001.065 189.04 8001.345 328.55 ;
      RECT 8000.505 189.04 8000.785 328.79 ;
      RECT 7999.945 189.04 8000.225 329.03 ;
      RECT 7999.385 189.04 7999.665 329.27 ;
      RECT 7998.825 187.94 7999.105 329.51 ;
      RECT 7998.265 189.04 7998.545 329.75 ;
      RECT 7997.705 187.94 7997.985 329.99 ;
      RECT 7997.145 189.04 7997.425 330.23 ;
      RECT 7996.585 189.04 7996.865 330.47 ;
      RECT 7996.025 189.04 7996.305 330.71 ;
      RECT 7995.465 189.04 7995.745 330.95 ;
      RECT 7994.905 189.04 7995.185 331.19 ;
      RECT 7994.345 189.04 7994.625 331.43 ;
      RECT 7993.785 189.04 7994.065 331.67 ;
      RECT 7993.225 189.04 7993.505 331.67 ;
      RECT 7992.665 189.04 7992.945 331.43 ;
      RECT 7992.105 189.04 7992.385 331.19 ;
      RECT 7991.545 189.04 7991.825 330.95 ;
      RECT 7990.985 189.04 7991.265 330.705 ;
      RECT 7990.425 189.04 7990.705 330.465 ;
      RECT 7989.865 189.04 7990.145 330.225 ;
      RECT 7989.305 187.94 7989.585 329.985 ;
      RECT 7988.745 189.04 7989.025 329.745 ;
      RECT 7975.305 187.94 7975.585 327.225 ;
      RECT 7974.745 189.04 7975.025 326.985 ;
      RECT 7974.185 189.04 7974.465 326.745 ;
      RECT 7973.625 189.04 7973.905 326.505 ;
      RECT 7973.065 187.94 7973.345 326.265 ;
      RECT 7972.505 189.04 7972.785 326.025 ;
      RECT 7971.945 187.94 7972.225 325.785 ;
      RECT 7971.385 189.04 7971.665 325.545 ;
      RECT 7970.825 187.94 7971.105 325.305 ;
      RECT 7970.265 189.04 7970.545 325.065 ;
      RECT 7969.705 189.04 7969.985 324.825 ;
      RECT 7969.145 189.04 7969.425 324.585 ;
      RECT 7968.585 189.04 7968.865 324.345 ;
      RECT 7968.025 189.04 7968.305 324.105 ;
      RECT 7967.465 189.04 7967.745 323.865 ;
      RECT 7966.905 189.04 7967.185 323.625 ;
      RECT 7966.345 189.04 7966.625 323.385 ;
      RECT 7965.785 189.04 7966.065 323.145 ;
      RECT 7965.225 189.04 7965.505 322.905 ;
      RECT 7964.665 189.04 7964.945 322.665 ;
      RECT 7964.105 189.04 7964.385 322.425 ;
      RECT 7963.545 187.94 7963.825 322.185 ;
      RECT 7962.985 189.04 7963.265 321.945 ;
      RECT 7962.425 187.94 7962.705 321.705 ;
      RECT 7922.665 189.04 7922.945 332.175 ;
      RECT 7922.105 187.94 7922.385 332.415 ;
      RECT 7921.545 189.04 7921.825 332.655 ;
      RECT 7920.985 189.04 7921.265 332.895 ;
      RECT 7920.425 189.04 7920.705 333.135 ;
      RECT 7919.865 189.04 7920.145 333.375 ;
      RECT 7919.305 189.04 7919.585 333.615 ;
      RECT 7918.745 189.04 7919.025 333.86 ;
      RECT 7918.185 189.04 7918.465 334.1 ;
      RECT 7917.625 189.04 7917.905 334.34 ;
      RECT 7917.065 187.94 7917.345 334.58 ;
      RECT 7916.505 189.04 7916.785 334.82 ;
      RECT 7915.945 187.94 7916.225 335.06 ;
      RECT 7915.385 189.04 7915.665 335.3 ;
      RECT 7914.825 189.04 7915.105 335.54 ;
      RECT 7914.265 189.04 7914.545 335.78 ;
      RECT 7913.705 189.04 7913.985 336.02 ;
      RECT 7913.145 189.04 7913.425 336.26 ;
      RECT 7912.585 189.04 7912.865 336.5 ;
      RECT 7912.025 189.04 7912.305 336.74 ;
      RECT 7911.465 189.04 7911.745 336.98 ;
      RECT 7910.905 189.04 7911.185 337.22 ;
      RECT 7910.345 189.04 7910.625 337.46 ;
      RECT 7909.785 189.04 7910.065 337.7 ;
      RECT 7900.825 189.04 7901.105 333.285 ;
      RECT 7900.265 189.04 7900.545 333.045 ;
      RECT 7899.705 189.04 7899.985 332.805 ;
      RECT 7899.145 187.94 7899.425 332.565 ;
      RECT 7898.585 189.04 7898.865 332.325 ;
      RECT 7898.025 187.94 7898.305 332.085 ;
      RECT 7897.465 189.04 7897.745 331.845 ;
      RECT 7896.905 189.04 7897.185 331.605 ;
      RECT 7896.345 189.04 7896.625 331.365 ;
      RECT 7895.785 187.94 7896.065 331.125 ;
      RECT 7895.225 189.04 7895.505 330.885 ;
      RECT 7894.665 187.94 7894.945 330.645 ;
      RECT 7894.105 189.04 7894.385 330.405 ;
      RECT 7893.545 187.94 7893.825 330.165 ;
      RECT 7891.025 189.04 7891.305 322.565 ;
      RECT 7890.465 189.04 7890.745 322.325 ;
      RECT 7889.905 189.04 7890.185 322.085 ;
      RECT 7889.345 189.04 7889.625 321.845 ;
      RECT 7888.785 189.04 7889.065 321.605 ;
      RECT 7888.225 189.04 7888.505 321.365 ;
      RECT 7887.665 189.04 7887.945 321.125 ;
      RECT 7861.625 189.04 7861.905 335 ;
      RECT 7861.065 189.04 7861.345 335.24 ;
      RECT 7860.505 189.04 7860.785 335.48 ;
      RECT 7859.945 189.04 7860.225 335.72 ;
      RECT 7859.385 189.04 7859.665 335.96 ;
      RECT 7858.825 187.94 7859.105 335.96 ;
      RECT 7858.265 189.04 7858.545 335.72 ;
      RECT 7857.705 187.94 7857.985 335.475 ;
      RECT 7857.145 189.04 7857.425 335.235 ;
      RECT 7856.585 187.94 7856.865 334.995 ;
      RECT 7856.025 189.04 7856.305 334.755 ;
      RECT 7855.465 189.04 7855.745 334.515 ;
      RECT 7854.905 189.04 7855.185 334.275 ;
      RECT 7854.345 189.04 7854.625 334.035 ;
      RECT 7853.785 189.04 7854.065 333.795 ;
      RECT 7853.225 189.04 7853.505 333.555 ;
      RECT 7852.665 189.04 7852.945 333.315 ;
      RECT 7852.105 189.04 7852.385 333.075 ;
      RECT 7851.545 187.94 7851.825 332.835 ;
      RECT 7850.985 189.04 7851.265 332.595 ;
      RECT 7850.425 187.94 7850.705 332.355 ;
      RECT 7849.865 189.04 7850.145 332.115 ;
      RECT 7849.305 189.04 7849.585 331.875 ;
      RECT 7848.745 189.04 7849.025 331.635 ;
      RECT 7835.305 189.04 7835.585 335.035 ;
      RECT 7834.745 189.04 7835.025 335.275 ;
      RECT 7834.185 189.04 7834.465 335.52 ;
      RECT 7833.625 189.04 7833.905 335.76 ;
      RECT 7833.065 189.04 7833.345 336 ;
      RECT 7832.505 189.04 7832.785 336 ;
      RECT 7831.945 189.04 7832.225 335.76 ;
      RECT 7831.385 189.04 7831.665 335.52 ;
      RECT 7830.825 189.04 7831.105 328.505 ;
      RECT 7830.265 189.04 7830.545 328.265 ;
      RECT 7829.705 189.04 7829.985 328.025 ;
      RECT 7829.145 187.94 7829.425 327.785 ;
      RECT 7828.585 189.04 7828.865 327.545 ;
      RECT 7828.025 187.94 7828.305 327.305 ;
      RECT 7827.465 189.04 7827.745 327.065 ;
      RECT 7826.905 189.04 7827.185 326.825 ;
      RECT 7826.345 189.04 7826.625 326.585 ;
      RECT 7825.785 187.94 7826.065 326.345 ;
      RECT 7825.225 189.04 7825.505 326.105 ;
      RECT 7824.665 187.94 7824.945 325.865 ;
      RECT 7824.105 189.04 7824.385 325.625 ;
      RECT 7823.545 187.94 7823.825 325.385 ;
      RECT 7822.985 189.04 7823.265 325.145 ;
      RECT 7822.425 189.04 7822.705 324.905 ;
      RECT 7782.105 189.04 7782.385 333.8 ;
      RECT 7781.545 189.04 7781.825 334.04 ;
      RECT 7780.985 189.04 7781.265 334.285 ;
      RECT 7780.425 189.04 7780.705 334.525 ;
      RECT 7779.865 189.04 7780.145 334.765 ;
      RECT 7779.305 189.04 7779.585 335.005 ;
      RECT 7778.745 189.04 7779.025 335.245 ;
      RECT 7778.185 189.04 7778.465 335.485 ;
      RECT 7777.625 189.04 7777.905 335.725 ;
      RECT 7777.065 189.04 7777.345 335.965 ;
      RECT 7776.505 187.94 7776.785 336.205 ;
      RECT 7775.945 189.04 7776.225 336.445 ;
      RECT 7775.385 187.94 7775.665 336.685 ;
      RECT 7774.825 189.04 7775.105 336.925 ;
      RECT 7774.265 187.94 7774.545 337.165 ;
      RECT 7773.705 189.04 7773.985 337.165 ;
      RECT 7773.145 189.04 7773.425 336.925 ;
      RECT 7772.585 189.04 7772.865 336.685 ;
      RECT 7772.025 189.04 7772.305 336.445 ;
      RECT 7771.465 189.04 7771.745 336.205 ;
      RECT 7770.905 189.04 7771.185 335.965 ;
      RECT 7770.345 189.04 7770.625 335.725 ;
      RECT 7769.785 189.04 7770.065 335.485 ;
      RECT 7760.825 187.94 7761.105 335.515 ;
      RECT 7760.265 189.04 7760.545 335.755 ;
      RECT 7759.705 187.94 7759.985 335.995 ;
      RECT 7759.145 189.04 7759.425 336.21 ;
      RECT 7758.585 189.04 7758.865 335.785 ;
      RECT 7758.025 189.04 7758.305 335.545 ;
      RECT 7757.465 189.04 7757.745 335.305 ;
      RECT 7756.905 189.04 7757.185 335.065 ;
      RECT 7756.345 189.04 7756.625 334.825 ;
      RECT 7755.785 189.04 7756.065 334.585 ;
      RECT 7755.225 189.04 7755.505 334.345 ;
      RECT 7754.665 189.04 7754.945 334.105 ;
      RECT 7754.105 189.04 7754.385 333.865 ;
      RECT 7753.545 189.04 7753.825 333.625 ;
      RECT 7751.025 189.04 7751.305 332.8 ;
      RECT 7750.465 189.04 7750.745 332.56 ;
      RECT 7749.905 189.04 7750.185 332.32 ;
      RECT 7749.345 187.94 7749.625 332.08 ;
      RECT 7748.785 189.04 7749.065 331.84 ;
      RECT 7748.225 187.94 7748.505 331.6 ;
      RECT 7747.665 189.04 7747.945 331.36 ;
      RECT 7747.105 189.04 7747.385 331.12 ;
      RECT 7720.505 189.04 7720.785 342.165 ;
      RECT 7719.945 187.94 7720.225 342.405 ;
      RECT 7719.385 189.04 7719.665 342.645 ;
      RECT 7718.825 187.94 7719.105 342.89 ;
      RECT 7718.265 189.04 7718.545 343.13 ;
      RECT 7717.705 187.94 7717.985 343.37 ;
      RECT 7717.145 189.04 7717.425 343.61 ;
      RECT 7716.585 189.04 7716.865 343.85 ;
      RECT 7716.025 189.04 7716.305 329.47 ;
      RECT 7715.465 189.04 7715.745 329.23 ;
      RECT 7714.905 189.04 7715.185 328.99 ;
      RECT 7714.345 189.04 7714.625 328.75 ;
      RECT 7713.785 189.04 7714.065 328.51 ;
      RECT 7713.225 189.04 7713.505 328.27 ;
      RECT 7712.665 189.04 7712.945 328.03 ;
      RECT 7712.105 189.04 7712.385 327.79 ;
      RECT 7711.545 189.04 7711.825 327.55 ;
      RECT 7710.985 189.04 7711.265 327.31 ;
      RECT 7710.425 187.94 7710.705 327.07 ;
      RECT 7709.865 189.04 7710.145 326.83 ;
      RECT 7709.305 187.94 7709.585 326.59 ;
      RECT 7708.745 189.04 7709.025 326.35 ;
      RECT 7694.745 187.94 7695.025 332.47 ;
      RECT 7694.185 189.04 7694.465 332.23 ;
      RECT 7693.625 189.04 7693.905 331.99 ;
      RECT 7693.065 189.04 7693.345 331.75 ;
      RECT 7692.505 189.04 7692.785 331.51 ;
      RECT 7691.945 189.04 7692.225 331.27 ;
      RECT 7691.385 189.04 7691.665 331.03 ;
      RECT 7690.825 189.04 7691.105 330.79 ;
      RECT 7690.265 189.04 7690.545 330.55 ;
      RECT 7689.705 187.94 7689.985 330.31 ;
      RECT 7689.145 189.04 7689.425 330.07 ;
      RECT 7688.585 187.94 7688.865 329.83 ;
      RECT 7688.025 189.04 7688.305 329.59 ;
      RECT 7687.465 189.04 7687.745 329.35 ;
      RECT 7686.905 189.04 7687.185 329.11 ;
      RECT 7686.345 189.04 7686.625 328.87 ;
      RECT 7685.785 189.04 7686.065 328.63 ;
      RECT 7685.225 189.04 7685.505 328.39 ;
      RECT 7684.665 189.04 7684.945 328.15 ;
      RECT 7684.105 189.04 7684.385 327.91 ;
      RECT 7683.545 189.04 7683.825 327.67 ;
      RECT 7682.985 189.04 7683.265 327.43 ;
      RECT 7682.425 189.04 7682.705 327.19 ;
      RECT 7643.225 189.04 7643.505 334.095 ;
      RECT 7642.665 189.04 7642.945 334.335 ;
      RECT 7642.105 189.04 7642.385 334.575 ;
      RECT 7641.545 187.94 7641.825 334.815 ;
      RECT 7640.985 189.04 7641.265 335.055 ;
      RECT 7640.425 187.94 7640.705 335.295 ;
      RECT 7639.865 189.04 7640.145 335.535 ;
      RECT 7639.305 189.04 7639.585 335.775 ;
      RECT 7638.745 189.04 7639.025 336.015 ;
      RECT 7638.185 187.94 7638.465 336.255 ;
      RECT 7637.625 189.04 7637.905 336.495 ;
      RECT 7637.065 187.94 7637.345 336.735 ;
      RECT 7636.505 189.04 7636.785 336.975 ;
      RECT 7635.945 187.94 7636.225 337.215 ;
      RECT 7635.385 189.04 7635.665 337.455 ;
      RECT 7634.825 189.04 7635.105 337.695 ;
      RECT 7634.265 189.04 7634.545 337.695 ;
      RECT 7633.705 189.04 7633.985 337.455 ;
      RECT 7633.145 189.04 7633.425 337.215 ;
      RECT 7632.585 189.04 7632.865 336.975 ;
      RECT 7632.025 189.04 7632.305 336.735 ;
      RECT 7631.465 189.04 7631.745 336.495 ;
      RECT 7630.905 189.04 7631.185 336.255 ;
      RECT 7630.345 189.04 7630.625 336.015 ;
      RECT 7629.785 189.04 7630.065 335.775 ;
      RECT 7620.825 189.04 7621.105 335.29 ;
      RECT 7620.265 187.94 7620.545 335.05 ;
      RECT 7619.705 189.04 7619.985 334.81 ;
      RECT 7619.145 187.94 7619.425 334.57 ;
      RECT 7618.585 189.04 7618.865 334.33 ;
      RECT 7618.025 187.94 7618.305 334.09 ;
      RECT 7617.465 189.04 7617.745 333.85 ;
      RECT 7616.905 189.04 7617.185 333.61 ;
      RECT 7616.345 189.04 7616.625 333.37 ;
      RECT 7615.785 189.04 7616.065 333.13 ;
      RECT 7615.225 189.04 7615.505 332.89 ;
      RECT 7614.665 189.04 7614.945 332.65 ;
      RECT 7614.105 189.04 7614.385 332.41 ;
      RECT 7613.545 189.04 7613.825 332.17 ;
      RECT 7611.025 187.94 7611.305 333.89 ;
      RECT 7610.465 189.04 7610.745 333.65 ;
      RECT 7609.905 187.94 7610.185 333.41 ;
      RECT 7609.345 189.04 7609.625 333.17 ;
      RECT 7608.785 189.04 7609.065 332.93 ;
      RECT 7608.225 189.04 7608.505 332.69 ;
      RECT 7607.665 189.04 7607.945 332.45 ;
      RECT 7607.105 189.04 7607.385 332.21 ;
      RECT 7581.065 189.04 7581.345 329.86 ;
      RECT 7580.505 189.04 7580.785 330.1 ;
      RECT 7579.945 189.04 7580.225 330.34 ;
      RECT 7579.385 189.04 7579.665 330.585 ;
      RECT 7578.825 189.04 7579.105 330.825 ;
      RECT 7578.265 189.04 7578.545 331.065 ;
      RECT 7577.705 189.04 7577.985 331.065 ;
      RECT 7577.145 189.04 7577.425 330.825 ;
      RECT 7576.585 189.04 7576.865 330.585 ;
      RECT 7576.025 187.94 7576.305 330.345 ;
      RECT 7575.465 189.04 7575.745 330.105 ;
      RECT 7574.905 187.94 7575.185 329.865 ;
      RECT 7574.345 189.04 7574.625 329.625 ;
      RECT 7573.785 189.04 7574.065 329.385 ;
      RECT 7573.225 189.04 7573.505 329.145 ;
      RECT 7572.665 187.94 7572.945 328.905 ;
      RECT 7572.105 189.04 7572.385 328.665 ;
      RECT 7571.545 187.94 7571.825 328.425 ;
      RECT 7570.985 189.04 7571.265 328.185 ;
      RECT 7570.425 187.94 7570.705 327.945 ;
      RECT 7569.865 189.04 7570.145 327.705 ;
      RECT 7569.305 189.04 7569.585 327.465 ;
      RECT 7568.745 189.04 7569.025 327.225 ;
      RECT 7568.185 189.04 7568.465 326.985 ;
      RECT 7554.745 189.04 7555.025 332.785 ;
      RECT 7554.185 189.04 7554.465 332.545 ;
      RECT 7553.625 189.04 7553.905 332.305 ;
      RECT 7553.065 189.04 7553.345 332.065 ;
      RECT 7552.505 189.04 7552.785 331.825 ;
      RECT 7551.945 189.04 7552.225 331.585 ;
      RECT 7551.385 189.04 7551.665 331.345 ;
      RECT 7550.825 189.04 7551.105 331.105 ;
      RECT 7550.265 187.94 7550.545 330.865 ;
      RECT 7549.705 189.04 7549.985 330.625 ;
      RECT 7549.145 187.94 7549.425 330.305 ;
      RECT 7548.585 189.04 7548.865 330.145 ;
      RECT 7548.025 187.94 7548.305 329.905 ;
      RECT 7547.465 189.04 7547.745 329.665 ;
      RECT 7546.905 189.04 7547.185 329.425 ;
      RECT 7546.345 189.04 7546.625 329.185 ;
      RECT 7545.785 189.04 7546.065 328.945 ;
      RECT 7545.225 189.04 7545.505 328.705 ;
      RECT 7544.665 189.04 7544.945 328.465 ;
      RECT 7544.105 189.04 7544.385 328.225 ;
      RECT 7543.545 189.04 7543.825 327.985 ;
      RECT 7542.985 187.94 7543.265 327.745 ;
      RECT 7542.425 189.04 7542.705 327.505 ;
      RECT 7541.865 187.94 7542.145 327.265 ;
      RECT 7502.665 189.04 7502.945 332.875 ;
      RECT 7502.105 189.04 7502.385 333.115 ;
      RECT 7501.545 189.04 7501.825 333.355 ;
      RECT 7500.985 189.04 7501.265 333.595 ;
      RECT 7500.425 189.04 7500.705 333.835 ;
      RECT 7499.865 189.04 7500.145 334.075 ;
      RECT 7499.305 189.04 7499.585 334.315 ;
      RECT 7498.745 189.04 7499.025 334.555 ;
      RECT 7498.185 189.04 7498.465 334.795 ;
      RECT 7497.625 189.04 7497.905 335.035 ;
      RECT 7497.065 189.04 7497.345 335.275 ;
      RECT 7496.505 189.04 7496.785 335.515 ;
      RECT 7495.945 189.04 7496.225 335.755 ;
      RECT 7495.385 189.04 7495.665 335.755 ;
      RECT 7494.825 187.94 7495.105 335.515 ;
      RECT 7494.265 189.04 7494.545 335.275 ;
      RECT 7493.705 187.94 7493.985 335.035 ;
      RECT 7493.145 189.04 7493.425 334.795 ;
      RECT 7492.585 189.04 7492.865 334.555 ;
      RECT 7492.025 189.04 7492.305 334.315 ;
      RECT 7491.465 187.94 7491.745 334.05 ;
      RECT 7490.905 189.04 7491.185 333.81 ;
      RECT 7490.345 187.94 7490.625 333.57 ;
      RECT 7489.785 189.04 7490.065 333.33 ;
      RECT 7480.825 187.94 7481.105 327.165 ;
      RECT 7480.265 189.04 7480.545 327.405 ;
      RECT 7479.705 189.04 7479.985 327.645 ;
      RECT 7479.145 189.04 7479.425 327.645 ;
      RECT 7478.585 189.04 7478.865 327.405 ;
      RECT 7478.025 189.04 7478.305 327.165 ;
      RECT 7477.465 189.04 7477.745 326.925 ;
      RECT 7476.905 189.04 7477.185 326.685 ;
      RECT 7476.345 189.04 7476.625 326.445 ;
      RECT 7475.785 189.04 7476.065 326.205 ;
      RECT 7475.225 189.04 7475.505 325.965 ;
      RECT 7474.665 189.04 7474.945 325.725 ;
      RECT 7474.105 189.04 7474.385 325.485 ;
      RECT 7473.545 187.94 7473.825 325.245 ;
      RECT 7471.025 189.04 7471.305 326.965 ;
      RECT 7470.465 187.94 7470.745 326.725 ;
      RECT 7469.905 189.04 7470.185 326.485 ;
      RECT 7469.345 187.94 7469.625 326.245 ;
      RECT 7468.785 189.04 7469.065 326.005 ;
      RECT 7468.225 189.04 7468.505 325.765 ;
      RECT 7467.665 189.04 7467.945 325.525 ;
      RECT 7441.625 189.04 7441.905 328.31 ;
      RECT 7441.065 189.04 7441.345 328.55 ;
      RECT 7440.505 189.04 7440.785 328.79 ;
      RECT 7439.945 189.04 7440.225 329.03 ;
      RECT 7439.385 189.04 7439.665 329.27 ;
      RECT 7438.825 187.94 7439.105 329.51 ;
      RECT 7438.265 189.04 7438.545 329.75 ;
      RECT 7437.705 187.94 7437.985 329.99 ;
      RECT 7437.145 189.04 7437.425 330.23 ;
      RECT 7436.585 189.04 7436.865 330.47 ;
      RECT 7436.025 189.04 7436.305 330.71 ;
      RECT 7435.465 189.04 7435.745 330.95 ;
      RECT 7434.905 189.04 7435.185 331.19 ;
      RECT 7434.345 189.04 7434.625 331.43 ;
      RECT 7433.785 189.04 7434.065 331.67 ;
      RECT 7433.225 189.04 7433.505 331.67 ;
      RECT 7432.665 189.04 7432.945 331.43 ;
      RECT 7432.105 189.04 7432.385 331.19 ;
      RECT 7431.545 189.04 7431.825 330.95 ;
      RECT 7430.985 189.04 7431.265 330.705 ;
      RECT 7430.425 189.04 7430.705 330.465 ;
      RECT 7429.865 189.04 7430.145 330.225 ;
      RECT 7429.305 187.94 7429.585 329.985 ;
      RECT 7428.745 189.04 7429.025 329.745 ;
      RECT 7415.305 187.94 7415.585 327.225 ;
      RECT 7414.745 189.04 7415.025 326.985 ;
      RECT 7414.185 189.04 7414.465 326.745 ;
      RECT 7413.625 189.04 7413.905 326.505 ;
      RECT 7413.065 187.94 7413.345 326.265 ;
      RECT 7412.505 189.04 7412.785 326.025 ;
      RECT 7411.945 187.94 7412.225 325.785 ;
      RECT 7411.385 189.04 7411.665 325.545 ;
      RECT 7410.825 187.94 7411.105 325.305 ;
      RECT 7410.265 189.04 7410.545 325.065 ;
      RECT 7409.705 189.04 7409.985 324.825 ;
      RECT 7409.145 189.04 7409.425 324.585 ;
      RECT 7408.585 189.04 7408.865 324.345 ;
      RECT 7408.025 189.04 7408.305 324.105 ;
      RECT 7407.465 189.04 7407.745 323.865 ;
      RECT 7406.905 189.04 7407.185 323.625 ;
      RECT 7406.345 189.04 7406.625 323.385 ;
      RECT 7405.785 189.04 7406.065 323.145 ;
      RECT 7405.225 189.04 7405.505 322.905 ;
      RECT 7404.665 189.04 7404.945 322.665 ;
      RECT 7404.105 189.04 7404.385 322.425 ;
      RECT 7403.545 187.94 7403.825 322.185 ;
      RECT 7402.985 189.04 7403.265 321.945 ;
      RECT 7402.425 187.94 7402.705 321.705 ;
      RECT 7362.665 189.04 7362.945 332.175 ;
      RECT 7362.105 187.94 7362.385 332.415 ;
      RECT 7361.545 189.04 7361.825 332.655 ;
      RECT 7360.985 189.04 7361.265 332.895 ;
      RECT 7360.425 189.04 7360.705 333.135 ;
      RECT 7359.865 189.04 7360.145 333.375 ;
      RECT 7359.305 189.04 7359.585 333.615 ;
      RECT 7358.745 189.04 7359.025 333.86 ;
      RECT 7358.185 189.04 7358.465 334.1 ;
      RECT 7357.625 189.04 7357.905 334.34 ;
      RECT 7357.065 187.94 7357.345 334.58 ;
      RECT 7356.505 189.04 7356.785 334.82 ;
      RECT 7355.945 187.94 7356.225 335.06 ;
      RECT 7355.385 189.04 7355.665 335.3 ;
      RECT 7354.825 189.04 7355.105 335.54 ;
      RECT 7354.265 189.04 7354.545 335.78 ;
      RECT 7353.705 189.04 7353.985 336.02 ;
      RECT 7353.145 189.04 7353.425 336.26 ;
      RECT 7352.585 189.04 7352.865 336.5 ;
      RECT 7352.025 189.04 7352.305 336.74 ;
      RECT 7351.465 189.04 7351.745 336.98 ;
      RECT 7350.905 189.04 7351.185 337.22 ;
      RECT 7350.345 189.04 7350.625 337.46 ;
      RECT 7349.785 189.04 7350.065 337.7 ;
      RECT 7340.825 189.04 7341.105 333.285 ;
      RECT 7340.265 189.04 7340.545 333.045 ;
      RECT 7339.705 189.04 7339.985 332.805 ;
      RECT 7339.145 187.94 7339.425 332.565 ;
      RECT 7338.585 189.04 7338.865 332.325 ;
      RECT 7338.025 187.94 7338.305 332.085 ;
      RECT 7337.465 189.04 7337.745 331.845 ;
      RECT 7336.905 189.04 7337.185 331.605 ;
      RECT 7336.345 189.04 7336.625 331.365 ;
      RECT 7335.785 187.94 7336.065 331.125 ;
      RECT 7335.225 189.04 7335.505 330.885 ;
      RECT 7334.665 187.94 7334.945 330.645 ;
      RECT 7334.105 189.04 7334.385 330.405 ;
      RECT 7333.545 187.94 7333.825 330.165 ;
      RECT 7331.025 189.04 7331.305 322.565 ;
      RECT 7330.465 189.04 7330.745 322.325 ;
      RECT 7329.905 189.04 7330.185 322.085 ;
      RECT 7329.345 189.04 7329.625 321.845 ;
      RECT 7328.785 189.04 7329.065 321.605 ;
      RECT 7328.225 189.04 7328.505 321.365 ;
      RECT 7327.665 189.04 7327.945 321.125 ;
      RECT 7301.625 189.04 7301.905 335 ;
      RECT 7301.065 189.04 7301.345 335.24 ;
      RECT 7300.505 189.04 7300.785 335.48 ;
      RECT 7299.945 189.04 7300.225 335.72 ;
      RECT 7299.385 189.04 7299.665 335.96 ;
      RECT 7298.825 187.94 7299.105 335.96 ;
      RECT 7298.265 189.04 7298.545 335.72 ;
      RECT 7297.705 187.94 7297.985 335.475 ;
      RECT 7297.145 189.04 7297.425 335.235 ;
      RECT 7296.585 187.94 7296.865 334.995 ;
      RECT 7296.025 189.04 7296.305 334.755 ;
      RECT 7295.465 189.04 7295.745 334.515 ;
      RECT 7294.905 189.04 7295.185 334.275 ;
      RECT 7294.345 189.04 7294.625 334.035 ;
      RECT 7293.785 189.04 7294.065 333.795 ;
      RECT 7293.225 189.04 7293.505 333.555 ;
      RECT 7292.665 189.04 7292.945 333.315 ;
      RECT 7292.105 189.04 7292.385 333.075 ;
      RECT 7291.545 187.94 7291.825 332.835 ;
      RECT 7290.985 189.04 7291.265 332.595 ;
      RECT 7290.425 187.94 7290.705 332.355 ;
      RECT 7289.865 189.04 7290.145 332.115 ;
      RECT 7289.305 189.04 7289.585 331.875 ;
      RECT 7288.745 189.04 7289.025 331.635 ;
      RECT 7275.305 189.04 7275.585 335.035 ;
      RECT 7274.745 189.04 7275.025 335.275 ;
      RECT 7274.185 189.04 7274.465 335.52 ;
      RECT 7273.625 189.04 7273.905 335.76 ;
      RECT 7273.065 189.04 7273.345 336 ;
      RECT 7272.505 189.04 7272.785 336 ;
      RECT 7271.945 189.04 7272.225 335.76 ;
      RECT 7271.385 189.04 7271.665 335.52 ;
      RECT 7270.825 189.04 7271.105 328.505 ;
      RECT 7270.265 189.04 7270.545 328.265 ;
      RECT 7269.705 189.04 7269.985 328.025 ;
      RECT 7269.145 187.94 7269.425 327.785 ;
      RECT 7268.585 189.04 7268.865 327.545 ;
      RECT 7268.025 187.94 7268.305 327.305 ;
      RECT 7267.465 189.04 7267.745 327.065 ;
      RECT 7266.905 189.04 7267.185 326.825 ;
      RECT 7266.345 189.04 7266.625 326.585 ;
      RECT 7265.785 187.94 7266.065 326.345 ;
      RECT 7265.225 189.04 7265.505 326.105 ;
      RECT 7264.665 187.94 7264.945 325.865 ;
      RECT 7264.105 189.04 7264.385 325.625 ;
      RECT 7263.545 187.94 7263.825 325.385 ;
      RECT 7262.985 189.04 7263.265 325.145 ;
      RECT 7262.425 189.04 7262.705 324.905 ;
      RECT 7222.105 189.04 7222.385 333.8 ;
      RECT 7221.545 189.04 7221.825 334.04 ;
      RECT 7220.985 189.04 7221.265 334.285 ;
      RECT 7220.425 189.04 7220.705 334.525 ;
      RECT 7219.865 189.04 7220.145 334.765 ;
      RECT 7219.305 189.04 7219.585 335.005 ;
      RECT 7218.745 189.04 7219.025 335.245 ;
      RECT 7218.185 189.04 7218.465 335.485 ;
      RECT 7217.625 189.04 7217.905 335.725 ;
      RECT 7217.065 189.04 7217.345 335.965 ;
      RECT 7216.505 187.94 7216.785 336.205 ;
      RECT 7215.945 189.04 7216.225 336.445 ;
      RECT 7215.385 187.94 7215.665 336.685 ;
      RECT 7214.825 189.04 7215.105 336.925 ;
      RECT 7214.265 187.94 7214.545 337.165 ;
      RECT 7213.705 189.04 7213.985 337.165 ;
      RECT 7213.145 189.04 7213.425 336.925 ;
      RECT 7212.585 189.04 7212.865 336.685 ;
      RECT 7212.025 189.04 7212.305 336.445 ;
      RECT 7211.465 189.04 7211.745 336.205 ;
      RECT 7210.905 189.04 7211.185 335.965 ;
      RECT 7210.345 189.04 7210.625 335.725 ;
      RECT 7209.785 189.04 7210.065 335.485 ;
      RECT 7200.825 187.94 7201.105 335.515 ;
      RECT 7200.265 189.04 7200.545 335.755 ;
      RECT 7199.705 187.94 7199.985 335.995 ;
      RECT 7199.145 189.04 7199.425 336.21 ;
      RECT 7198.585 189.04 7198.865 335.785 ;
      RECT 7198.025 189.04 7198.305 335.545 ;
      RECT 7197.465 189.04 7197.745 335.305 ;
      RECT 7196.905 189.04 7197.185 335.065 ;
      RECT 7196.345 189.04 7196.625 334.825 ;
      RECT 7195.785 189.04 7196.065 334.585 ;
      RECT 7195.225 189.04 7195.505 334.345 ;
      RECT 7194.665 189.04 7194.945 334.105 ;
      RECT 7194.105 189.04 7194.385 333.865 ;
      RECT 7193.545 189.04 7193.825 333.625 ;
      RECT 7191.025 189.04 7191.305 332.8 ;
      RECT 7190.465 189.04 7190.745 332.56 ;
      RECT 7189.905 189.04 7190.185 332.32 ;
      RECT 7189.345 187.94 7189.625 332.08 ;
      RECT 7188.785 189.04 7189.065 331.84 ;
      RECT 7188.225 187.94 7188.505 331.6 ;
      RECT 7187.665 189.04 7187.945 331.36 ;
      RECT 7187.105 189.04 7187.385 331.12 ;
      RECT 7160.505 189.04 7160.785 342.165 ;
      RECT 7159.945 187.94 7160.225 342.405 ;
      RECT 7159.385 189.04 7159.665 342.645 ;
      RECT 7158.825 187.94 7159.105 342.89 ;
      RECT 7158.265 189.04 7158.545 343.13 ;
      RECT 7157.705 187.94 7157.985 343.37 ;
      RECT 7157.145 189.04 7157.425 343.61 ;
      RECT 7156.585 189.04 7156.865 343.85 ;
      RECT 7156.025 189.04 7156.305 329.47 ;
      RECT 7155.465 189.04 7155.745 329.23 ;
      RECT 7154.905 189.04 7155.185 328.99 ;
      RECT 7154.345 189.04 7154.625 328.75 ;
      RECT 7153.785 189.04 7154.065 328.51 ;
      RECT 7153.225 189.04 7153.505 328.27 ;
      RECT 7152.665 189.04 7152.945 328.03 ;
      RECT 7152.105 189.04 7152.385 327.79 ;
      RECT 7151.545 189.04 7151.825 327.55 ;
      RECT 7150.985 189.04 7151.265 327.31 ;
      RECT 7150.425 187.94 7150.705 327.07 ;
      RECT 7149.865 189.04 7150.145 326.83 ;
      RECT 7149.305 187.94 7149.585 326.59 ;
      RECT 7148.745 189.04 7149.025 326.35 ;
      RECT 7134.745 187.94 7135.025 332.47 ;
      RECT 7134.185 189.04 7134.465 332.23 ;
      RECT 7133.625 189.04 7133.905 331.99 ;
      RECT 7133.065 189.04 7133.345 331.75 ;
      RECT 7132.505 189.04 7132.785 331.51 ;
      RECT 7131.945 189.04 7132.225 331.27 ;
      RECT 7131.385 189.04 7131.665 331.03 ;
      RECT 7130.825 189.04 7131.105 330.79 ;
      RECT 7130.265 189.04 7130.545 330.55 ;
      RECT 7129.705 187.94 7129.985 330.31 ;
      RECT 7129.145 189.04 7129.425 330.07 ;
      RECT 7128.585 187.94 7128.865 329.83 ;
      RECT 7128.025 189.04 7128.305 329.59 ;
      RECT 7127.465 189.04 7127.745 329.35 ;
      RECT 7126.905 189.04 7127.185 329.11 ;
      RECT 7126.345 189.04 7126.625 328.87 ;
      RECT 7125.785 189.04 7126.065 328.63 ;
      RECT 7125.225 189.04 7125.505 328.39 ;
      RECT 7124.665 189.04 7124.945 328.15 ;
      RECT 7124.105 189.04 7124.385 327.91 ;
      RECT 7123.545 189.04 7123.825 327.67 ;
      RECT 7122.985 189.04 7123.265 327.43 ;
      RECT 7122.425 189.04 7122.705 327.19 ;
      RECT 7083.225 189.04 7083.505 334.095 ;
      RECT 7082.665 189.04 7082.945 334.335 ;
      RECT 7082.105 189.04 7082.385 334.575 ;
      RECT 7081.545 187.94 7081.825 334.815 ;
      RECT 7080.985 189.04 7081.265 335.055 ;
      RECT 7080.425 187.94 7080.705 335.295 ;
      RECT 7079.865 189.04 7080.145 335.535 ;
      RECT 7079.305 189.04 7079.585 335.775 ;
      RECT 7078.745 189.04 7079.025 336.015 ;
      RECT 7078.185 187.94 7078.465 336.255 ;
      RECT 7077.625 189.04 7077.905 336.495 ;
      RECT 7077.065 187.94 7077.345 336.735 ;
      RECT 7076.505 189.04 7076.785 336.975 ;
      RECT 7075.945 187.94 7076.225 337.215 ;
      RECT 7075.385 189.04 7075.665 337.455 ;
      RECT 7074.825 189.04 7075.105 337.695 ;
      RECT 7074.265 189.04 7074.545 337.695 ;
      RECT 7073.705 189.04 7073.985 337.455 ;
      RECT 7073.145 189.04 7073.425 337.215 ;
      RECT 7072.585 189.04 7072.865 336.975 ;
      RECT 7072.025 189.04 7072.305 336.735 ;
      RECT 7071.465 189.04 7071.745 336.495 ;
      RECT 7070.905 189.04 7071.185 336.255 ;
      RECT 7070.345 189.04 7070.625 336.015 ;
      RECT 7069.785 189.04 7070.065 335.775 ;
      RECT 7060.825 189.04 7061.105 335.29 ;
      RECT 7060.265 187.94 7060.545 335.05 ;
      RECT 7059.705 189.04 7059.985 334.81 ;
      RECT 7059.145 187.94 7059.425 334.57 ;
      RECT 7058.585 189.04 7058.865 334.33 ;
      RECT 7058.025 187.94 7058.305 334.09 ;
      RECT 7057.465 189.04 7057.745 333.85 ;
      RECT 7056.905 189.04 7057.185 333.61 ;
      RECT 7056.345 189.04 7056.625 333.37 ;
      RECT 7055.785 189.04 7056.065 333.13 ;
      RECT 7055.225 189.04 7055.505 332.89 ;
      RECT 7054.665 189.04 7054.945 332.65 ;
      RECT 7054.105 189.04 7054.385 332.41 ;
      RECT 7053.545 189.04 7053.825 332.17 ;
      RECT 7051.025 187.94 7051.305 333.89 ;
      RECT 7050.465 189.04 7050.745 333.65 ;
      RECT 7049.905 187.94 7050.185 333.41 ;
      RECT 7049.345 189.04 7049.625 333.17 ;
      RECT 7048.785 189.04 7049.065 332.93 ;
      RECT 7048.225 189.04 7048.505 332.69 ;
      RECT 7047.665 189.04 7047.945 332.45 ;
      RECT 7047.105 189.04 7047.385 332.21 ;
      RECT 7021.065 189.04 7021.345 329.86 ;
      RECT 7020.505 189.04 7020.785 330.1 ;
      RECT 7019.945 189.04 7020.225 330.34 ;
      RECT 7019.385 189.04 7019.665 330.585 ;
      RECT 7018.825 189.04 7019.105 330.825 ;
      RECT 7018.265 189.04 7018.545 331.065 ;
      RECT 7017.705 189.04 7017.985 331.065 ;
      RECT 7017.145 189.04 7017.425 330.825 ;
      RECT 7016.585 189.04 7016.865 330.585 ;
      RECT 7016.025 187.94 7016.305 330.345 ;
      RECT 7015.465 189.04 7015.745 330.105 ;
      RECT 7014.905 187.94 7015.185 329.865 ;
      RECT 7014.345 189.04 7014.625 329.625 ;
      RECT 7013.785 189.04 7014.065 329.385 ;
      RECT 7013.225 189.04 7013.505 329.145 ;
      RECT 7012.665 187.94 7012.945 328.905 ;
      RECT 7012.105 189.04 7012.385 328.665 ;
      RECT 7011.545 187.94 7011.825 328.425 ;
      RECT 7010.985 189.04 7011.265 328.185 ;
      RECT 7010.425 187.94 7010.705 327.945 ;
      RECT 7009.865 189.04 7010.145 327.705 ;
      RECT 7009.305 189.04 7009.585 327.465 ;
      RECT 7008.745 189.04 7009.025 327.225 ;
      RECT 7008.185 189.04 7008.465 326.985 ;
      RECT 6994.745 189.04 6995.025 332.785 ;
      RECT 6994.185 189.04 6994.465 332.545 ;
      RECT 6993.625 189.04 6993.905 332.305 ;
      RECT 6993.065 189.04 6993.345 332.065 ;
      RECT 6992.505 189.04 6992.785 331.825 ;
      RECT 6991.945 189.04 6992.225 331.585 ;
      RECT 6991.385 189.04 6991.665 331.345 ;
      RECT 6990.825 189.04 6991.105 331.105 ;
      RECT 6990.265 187.94 6990.545 330.865 ;
      RECT 6989.705 189.04 6989.985 330.625 ;
      RECT 6989.145 187.94 6989.425 330.305 ;
      RECT 6988.585 189.04 6988.865 330.145 ;
      RECT 6988.025 187.94 6988.305 329.905 ;
      RECT 6987.465 189.04 6987.745 329.665 ;
      RECT 6986.905 189.04 6987.185 329.425 ;
      RECT 6986.345 189.04 6986.625 329.185 ;
      RECT 6985.785 189.04 6986.065 328.945 ;
      RECT 6985.225 189.04 6985.505 328.705 ;
      RECT 6984.665 189.04 6984.945 328.465 ;
      RECT 6984.105 189.04 6984.385 328.225 ;
      RECT 6983.545 189.04 6983.825 327.985 ;
      RECT 6982.985 187.94 6983.265 327.745 ;
      RECT 6982.425 189.04 6982.705 327.505 ;
      RECT 6981.865 187.94 6982.145 327.265 ;
      RECT 6942.665 189.04 6942.945 332.875 ;
      RECT 6942.105 189.04 6942.385 333.115 ;
      RECT 6941.545 189.04 6941.825 333.355 ;
      RECT 6940.985 189.04 6941.265 333.595 ;
      RECT 6940.425 189.04 6940.705 333.835 ;
      RECT 6939.865 189.04 6940.145 334.075 ;
      RECT 6939.305 189.04 6939.585 334.315 ;
      RECT 6938.745 189.04 6939.025 334.555 ;
      RECT 6938.185 189.04 6938.465 334.795 ;
      RECT 6937.625 189.04 6937.905 335.035 ;
      RECT 6937.065 189.04 6937.345 335.275 ;
      RECT 6936.505 189.04 6936.785 335.515 ;
      RECT 6935.945 189.04 6936.225 335.755 ;
      RECT 6935.385 189.04 6935.665 335.755 ;
      RECT 6934.825 187.94 6935.105 335.515 ;
      RECT 6934.265 189.04 6934.545 335.275 ;
      RECT 6933.705 187.94 6933.985 335.035 ;
      RECT 6933.145 189.04 6933.425 334.795 ;
      RECT 6932.585 189.04 6932.865 334.555 ;
      RECT 6932.025 189.04 6932.305 334.315 ;
      RECT 6931.465 187.94 6931.745 334.05 ;
      RECT 6930.905 189.04 6931.185 333.81 ;
      RECT 6930.345 187.94 6930.625 333.57 ;
      RECT 6929.785 189.04 6930.065 333.33 ;
      RECT 6920.825 187.94 6921.105 327.165 ;
      RECT 6920.265 189.04 6920.545 327.405 ;
      RECT 6919.705 189.04 6919.985 327.645 ;
      RECT 6919.145 189.04 6919.425 327.645 ;
      RECT 6918.585 189.04 6918.865 327.405 ;
      RECT 6918.025 189.04 6918.305 327.165 ;
      RECT 6917.465 189.04 6917.745 326.925 ;
      RECT 6916.905 189.04 6917.185 326.685 ;
      RECT 6916.345 189.04 6916.625 326.445 ;
      RECT 6915.785 189.04 6916.065 326.205 ;
      RECT 6915.225 189.04 6915.505 325.965 ;
      RECT 6914.665 189.04 6914.945 325.725 ;
      RECT 6914.105 189.04 6914.385 325.485 ;
      RECT 6913.545 187.94 6913.825 325.245 ;
      RECT 6911.025 189.04 6911.305 326.965 ;
      RECT 6910.465 187.94 6910.745 326.725 ;
      RECT 6909.905 189.04 6910.185 326.485 ;
      RECT 6909.345 187.94 6909.625 326.245 ;
      RECT 6908.785 189.04 6909.065 326.005 ;
      RECT 6908.225 189.04 6908.505 325.765 ;
      RECT 6907.665 189.04 6907.945 325.525 ;
      RECT 6881.625 189.04 6881.905 328.31 ;
      RECT 6881.065 189.04 6881.345 328.55 ;
      RECT 6880.505 189.04 6880.785 328.79 ;
      RECT 6879.945 189.04 6880.225 329.03 ;
      RECT 6879.385 189.04 6879.665 329.27 ;
      RECT 6878.825 187.94 6879.105 329.51 ;
      RECT 6878.265 189.04 6878.545 329.75 ;
      RECT 6877.705 187.94 6877.985 329.99 ;
      RECT 6877.145 189.04 6877.425 330.23 ;
      RECT 6876.585 189.04 6876.865 330.47 ;
      RECT 6876.025 189.04 6876.305 330.71 ;
      RECT 6875.465 189.04 6875.745 330.95 ;
      RECT 6874.905 189.04 6875.185 331.19 ;
      RECT 6874.345 189.04 6874.625 331.43 ;
      RECT 6873.785 189.04 6874.065 331.67 ;
      RECT 6873.225 189.04 6873.505 331.67 ;
      RECT 6872.665 189.04 6872.945 331.43 ;
      RECT 6872.105 189.04 6872.385 331.19 ;
      RECT 6871.545 189.04 6871.825 330.95 ;
      RECT 6870.985 189.04 6871.265 330.705 ;
      RECT 6870.425 189.04 6870.705 330.465 ;
      RECT 6869.865 189.04 6870.145 330.225 ;
      RECT 6869.305 187.94 6869.585 329.985 ;
      RECT 6868.745 189.04 6869.025 329.745 ;
      RECT 6855.305 187.94 6855.585 327.225 ;
      RECT 6854.745 189.04 6855.025 326.985 ;
      RECT 6854.185 189.04 6854.465 326.745 ;
      RECT 6853.625 189.04 6853.905 326.505 ;
      RECT 6853.065 187.94 6853.345 326.265 ;
      RECT 6852.505 189.04 6852.785 326.025 ;
      RECT 6851.945 187.94 6852.225 325.785 ;
      RECT 6851.385 189.04 6851.665 325.545 ;
      RECT 6850.825 187.94 6851.105 325.305 ;
      RECT 6850.265 189.04 6850.545 325.065 ;
      RECT 6849.705 189.04 6849.985 324.825 ;
      RECT 6849.145 189.04 6849.425 324.585 ;
      RECT 6848.585 189.04 6848.865 324.345 ;
      RECT 6848.025 189.04 6848.305 324.105 ;
      RECT 6847.465 189.04 6847.745 323.865 ;
      RECT 6846.905 189.04 6847.185 323.625 ;
      RECT 6846.345 189.04 6846.625 323.385 ;
      RECT 6845.785 189.04 6846.065 323.145 ;
      RECT 6845.225 189.04 6845.505 322.905 ;
      RECT 6844.665 189.04 6844.945 322.665 ;
      RECT 6844.105 189.04 6844.385 322.425 ;
      RECT 6843.545 187.94 6843.825 322.185 ;
      RECT 6842.985 189.04 6843.265 321.945 ;
      RECT 6842.425 187.94 6842.705 321.705 ;
      RECT 6802.665 189.04 6802.945 332.175 ;
      RECT 6802.105 187.94 6802.385 332.415 ;
      RECT 6801.545 189.04 6801.825 332.655 ;
      RECT 6800.985 189.04 6801.265 332.895 ;
      RECT 6800.425 189.04 6800.705 333.135 ;
      RECT 6799.865 189.04 6800.145 333.375 ;
      RECT 6799.305 189.04 6799.585 333.615 ;
      RECT 6798.745 189.04 6799.025 333.86 ;
      RECT 6798.185 189.04 6798.465 334.1 ;
      RECT 6797.625 189.04 6797.905 334.34 ;
      RECT 6797.065 187.94 6797.345 334.58 ;
      RECT 6796.505 189.04 6796.785 334.82 ;
      RECT 6795.945 187.94 6796.225 335.06 ;
      RECT 6795.385 189.04 6795.665 335.3 ;
      RECT 6794.825 189.04 6795.105 335.54 ;
      RECT 6794.265 189.04 6794.545 335.78 ;
      RECT 6793.705 189.04 6793.985 336.02 ;
      RECT 6793.145 189.04 6793.425 336.26 ;
      RECT 6792.585 189.04 6792.865 336.5 ;
      RECT 6792.025 189.04 6792.305 336.74 ;
      RECT 6791.465 189.04 6791.745 336.98 ;
      RECT 6790.905 189.04 6791.185 337.22 ;
      RECT 6790.345 189.04 6790.625 337.46 ;
      RECT 6789.785 189.04 6790.065 337.7 ;
      RECT 6780.825 189.04 6781.105 333.285 ;
      RECT 6780.265 189.04 6780.545 333.045 ;
      RECT 6779.705 189.04 6779.985 332.805 ;
      RECT 6779.145 187.94 6779.425 332.565 ;
      RECT 6778.585 189.04 6778.865 332.325 ;
      RECT 6778.025 187.94 6778.305 332.085 ;
      RECT 6777.465 189.04 6777.745 331.845 ;
      RECT 6776.905 189.04 6777.185 331.605 ;
      RECT 6776.345 189.04 6776.625 331.365 ;
      RECT 6775.785 187.94 6776.065 331.125 ;
      RECT 6775.225 189.04 6775.505 330.885 ;
      RECT 6774.665 187.94 6774.945 330.645 ;
      RECT 6774.105 189.04 6774.385 330.405 ;
      RECT 6773.545 187.94 6773.825 330.165 ;
      RECT 6771.025 189.04 6771.305 322.565 ;
      RECT 6770.465 189.04 6770.745 322.325 ;
      RECT 6769.905 189.04 6770.185 322.085 ;
      RECT 6769.345 189.04 6769.625 321.845 ;
      RECT 6768.785 189.04 6769.065 321.605 ;
      RECT 6768.225 189.04 6768.505 321.365 ;
      RECT 6767.665 189.04 6767.945 321.125 ;
      RECT 6741.625 189.04 6741.905 335 ;
      RECT 6741.065 189.04 6741.345 335.24 ;
      RECT 6740.505 189.04 6740.785 335.48 ;
      RECT 6739.945 189.04 6740.225 335.72 ;
      RECT 6739.385 189.04 6739.665 335.96 ;
      RECT 6738.825 187.94 6739.105 335.96 ;
      RECT 6738.265 189.04 6738.545 335.72 ;
      RECT 6737.705 187.94 6737.985 335.475 ;
      RECT 6737.145 189.04 6737.425 335.235 ;
      RECT 6736.585 187.94 6736.865 334.995 ;
      RECT 6736.025 189.04 6736.305 334.755 ;
      RECT 6735.465 189.04 6735.745 334.515 ;
      RECT 6734.905 189.04 6735.185 334.275 ;
      RECT 6734.345 189.04 6734.625 334.035 ;
      RECT 6733.785 189.04 6734.065 333.795 ;
      RECT 6733.225 189.04 6733.505 333.555 ;
      RECT 6732.665 189.04 6732.945 333.315 ;
      RECT 6732.105 189.04 6732.385 333.075 ;
      RECT 6731.545 187.94 6731.825 332.835 ;
      RECT 6730.985 189.04 6731.265 332.595 ;
      RECT 6730.425 187.94 6730.705 332.355 ;
      RECT 6729.865 189.04 6730.145 332.115 ;
      RECT 6729.305 189.04 6729.585 331.875 ;
      RECT 6728.745 189.04 6729.025 331.635 ;
      RECT 6715.305 189.04 6715.585 335.035 ;
      RECT 6714.745 189.04 6715.025 335.275 ;
      RECT 6714.185 189.04 6714.465 335.52 ;
      RECT 6713.625 189.04 6713.905 335.76 ;
      RECT 6713.065 189.04 6713.345 336 ;
      RECT 6712.505 189.04 6712.785 336 ;
      RECT 6711.945 189.04 6712.225 335.76 ;
      RECT 6711.385 189.04 6711.665 335.52 ;
      RECT 6710.825 189.04 6711.105 328.505 ;
      RECT 6710.265 189.04 6710.545 328.265 ;
      RECT 6709.705 189.04 6709.985 328.025 ;
      RECT 6709.145 187.94 6709.425 327.785 ;
      RECT 6708.585 189.04 6708.865 327.545 ;
      RECT 6708.025 187.94 6708.305 327.305 ;
      RECT 6707.465 189.04 6707.745 327.065 ;
      RECT 6706.905 189.04 6707.185 326.825 ;
      RECT 6706.345 189.04 6706.625 326.585 ;
      RECT 6705.785 187.94 6706.065 326.345 ;
      RECT 6705.225 189.04 6705.505 326.105 ;
      RECT 6704.665 187.94 6704.945 325.865 ;
      RECT 6704.105 189.04 6704.385 325.625 ;
      RECT 6703.545 187.94 6703.825 325.385 ;
      RECT 6702.985 189.04 6703.265 325.145 ;
      RECT 6702.425 189.04 6702.705 324.905 ;
      RECT 6662.105 189.04 6662.385 333.8 ;
      RECT 6661.545 189.04 6661.825 334.04 ;
      RECT 6660.985 189.04 6661.265 334.285 ;
      RECT 6660.425 189.04 6660.705 334.525 ;
      RECT 6659.865 189.04 6660.145 334.765 ;
      RECT 6659.305 189.04 6659.585 335.005 ;
      RECT 6658.745 189.04 6659.025 335.245 ;
      RECT 6658.185 189.04 6658.465 335.485 ;
      RECT 6657.625 189.04 6657.905 335.725 ;
      RECT 6657.065 189.04 6657.345 335.965 ;
      RECT 6656.505 187.94 6656.785 336.205 ;
      RECT 6655.945 189.04 6656.225 336.445 ;
      RECT 6655.385 187.94 6655.665 336.685 ;
      RECT 6654.825 189.04 6655.105 336.925 ;
      RECT 6654.265 187.94 6654.545 337.165 ;
      RECT 6653.705 189.04 6653.985 337.165 ;
      RECT 6653.145 189.04 6653.425 336.925 ;
      RECT 6652.585 189.04 6652.865 336.685 ;
      RECT 6652.025 189.04 6652.305 336.445 ;
      RECT 6651.465 189.04 6651.745 336.205 ;
      RECT 6650.905 189.04 6651.185 335.965 ;
      RECT 6650.345 189.04 6650.625 335.725 ;
      RECT 6649.785 189.04 6650.065 335.485 ;
      RECT 6640.825 187.94 6641.105 335.515 ;
      RECT 6640.265 189.04 6640.545 335.755 ;
      RECT 6639.705 187.94 6639.985 335.995 ;
      RECT 6639.145 189.04 6639.425 336.21 ;
      RECT 6638.585 189.04 6638.865 335.785 ;
      RECT 6638.025 189.04 6638.305 335.545 ;
      RECT 6637.465 189.04 6637.745 335.305 ;
      RECT 6636.905 189.04 6637.185 335.065 ;
      RECT 6636.345 189.04 6636.625 334.825 ;
      RECT 6635.785 189.04 6636.065 334.585 ;
      RECT 6635.225 189.04 6635.505 334.345 ;
      RECT 6634.665 189.04 6634.945 334.105 ;
      RECT 6634.105 189.04 6634.385 333.865 ;
      RECT 6633.545 189.04 6633.825 333.625 ;
      RECT 6631.025 189.04 6631.305 332.8 ;
      RECT 6630.465 189.04 6630.745 332.56 ;
      RECT 6629.905 189.04 6630.185 332.32 ;
      RECT 6629.345 187.94 6629.625 332.08 ;
      RECT 6628.785 189.04 6629.065 331.84 ;
      RECT 6628.225 187.94 6628.505 331.6 ;
      RECT 6627.665 189.04 6627.945 331.36 ;
      RECT 6627.105 189.04 6627.385 331.12 ;
      RECT 6600.505 189.04 6600.785 342.165 ;
      RECT 6599.945 187.94 6600.225 342.405 ;
      RECT 6599.385 189.04 6599.665 342.645 ;
      RECT 6598.825 187.94 6599.105 342.89 ;
      RECT 6598.265 189.04 6598.545 343.13 ;
      RECT 6597.705 187.94 6597.985 343.37 ;
      RECT 6597.145 189.04 6597.425 343.61 ;
      RECT 6596.585 189.04 6596.865 343.85 ;
      RECT 6596.025 189.04 6596.305 329.47 ;
      RECT 6595.465 189.04 6595.745 329.23 ;
      RECT 6594.905 189.04 6595.185 328.99 ;
      RECT 6594.345 189.04 6594.625 328.75 ;
      RECT 6593.785 189.04 6594.065 328.51 ;
      RECT 6593.225 189.04 6593.505 328.27 ;
      RECT 6592.665 189.04 6592.945 328.03 ;
      RECT 6592.105 189.04 6592.385 327.79 ;
      RECT 6591.545 189.04 6591.825 327.55 ;
      RECT 6590.985 189.04 6591.265 327.31 ;
      RECT 6590.425 187.94 6590.705 327.07 ;
      RECT 6589.865 189.04 6590.145 326.83 ;
      RECT 6589.305 187.94 6589.585 326.59 ;
      RECT 6588.745 189.04 6589.025 326.35 ;
      RECT 6574.745 187.94 6575.025 332.47 ;
      RECT 6574.185 189.04 6574.465 332.23 ;
      RECT 6573.625 189.04 6573.905 331.99 ;
      RECT 6573.065 189.04 6573.345 331.75 ;
      RECT 6572.505 189.04 6572.785 331.51 ;
      RECT 6571.945 189.04 6572.225 331.27 ;
      RECT 6571.385 189.04 6571.665 331.03 ;
      RECT 6570.825 189.04 6571.105 330.79 ;
      RECT 6570.265 189.04 6570.545 330.55 ;
      RECT 6569.705 187.94 6569.985 330.31 ;
      RECT 6569.145 189.04 6569.425 330.07 ;
      RECT 6568.585 187.94 6568.865 329.83 ;
      RECT 6568.025 189.04 6568.305 329.59 ;
      RECT 6567.465 189.04 6567.745 329.35 ;
      RECT 6566.905 189.04 6567.185 329.11 ;
      RECT 6566.345 189.04 6566.625 328.87 ;
      RECT 6565.785 189.04 6566.065 328.63 ;
      RECT 6565.225 189.04 6565.505 328.39 ;
      RECT 6564.665 189.04 6564.945 328.15 ;
      RECT 6564.105 189.04 6564.385 327.91 ;
      RECT 6563.545 189.04 6563.825 327.67 ;
      RECT 6562.985 189.04 6563.265 327.43 ;
      RECT 6562.425 189.04 6562.705 327.19 ;
      RECT 6523.225 189.04 6523.505 334.095 ;
      RECT 6522.665 189.04 6522.945 334.335 ;
      RECT 6522.105 189.04 6522.385 334.575 ;
      RECT 6521.545 187.94 6521.825 334.815 ;
      RECT 6520.985 189.04 6521.265 335.055 ;
      RECT 6520.425 187.94 6520.705 335.295 ;
      RECT 6519.865 189.04 6520.145 335.535 ;
      RECT 6519.305 189.04 6519.585 335.775 ;
      RECT 6518.745 189.04 6519.025 336.015 ;
      RECT 6518.185 187.94 6518.465 336.255 ;
      RECT 6517.625 189.04 6517.905 336.495 ;
      RECT 6517.065 187.94 6517.345 336.735 ;
      RECT 6516.505 189.04 6516.785 336.975 ;
      RECT 6515.945 187.94 6516.225 337.215 ;
      RECT 6515.385 189.04 6515.665 337.455 ;
      RECT 6514.825 189.04 6515.105 337.695 ;
      RECT 6514.265 189.04 6514.545 337.695 ;
      RECT 6513.705 189.04 6513.985 337.455 ;
      RECT 6513.145 189.04 6513.425 337.215 ;
      RECT 6512.585 189.04 6512.865 336.975 ;
      RECT 6512.025 189.04 6512.305 336.735 ;
      RECT 6511.465 189.04 6511.745 336.495 ;
      RECT 6510.905 189.04 6511.185 336.255 ;
      RECT 6510.345 189.04 6510.625 336.015 ;
      RECT 6509.785 189.04 6510.065 335.775 ;
      RECT 6500.825 189.04 6501.105 335.29 ;
      RECT 6500.265 187.94 6500.545 335.05 ;
      RECT 6499.705 189.04 6499.985 334.81 ;
      RECT 6499.145 187.94 6499.425 334.57 ;
      RECT 6498.585 189.04 6498.865 334.33 ;
      RECT 6498.025 187.94 6498.305 334.09 ;
      RECT 6497.465 189.04 6497.745 333.85 ;
      RECT 6496.905 189.04 6497.185 333.61 ;
      RECT 6496.345 189.04 6496.625 333.37 ;
      RECT 6495.785 189.04 6496.065 333.13 ;
      RECT 6495.225 189.04 6495.505 332.89 ;
      RECT 6494.665 189.04 6494.945 332.65 ;
      RECT 6494.105 189.04 6494.385 332.41 ;
      RECT 6493.545 189.04 6493.825 332.17 ;
      RECT 6491.025 187.94 6491.305 333.89 ;
      RECT 6490.465 189.04 6490.745 333.65 ;
      RECT 6489.905 187.94 6490.185 333.41 ;
      RECT 6489.345 189.04 6489.625 333.17 ;
      RECT 6488.785 189.04 6489.065 332.93 ;
      RECT 6488.225 189.04 6488.505 332.69 ;
      RECT 6487.665 189.04 6487.945 332.45 ;
      RECT 6487.105 189.04 6487.385 332.21 ;
      RECT 6461.065 189.04 6461.345 329.86 ;
      RECT 6460.505 189.04 6460.785 330.1 ;
      RECT 6459.945 189.04 6460.225 330.34 ;
      RECT 6459.385 189.04 6459.665 330.585 ;
      RECT 6458.825 189.04 6459.105 330.825 ;
      RECT 6458.265 189.04 6458.545 331.065 ;
      RECT 6457.705 189.04 6457.985 331.065 ;
      RECT 6457.145 189.04 6457.425 330.825 ;
      RECT 6456.585 189.04 6456.865 330.585 ;
      RECT 6456.025 187.94 6456.305 330.345 ;
      RECT 6455.465 189.04 6455.745 330.105 ;
      RECT 6454.905 187.94 6455.185 329.865 ;
      RECT 6454.345 189.04 6454.625 329.625 ;
      RECT 6453.785 189.04 6454.065 329.385 ;
      RECT 6453.225 189.04 6453.505 329.145 ;
      RECT 6452.665 187.94 6452.945 328.905 ;
      RECT 6452.105 189.04 6452.385 328.665 ;
      RECT 6451.545 187.94 6451.825 328.425 ;
      RECT 6450.985 189.04 6451.265 328.185 ;
      RECT 6450.425 187.94 6450.705 327.945 ;
      RECT 6449.865 189.04 6450.145 327.705 ;
      RECT 6449.305 189.04 6449.585 327.465 ;
      RECT 6448.745 189.04 6449.025 327.225 ;
      RECT 6448.185 189.04 6448.465 326.985 ;
      RECT 6434.745 189.04 6435.025 332.785 ;
      RECT 6434.185 189.04 6434.465 332.545 ;
      RECT 6433.625 189.04 6433.905 332.305 ;
      RECT 6433.065 189.04 6433.345 332.065 ;
      RECT 6432.505 189.04 6432.785 331.825 ;
      RECT 6431.945 189.04 6432.225 331.585 ;
      RECT 6431.385 189.04 6431.665 331.345 ;
      RECT 6430.825 189.04 6431.105 331.105 ;
      RECT 6430.265 187.94 6430.545 330.865 ;
      RECT 6429.705 189.04 6429.985 330.625 ;
      RECT 6429.145 187.94 6429.425 330.305 ;
      RECT 6428.585 189.04 6428.865 330.145 ;
      RECT 6428.025 187.94 6428.305 329.905 ;
      RECT 6427.465 189.04 6427.745 329.665 ;
      RECT 6426.905 189.04 6427.185 329.425 ;
      RECT 6426.345 189.04 6426.625 329.185 ;
      RECT 6425.785 189.04 6426.065 328.945 ;
      RECT 6425.225 189.04 6425.505 328.705 ;
      RECT 6424.665 189.04 6424.945 328.465 ;
      RECT 6424.105 189.04 6424.385 328.225 ;
      RECT 6423.545 189.04 6423.825 327.985 ;
      RECT 6422.985 187.94 6423.265 327.745 ;
      RECT 6422.425 189.04 6422.705 327.505 ;
      RECT 6421.865 187.94 6422.145 327.265 ;
      RECT 6382.665 189.04 6382.945 332.875 ;
      RECT 6382.105 189.04 6382.385 333.115 ;
      RECT 6381.545 189.04 6381.825 333.355 ;
      RECT 6380.985 189.04 6381.265 333.595 ;
      RECT 6380.425 189.04 6380.705 333.835 ;
      RECT 6379.865 189.04 6380.145 334.075 ;
      RECT 6379.305 189.04 6379.585 334.315 ;
      RECT 6378.745 189.04 6379.025 334.555 ;
      RECT 6378.185 189.04 6378.465 334.795 ;
      RECT 6377.625 189.04 6377.905 335.035 ;
      RECT 6377.065 189.04 6377.345 335.275 ;
      RECT 6376.505 189.04 6376.785 335.515 ;
      RECT 6375.945 189.04 6376.225 335.755 ;
      RECT 6375.385 189.04 6375.665 335.755 ;
      RECT 6374.825 187.94 6375.105 335.515 ;
      RECT 6374.265 189.04 6374.545 335.275 ;
      RECT 6373.705 187.94 6373.985 335.035 ;
      RECT 6373.145 189.04 6373.425 334.795 ;
      RECT 6372.585 189.04 6372.865 334.555 ;
      RECT 6372.025 189.04 6372.305 334.315 ;
      RECT 6371.465 187.94 6371.745 334.05 ;
      RECT 6370.905 189.04 6371.185 333.81 ;
      RECT 6370.345 187.94 6370.625 333.57 ;
      RECT 6369.785 189.04 6370.065 333.33 ;
      RECT 6360.825 187.94 6361.105 327.165 ;
      RECT 6360.265 189.04 6360.545 327.405 ;
      RECT 6359.705 189.04 6359.985 327.645 ;
      RECT 6359.145 189.04 6359.425 327.645 ;
      RECT 6358.585 189.04 6358.865 327.405 ;
      RECT 6358.025 189.04 6358.305 327.165 ;
      RECT 6357.465 189.04 6357.745 326.925 ;
      RECT 6356.905 189.04 6357.185 326.685 ;
      RECT 6356.345 189.04 6356.625 326.445 ;
      RECT 6355.785 189.04 6356.065 326.205 ;
      RECT 6355.225 189.04 6355.505 325.965 ;
      RECT 6354.665 189.04 6354.945 325.725 ;
      RECT 6354.105 189.04 6354.385 325.485 ;
      RECT 6353.545 187.94 6353.825 325.245 ;
      RECT 6351.025 189.04 6351.305 326.965 ;
      RECT 6350.465 187.94 6350.745 326.725 ;
      RECT 6349.905 189.04 6350.185 326.485 ;
      RECT 6349.345 187.94 6349.625 326.245 ;
      RECT 6348.785 189.04 6349.065 326.005 ;
      RECT 6348.225 189.04 6348.505 325.765 ;
      RECT 6347.665 189.04 6347.945 325.525 ;
      RECT 6321.625 189.04 6321.905 328.31 ;
      RECT 6321.065 189.04 6321.345 328.55 ;
      RECT 6320.505 189.04 6320.785 328.79 ;
      RECT 6319.945 189.04 6320.225 329.03 ;
      RECT 6319.385 189.04 6319.665 329.27 ;
      RECT 6318.825 187.94 6319.105 329.51 ;
      RECT 6318.265 189.04 6318.545 329.75 ;
      RECT 6317.705 187.94 6317.985 329.99 ;
      RECT 6317.145 189.04 6317.425 330.23 ;
      RECT 6316.585 189.04 6316.865 330.47 ;
      RECT 6316.025 189.04 6316.305 330.71 ;
      RECT 6315.465 189.04 6315.745 330.95 ;
      RECT 6314.905 189.04 6315.185 331.19 ;
      RECT 6314.345 189.04 6314.625 331.43 ;
      RECT 6313.785 189.04 6314.065 331.67 ;
      RECT 6313.225 189.04 6313.505 331.67 ;
      RECT 6312.665 189.04 6312.945 331.43 ;
      RECT 6312.105 189.04 6312.385 331.19 ;
      RECT 6311.545 189.04 6311.825 330.95 ;
      RECT 6310.985 189.04 6311.265 330.705 ;
      RECT 6310.425 189.04 6310.705 330.465 ;
      RECT 6309.865 189.04 6310.145 330.225 ;
      RECT 6309.305 187.94 6309.585 329.985 ;
      RECT 6308.745 189.04 6309.025 329.745 ;
      RECT 6295.305 187.94 6295.585 327.225 ;
      RECT 6294.745 189.04 6295.025 326.985 ;
      RECT 6294.185 189.04 6294.465 326.745 ;
      RECT 6293.625 189.04 6293.905 326.505 ;
      RECT 6293.065 187.94 6293.345 326.265 ;
      RECT 6292.505 189.04 6292.785 326.025 ;
      RECT 6291.945 187.94 6292.225 325.785 ;
      RECT 6291.385 189.04 6291.665 325.545 ;
      RECT 6290.825 187.94 6291.105 325.305 ;
      RECT 6290.265 189.04 6290.545 325.065 ;
      RECT 6289.705 189.04 6289.985 324.825 ;
      RECT 6289.145 189.04 6289.425 324.585 ;
      RECT 6288.585 189.04 6288.865 324.345 ;
      RECT 6288.025 189.04 6288.305 324.105 ;
      RECT 6287.465 189.04 6287.745 323.865 ;
      RECT 6286.905 189.04 6287.185 323.625 ;
      RECT 6286.345 189.04 6286.625 323.385 ;
      RECT 6285.785 189.04 6286.065 323.145 ;
      RECT 6285.225 189.04 6285.505 322.905 ;
      RECT 6284.665 189.04 6284.945 322.665 ;
      RECT 6284.105 189.04 6284.385 322.425 ;
      RECT 6283.545 187.94 6283.825 322.185 ;
      RECT 6282.985 189.04 6283.265 321.945 ;
      RECT 6282.425 187.94 6282.705 321.705 ;
      RECT 6242.665 189.04 6242.945 332.175 ;
      RECT 6242.105 187.94 6242.385 332.415 ;
      RECT 6241.545 189.04 6241.825 332.655 ;
      RECT 6240.985 189.04 6241.265 332.895 ;
      RECT 6240.425 189.04 6240.705 333.135 ;
      RECT 6239.865 189.04 6240.145 333.375 ;
      RECT 6239.305 189.04 6239.585 333.615 ;
      RECT 6238.745 189.04 6239.025 333.86 ;
      RECT 6238.185 189.04 6238.465 334.1 ;
      RECT 6237.625 189.04 6237.905 334.34 ;
      RECT 6237.065 187.94 6237.345 334.58 ;
      RECT 6236.505 189.04 6236.785 334.82 ;
      RECT 6235.945 187.94 6236.225 335.06 ;
      RECT 6235.385 189.04 6235.665 335.3 ;
      RECT 6234.825 189.04 6235.105 335.54 ;
      RECT 6234.265 189.04 6234.545 335.78 ;
      RECT 6233.705 189.04 6233.985 336.02 ;
      RECT 6233.145 189.04 6233.425 336.26 ;
      RECT 6232.585 189.04 6232.865 336.5 ;
      RECT 6232.025 189.04 6232.305 336.74 ;
      RECT 6231.465 189.04 6231.745 336.98 ;
      RECT 6230.905 189.04 6231.185 337.22 ;
      RECT 6230.345 189.04 6230.625 337.46 ;
      RECT 6229.785 189.04 6230.065 337.7 ;
      RECT 6220.825 189.04 6221.105 333.285 ;
      RECT 6220.265 189.04 6220.545 333.045 ;
      RECT 6219.705 189.04 6219.985 332.805 ;
      RECT 6219.145 187.94 6219.425 332.565 ;
      RECT 6218.585 189.04 6218.865 332.325 ;
      RECT 6218.025 187.94 6218.305 332.085 ;
      RECT 6217.465 189.04 6217.745 331.845 ;
      RECT 6216.905 189.04 6217.185 331.605 ;
      RECT 6216.345 189.04 6216.625 331.365 ;
      RECT 6215.785 187.94 6216.065 331.125 ;
      RECT 6215.225 189.04 6215.505 330.885 ;
      RECT 6214.665 187.94 6214.945 330.645 ;
      RECT 6214.105 189.04 6214.385 330.405 ;
      RECT 6213.545 187.94 6213.825 330.165 ;
      RECT 6211.025 189.04 6211.305 322.565 ;
      RECT 6210.465 189.04 6210.745 322.325 ;
      RECT 6209.905 189.04 6210.185 322.085 ;
      RECT 6209.345 189.04 6209.625 321.845 ;
      RECT 6208.785 189.04 6209.065 321.605 ;
      RECT 6208.225 189.04 6208.505 321.365 ;
      RECT 6207.665 189.04 6207.945 321.125 ;
      RECT 6181.625 189.04 6181.905 335 ;
      RECT 6181.065 189.04 6181.345 335.24 ;
      RECT 6180.505 189.04 6180.785 335.48 ;
      RECT 6179.945 189.04 6180.225 335.72 ;
      RECT 6179.385 189.04 6179.665 335.96 ;
      RECT 6178.825 187.94 6179.105 335.96 ;
      RECT 6178.265 189.04 6178.545 335.72 ;
      RECT 6177.705 187.94 6177.985 335.475 ;
      RECT 6177.145 189.04 6177.425 335.235 ;
      RECT 6176.585 187.94 6176.865 334.995 ;
      RECT 6176.025 189.04 6176.305 334.755 ;
      RECT 6175.465 189.04 6175.745 334.515 ;
      RECT 6174.905 189.04 6175.185 334.275 ;
      RECT 6174.345 189.04 6174.625 334.035 ;
      RECT 6173.785 189.04 6174.065 333.795 ;
      RECT 6173.225 189.04 6173.505 333.555 ;
      RECT 6172.665 189.04 6172.945 333.315 ;
      RECT 6172.105 189.04 6172.385 333.075 ;
      RECT 6171.545 187.94 6171.825 332.835 ;
      RECT 6170.985 189.04 6171.265 332.595 ;
      RECT 6170.425 187.94 6170.705 332.355 ;
      RECT 6169.865 189.04 6170.145 332.115 ;
      RECT 6169.305 189.04 6169.585 331.875 ;
      RECT 6168.745 189.04 6169.025 331.635 ;
      RECT 6155.305 189.04 6155.585 335.035 ;
      RECT 6154.745 189.04 6155.025 335.275 ;
      RECT 6154.185 189.04 6154.465 335.52 ;
      RECT 6153.625 189.04 6153.905 335.76 ;
      RECT 6153.065 189.04 6153.345 336 ;
      RECT 6152.505 189.04 6152.785 336 ;
      RECT 6151.945 189.04 6152.225 335.76 ;
      RECT 6151.385 189.04 6151.665 335.52 ;
      RECT 6150.825 189.04 6151.105 328.505 ;
      RECT 6150.265 189.04 6150.545 328.265 ;
      RECT 6149.705 189.04 6149.985 328.025 ;
      RECT 6149.145 187.94 6149.425 327.785 ;
      RECT 6148.585 189.04 6148.865 327.545 ;
      RECT 6148.025 187.94 6148.305 327.305 ;
      RECT 6147.465 189.04 6147.745 327.065 ;
      RECT 6146.905 189.04 6147.185 326.825 ;
      RECT 6146.345 189.04 6146.625 326.585 ;
      RECT 6145.785 187.94 6146.065 326.345 ;
      RECT 6145.225 189.04 6145.505 326.105 ;
      RECT 6144.665 187.94 6144.945 325.865 ;
      RECT 6144.105 189.04 6144.385 325.625 ;
      RECT 6143.545 187.94 6143.825 325.385 ;
      RECT 6142.985 189.04 6143.265 325.145 ;
      RECT 6142.425 189.04 6142.705 324.905 ;
      RECT 6102.105 189.04 6102.385 333.8 ;
      RECT 6101.545 189.04 6101.825 334.04 ;
      RECT 6100.985 189.04 6101.265 334.285 ;
      RECT 6100.425 189.04 6100.705 334.525 ;
      RECT 6099.865 189.04 6100.145 334.765 ;
      RECT 6099.305 189.04 6099.585 335.005 ;
      RECT 6098.745 189.04 6099.025 335.245 ;
      RECT 6098.185 189.04 6098.465 335.485 ;
      RECT 6097.625 189.04 6097.905 335.725 ;
      RECT 6097.065 189.04 6097.345 335.965 ;
      RECT 6096.505 187.94 6096.785 336.205 ;
      RECT 6095.945 189.04 6096.225 336.445 ;
      RECT 6095.385 187.94 6095.665 336.685 ;
      RECT 6094.825 189.04 6095.105 336.925 ;
      RECT 6094.265 187.94 6094.545 337.165 ;
      RECT 6093.705 189.04 6093.985 337.165 ;
      RECT 6093.145 189.04 6093.425 336.925 ;
      RECT 6092.585 189.04 6092.865 336.685 ;
      RECT 6092.025 189.04 6092.305 336.445 ;
      RECT 6091.465 189.04 6091.745 336.205 ;
      RECT 6090.905 189.04 6091.185 335.965 ;
      RECT 6090.345 189.04 6090.625 335.725 ;
      RECT 6089.785 189.04 6090.065 335.485 ;
      RECT 6080.825 187.94 6081.105 335.515 ;
      RECT 6080.265 189.04 6080.545 335.755 ;
      RECT 6079.705 187.94 6079.985 335.995 ;
      RECT 6079.145 189.04 6079.425 336.21 ;
      RECT 6078.585 189.04 6078.865 335.785 ;
      RECT 6078.025 189.04 6078.305 335.545 ;
      RECT 6077.465 189.04 6077.745 335.305 ;
      RECT 6076.905 189.04 6077.185 335.065 ;
      RECT 6076.345 189.04 6076.625 334.825 ;
      RECT 6075.785 189.04 6076.065 334.585 ;
      RECT 6075.225 189.04 6075.505 334.345 ;
      RECT 6074.665 189.04 6074.945 334.105 ;
      RECT 6074.105 189.04 6074.385 333.865 ;
      RECT 6073.545 189.04 6073.825 333.625 ;
      RECT 6071.025 189.04 6071.305 332.8 ;
      RECT 6070.465 189.04 6070.745 332.56 ;
      RECT 6069.905 189.04 6070.185 332.32 ;
      RECT 6069.345 187.94 6069.625 332.08 ;
      RECT 6068.785 189.04 6069.065 331.84 ;
      RECT 6068.225 187.94 6068.505 331.6 ;
      RECT 6067.665 189.04 6067.945 331.36 ;
      RECT 6067.105 189.04 6067.385 331.12 ;
      RECT 6040.505 189.04 6040.785 342.165 ;
      RECT 6039.945 187.94 6040.225 342.405 ;
      RECT 6039.385 189.04 6039.665 342.645 ;
      RECT 6038.825 187.94 6039.105 342.89 ;
      RECT 6038.265 189.04 6038.545 343.13 ;
      RECT 6037.705 187.94 6037.985 343.37 ;
      RECT 6037.145 189.04 6037.425 343.61 ;
      RECT 6036.585 189.04 6036.865 343.85 ;
      RECT 6036.025 189.04 6036.305 329.47 ;
      RECT 6035.465 189.04 6035.745 329.23 ;
      RECT 6034.905 189.04 6035.185 328.99 ;
      RECT 6034.345 189.04 6034.625 328.75 ;
      RECT 6033.785 189.04 6034.065 328.51 ;
      RECT 6033.225 189.04 6033.505 328.27 ;
      RECT 6032.665 189.04 6032.945 328.03 ;
      RECT 6032.105 189.04 6032.385 327.79 ;
      RECT 6031.545 189.04 6031.825 327.55 ;
      RECT 6030.985 189.04 6031.265 327.31 ;
      RECT 6030.425 187.94 6030.705 327.07 ;
      RECT 6029.865 189.04 6030.145 326.83 ;
      RECT 6029.305 187.94 6029.585 326.59 ;
      RECT 6028.745 189.04 6029.025 326.35 ;
      RECT 6014.745 187.94 6015.025 332.47 ;
      RECT 6014.185 189.04 6014.465 332.23 ;
      RECT 6013.625 189.04 6013.905 331.99 ;
      RECT 6013.065 189.04 6013.345 331.75 ;
      RECT 6012.505 189.04 6012.785 331.51 ;
      RECT 6011.945 189.04 6012.225 331.27 ;
      RECT 6011.385 189.04 6011.665 331.03 ;
      RECT 6010.825 189.04 6011.105 330.79 ;
      RECT 6010.265 189.04 6010.545 330.55 ;
      RECT 6009.705 187.94 6009.985 330.31 ;
      RECT 6009.145 189.04 6009.425 330.07 ;
      RECT 6008.585 187.94 6008.865 329.83 ;
      RECT 6008.025 189.04 6008.305 329.59 ;
      RECT 6007.465 189.04 6007.745 329.35 ;
      RECT 6006.905 189.04 6007.185 329.11 ;
      RECT 6006.345 189.04 6006.625 328.87 ;
      RECT 6005.785 189.04 6006.065 328.63 ;
      RECT 6005.225 189.04 6005.505 328.39 ;
      RECT 6004.665 189.04 6004.945 328.15 ;
      RECT 6004.105 189.04 6004.385 327.91 ;
      RECT 6003.545 189.04 6003.825 327.67 ;
      RECT 6002.985 189.04 6003.265 327.43 ;
      RECT 6002.425 189.04 6002.705 327.19 ;
      RECT 5963.225 189.04 5963.505 334.095 ;
      RECT 5962.665 189.04 5962.945 334.335 ;
      RECT 5962.105 189.04 5962.385 334.575 ;
      RECT 5961.545 187.94 5961.825 334.815 ;
      RECT 5960.985 189.04 5961.265 335.055 ;
      RECT 5960.425 187.94 5960.705 335.295 ;
      RECT 5959.865 189.04 5960.145 335.535 ;
      RECT 5959.305 189.04 5959.585 335.775 ;
      RECT 5958.745 189.04 5959.025 336.015 ;
      RECT 5958.185 187.94 5958.465 336.255 ;
      RECT 5957.625 189.04 5957.905 336.495 ;
      RECT 5957.065 187.94 5957.345 336.735 ;
      RECT 5956.505 189.04 5956.785 336.975 ;
      RECT 5955.945 187.94 5956.225 337.215 ;
      RECT 5955.385 189.04 5955.665 337.455 ;
      RECT 5954.825 189.04 5955.105 337.695 ;
      RECT 5954.265 189.04 5954.545 337.695 ;
      RECT 5953.705 189.04 5953.985 337.455 ;
      RECT 5953.145 189.04 5953.425 337.215 ;
      RECT 5952.585 189.04 5952.865 336.975 ;
      RECT 5952.025 189.04 5952.305 336.735 ;
      RECT 5951.465 189.04 5951.745 336.495 ;
      RECT 5950.905 189.04 5951.185 336.255 ;
      RECT 5950.345 189.04 5950.625 336.015 ;
      RECT 5949.785 189.04 5950.065 335.775 ;
      RECT 5940.825 189.04 5941.105 335.29 ;
      RECT 5940.265 187.94 5940.545 335.05 ;
      RECT 5939.705 189.04 5939.985 334.81 ;
      RECT 5939.145 187.94 5939.425 334.57 ;
      RECT 5938.585 189.04 5938.865 334.33 ;
      RECT 5938.025 187.94 5938.305 334.09 ;
      RECT 5937.465 189.04 5937.745 333.85 ;
      RECT 5936.905 189.04 5937.185 333.61 ;
      RECT 5936.345 189.04 5936.625 333.37 ;
      RECT 5935.785 189.04 5936.065 333.13 ;
      RECT 5935.225 189.04 5935.505 332.89 ;
      RECT 5934.665 189.04 5934.945 332.65 ;
      RECT 5934.105 189.04 5934.385 332.41 ;
      RECT 5933.545 189.04 5933.825 332.17 ;
      RECT 5931.025 187.94 5931.305 333.89 ;
      RECT 5930.465 189.04 5930.745 333.65 ;
      RECT 5929.905 187.94 5930.185 333.41 ;
      RECT 5929.345 189.04 5929.625 333.17 ;
      RECT 5928.785 189.04 5929.065 332.93 ;
      RECT 5928.225 189.04 5928.505 332.69 ;
      RECT 5927.665 189.04 5927.945 332.45 ;
      RECT 5927.105 189.04 5927.385 332.21 ;
      RECT 5901.065 189.04 5901.345 329.86 ;
      RECT 5900.505 189.04 5900.785 330.1 ;
      RECT 5899.945 189.04 5900.225 330.34 ;
      RECT 5899.385 189.04 5899.665 330.585 ;
      RECT 5898.825 189.04 5899.105 330.825 ;
      RECT 5898.265 189.04 5898.545 331.065 ;
      RECT 5897.705 189.04 5897.985 331.065 ;
      RECT 5897.145 189.04 5897.425 330.825 ;
      RECT 5896.585 189.04 5896.865 330.585 ;
      RECT 5896.025 187.94 5896.305 330.345 ;
      RECT 5895.465 189.04 5895.745 330.105 ;
      RECT 5894.905 187.94 5895.185 329.865 ;
      RECT 5894.345 189.04 5894.625 329.625 ;
      RECT 5893.785 189.04 5894.065 329.385 ;
      RECT 5893.225 189.04 5893.505 329.145 ;
      RECT 5892.665 187.94 5892.945 328.905 ;
      RECT 5892.105 189.04 5892.385 328.665 ;
      RECT 5891.545 187.94 5891.825 328.425 ;
      RECT 5890.985 189.04 5891.265 328.185 ;
      RECT 5890.425 187.94 5890.705 327.945 ;
      RECT 5889.865 189.04 5890.145 327.705 ;
      RECT 5889.305 189.04 5889.585 327.465 ;
      RECT 5888.745 189.04 5889.025 327.225 ;
      RECT 5888.185 189.04 5888.465 326.985 ;
      RECT 5874.745 189.04 5875.025 332.785 ;
      RECT 5874.185 189.04 5874.465 332.545 ;
      RECT 5873.625 189.04 5873.905 332.305 ;
      RECT 5873.065 189.04 5873.345 332.065 ;
      RECT 5872.505 189.04 5872.785 331.825 ;
      RECT 5871.945 189.04 5872.225 331.585 ;
      RECT 5871.385 189.04 5871.665 331.345 ;
      RECT 5870.825 189.04 5871.105 331.105 ;
      RECT 5870.265 187.94 5870.545 330.865 ;
      RECT 5869.705 189.04 5869.985 330.625 ;
      RECT 5869.145 187.94 5869.425 330.305 ;
      RECT 5868.585 189.04 5868.865 330.145 ;
      RECT 5868.025 187.94 5868.305 329.905 ;
      RECT 5867.465 189.04 5867.745 329.665 ;
      RECT 5866.905 189.04 5867.185 329.425 ;
      RECT 5866.345 189.04 5866.625 329.185 ;
      RECT 5865.785 189.04 5866.065 328.945 ;
      RECT 5865.225 189.04 5865.505 328.705 ;
      RECT 5864.665 189.04 5864.945 328.465 ;
      RECT 5864.105 189.04 5864.385 328.225 ;
      RECT 5863.545 189.04 5863.825 327.985 ;
      RECT 5862.985 187.94 5863.265 327.745 ;
      RECT 5862.425 189.04 5862.705 327.505 ;
      RECT 5861.865 187.94 5862.145 327.265 ;
      RECT 5822.665 189.04 5822.945 332.875 ;
      RECT 5822.105 189.04 5822.385 333.115 ;
      RECT 5821.545 189.04 5821.825 333.355 ;
      RECT 5820.985 189.04 5821.265 333.595 ;
      RECT 5820.425 189.04 5820.705 333.835 ;
      RECT 5819.865 189.04 5820.145 334.075 ;
      RECT 5819.305 189.04 5819.585 334.315 ;
      RECT 5818.745 189.04 5819.025 334.555 ;
      RECT 5818.185 189.04 5818.465 334.795 ;
      RECT 5817.625 189.04 5817.905 335.035 ;
      RECT 5817.065 189.04 5817.345 335.275 ;
      RECT 5816.505 189.04 5816.785 335.515 ;
      RECT 5815.945 189.04 5816.225 335.755 ;
      RECT 5815.385 189.04 5815.665 335.755 ;
      RECT 5814.825 187.94 5815.105 335.515 ;
      RECT 5814.265 189.04 5814.545 335.275 ;
      RECT 5813.705 187.94 5813.985 335.035 ;
      RECT 5813.145 189.04 5813.425 334.795 ;
      RECT 5812.585 189.04 5812.865 334.555 ;
      RECT 5812.025 189.04 5812.305 334.315 ;
      RECT 5811.465 187.94 5811.745 334.05 ;
      RECT 5810.905 189.04 5811.185 333.81 ;
      RECT 5810.345 187.94 5810.625 333.57 ;
      RECT 5809.785 189.04 5810.065 333.33 ;
      RECT 5800.825 187.94 5801.105 327.165 ;
      RECT 5800.265 189.04 5800.545 327.405 ;
      RECT 5799.705 189.04 5799.985 327.645 ;
      RECT 5799.145 189.04 5799.425 327.645 ;
      RECT 5798.585 189.04 5798.865 327.405 ;
      RECT 5798.025 189.04 5798.305 327.165 ;
      RECT 5797.465 189.04 5797.745 326.925 ;
      RECT 5796.905 189.04 5797.185 326.685 ;
      RECT 5796.345 189.04 5796.625 326.445 ;
      RECT 5795.785 189.04 5796.065 326.205 ;
      RECT 5795.225 189.04 5795.505 325.965 ;
      RECT 5794.665 189.04 5794.945 325.725 ;
      RECT 5794.105 189.04 5794.385 325.485 ;
      RECT 5793.545 187.94 5793.825 325.245 ;
      RECT 5791.025 189.04 5791.305 326.965 ;
      RECT 5790.465 187.94 5790.745 326.725 ;
      RECT 5789.905 189.04 5790.185 326.485 ;
      RECT 5789.345 187.94 5789.625 326.245 ;
      RECT 5788.785 189.04 5789.065 326.005 ;
      RECT 5788.225 189.04 5788.505 325.765 ;
      RECT 5787.665 189.04 5787.945 325.525 ;
      RECT 5761.625 189.04 5761.905 328.31 ;
      RECT 5761.065 189.04 5761.345 328.55 ;
      RECT 5760.505 189.04 5760.785 328.79 ;
      RECT 5759.945 189.04 5760.225 329.03 ;
      RECT 5759.385 189.04 5759.665 329.27 ;
      RECT 5758.825 187.94 5759.105 329.51 ;
      RECT 5758.265 189.04 5758.545 329.75 ;
      RECT 5757.705 187.94 5757.985 329.99 ;
      RECT 5757.145 189.04 5757.425 330.23 ;
      RECT 5756.585 189.04 5756.865 330.47 ;
      RECT 5756.025 189.04 5756.305 330.71 ;
      RECT 5755.465 189.04 5755.745 330.95 ;
      RECT 5754.905 189.04 5755.185 331.19 ;
      RECT 5754.345 189.04 5754.625 331.43 ;
      RECT 5753.785 189.04 5754.065 331.67 ;
      RECT 5753.225 189.04 5753.505 331.67 ;
      RECT 5752.665 189.04 5752.945 331.43 ;
      RECT 5752.105 189.04 5752.385 331.19 ;
      RECT 5751.545 189.04 5751.825 330.95 ;
      RECT 5750.985 189.04 5751.265 330.705 ;
      RECT 5750.425 189.04 5750.705 330.465 ;
      RECT 5749.865 189.04 5750.145 330.225 ;
      RECT 5749.305 187.94 5749.585 329.985 ;
      RECT 5748.745 189.04 5749.025 329.745 ;
      RECT 5735.305 187.94 5735.585 327.225 ;
      RECT 5734.745 189.04 5735.025 326.985 ;
      RECT 5734.185 189.04 5734.465 326.745 ;
      RECT 5733.625 189.04 5733.905 326.505 ;
      RECT 5733.065 187.94 5733.345 326.265 ;
      RECT 5732.505 189.04 5732.785 326.025 ;
      RECT 5731.945 187.94 5732.225 325.785 ;
      RECT 5731.385 189.04 5731.665 325.545 ;
      RECT 5730.825 187.94 5731.105 325.305 ;
      RECT 5730.265 189.04 5730.545 325.065 ;
      RECT 5729.705 189.04 5729.985 324.825 ;
      RECT 5729.145 189.04 5729.425 324.585 ;
      RECT 5728.585 189.04 5728.865 324.345 ;
      RECT 5728.025 189.04 5728.305 324.105 ;
      RECT 5727.465 189.04 5727.745 323.865 ;
      RECT 5726.905 189.04 5727.185 323.625 ;
      RECT 5726.345 189.04 5726.625 323.385 ;
      RECT 5725.785 189.04 5726.065 323.145 ;
      RECT 5725.225 189.04 5725.505 322.905 ;
      RECT 5724.665 189.04 5724.945 322.665 ;
      RECT 5724.105 189.04 5724.385 322.425 ;
      RECT 5723.545 187.94 5723.825 322.185 ;
      RECT 5722.985 189.04 5723.265 321.945 ;
      RECT 5722.425 187.94 5722.705 321.705 ;
      RECT 5682.665 189.04 5682.945 332.175 ;
      RECT 5682.105 187.94 5682.385 332.415 ;
      RECT 5681.545 189.04 5681.825 332.655 ;
      RECT 5680.985 189.04 5681.265 332.895 ;
      RECT 5680.425 189.04 5680.705 333.135 ;
      RECT 5679.865 189.04 5680.145 333.375 ;
      RECT 5679.305 189.04 5679.585 333.615 ;
      RECT 5678.745 189.04 5679.025 333.86 ;
      RECT 5678.185 189.04 5678.465 334.1 ;
      RECT 5677.625 189.04 5677.905 334.34 ;
      RECT 5677.065 187.94 5677.345 334.58 ;
      RECT 5676.505 189.04 5676.785 334.82 ;
      RECT 5675.945 187.94 5676.225 335.06 ;
      RECT 5675.385 189.04 5675.665 335.3 ;
      RECT 5674.825 189.04 5675.105 335.54 ;
      RECT 5674.265 189.04 5674.545 335.78 ;
      RECT 5673.705 189.04 5673.985 336.02 ;
      RECT 5673.145 189.04 5673.425 336.26 ;
      RECT 5672.585 189.04 5672.865 336.5 ;
      RECT 5672.025 189.04 5672.305 336.74 ;
      RECT 5671.465 189.04 5671.745 336.98 ;
      RECT 5670.905 189.04 5671.185 337.22 ;
      RECT 5670.345 189.04 5670.625 337.46 ;
      RECT 5669.785 189.04 5670.065 337.7 ;
      RECT 5660.825 189.04 5661.105 333.285 ;
      RECT 5660.265 189.04 5660.545 333.045 ;
      RECT 5659.705 189.04 5659.985 332.805 ;
      RECT 5659.145 187.94 5659.425 332.565 ;
      RECT 5658.585 189.04 5658.865 332.325 ;
      RECT 5658.025 187.94 5658.305 332.085 ;
      RECT 5657.465 189.04 5657.745 331.845 ;
      RECT 5656.905 189.04 5657.185 331.605 ;
      RECT 5656.345 189.04 5656.625 331.365 ;
      RECT 5655.785 187.94 5656.065 331.125 ;
      RECT 5655.225 189.04 5655.505 330.885 ;
      RECT 5654.665 187.94 5654.945 330.645 ;
      RECT 5654.105 189.04 5654.385 330.405 ;
      RECT 5653.545 187.94 5653.825 330.165 ;
      RECT 5651.025 189.04 5651.305 322.565 ;
      RECT 5650.465 189.04 5650.745 322.325 ;
      RECT 5649.905 189.04 5650.185 322.085 ;
      RECT 5649.345 189.04 5649.625 321.845 ;
      RECT 5648.785 189.04 5649.065 321.605 ;
      RECT 5648.225 189.04 5648.505 321.365 ;
      RECT 5647.665 189.04 5647.945 321.125 ;
      RECT 5621.625 189.04 5621.905 335 ;
      RECT 5621.065 189.04 5621.345 335.24 ;
      RECT 5620.505 189.04 5620.785 335.48 ;
      RECT 5619.945 189.04 5620.225 335.72 ;
      RECT 5619.385 189.04 5619.665 335.96 ;
      RECT 5618.825 187.94 5619.105 335.96 ;
      RECT 5618.265 189.04 5618.545 335.72 ;
      RECT 5617.705 187.94 5617.985 335.475 ;
      RECT 5617.145 189.04 5617.425 335.235 ;
      RECT 5616.585 187.94 5616.865 334.995 ;
      RECT 5616.025 189.04 5616.305 334.755 ;
      RECT 5615.465 189.04 5615.745 334.515 ;
      RECT 5614.905 189.04 5615.185 334.275 ;
      RECT 5614.345 189.04 5614.625 334.035 ;
      RECT 5613.785 189.04 5614.065 333.795 ;
      RECT 5613.225 189.04 5613.505 333.555 ;
      RECT 5612.665 189.04 5612.945 333.315 ;
      RECT 5612.105 189.04 5612.385 333.075 ;
      RECT 5611.545 187.94 5611.825 332.835 ;
      RECT 5610.985 189.04 5611.265 332.595 ;
      RECT 5610.425 187.94 5610.705 332.355 ;
      RECT 5609.865 189.04 5610.145 332.115 ;
      RECT 5609.305 189.04 5609.585 331.875 ;
      RECT 5608.745 189.04 5609.025 331.635 ;
      RECT 5595.305 189.04 5595.585 335.035 ;
      RECT 5594.745 189.04 5595.025 335.275 ;
      RECT 5594.185 189.04 5594.465 335.52 ;
      RECT 5593.625 189.04 5593.905 335.76 ;
      RECT 5593.065 189.04 5593.345 336 ;
      RECT 5592.505 189.04 5592.785 336 ;
      RECT 5591.945 189.04 5592.225 335.76 ;
      RECT 5591.385 189.04 5591.665 335.52 ;
      RECT 5590.825 189.04 5591.105 328.505 ;
      RECT 5590.265 189.04 5590.545 328.265 ;
      RECT 5589.705 189.04 5589.985 328.025 ;
      RECT 5589.145 187.94 5589.425 327.785 ;
      RECT 5588.585 189.04 5588.865 327.545 ;
      RECT 5588.025 187.94 5588.305 327.305 ;
      RECT 5587.465 189.04 5587.745 327.065 ;
      RECT 5586.905 189.04 5587.185 326.825 ;
      RECT 5586.345 189.04 5586.625 326.585 ;
      RECT 5585.785 187.94 5586.065 326.345 ;
      RECT 5585.225 189.04 5585.505 326.105 ;
      RECT 5584.665 187.94 5584.945 325.865 ;
      RECT 5584.105 189.04 5584.385 325.625 ;
      RECT 5583.545 187.94 5583.825 325.385 ;
      RECT 5582.985 189.04 5583.265 325.145 ;
      RECT 5582.425 189.04 5582.705 324.905 ;
      RECT 5542.105 189.04 5542.385 333.8 ;
      RECT 5541.545 189.04 5541.825 334.04 ;
      RECT 5540.985 189.04 5541.265 334.285 ;
      RECT 5540.425 189.04 5540.705 334.525 ;
      RECT 5539.865 189.04 5540.145 334.765 ;
      RECT 5539.305 189.04 5539.585 335.005 ;
      RECT 5538.745 189.04 5539.025 335.245 ;
      RECT 5538.185 189.04 5538.465 335.485 ;
      RECT 5537.625 189.04 5537.905 335.725 ;
      RECT 5537.065 189.04 5537.345 335.965 ;
      RECT 5536.505 187.94 5536.785 336.205 ;
      RECT 5535.945 189.04 5536.225 336.445 ;
      RECT 5535.385 187.94 5535.665 336.685 ;
      RECT 5534.825 189.04 5535.105 336.925 ;
      RECT 5534.265 187.94 5534.545 337.165 ;
      RECT 5533.705 189.04 5533.985 337.165 ;
      RECT 5533.145 189.04 5533.425 336.925 ;
      RECT 5532.585 189.04 5532.865 336.685 ;
      RECT 5532.025 189.04 5532.305 336.445 ;
      RECT 5531.465 189.04 5531.745 336.205 ;
      RECT 5530.905 189.04 5531.185 335.965 ;
      RECT 5530.345 189.04 5530.625 335.725 ;
      RECT 5529.785 189.04 5530.065 335.485 ;
      RECT 5520.825 187.94 5521.105 335.515 ;
      RECT 5520.265 189.04 5520.545 335.755 ;
      RECT 5519.705 187.94 5519.985 335.995 ;
      RECT 5519.145 189.04 5519.425 336.21 ;
      RECT 5518.585 189.04 5518.865 335.785 ;
      RECT 5518.025 189.04 5518.305 335.545 ;
      RECT 5517.465 189.04 5517.745 335.305 ;
      RECT 5516.905 189.04 5517.185 335.065 ;
      RECT 5516.345 189.04 5516.625 334.825 ;
      RECT 5515.785 189.04 5516.065 334.585 ;
      RECT 5515.225 189.04 5515.505 334.345 ;
      RECT 5514.665 189.04 5514.945 334.105 ;
      RECT 5514.105 189.04 5514.385 333.865 ;
      RECT 5513.545 189.04 5513.825 333.625 ;
      RECT 5511.025 189.04 5511.305 332.8 ;
      RECT 5510.465 189.04 5510.745 332.56 ;
      RECT 5509.905 189.04 5510.185 332.32 ;
      RECT 5509.345 187.94 5509.625 332.08 ;
      RECT 5508.785 189.04 5509.065 331.84 ;
      RECT 5508.225 187.94 5508.505 331.6 ;
      RECT 5507.665 189.04 5507.945 331.36 ;
      RECT 5507.105 189.04 5507.385 331.12 ;
      RECT 5480.505 189.04 5480.785 342.165 ;
      RECT 5479.945 187.94 5480.225 342.405 ;
      RECT 5479.385 189.04 5479.665 342.645 ;
      RECT 5478.825 187.94 5479.105 342.89 ;
      RECT 5478.265 189.04 5478.545 343.13 ;
      RECT 5477.705 187.94 5477.985 343.37 ;
      RECT 5477.145 189.04 5477.425 343.61 ;
      RECT 5476.585 189.04 5476.865 343.85 ;
      RECT 5476.025 189.04 5476.305 329.47 ;
      RECT 5475.465 189.04 5475.745 329.23 ;
      RECT 5474.905 189.04 5475.185 328.99 ;
      RECT 5474.345 189.04 5474.625 328.75 ;
      RECT 5473.785 189.04 5474.065 328.51 ;
      RECT 5473.225 189.04 5473.505 328.27 ;
      RECT 5472.665 189.04 5472.945 328.03 ;
      RECT 5472.105 189.04 5472.385 327.79 ;
      RECT 5471.545 189.04 5471.825 327.55 ;
      RECT 5470.985 189.04 5471.265 327.31 ;
      RECT 5470.425 187.94 5470.705 327.07 ;
      RECT 5469.865 189.04 5470.145 326.83 ;
      RECT 5469.305 187.94 5469.585 326.59 ;
      RECT 5468.745 189.04 5469.025 326.35 ;
      RECT 5454.745 187.94 5455.025 332.47 ;
      RECT 5454.185 189.04 5454.465 332.23 ;
      RECT 5453.625 189.04 5453.905 331.99 ;
      RECT 5453.065 189.04 5453.345 331.75 ;
      RECT 5452.505 189.04 5452.785 331.51 ;
      RECT 5451.945 189.04 5452.225 331.27 ;
      RECT 5451.385 189.04 5451.665 331.03 ;
      RECT 5450.825 189.04 5451.105 330.79 ;
      RECT 5450.265 189.04 5450.545 330.55 ;
      RECT 5449.705 187.94 5449.985 330.31 ;
      RECT 5449.145 189.04 5449.425 330.07 ;
      RECT 5448.585 187.94 5448.865 329.83 ;
      RECT 5448.025 189.04 5448.305 329.59 ;
      RECT 5447.465 189.04 5447.745 329.35 ;
      RECT 5446.905 189.04 5447.185 329.11 ;
      RECT 5446.345 189.04 5446.625 328.87 ;
      RECT 5445.785 189.04 5446.065 328.63 ;
      RECT 5445.225 189.04 5445.505 328.39 ;
      RECT 5444.665 189.04 5444.945 328.15 ;
      RECT 5444.105 189.04 5444.385 327.91 ;
      RECT 5443.545 189.04 5443.825 327.67 ;
      RECT 5442.985 189.04 5443.265 327.43 ;
      RECT 5442.425 189.04 5442.705 327.19 ;
      RECT 5403.225 189.04 5403.505 334.095 ;
      RECT 5402.665 189.04 5402.945 334.335 ;
      RECT 5402.105 189.04 5402.385 334.575 ;
      RECT 5401.545 187.94 5401.825 334.815 ;
      RECT 5400.985 189.04 5401.265 335.055 ;
      RECT 5400.425 187.94 5400.705 335.295 ;
      RECT 5399.865 189.04 5400.145 335.535 ;
      RECT 5399.305 189.04 5399.585 335.775 ;
      RECT 5398.745 189.04 5399.025 336.015 ;
      RECT 5398.185 187.94 5398.465 336.255 ;
      RECT 5397.625 189.04 5397.905 336.495 ;
      RECT 5397.065 187.94 5397.345 336.735 ;
      RECT 5396.505 189.04 5396.785 336.975 ;
      RECT 5395.945 187.94 5396.225 337.215 ;
      RECT 5395.385 189.04 5395.665 337.455 ;
      RECT 5394.825 189.04 5395.105 337.695 ;
      RECT 5394.265 189.04 5394.545 337.695 ;
      RECT 5393.705 189.04 5393.985 337.455 ;
      RECT 5393.145 189.04 5393.425 337.215 ;
      RECT 5392.585 189.04 5392.865 336.975 ;
      RECT 5392.025 189.04 5392.305 336.735 ;
      RECT 5391.465 189.04 5391.745 336.495 ;
      RECT 5390.905 189.04 5391.185 336.255 ;
      RECT 5390.345 189.04 5390.625 336.015 ;
      RECT 5389.785 189.04 5390.065 335.775 ;
      RECT 5380.825 189.04 5381.105 335.29 ;
      RECT 5380.265 187.94 5380.545 335.05 ;
      RECT 5379.705 189.04 5379.985 334.81 ;
      RECT 5379.145 187.94 5379.425 334.57 ;
      RECT 5378.585 189.04 5378.865 334.33 ;
      RECT 5378.025 187.94 5378.305 334.09 ;
      RECT 5377.465 189.04 5377.745 333.85 ;
      RECT 5376.905 189.04 5377.185 333.61 ;
      RECT 5376.345 189.04 5376.625 333.37 ;
      RECT 5375.785 189.04 5376.065 333.13 ;
      RECT 5375.225 189.04 5375.505 332.89 ;
      RECT 5374.665 189.04 5374.945 332.65 ;
      RECT 5374.105 189.04 5374.385 332.41 ;
      RECT 5373.545 189.04 5373.825 332.17 ;
      RECT 5371.025 187.94 5371.305 333.89 ;
      RECT 5370.465 189.04 5370.745 333.65 ;
      RECT 5369.905 187.94 5370.185 333.41 ;
      RECT 5369.345 189.04 5369.625 333.17 ;
      RECT 5368.785 189.04 5369.065 332.93 ;
      RECT 5368.225 189.04 5368.505 332.69 ;
      RECT 5367.665 189.04 5367.945 332.45 ;
      RECT 5367.105 189.04 5367.385 332.21 ;
      RECT 5341.065 189.04 5341.345 329.86 ;
      RECT 5340.505 189.04 5340.785 330.1 ;
      RECT 5339.945 189.04 5340.225 330.34 ;
      RECT 5339.385 189.04 5339.665 330.585 ;
      RECT 5338.825 189.04 5339.105 330.825 ;
      RECT 5338.265 189.04 5338.545 331.065 ;
      RECT 5337.705 189.04 5337.985 331.065 ;
      RECT 5337.145 189.04 5337.425 330.825 ;
      RECT 5336.585 189.04 5336.865 330.585 ;
      RECT 5336.025 187.94 5336.305 330.345 ;
      RECT 5335.465 189.04 5335.745 330.105 ;
      RECT 5334.905 187.94 5335.185 329.865 ;
      RECT 5334.345 189.04 5334.625 329.625 ;
      RECT 5333.785 189.04 5334.065 329.385 ;
      RECT 5333.225 189.04 5333.505 329.145 ;
      RECT 5332.665 187.94 5332.945 328.905 ;
      RECT 5332.105 189.04 5332.385 328.665 ;
      RECT 5331.545 187.94 5331.825 328.425 ;
      RECT 5330.985 189.04 5331.265 328.185 ;
      RECT 5330.425 187.94 5330.705 327.945 ;
      RECT 5329.865 189.04 5330.145 327.705 ;
      RECT 5329.305 189.04 5329.585 327.465 ;
      RECT 5328.745 189.04 5329.025 327.225 ;
      RECT 5328.185 189.04 5328.465 326.985 ;
      RECT 5314.745 189.04 5315.025 332.785 ;
      RECT 5314.185 189.04 5314.465 332.545 ;
      RECT 5313.625 189.04 5313.905 332.305 ;
      RECT 5313.065 189.04 5313.345 332.065 ;
      RECT 5312.505 189.04 5312.785 331.825 ;
      RECT 5311.945 189.04 5312.225 331.585 ;
      RECT 5311.385 189.04 5311.665 331.345 ;
      RECT 5310.825 189.04 5311.105 331.105 ;
      RECT 5310.265 187.94 5310.545 330.865 ;
      RECT 5309.705 189.04 5309.985 330.625 ;
      RECT 5309.145 187.94 5309.425 330.305 ;
      RECT 5308.585 189.04 5308.865 330.145 ;
      RECT 5308.025 187.94 5308.305 329.905 ;
      RECT 5307.465 189.04 5307.745 329.665 ;
      RECT 5306.905 189.04 5307.185 329.425 ;
      RECT 5306.345 189.04 5306.625 329.185 ;
      RECT 5305.785 189.04 5306.065 328.945 ;
      RECT 5305.225 189.04 5305.505 328.705 ;
      RECT 5304.665 189.04 5304.945 328.465 ;
      RECT 5304.105 189.04 5304.385 328.225 ;
      RECT 5303.545 189.04 5303.825 327.985 ;
      RECT 5302.985 187.94 5303.265 327.745 ;
      RECT 5302.425 189.04 5302.705 327.505 ;
      RECT 5301.865 187.94 5302.145 327.265 ;
      RECT 5262.665 189.04 5262.945 332.875 ;
      RECT 5262.105 189.04 5262.385 333.115 ;
      RECT 5261.545 189.04 5261.825 333.355 ;
      RECT 5260.985 189.04 5261.265 333.595 ;
      RECT 5260.425 189.04 5260.705 333.835 ;
      RECT 5259.865 189.04 5260.145 334.075 ;
      RECT 5259.305 189.04 5259.585 334.315 ;
      RECT 5258.745 189.04 5259.025 334.555 ;
      RECT 5258.185 189.04 5258.465 334.795 ;
      RECT 5257.625 189.04 5257.905 335.035 ;
      RECT 5257.065 189.04 5257.345 335.275 ;
      RECT 5256.505 189.04 5256.785 335.515 ;
      RECT 5255.945 189.04 5256.225 335.755 ;
      RECT 5255.385 189.04 5255.665 335.755 ;
      RECT 5254.825 187.94 5255.105 335.515 ;
      RECT 5254.265 189.04 5254.545 335.275 ;
      RECT 5253.705 187.94 5253.985 335.035 ;
      RECT 5253.145 189.04 5253.425 334.795 ;
      RECT 5252.585 189.04 5252.865 334.555 ;
      RECT 5252.025 189.04 5252.305 334.315 ;
      RECT 5251.465 187.94 5251.745 334.05 ;
      RECT 5250.905 189.04 5251.185 333.81 ;
      RECT 5250.345 187.94 5250.625 333.57 ;
      RECT 5249.785 189.04 5250.065 333.33 ;
      RECT 5240.825 187.94 5241.105 327.165 ;
      RECT 5240.265 189.04 5240.545 327.405 ;
      RECT 5239.705 189.04 5239.985 327.645 ;
      RECT 5239.145 189.04 5239.425 327.645 ;
      RECT 5238.585 189.04 5238.865 327.405 ;
      RECT 5238.025 189.04 5238.305 327.165 ;
      RECT 5237.465 189.04 5237.745 326.925 ;
      RECT 5236.905 189.04 5237.185 326.685 ;
      RECT 5236.345 189.04 5236.625 326.445 ;
      RECT 5235.785 189.04 5236.065 326.205 ;
      RECT 5235.225 189.04 5235.505 325.965 ;
      RECT 5234.665 189.04 5234.945 325.725 ;
      RECT 5234.105 189.04 5234.385 325.485 ;
      RECT 5233.545 187.94 5233.825 325.245 ;
      RECT 5231.025 189.04 5231.305 326.965 ;
      RECT 5230.465 187.94 5230.745 326.725 ;
      RECT 5229.905 189.04 5230.185 326.485 ;
      RECT 5229.345 187.94 5229.625 326.245 ;
      RECT 5228.785 189.04 5229.065 326.005 ;
      RECT 5228.225 189.04 5228.505 325.765 ;
      RECT 5227.665 189.04 5227.945 325.525 ;
      RECT 5201.625 189.04 5201.905 328.31 ;
      RECT 5201.065 189.04 5201.345 328.55 ;
      RECT 5200.505 189.04 5200.785 328.79 ;
      RECT 5199.945 189.04 5200.225 329.03 ;
      RECT 5199.385 189.04 5199.665 329.27 ;
      RECT 5198.825 187.94 5199.105 329.51 ;
      RECT 5198.265 189.04 5198.545 329.75 ;
      RECT 5197.705 187.94 5197.985 329.99 ;
      RECT 5197.145 189.04 5197.425 330.23 ;
      RECT 5196.585 189.04 5196.865 330.47 ;
      RECT 5196.025 189.04 5196.305 330.71 ;
      RECT 5195.465 189.04 5195.745 330.95 ;
      RECT 5194.905 189.04 5195.185 331.19 ;
      RECT 5194.345 189.04 5194.625 331.43 ;
      RECT 5193.785 189.04 5194.065 331.67 ;
      RECT 5193.225 189.04 5193.505 331.67 ;
      RECT 5192.665 189.04 5192.945 331.43 ;
      RECT 5192.105 189.04 5192.385 331.19 ;
      RECT 5191.545 189.04 5191.825 330.95 ;
      RECT 5190.985 189.04 5191.265 330.705 ;
      RECT 5190.425 189.04 5190.705 330.465 ;
      RECT 5189.865 189.04 5190.145 330.225 ;
      RECT 5189.305 187.94 5189.585 329.985 ;
      RECT 5188.745 189.04 5189.025 329.745 ;
      RECT 5175.305 187.94 5175.585 327.225 ;
      RECT 5174.745 189.04 5175.025 326.985 ;
      RECT 5174.185 189.04 5174.465 326.745 ;
      RECT 5173.625 189.04 5173.905 326.505 ;
      RECT 5173.065 187.94 5173.345 326.265 ;
      RECT 5172.505 189.04 5172.785 326.025 ;
      RECT 5171.945 187.94 5172.225 325.785 ;
      RECT 5171.385 189.04 5171.665 325.545 ;
      RECT 5170.825 187.94 5171.105 325.305 ;
      RECT 5170.265 189.04 5170.545 325.065 ;
      RECT 5169.705 189.04 5169.985 324.825 ;
      RECT 5169.145 189.04 5169.425 324.585 ;
      RECT 5168.585 189.04 5168.865 324.345 ;
      RECT 5168.025 189.04 5168.305 324.105 ;
      RECT 5167.465 189.04 5167.745 323.865 ;
      RECT 5166.905 189.04 5167.185 323.625 ;
      RECT 5166.345 189.04 5166.625 323.385 ;
      RECT 5165.785 189.04 5166.065 323.145 ;
      RECT 5165.225 189.04 5165.505 322.905 ;
      RECT 5164.665 189.04 5164.945 322.665 ;
      RECT 5164.105 189.04 5164.385 322.425 ;
      RECT 5163.545 187.94 5163.825 322.185 ;
      RECT 5162.985 189.04 5163.265 321.945 ;
      RECT 5162.425 187.94 5162.705 321.705 ;
      RECT 5122.665 189.04 5122.945 332.175 ;
      RECT 5122.105 187.94 5122.385 332.415 ;
      RECT 5121.545 189.04 5121.825 332.655 ;
      RECT 5120.985 189.04 5121.265 332.895 ;
      RECT 5120.425 189.04 5120.705 333.135 ;
      RECT 5119.865 189.04 5120.145 333.375 ;
      RECT 5119.305 189.04 5119.585 333.615 ;
      RECT 5118.745 189.04 5119.025 333.86 ;
      RECT 5118.185 189.04 5118.465 334.1 ;
      RECT 5117.625 189.04 5117.905 334.34 ;
      RECT 5117.065 187.94 5117.345 334.58 ;
      RECT 5116.505 189.04 5116.785 334.82 ;
      RECT 5115.945 187.94 5116.225 335.06 ;
      RECT 5115.385 189.04 5115.665 335.3 ;
      RECT 5114.825 189.04 5115.105 335.54 ;
      RECT 5114.265 189.04 5114.545 335.78 ;
      RECT 5113.705 189.04 5113.985 336.02 ;
      RECT 5113.145 189.04 5113.425 336.26 ;
      RECT 5112.585 189.04 5112.865 336.5 ;
      RECT 5112.025 189.04 5112.305 336.74 ;
      RECT 5111.465 189.04 5111.745 336.98 ;
      RECT 5110.905 189.04 5111.185 337.22 ;
      RECT 5110.345 189.04 5110.625 337.46 ;
      RECT 5109.785 189.04 5110.065 337.7 ;
      RECT 5100.825 189.04 5101.105 333.285 ;
      RECT 5100.265 189.04 5100.545 333.045 ;
      RECT 5099.705 189.04 5099.985 332.805 ;
      RECT 5099.145 187.94 5099.425 332.565 ;
      RECT 5098.585 189.04 5098.865 332.325 ;
      RECT 5098.025 187.94 5098.305 332.085 ;
      RECT 5097.465 189.04 5097.745 331.845 ;
      RECT 5096.905 189.04 5097.185 331.605 ;
      RECT 5096.345 189.04 5096.625 331.365 ;
      RECT 5095.785 187.94 5096.065 331.125 ;
      RECT 5095.225 189.04 5095.505 330.885 ;
      RECT 5094.665 187.94 5094.945 330.645 ;
      RECT 5094.105 189.04 5094.385 330.405 ;
      RECT 5093.545 187.94 5093.825 330.165 ;
      RECT 5091.025 189.04 5091.305 322.565 ;
      RECT 5090.465 189.04 5090.745 322.325 ;
      RECT 5089.905 189.04 5090.185 322.085 ;
      RECT 5089.345 189.04 5089.625 321.845 ;
      RECT 5088.785 189.04 5089.065 321.605 ;
      RECT 5088.225 189.04 5088.505 321.365 ;
      RECT 5087.665 189.04 5087.945 321.125 ;
      RECT 5061.625 189.04 5061.905 335 ;
      RECT 5061.065 189.04 5061.345 335.24 ;
      RECT 5060.505 189.04 5060.785 335.48 ;
      RECT 5059.945 189.04 5060.225 335.72 ;
      RECT 5059.385 189.04 5059.665 335.96 ;
      RECT 5058.825 187.94 5059.105 335.96 ;
      RECT 5058.265 189.04 5058.545 335.72 ;
      RECT 5057.705 187.94 5057.985 335.475 ;
      RECT 5057.145 189.04 5057.425 335.235 ;
      RECT 5056.585 187.94 5056.865 334.995 ;
      RECT 5056.025 189.04 5056.305 334.755 ;
      RECT 5055.465 189.04 5055.745 334.515 ;
      RECT 5054.905 189.04 5055.185 334.275 ;
      RECT 5054.345 189.04 5054.625 334.035 ;
      RECT 5053.785 189.04 5054.065 333.795 ;
      RECT 5053.225 189.04 5053.505 333.555 ;
      RECT 5052.665 189.04 5052.945 333.315 ;
      RECT 5052.105 189.04 5052.385 333.075 ;
      RECT 5051.545 187.94 5051.825 332.835 ;
      RECT 5050.985 189.04 5051.265 332.595 ;
      RECT 5050.425 187.94 5050.705 332.355 ;
      RECT 5049.865 189.04 5050.145 332.115 ;
      RECT 5049.305 189.04 5049.585 331.875 ;
      RECT 5048.745 189.04 5049.025 331.635 ;
      RECT 5035.305 189.04 5035.585 335.035 ;
      RECT 5034.745 189.04 5035.025 335.275 ;
      RECT 5034.185 189.04 5034.465 335.52 ;
      RECT 5033.625 189.04 5033.905 335.76 ;
      RECT 5033.065 189.04 5033.345 336 ;
      RECT 5032.505 189.04 5032.785 336 ;
      RECT 5031.945 189.04 5032.225 335.76 ;
      RECT 5031.385 189.04 5031.665 335.52 ;
      RECT 5030.825 189.04 5031.105 328.505 ;
      RECT 5030.265 189.04 5030.545 328.265 ;
      RECT 5029.705 189.04 5029.985 328.025 ;
      RECT 5029.145 187.94 5029.425 327.785 ;
      RECT 5028.585 189.04 5028.865 327.545 ;
      RECT 5028.025 187.94 5028.305 327.305 ;
      RECT 5027.465 189.04 5027.745 327.065 ;
      RECT 5026.905 189.04 5027.185 326.825 ;
      RECT 5026.345 189.04 5026.625 326.585 ;
      RECT 5025.785 187.94 5026.065 326.345 ;
      RECT 5025.225 189.04 5025.505 326.105 ;
      RECT 5024.665 187.94 5024.945 325.865 ;
      RECT 5024.105 189.04 5024.385 325.625 ;
      RECT 5023.545 187.94 5023.825 325.385 ;
      RECT 5022.985 189.04 5023.265 325.145 ;
      RECT 5022.425 189.04 5022.705 324.905 ;
      RECT 4982.105 189.04 4982.385 333.8 ;
      RECT 4981.545 189.04 4981.825 334.04 ;
      RECT 4980.985 189.04 4981.265 334.285 ;
      RECT 4980.425 189.04 4980.705 334.525 ;
      RECT 4979.865 189.04 4980.145 334.765 ;
      RECT 4979.305 189.04 4979.585 335.005 ;
      RECT 4978.745 189.04 4979.025 335.245 ;
      RECT 4978.185 189.04 4978.465 335.485 ;
      RECT 4977.625 189.04 4977.905 335.725 ;
      RECT 4977.065 189.04 4977.345 335.965 ;
      RECT 4976.505 187.94 4976.785 336.205 ;
      RECT 4975.945 189.04 4976.225 336.445 ;
      RECT 4975.385 187.94 4975.665 336.685 ;
      RECT 4974.825 189.04 4975.105 336.925 ;
      RECT 4974.265 187.94 4974.545 337.165 ;
      RECT 4973.705 189.04 4973.985 337.165 ;
      RECT 4973.145 189.04 4973.425 336.925 ;
      RECT 4972.585 189.04 4972.865 336.685 ;
      RECT 4972.025 189.04 4972.305 336.445 ;
      RECT 4971.465 189.04 4971.745 336.205 ;
      RECT 4970.905 189.04 4971.185 335.965 ;
      RECT 4970.345 189.04 4970.625 335.725 ;
      RECT 4969.785 189.04 4970.065 335.485 ;
      RECT 4960.825 187.94 4961.105 335.515 ;
      RECT 4960.265 189.04 4960.545 335.755 ;
      RECT 4959.705 187.94 4959.985 335.995 ;
      RECT 4959.145 189.04 4959.425 336.21 ;
      RECT 4958.585 189.04 4958.865 335.785 ;
      RECT 4958.025 189.04 4958.305 335.545 ;
      RECT 4957.465 189.04 4957.745 335.305 ;
      RECT 4956.905 189.04 4957.185 335.065 ;
      RECT 4956.345 189.04 4956.625 334.825 ;
      RECT 4955.785 189.04 4956.065 334.585 ;
      RECT 4955.225 189.04 4955.505 334.345 ;
      RECT 4954.665 189.04 4954.945 334.105 ;
      RECT 4954.105 189.04 4954.385 333.865 ;
      RECT 4953.545 189.04 4953.825 333.625 ;
      RECT 4951.025 189.04 4951.305 332.8 ;
      RECT 4950.465 189.04 4950.745 332.56 ;
      RECT 4949.905 189.04 4950.185 332.32 ;
      RECT 4949.345 187.94 4949.625 332.08 ;
      RECT 4948.785 189.04 4949.065 331.84 ;
      RECT 4948.225 187.94 4948.505 331.6 ;
      RECT 4947.665 189.04 4947.945 331.36 ;
      RECT 4947.105 189.04 4947.385 331.12 ;
      RECT 4920.505 189.04 4920.785 342.165 ;
      RECT 4919.945 187.94 4920.225 342.405 ;
      RECT 4919.385 189.04 4919.665 342.645 ;
      RECT 4918.825 187.94 4919.105 342.89 ;
      RECT 4918.265 189.04 4918.545 343.13 ;
      RECT 4917.705 187.94 4917.985 343.37 ;
      RECT 4917.145 189.04 4917.425 343.61 ;
      RECT 4916.585 189.04 4916.865 343.85 ;
      RECT 4916.025 189.04 4916.305 329.47 ;
      RECT 4915.465 189.04 4915.745 329.23 ;
      RECT 4914.905 189.04 4915.185 328.99 ;
      RECT 4914.345 189.04 4914.625 328.75 ;
      RECT 4913.785 189.04 4914.065 328.51 ;
      RECT 4913.225 189.04 4913.505 328.27 ;
      RECT 4912.665 189.04 4912.945 328.03 ;
      RECT 4912.105 189.04 4912.385 327.79 ;
      RECT 4911.545 189.04 4911.825 327.55 ;
      RECT 4910.985 189.04 4911.265 327.31 ;
      RECT 4910.425 187.94 4910.705 327.07 ;
      RECT 4909.865 189.04 4910.145 326.83 ;
      RECT 4909.305 187.94 4909.585 326.59 ;
      RECT 4908.745 189.04 4909.025 326.35 ;
      RECT 4894.745 187.94 4895.025 332.47 ;
      RECT 4894.185 189.04 4894.465 332.23 ;
      RECT 4893.625 189.04 4893.905 331.99 ;
      RECT 4893.065 189.04 4893.345 331.75 ;
      RECT 4892.505 189.04 4892.785 331.51 ;
      RECT 4891.945 189.04 4892.225 331.27 ;
      RECT 4891.385 189.04 4891.665 331.03 ;
      RECT 4890.825 189.04 4891.105 330.79 ;
      RECT 4890.265 189.04 4890.545 330.55 ;
      RECT 4889.705 187.94 4889.985 330.31 ;
      RECT 4889.145 189.04 4889.425 330.07 ;
      RECT 4888.585 187.94 4888.865 329.83 ;
      RECT 4888.025 189.04 4888.305 329.59 ;
      RECT 4887.465 189.04 4887.745 329.35 ;
      RECT 4886.905 189.04 4887.185 329.11 ;
      RECT 4886.345 189.04 4886.625 328.87 ;
      RECT 4885.785 189.04 4886.065 328.63 ;
      RECT 4885.225 189.04 4885.505 328.39 ;
      RECT 4884.665 189.04 4884.945 328.15 ;
      RECT 4884.105 189.04 4884.385 327.91 ;
      RECT 4883.545 189.04 4883.825 327.67 ;
      RECT 4882.985 189.04 4883.265 327.43 ;
      RECT 4882.425 189.04 4882.705 327.19 ;
      RECT 4843.225 189.04 4843.505 334.095 ;
      RECT 4842.665 189.04 4842.945 334.335 ;
      RECT 4842.105 189.04 4842.385 334.575 ;
      RECT 4841.545 187.94 4841.825 334.815 ;
      RECT 4840.985 189.04 4841.265 335.055 ;
      RECT 4840.425 187.94 4840.705 335.295 ;
      RECT 4839.865 189.04 4840.145 335.535 ;
      RECT 4839.305 189.04 4839.585 335.775 ;
      RECT 4838.745 189.04 4839.025 336.015 ;
      RECT 4838.185 187.94 4838.465 336.255 ;
      RECT 4837.625 189.04 4837.905 336.495 ;
      RECT 4837.065 187.94 4837.345 336.735 ;
      RECT 4836.505 189.04 4836.785 336.975 ;
      RECT 4835.945 187.94 4836.225 337.215 ;
      RECT 4835.385 189.04 4835.665 337.455 ;
      RECT 4834.825 189.04 4835.105 337.695 ;
      RECT 4834.265 189.04 4834.545 337.695 ;
      RECT 4833.705 189.04 4833.985 337.455 ;
      RECT 4833.145 189.04 4833.425 337.215 ;
      RECT 4832.585 189.04 4832.865 336.975 ;
      RECT 4832.025 189.04 4832.305 336.735 ;
      RECT 4831.465 189.04 4831.745 336.495 ;
      RECT 4830.905 189.04 4831.185 336.255 ;
      RECT 4830.345 189.04 4830.625 336.015 ;
      RECT 4829.785 189.04 4830.065 335.775 ;
      RECT 4820.825 189.04 4821.105 335.29 ;
      RECT 4820.265 187.94 4820.545 335.05 ;
      RECT 4819.705 189.04 4819.985 334.81 ;
      RECT 4819.145 187.94 4819.425 334.57 ;
      RECT 4818.585 189.04 4818.865 334.33 ;
      RECT 4818.025 187.94 4818.305 334.09 ;
      RECT 4817.465 189.04 4817.745 333.85 ;
      RECT 4816.905 189.04 4817.185 333.61 ;
      RECT 4816.345 189.04 4816.625 333.37 ;
      RECT 4815.785 189.04 4816.065 333.13 ;
      RECT 4815.225 189.04 4815.505 332.89 ;
      RECT 4814.665 189.04 4814.945 332.65 ;
      RECT 4814.105 189.04 4814.385 332.41 ;
      RECT 4813.545 189.04 4813.825 332.17 ;
      RECT 4811.025 187.94 4811.305 333.89 ;
      RECT 4810.465 189.04 4810.745 333.65 ;
      RECT 4809.905 187.94 4810.185 333.41 ;
      RECT 4809.345 189.04 4809.625 333.17 ;
      RECT 4808.785 189.04 4809.065 332.93 ;
      RECT 4808.225 189.04 4808.505 332.69 ;
      RECT 4807.665 189.04 4807.945 332.45 ;
      RECT 4807.105 189.04 4807.385 332.21 ;
      RECT 4781.065 189.04 4781.345 329.86 ;
      RECT 4780.505 189.04 4780.785 330.1 ;
      RECT 4779.945 189.04 4780.225 330.34 ;
      RECT 4779.385 189.04 4779.665 330.585 ;
      RECT 4778.825 189.04 4779.105 330.825 ;
      RECT 4778.265 189.04 4778.545 331.065 ;
      RECT 4777.705 189.04 4777.985 331.065 ;
      RECT 4777.145 189.04 4777.425 330.825 ;
      RECT 4776.585 189.04 4776.865 330.585 ;
      RECT 4776.025 187.94 4776.305 330.345 ;
      RECT 4775.465 189.04 4775.745 330.105 ;
      RECT 4774.905 187.94 4775.185 329.865 ;
      RECT 4774.345 189.04 4774.625 329.625 ;
      RECT 4773.785 189.04 4774.065 329.385 ;
      RECT 4773.225 189.04 4773.505 329.145 ;
      RECT 4772.665 187.94 4772.945 328.905 ;
      RECT 4772.105 189.04 4772.385 328.665 ;
      RECT 4771.545 187.94 4771.825 328.425 ;
      RECT 4770.985 189.04 4771.265 328.185 ;
      RECT 4770.425 187.94 4770.705 327.945 ;
      RECT 4769.865 189.04 4770.145 327.705 ;
      RECT 4769.305 189.04 4769.585 327.465 ;
      RECT 4768.745 189.04 4769.025 327.225 ;
      RECT 4768.185 189.04 4768.465 326.985 ;
      RECT 4754.745 189.04 4755.025 332.785 ;
      RECT 4754.185 189.04 4754.465 332.545 ;
      RECT 4753.625 189.04 4753.905 332.305 ;
      RECT 4753.065 189.04 4753.345 332.065 ;
      RECT 4752.505 189.04 4752.785 331.825 ;
      RECT 4751.945 189.04 4752.225 331.585 ;
      RECT 4751.385 189.04 4751.665 331.345 ;
      RECT 4750.825 189.04 4751.105 331.105 ;
      RECT 4750.265 187.94 4750.545 330.865 ;
      RECT 4749.705 189.04 4749.985 330.625 ;
      RECT 4749.145 187.94 4749.425 330.305 ;
      RECT 4748.585 189.04 4748.865 330.145 ;
      RECT 4748.025 187.94 4748.305 329.905 ;
      RECT 4747.465 189.04 4747.745 329.665 ;
      RECT 4746.905 189.04 4747.185 329.425 ;
      RECT 4746.345 189.04 4746.625 329.185 ;
      RECT 4745.785 189.04 4746.065 328.945 ;
      RECT 4745.225 189.04 4745.505 328.705 ;
      RECT 4744.665 189.04 4744.945 328.465 ;
      RECT 4744.105 189.04 4744.385 328.225 ;
      RECT 4743.545 189.04 4743.825 327.985 ;
      RECT 4742.985 187.94 4743.265 327.745 ;
      RECT 4742.425 189.04 4742.705 327.505 ;
      RECT 4741.865 187.94 4742.145 327.265 ;
      RECT 4702.665 189.04 4702.945 332.875 ;
      RECT 4702.105 189.04 4702.385 333.115 ;
      RECT 4701.545 189.04 4701.825 333.355 ;
      RECT 4700.985 189.04 4701.265 333.595 ;
      RECT 4700.425 189.04 4700.705 333.835 ;
      RECT 4699.865 189.04 4700.145 334.075 ;
      RECT 4699.305 189.04 4699.585 334.315 ;
      RECT 4698.745 189.04 4699.025 334.555 ;
      RECT 4698.185 189.04 4698.465 334.795 ;
      RECT 4697.625 189.04 4697.905 335.035 ;
      RECT 4697.065 189.04 4697.345 335.275 ;
      RECT 4696.505 189.04 4696.785 335.515 ;
      RECT 4695.945 189.04 4696.225 335.755 ;
      RECT 4695.385 189.04 4695.665 335.755 ;
      RECT 4694.825 187.94 4695.105 335.515 ;
      RECT 4694.265 189.04 4694.545 335.275 ;
      RECT 4693.705 187.94 4693.985 335.035 ;
      RECT 4693.145 189.04 4693.425 334.795 ;
      RECT 4692.585 189.04 4692.865 334.555 ;
      RECT 4692.025 189.04 4692.305 334.315 ;
      RECT 4691.465 187.94 4691.745 334.05 ;
      RECT 4690.905 189.04 4691.185 333.81 ;
      RECT 4690.345 187.94 4690.625 333.57 ;
      RECT 4689.785 189.04 4690.065 333.33 ;
      RECT 4680.825 187.94 4681.105 327.165 ;
      RECT 4680.265 189.04 4680.545 327.405 ;
      RECT 4679.705 189.04 4679.985 327.645 ;
      RECT 4679.145 189.04 4679.425 327.645 ;
      RECT 4678.585 189.04 4678.865 327.405 ;
      RECT 4678.025 189.04 4678.305 327.165 ;
      RECT 4677.465 189.04 4677.745 326.925 ;
      RECT 4676.905 189.04 4677.185 326.685 ;
      RECT 4676.345 189.04 4676.625 326.445 ;
      RECT 4675.785 189.04 4676.065 326.205 ;
      RECT 4675.225 189.04 4675.505 325.965 ;
      RECT 4674.665 189.04 4674.945 325.725 ;
      RECT 4674.105 189.04 4674.385 325.485 ;
      RECT 4673.545 187.94 4673.825 325.245 ;
      RECT 4671.025 189.04 4671.305 326.965 ;
      RECT 4670.465 187.94 4670.745 326.725 ;
      RECT 4669.905 189.04 4670.185 326.485 ;
      RECT 4669.345 187.94 4669.625 326.245 ;
      RECT 4668.785 189.04 4669.065 326.005 ;
      RECT 4668.225 189.04 4668.505 325.765 ;
      RECT 4667.665 189.04 4667.945 325.525 ;
      RECT 4641.625 189.04 4641.905 328.31 ;
      RECT 4641.065 189.04 4641.345 328.55 ;
      RECT 4640.505 189.04 4640.785 328.79 ;
      RECT 4639.945 189.04 4640.225 329.03 ;
      RECT 4639.385 189.04 4639.665 329.27 ;
      RECT 4638.825 187.94 4639.105 329.51 ;
      RECT 4638.265 189.04 4638.545 329.75 ;
      RECT 4637.705 187.94 4637.985 329.99 ;
      RECT 4637.145 189.04 4637.425 330.23 ;
      RECT 4636.585 189.04 4636.865 330.47 ;
      RECT 4636.025 189.04 4636.305 330.71 ;
      RECT 4635.465 189.04 4635.745 330.95 ;
      RECT 4634.905 189.04 4635.185 331.19 ;
      RECT 4634.345 189.04 4634.625 331.43 ;
      RECT 4633.785 189.04 4634.065 331.67 ;
      RECT 4633.225 189.04 4633.505 331.67 ;
      RECT 4632.665 189.04 4632.945 331.43 ;
      RECT 4632.105 189.04 4632.385 331.19 ;
      RECT 4631.545 189.04 4631.825 330.95 ;
      RECT 4630.985 189.04 4631.265 330.705 ;
      RECT 4630.425 189.04 4630.705 330.465 ;
      RECT 4629.865 189.04 4630.145 330.225 ;
      RECT 4629.305 187.94 4629.585 329.985 ;
      RECT 4628.745 189.04 4629.025 329.745 ;
      RECT 4615.305 187.94 4615.585 327.225 ;
      RECT 4614.745 189.04 4615.025 326.985 ;
      RECT 4614.185 189.04 4614.465 326.745 ;
      RECT 4613.625 189.04 4613.905 326.505 ;
      RECT 4613.065 187.94 4613.345 326.265 ;
      RECT 4612.505 189.04 4612.785 326.025 ;
      RECT 4611.945 187.94 4612.225 325.785 ;
      RECT 4611.385 189.04 4611.665 325.545 ;
      RECT 4610.825 187.94 4611.105 325.305 ;
      RECT 4610.265 189.04 4610.545 325.065 ;
      RECT 4609.705 189.04 4609.985 324.825 ;
      RECT 4609.145 189.04 4609.425 324.585 ;
      RECT 4608.585 189.04 4608.865 324.345 ;
      RECT 4608.025 189.04 4608.305 324.105 ;
      RECT 4607.465 189.04 4607.745 323.865 ;
      RECT 4606.905 189.04 4607.185 323.625 ;
      RECT 4606.345 189.04 4606.625 323.385 ;
      RECT 4605.785 189.04 4606.065 323.145 ;
      RECT 4605.225 189.04 4605.505 322.905 ;
      RECT 4604.665 189.04 4604.945 322.665 ;
      RECT 4604.105 189.04 4604.385 322.425 ;
      RECT 4603.545 187.94 4603.825 322.185 ;
      RECT 4602.985 189.04 4603.265 321.945 ;
      RECT 4602.425 187.94 4602.705 321.705 ;
      RECT 4562.665 189.04 4562.945 332.175 ;
      RECT 4562.105 187.94 4562.385 332.415 ;
      RECT 4561.545 189.04 4561.825 332.655 ;
      RECT 4560.985 189.04 4561.265 332.895 ;
      RECT 4560.425 189.04 4560.705 333.135 ;
      RECT 4559.865 189.04 4560.145 333.375 ;
      RECT 4559.305 189.04 4559.585 333.615 ;
      RECT 4558.745 189.04 4559.025 333.86 ;
      RECT 4558.185 189.04 4558.465 334.1 ;
      RECT 4557.625 189.04 4557.905 334.34 ;
      RECT 4557.065 187.94 4557.345 334.58 ;
      RECT 4556.505 189.04 4556.785 334.82 ;
      RECT 4555.945 187.94 4556.225 335.06 ;
      RECT 4555.385 189.04 4555.665 335.3 ;
      RECT 4554.825 189.04 4555.105 335.54 ;
      RECT 4554.265 189.04 4554.545 335.78 ;
      RECT 4553.705 189.04 4553.985 336.02 ;
      RECT 4553.145 189.04 4553.425 336.26 ;
      RECT 4552.585 189.04 4552.865 336.5 ;
      RECT 4552.025 189.04 4552.305 336.74 ;
      RECT 4551.465 189.04 4551.745 336.98 ;
      RECT 4550.905 189.04 4551.185 337.22 ;
      RECT 4550.345 189.04 4550.625 337.46 ;
      RECT 4549.785 189.04 4550.065 337.7 ;
      RECT 4540.825 189.04 4541.105 333.285 ;
      RECT 4540.265 189.04 4540.545 333.045 ;
      RECT 4539.705 189.04 4539.985 332.805 ;
      RECT 4539.145 187.94 4539.425 332.565 ;
      RECT 4538.585 189.04 4538.865 332.325 ;
      RECT 4538.025 187.94 4538.305 332.085 ;
      RECT 4537.465 189.04 4537.745 331.845 ;
      RECT 4536.905 189.04 4537.185 331.605 ;
      RECT 4536.345 189.04 4536.625 331.365 ;
      RECT 4535.785 187.94 4536.065 331.125 ;
      RECT 4535.225 189.04 4535.505 330.885 ;
      RECT 4534.665 187.94 4534.945 330.645 ;
      RECT 4534.105 189.04 4534.385 330.405 ;
      RECT 4533.545 187.94 4533.825 330.165 ;
      RECT 4531.025 189.04 4531.305 322.565 ;
      RECT 4530.465 189.04 4530.745 322.325 ;
      RECT 4529.905 189.04 4530.185 322.085 ;
      RECT 4529.345 189.04 4529.625 321.845 ;
      RECT 4528.785 189.04 4529.065 321.605 ;
      RECT 4528.225 189.04 4528.505 321.365 ;
      RECT 4527.665 189.04 4527.945 321.125 ;
      RECT 4501.625 189.04 4501.905 335 ;
      RECT 4501.065 189.04 4501.345 335.24 ;
      RECT 4500.505 189.04 4500.785 335.48 ;
      RECT 4499.945 189.04 4500.225 335.72 ;
      RECT 4499.385 189.04 4499.665 335.96 ;
      RECT 4498.825 187.94 4499.105 335.96 ;
      RECT 4498.265 189.04 4498.545 335.72 ;
      RECT 4497.705 187.94 4497.985 335.475 ;
      RECT 4497.145 189.04 4497.425 335.235 ;
      RECT 4496.585 187.94 4496.865 334.995 ;
      RECT 4496.025 189.04 4496.305 334.755 ;
      RECT 4495.465 189.04 4495.745 334.515 ;
      RECT 4494.905 189.04 4495.185 334.275 ;
      RECT 4494.345 189.04 4494.625 334.035 ;
      RECT 4493.785 189.04 4494.065 333.795 ;
      RECT 4493.225 189.04 4493.505 333.555 ;
      RECT 4492.665 189.04 4492.945 333.315 ;
      RECT 4492.105 189.04 4492.385 333.075 ;
      RECT 4491.545 187.94 4491.825 332.835 ;
      RECT 4490.985 189.04 4491.265 332.595 ;
      RECT 4490.425 187.94 4490.705 332.355 ;
      RECT 4489.865 189.04 4490.145 332.115 ;
      RECT 4489.305 189.04 4489.585 331.875 ;
      RECT 4488.745 189.04 4489.025 331.635 ;
      RECT 4475.305 189.04 4475.585 335.035 ;
      RECT 4474.745 189.04 4475.025 335.275 ;
      RECT 4474.185 189.04 4474.465 335.52 ;
      RECT 4473.625 189.04 4473.905 335.76 ;
      RECT 4473.065 189.04 4473.345 336 ;
      RECT 4472.505 189.04 4472.785 336 ;
      RECT 4471.945 189.04 4472.225 335.76 ;
      RECT 4471.385 189.04 4471.665 335.52 ;
      RECT 4470.825 189.04 4471.105 328.505 ;
      RECT 4470.265 189.04 4470.545 328.265 ;
      RECT 4469.705 189.04 4469.985 328.025 ;
      RECT 4469.145 187.94 4469.425 327.785 ;
      RECT 4468.585 189.04 4468.865 327.545 ;
      RECT 4468.025 187.94 4468.305 327.305 ;
      RECT 4467.465 189.04 4467.745 327.065 ;
      RECT 4466.905 189.04 4467.185 326.825 ;
      RECT 4466.345 189.04 4466.625 326.585 ;
      RECT 4465.785 187.94 4466.065 326.345 ;
      RECT 4465.225 189.04 4465.505 326.105 ;
      RECT 4464.665 187.94 4464.945 325.865 ;
      RECT 4464.105 189.04 4464.385 325.625 ;
      RECT 4463.545 187.94 4463.825 325.385 ;
      RECT 4462.985 189.04 4463.265 325.145 ;
      RECT 4462.425 189.04 4462.705 324.905 ;
      RECT 4422.105 189.04 4422.385 333.8 ;
      RECT 4421.545 189.04 4421.825 334.04 ;
      RECT 4420.985 189.04 4421.265 334.285 ;
      RECT 4420.425 189.04 4420.705 334.525 ;
      RECT 4419.865 189.04 4420.145 334.765 ;
      RECT 4419.305 189.04 4419.585 335.005 ;
      RECT 4418.745 189.04 4419.025 335.245 ;
      RECT 4418.185 189.04 4418.465 335.485 ;
      RECT 4417.625 189.04 4417.905 335.725 ;
      RECT 4417.065 189.04 4417.345 335.965 ;
      RECT 4416.505 187.94 4416.785 336.205 ;
      RECT 4415.945 189.04 4416.225 336.445 ;
      RECT 4415.385 187.94 4415.665 336.685 ;
      RECT 4414.825 189.04 4415.105 336.925 ;
      RECT 4414.265 187.94 4414.545 337.165 ;
      RECT 4413.705 189.04 4413.985 337.165 ;
      RECT 4413.145 189.04 4413.425 336.925 ;
      RECT 4412.585 189.04 4412.865 336.685 ;
      RECT 4412.025 189.04 4412.305 336.445 ;
      RECT 4411.465 189.04 4411.745 336.205 ;
      RECT 4410.905 189.04 4411.185 335.965 ;
      RECT 4410.345 189.04 4410.625 335.725 ;
      RECT 4409.785 189.04 4410.065 335.485 ;
      RECT 4400.825 187.94 4401.105 335.515 ;
      RECT 4400.265 189.04 4400.545 335.755 ;
      RECT 4399.705 187.94 4399.985 335.995 ;
      RECT 4399.145 189.04 4399.425 336.21 ;
      RECT 4398.585 189.04 4398.865 335.785 ;
      RECT 4398.025 189.04 4398.305 335.545 ;
      RECT 4397.465 189.04 4397.745 335.305 ;
      RECT 4396.905 189.04 4397.185 335.065 ;
      RECT 4396.345 189.04 4396.625 334.825 ;
      RECT 4395.785 189.04 4396.065 334.585 ;
      RECT 4395.225 189.04 4395.505 334.345 ;
      RECT 4394.665 189.04 4394.945 334.105 ;
      RECT 4394.105 189.04 4394.385 333.865 ;
      RECT 4393.545 189.04 4393.825 333.625 ;
      RECT 4391.025 189.04 4391.305 332.8 ;
      RECT 4390.465 189.04 4390.745 332.56 ;
      RECT 4389.905 189.04 4390.185 332.32 ;
      RECT 4389.345 187.94 4389.625 332.08 ;
      RECT 4388.785 189.04 4389.065 331.84 ;
      RECT 4388.225 187.94 4388.505 331.6 ;
      RECT 4387.665 189.04 4387.945 331.36 ;
      RECT 4387.105 189.04 4387.385 331.12 ;
      RECT 4360.505 189.04 4360.785 342.165 ;
      RECT 4359.945 187.94 4360.225 342.405 ;
      RECT 4359.385 189.04 4359.665 342.645 ;
      RECT 4358.825 187.94 4359.105 342.89 ;
      RECT 4358.265 189.04 4358.545 343.13 ;
      RECT 4357.705 187.94 4357.985 343.37 ;
      RECT 4357.145 189.04 4357.425 343.61 ;
      RECT 4356.585 189.04 4356.865 343.85 ;
      RECT 4356.025 189.04 4356.305 329.47 ;
      RECT 4355.465 189.04 4355.745 329.23 ;
      RECT 4354.905 189.04 4355.185 328.99 ;
      RECT 4354.345 189.04 4354.625 328.75 ;
      RECT 4353.785 189.04 4354.065 328.51 ;
      RECT 4353.225 189.04 4353.505 328.27 ;
      RECT 4352.665 189.04 4352.945 328.03 ;
      RECT 4352.105 189.04 4352.385 327.79 ;
      RECT 4351.545 189.04 4351.825 327.55 ;
      RECT 4350.985 189.04 4351.265 327.31 ;
      RECT 4350.425 187.94 4350.705 327.07 ;
      RECT 4349.865 189.04 4350.145 326.83 ;
      RECT 4349.305 187.94 4349.585 326.59 ;
      RECT 4348.745 189.04 4349.025 326.35 ;
      RECT 4334.745 187.94 4335.025 332.47 ;
      RECT 4334.185 189.04 4334.465 332.23 ;
      RECT 4333.625 189.04 4333.905 331.99 ;
      RECT 4333.065 189.04 4333.345 331.75 ;
      RECT 4332.505 189.04 4332.785 331.51 ;
      RECT 4331.945 189.04 4332.225 331.27 ;
      RECT 4331.385 189.04 4331.665 331.03 ;
      RECT 4330.825 189.04 4331.105 330.79 ;
      RECT 4330.265 189.04 4330.545 330.55 ;
      RECT 4329.705 187.94 4329.985 330.31 ;
      RECT 4329.145 189.04 4329.425 330.07 ;
      RECT 4328.585 187.94 4328.865 329.83 ;
      RECT 4328.025 189.04 4328.305 329.59 ;
      RECT 4327.465 189.04 4327.745 329.35 ;
      RECT 4326.905 189.04 4327.185 329.11 ;
      RECT 4326.345 189.04 4326.625 328.87 ;
      RECT 4325.785 189.04 4326.065 328.63 ;
      RECT 4325.225 189.04 4325.505 328.39 ;
      RECT 4324.665 189.04 4324.945 328.15 ;
      RECT 4324.105 189.04 4324.385 327.91 ;
      RECT 4323.545 189.04 4323.825 327.67 ;
      RECT 4322.985 189.04 4323.265 327.43 ;
      RECT 4322.425 189.04 4322.705 327.19 ;
      RECT 4283.225 189.04 4283.505 334.095 ;
      RECT 4282.665 189.04 4282.945 334.335 ;
      RECT 4282.105 189.04 4282.385 334.575 ;
      RECT 4281.545 187.94 4281.825 334.815 ;
      RECT 4280.985 189.04 4281.265 335.055 ;
      RECT 4280.425 187.94 4280.705 335.295 ;
      RECT 4279.865 189.04 4280.145 335.535 ;
      RECT 4279.305 189.04 4279.585 335.775 ;
      RECT 4278.745 189.04 4279.025 336.015 ;
      RECT 4278.185 187.94 4278.465 336.255 ;
      RECT 4277.625 189.04 4277.905 336.495 ;
      RECT 4277.065 187.94 4277.345 336.735 ;
      RECT 4276.505 189.04 4276.785 336.975 ;
      RECT 4275.945 187.94 4276.225 337.215 ;
      RECT 4275.385 189.04 4275.665 337.455 ;
      RECT 4274.825 189.04 4275.105 337.695 ;
      RECT 4274.265 189.04 4274.545 337.695 ;
      RECT 4273.705 189.04 4273.985 337.455 ;
      RECT 4273.145 189.04 4273.425 337.215 ;
      RECT 4272.585 189.04 4272.865 336.975 ;
      RECT 4272.025 189.04 4272.305 336.735 ;
      RECT 4271.465 189.04 4271.745 336.495 ;
      RECT 4270.905 189.04 4271.185 336.255 ;
      RECT 4270.345 189.04 4270.625 336.015 ;
      RECT 4269.785 189.04 4270.065 335.775 ;
      RECT 4260.825 189.04 4261.105 335.29 ;
      RECT 4260.265 187.94 4260.545 335.05 ;
      RECT 4259.705 189.04 4259.985 334.81 ;
      RECT 4259.145 187.94 4259.425 334.57 ;
      RECT 4258.585 189.04 4258.865 334.33 ;
      RECT 4258.025 187.94 4258.305 334.09 ;
      RECT 4257.465 189.04 4257.745 333.85 ;
      RECT 4256.905 189.04 4257.185 333.61 ;
      RECT 4256.345 189.04 4256.625 333.37 ;
      RECT 4255.785 189.04 4256.065 333.13 ;
      RECT 4255.225 189.04 4255.505 332.89 ;
      RECT 4254.665 189.04 4254.945 332.65 ;
      RECT 4254.105 189.04 4254.385 332.41 ;
      RECT 4253.545 189.04 4253.825 332.17 ;
      RECT 4251.025 187.94 4251.305 333.89 ;
      RECT 4250.465 189.04 4250.745 333.65 ;
      RECT 4249.905 187.94 4250.185 333.41 ;
      RECT 4249.345 189.04 4249.625 333.17 ;
      RECT 4248.785 189.04 4249.065 332.93 ;
      RECT 4248.225 189.04 4248.505 332.69 ;
      RECT 4247.665 189.04 4247.945 332.45 ;
      RECT 4247.105 189.04 4247.385 332.21 ;
      RECT 4221.065 189.04 4221.345 329.86 ;
      RECT 4220.505 189.04 4220.785 330.1 ;
      RECT 4219.945 189.04 4220.225 330.34 ;
      RECT 4219.385 189.04 4219.665 330.585 ;
      RECT 4218.825 189.04 4219.105 330.825 ;
      RECT 4218.265 189.04 4218.545 331.065 ;
      RECT 4217.705 189.04 4217.985 331.065 ;
      RECT 4217.145 189.04 4217.425 330.825 ;
      RECT 4216.585 189.04 4216.865 330.585 ;
      RECT 4216.025 187.94 4216.305 330.345 ;
      RECT 4215.465 189.04 4215.745 330.105 ;
      RECT 4214.905 187.94 4215.185 329.865 ;
      RECT 4214.345 189.04 4214.625 329.625 ;
      RECT 4213.785 189.04 4214.065 329.385 ;
      RECT 4213.225 189.04 4213.505 329.145 ;
      RECT 4212.665 187.94 4212.945 328.905 ;
      RECT 4212.105 189.04 4212.385 328.665 ;
      RECT 4211.545 187.94 4211.825 328.425 ;
      RECT 4210.985 189.04 4211.265 328.185 ;
      RECT 4210.425 187.94 4210.705 327.945 ;
      RECT 4209.865 189.04 4210.145 327.705 ;
      RECT 4209.305 189.04 4209.585 327.465 ;
      RECT 4208.745 189.04 4209.025 327.225 ;
      RECT 4208.185 189.04 4208.465 326.985 ;
      RECT 4194.745 189.04 4195.025 332.785 ;
      RECT 4194.185 189.04 4194.465 332.545 ;
      RECT 4193.625 189.04 4193.905 332.305 ;
      RECT 4193.065 189.04 4193.345 332.065 ;
      RECT 4192.505 189.04 4192.785 331.825 ;
      RECT 4191.945 189.04 4192.225 331.585 ;
      RECT 4191.385 189.04 4191.665 331.345 ;
      RECT 4190.825 189.04 4191.105 331.105 ;
      RECT 4190.265 187.94 4190.545 330.865 ;
      RECT 4189.705 189.04 4189.985 330.625 ;
      RECT 4189.145 187.94 4189.425 330.305 ;
      RECT 4188.585 189.04 4188.865 330.145 ;
      RECT 4188.025 187.94 4188.305 329.905 ;
      RECT 4187.465 189.04 4187.745 329.665 ;
      RECT 4186.905 189.04 4187.185 329.425 ;
      RECT 4186.345 189.04 4186.625 329.185 ;
      RECT 4185.785 189.04 4186.065 328.945 ;
      RECT 4185.225 189.04 4185.505 328.705 ;
      RECT 4184.665 189.04 4184.945 328.465 ;
      RECT 4184.105 189.04 4184.385 328.225 ;
      RECT 4183.545 189.04 4183.825 327.985 ;
      RECT 4182.985 187.94 4183.265 327.745 ;
      RECT 4182.425 189.04 4182.705 327.505 ;
      RECT 4181.865 187.94 4182.145 327.265 ;
      RECT 4142.665 189.04 4142.945 332.875 ;
      RECT 4142.105 189.04 4142.385 333.115 ;
      RECT 4141.545 189.04 4141.825 333.355 ;
      RECT 4140.985 189.04 4141.265 333.595 ;
      RECT 4140.425 189.04 4140.705 333.835 ;
      RECT 4139.865 189.04 4140.145 334.075 ;
      RECT 4139.305 189.04 4139.585 334.315 ;
      RECT 4138.745 189.04 4139.025 334.555 ;
      RECT 4138.185 189.04 4138.465 334.795 ;
      RECT 4137.625 189.04 4137.905 335.035 ;
      RECT 4137.065 189.04 4137.345 335.275 ;
      RECT 4136.505 189.04 4136.785 335.515 ;
      RECT 4135.945 189.04 4136.225 335.755 ;
      RECT 4135.385 189.04 4135.665 335.755 ;
      RECT 4134.825 187.94 4135.105 335.515 ;
      RECT 4134.265 189.04 4134.545 335.275 ;
      RECT 4133.705 187.94 4133.985 335.035 ;
      RECT 4133.145 189.04 4133.425 334.795 ;
      RECT 4132.585 189.04 4132.865 334.555 ;
      RECT 4132.025 189.04 4132.305 334.315 ;
      RECT 4131.465 187.94 4131.745 334.05 ;
      RECT 4130.905 189.04 4131.185 333.81 ;
      RECT 4130.345 187.94 4130.625 333.57 ;
      RECT 4129.785 189.04 4130.065 333.33 ;
      RECT 4120.825 187.94 4121.105 327.165 ;
      RECT 4120.265 189.04 4120.545 327.405 ;
      RECT 4119.705 189.04 4119.985 327.645 ;
      RECT 4119.145 189.04 4119.425 327.645 ;
      RECT 4118.585 189.04 4118.865 327.405 ;
      RECT 4118.025 189.04 4118.305 327.165 ;
      RECT 4117.465 189.04 4117.745 326.925 ;
      RECT 4116.905 189.04 4117.185 326.685 ;
      RECT 4116.345 189.04 4116.625 326.445 ;
      RECT 4115.785 189.04 4116.065 326.205 ;
      RECT 4115.225 189.04 4115.505 325.965 ;
      RECT 4114.665 189.04 4114.945 325.725 ;
      RECT 4114.105 189.04 4114.385 325.485 ;
      RECT 4113.545 187.94 4113.825 325.245 ;
      RECT 4111.025 189.04 4111.305 326.965 ;
      RECT 4110.465 187.94 4110.745 326.725 ;
      RECT 4109.905 189.04 4110.185 326.485 ;
      RECT 4109.345 187.94 4109.625 326.245 ;
      RECT 4108.785 189.04 4109.065 326.005 ;
      RECT 4108.225 189.04 4108.505 325.765 ;
      RECT 4107.665 189.04 4107.945 325.525 ;
      RECT 4081.625 189.04 4081.905 328.31 ;
      RECT 4081.065 189.04 4081.345 328.55 ;
      RECT 4080.505 189.04 4080.785 328.79 ;
      RECT 4079.945 189.04 4080.225 329.03 ;
      RECT 4079.385 189.04 4079.665 329.27 ;
      RECT 4078.825 187.94 4079.105 329.51 ;
      RECT 4078.265 189.04 4078.545 329.75 ;
      RECT 4077.705 187.94 4077.985 329.99 ;
      RECT 4077.145 189.04 4077.425 330.23 ;
      RECT 4076.585 189.04 4076.865 330.47 ;
      RECT 4076.025 189.04 4076.305 330.71 ;
      RECT 4075.465 189.04 4075.745 330.95 ;
      RECT 4074.905 189.04 4075.185 331.19 ;
      RECT 4074.345 189.04 4074.625 331.43 ;
      RECT 4073.785 189.04 4074.065 331.67 ;
      RECT 4073.225 189.04 4073.505 331.67 ;
      RECT 4072.665 189.04 4072.945 331.43 ;
      RECT 4072.105 189.04 4072.385 331.19 ;
      RECT 4071.545 189.04 4071.825 330.95 ;
      RECT 4070.985 189.04 4071.265 330.705 ;
      RECT 4070.425 189.04 4070.705 330.465 ;
      RECT 4069.865 189.04 4070.145 330.225 ;
      RECT 4069.305 187.94 4069.585 329.985 ;
      RECT 4068.745 189.04 4069.025 329.745 ;
      RECT 4055.305 187.94 4055.585 327.225 ;
      RECT 4054.745 189.04 4055.025 326.985 ;
      RECT 4054.185 189.04 4054.465 326.745 ;
      RECT 4053.625 189.04 4053.905 326.505 ;
      RECT 4053.065 187.94 4053.345 326.265 ;
      RECT 4052.505 189.04 4052.785 326.025 ;
      RECT 4051.945 187.94 4052.225 325.785 ;
      RECT 4051.385 189.04 4051.665 325.545 ;
      RECT 4050.825 187.94 4051.105 325.305 ;
      RECT 4050.265 189.04 4050.545 325.065 ;
      RECT 4049.705 189.04 4049.985 324.825 ;
      RECT 4049.145 189.04 4049.425 324.585 ;
      RECT 4048.585 189.04 4048.865 324.345 ;
      RECT 4048.025 189.04 4048.305 324.105 ;
      RECT 4047.465 189.04 4047.745 323.865 ;
      RECT 4046.905 189.04 4047.185 323.625 ;
      RECT 4046.345 189.04 4046.625 323.385 ;
      RECT 4045.785 189.04 4046.065 323.145 ;
      RECT 4045.225 189.04 4045.505 322.905 ;
      RECT 4044.665 189.04 4044.945 322.665 ;
      RECT 4044.105 189.04 4044.385 322.425 ;
      RECT 4043.545 187.94 4043.825 322.185 ;
      RECT 4042.985 189.04 4043.265 321.945 ;
      RECT 4042.425 187.94 4042.705 321.705 ;
      RECT 4002.665 189.04 4002.945 332.175 ;
      RECT 4002.105 187.94 4002.385 332.415 ;
      RECT 4001.545 189.04 4001.825 332.655 ;
      RECT 4000.985 189.04 4001.265 332.895 ;
      RECT 4000.425 189.04 4000.705 333.135 ;
      RECT 3999.865 189.04 4000.145 333.375 ;
      RECT 3999.305 189.04 3999.585 333.615 ;
      RECT 3998.745 189.04 3999.025 333.86 ;
      RECT 3998.185 189.04 3998.465 334.1 ;
      RECT 3997.625 189.04 3997.905 334.34 ;
      RECT 3997.065 187.94 3997.345 334.58 ;
      RECT 3996.505 189.04 3996.785 334.82 ;
      RECT 3995.945 187.94 3996.225 335.06 ;
      RECT 3995.385 189.04 3995.665 335.3 ;
      RECT 3994.825 189.04 3995.105 335.54 ;
      RECT 3994.265 189.04 3994.545 335.78 ;
      RECT 3993.705 189.04 3993.985 336.02 ;
      RECT 3993.145 189.04 3993.425 336.26 ;
      RECT 3992.585 189.04 3992.865 336.5 ;
      RECT 3992.025 189.04 3992.305 336.74 ;
      RECT 3991.465 189.04 3991.745 336.98 ;
      RECT 3990.905 189.04 3991.185 337.22 ;
      RECT 3990.345 189.04 3990.625 337.46 ;
      RECT 3989.785 189.04 3990.065 337.7 ;
      RECT 3980.825 189.04 3981.105 333.285 ;
      RECT 3980.265 189.04 3980.545 333.045 ;
      RECT 3979.705 189.04 3979.985 332.805 ;
      RECT 3979.145 187.94 3979.425 332.565 ;
      RECT 3978.585 189.04 3978.865 332.325 ;
      RECT 3978.025 187.94 3978.305 332.085 ;
      RECT 3977.465 189.04 3977.745 331.845 ;
      RECT 3976.905 189.04 3977.185 331.605 ;
      RECT 3976.345 189.04 3976.625 331.365 ;
      RECT 3975.785 187.94 3976.065 331.125 ;
      RECT 3975.225 189.04 3975.505 330.885 ;
      RECT 3974.665 187.94 3974.945 330.645 ;
      RECT 3974.105 189.04 3974.385 330.405 ;
      RECT 3973.545 187.94 3973.825 330.165 ;
      RECT 3971.025 189.04 3971.305 322.565 ;
      RECT 3970.465 189.04 3970.745 322.325 ;
      RECT 3969.905 189.04 3970.185 322.085 ;
      RECT 3969.345 189.04 3969.625 321.845 ;
      RECT 3968.785 189.04 3969.065 321.605 ;
      RECT 3968.225 189.04 3968.505 321.365 ;
      RECT 3967.665 189.04 3967.945 321.125 ;
      RECT 3941.625 189.04 3941.905 335 ;
      RECT 3941.065 189.04 3941.345 335.24 ;
      RECT 3940.505 189.04 3940.785 335.48 ;
      RECT 3939.945 189.04 3940.225 335.72 ;
      RECT 3939.385 189.04 3939.665 335.96 ;
      RECT 3938.825 187.94 3939.105 335.96 ;
      RECT 3938.265 189.04 3938.545 335.72 ;
      RECT 3937.705 187.94 3937.985 335.475 ;
      RECT 3937.145 189.04 3937.425 335.235 ;
      RECT 3936.585 187.94 3936.865 334.995 ;
      RECT 3936.025 189.04 3936.305 334.755 ;
      RECT 3935.465 189.04 3935.745 334.515 ;
      RECT 3934.905 189.04 3935.185 334.275 ;
      RECT 3934.345 189.04 3934.625 334.035 ;
      RECT 3933.785 189.04 3934.065 333.795 ;
      RECT 3933.225 189.04 3933.505 333.555 ;
      RECT 3932.665 189.04 3932.945 333.315 ;
      RECT 3932.105 189.04 3932.385 333.075 ;
      RECT 3931.545 187.94 3931.825 332.835 ;
      RECT 3930.985 189.04 3931.265 332.595 ;
      RECT 3930.425 187.94 3930.705 332.355 ;
      RECT 3929.865 189.04 3930.145 332.115 ;
      RECT 3929.305 189.04 3929.585 331.875 ;
      RECT 3928.745 189.04 3929.025 331.635 ;
      RECT 3915.305 189.04 3915.585 335.035 ;
      RECT 3914.745 189.04 3915.025 335.275 ;
      RECT 3914.185 189.04 3914.465 335.52 ;
      RECT 3913.625 189.04 3913.905 335.76 ;
      RECT 3913.065 189.04 3913.345 336 ;
      RECT 3912.505 189.04 3912.785 336 ;
      RECT 3911.945 189.04 3912.225 335.76 ;
      RECT 3911.385 189.04 3911.665 335.52 ;
      RECT 3910.825 189.04 3911.105 328.505 ;
      RECT 3910.265 189.04 3910.545 328.265 ;
      RECT 3909.705 189.04 3909.985 328.025 ;
      RECT 3909.145 187.94 3909.425 327.785 ;
      RECT 3908.585 189.04 3908.865 327.545 ;
      RECT 3908.025 187.94 3908.305 327.305 ;
      RECT 3907.465 189.04 3907.745 327.065 ;
      RECT 3906.905 189.04 3907.185 326.825 ;
      RECT 3906.345 189.04 3906.625 326.585 ;
      RECT 3905.785 187.94 3906.065 326.345 ;
      RECT 3905.225 189.04 3905.505 326.105 ;
      RECT 3904.665 187.94 3904.945 325.865 ;
      RECT 3904.105 189.04 3904.385 325.625 ;
      RECT 3903.545 187.94 3903.825 325.385 ;
      RECT 3902.985 189.04 3903.265 325.145 ;
      RECT 3902.425 189.04 3902.705 324.905 ;
      RECT 3862.105 189.04 3862.385 333.8 ;
      RECT 3861.545 189.04 3861.825 334.04 ;
      RECT 3860.985 189.04 3861.265 334.285 ;
      RECT 3860.425 189.04 3860.705 334.525 ;
      RECT 3859.865 189.04 3860.145 334.765 ;
      RECT 3859.305 189.04 3859.585 335.005 ;
      RECT 3858.745 189.04 3859.025 335.245 ;
      RECT 3858.185 189.04 3858.465 335.485 ;
      RECT 3857.625 189.04 3857.905 335.725 ;
      RECT 3857.065 189.04 3857.345 335.965 ;
      RECT 3856.505 187.94 3856.785 336.205 ;
      RECT 3855.945 189.04 3856.225 336.445 ;
      RECT 3855.385 187.94 3855.665 336.685 ;
      RECT 3854.825 189.04 3855.105 336.925 ;
      RECT 3854.265 187.94 3854.545 337.165 ;
      RECT 3853.705 189.04 3853.985 337.165 ;
      RECT 3853.145 189.04 3853.425 336.925 ;
      RECT 3852.585 189.04 3852.865 336.685 ;
      RECT 3852.025 189.04 3852.305 336.445 ;
      RECT 3851.465 189.04 3851.745 336.205 ;
      RECT 3850.905 189.04 3851.185 335.965 ;
      RECT 3850.345 189.04 3850.625 335.725 ;
      RECT 3849.785 189.04 3850.065 335.485 ;
      RECT 3840.825 187.94 3841.105 335.515 ;
      RECT 3840.265 189.04 3840.545 335.755 ;
      RECT 3839.705 187.94 3839.985 335.995 ;
      RECT 3839.145 189.04 3839.425 336.21 ;
      RECT 3838.585 189.04 3838.865 335.785 ;
      RECT 3838.025 189.04 3838.305 335.545 ;
      RECT 3837.465 189.04 3837.745 335.305 ;
      RECT 3836.905 189.04 3837.185 335.065 ;
      RECT 3836.345 189.04 3836.625 334.825 ;
      RECT 3835.785 189.04 3836.065 334.585 ;
      RECT 3835.225 189.04 3835.505 334.345 ;
      RECT 3834.665 189.04 3834.945 334.105 ;
      RECT 3834.105 189.04 3834.385 333.865 ;
      RECT 3833.545 189.04 3833.825 333.625 ;
      RECT 3831.025 189.04 3831.305 332.8 ;
      RECT 3830.465 189.04 3830.745 332.56 ;
      RECT 3829.905 189.04 3830.185 332.32 ;
      RECT 3829.345 187.94 3829.625 332.08 ;
      RECT 3828.785 189.04 3829.065 331.84 ;
      RECT 3828.225 187.94 3828.505 331.6 ;
      RECT 3827.665 189.04 3827.945 331.36 ;
      RECT 3827.105 189.04 3827.385 331.12 ;
      RECT 3800.505 189.04 3800.785 342.165 ;
      RECT 3799.945 187.94 3800.225 342.405 ;
      RECT 3799.385 189.04 3799.665 342.645 ;
      RECT 3798.825 187.94 3799.105 342.89 ;
      RECT 3798.265 189.04 3798.545 343.13 ;
      RECT 3797.705 187.94 3797.985 343.37 ;
      RECT 3797.145 189.04 3797.425 343.61 ;
      RECT 3796.585 189.04 3796.865 343.85 ;
      RECT 3796.025 189.04 3796.305 329.47 ;
      RECT 3795.465 189.04 3795.745 329.23 ;
      RECT 3794.905 189.04 3795.185 328.99 ;
      RECT 3794.345 189.04 3794.625 328.75 ;
      RECT 3793.785 189.04 3794.065 328.51 ;
      RECT 3793.225 189.04 3793.505 328.27 ;
      RECT 3792.665 189.04 3792.945 328.03 ;
      RECT 3792.105 189.04 3792.385 327.79 ;
      RECT 3791.545 189.04 3791.825 327.55 ;
      RECT 3790.985 189.04 3791.265 327.31 ;
      RECT 3790.425 187.94 3790.705 327.07 ;
      RECT 3789.865 189.04 3790.145 326.83 ;
      RECT 3789.305 187.94 3789.585 326.59 ;
      RECT 3788.745 189.04 3789.025 326.35 ;
      RECT 3774.745 187.94 3775.025 332.47 ;
      RECT 3774.185 189.04 3774.465 332.23 ;
      RECT 3773.625 189.04 3773.905 331.99 ;
      RECT 3773.065 189.04 3773.345 331.75 ;
      RECT 3772.505 189.04 3772.785 331.51 ;
      RECT 3771.945 189.04 3772.225 331.27 ;
      RECT 3771.385 189.04 3771.665 331.03 ;
      RECT 3770.825 189.04 3771.105 330.79 ;
      RECT 3770.265 189.04 3770.545 330.55 ;
      RECT 3769.705 187.94 3769.985 330.31 ;
      RECT 3769.145 189.04 3769.425 330.07 ;
      RECT 3768.585 187.94 3768.865 329.83 ;
      RECT 3768.025 189.04 3768.305 329.59 ;
      RECT 3767.465 189.04 3767.745 329.35 ;
      RECT 3766.905 189.04 3767.185 329.11 ;
      RECT 3766.345 189.04 3766.625 328.87 ;
      RECT 3765.785 189.04 3766.065 328.63 ;
      RECT 3765.225 189.04 3765.505 328.39 ;
      RECT 3764.665 189.04 3764.945 328.15 ;
      RECT 3764.105 189.04 3764.385 327.91 ;
      RECT 3763.545 189.04 3763.825 327.67 ;
      RECT 3762.985 189.04 3763.265 327.43 ;
      RECT 3762.425 189.04 3762.705 327.19 ;
      RECT 3723.225 189.04 3723.505 334.095 ;
      RECT 3722.665 189.04 3722.945 334.335 ;
      RECT 3722.105 189.04 3722.385 334.575 ;
      RECT 3721.545 187.94 3721.825 334.815 ;
      RECT 3720.985 189.04 3721.265 335.055 ;
      RECT 3720.425 187.94 3720.705 335.295 ;
      RECT 3719.865 189.04 3720.145 335.535 ;
      RECT 3719.305 189.04 3719.585 335.775 ;
      RECT 3718.745 189.04 3719.025 336.015 ;
      RECT 3718.185 187.94 3718.465 336.255 ;
      RECT 3717.625 189.04 3717.905 336.495 ;
      RECT 3717.065 187.94 3717.345 336.735 ;
      RECT 3716.505 189.04 3716.785 336.975 ;
      RECT 3715.945 187.94 3716.225 337.215 ;
      RECT 3715.385 189.04 3715.665 337.455 ;
      RECT 3714.825 189.04 3715.105 337.695 ;
      RECT 3714.265 189.04 3714.545 337.695 ;
      RECT 3713.705 189.04 3713.985 337.455 ;
      RECT 3713.145 189.04 3713.425 337.215 ;
      RECT 3712.585 189.04 3712.865 336.975 ;
      RECT 3712.025 189.04 3712.305 336.735 ;
      RECT 3711.465 189.04 3711.745 336.495 ;
      RECT 3710.905 189.04 3711.185 336.255 ;
      RECT 3710.345 189.04 3710.625 336.015 ;
      RECT 3709.785 189.04 3710.065 335.775 ;
      RECT 3700.825 189.04 3701.105 335.29 ;
      RECT 3700.265 187.94 3700.545 335.05 ;
      RECT 3699.705 189.04 3699.985 334.81 ;
      RECT 3699.145 187.94 3699.425 334.57 ;
      RECT 3698.585 189.04 3698.865 334.33 ;
      RECT 3698.025 187.94 3698.305 334.09 ;
      RECT 3697.465 189.04 3697.745 333.85 ;
      RECT 3696.905 189.04 3697.185 333.61 ;
      RECT 3696.345 189.04 3696.625 333.37 ;
      RECT 3695.785 189.04 3696.065 333.13 ;
      RECT 3695.225 189.04 3695.505 332.89 ;
      RECT 3694.665 189.04 3694.945 332.65 ;
      RECT 3694.105 189.04 3694.385 332.41 ;
      RECT 3693.545 189.04 3693.825 332.17 ;
      RECT 3691.025 187.94 3691.305 333.89 ;
      RECT 3690.465 189.04 3690.745 333.65 ;
      RECT 3689.905 187.94 3690.185 333.41 ;
      RECT 3689.345 189.04 3689.625 333.17 ;
      RECT 3688.785 189.04 3689.065 332.93 ;
      RECT 3688.225 189.04 3688.505 332.69 ;
      RECT 3687.665 189.04 3687.945 332.45 ;
      RECT 3687.105 189.04 3687.385 332.21 ;
      RECT 3661.065 189.04 3661.345 329.86 ;
      RECT 3660.505 189.04 3660.785 330.1 ;
      RECT 3659.945 189.04 3660.225 330.34 ;
      RECT 3659.385 189.04 3659.665 330.585 ;
      RECT 3658.825 189.04 3659.105 330.825 ;
      RECT 3658.265 189.04 3658.545 331.065 ;
      RECT 3657.705 189.04 3657.985 331.065 ;
      RECT 3657.145 189.04 3657.425 330.825 ;
      RECT 3656.585 189.04 3656.865 330.585 ;
      RECT 3656.025 187.94 3656.305 330.345 ;
      RECT 3655.465 189.04 3655.745 330.105 ;
      RECT 3654.905 187.94 3655.185 329.865 ;
      RECT 3654.345 189.04 3654.625 329.625 ;
      RECT 3653.785 189.04 3654.065 329.385 ;
      RECT 3653.225 189.04 3653.505 329.145 ;
      RECT 3652.665 187.94 3652.945 328.905 ;
      RECT 3652.105 189.04 3652.385 328.665 ;
      RECT 3651.545 187.94 3651.825 328.425 ;
      RECT 3650.985 189.04 3651.265 328.185 ;
      RECT 3650.425 187.94 3650.705 327.945 ;
      RECT 3649.865 189.04 3650.145 327.705 ;
      RECT 3649.305 189.04 3649.585 327.465 ;
      RECT 3648.745 189.04 3649.025 327.225 ;
      RECT 3648.185 189.04 3648.465 326.985 ;
      RECT 3634.745 189.04 3635.025 332.785 ;
      RECT 3634.185 189.04 3634.465 332.545 ;
      RECT 3633.625 189.04 3633.905 332.305 ;
      RECT 3633.065 189.04 3633.345 332.065 ;
      RECT 3632.505 189.04 3632.785 331.825 ;
      RECT 3631.945 189.04 3632.225 331.585 ;
      RECT 3631.385 189.04 3631.665 331.345 ;
      RECT 3630.825 189.04 3631.105 331.105 ;
      RECT 3630.265 187.94 3630.545 330.865 ;
      RECT 3629.705 189.04 3629.985 330.625 ;
      RECT 3629.145 187.94 3629.425 330.305 ;
      RECT 3628.585 189.04 3628.865 330.145 ;
      RECT 3628.025 187.94 3628.305 329.905 ;
      RECT 3627.465 189.04 3627.745 329.665 ;
      RECT 3626.905 189.04 3627.185 329.425 ;
      RECT 3626.345 189.04 3626.625 329.185 ;
      RECT 3625.785 189.04 3626.065 328.945 ;
      RECT 3625.225 189.04 3625.505 328.705 ;
      RECT 3624.665 189.04 3624.945 328.465 ;
      RECT 3624.105 189.04 3624.385 328.225 ;
      RECT 3623.545 189.04 3623.825 327.985 ;
      RECT 3622.985 187.94 3623.265 327.745 ;
      RECT 3622.425 189.04 3622.705 327.505 ;
      RECT 3621.865 187.94 3622.145 327.265 ;
      RECT 3582.665 189.04 3582.945 332.875 ;
      RECT 3582.105 189.04 3582.385 333.115 ;
      RECT 3581.545 189.04 3581.825 333.355 ;
      RECT 3580.985 189.04 3581.265 333.595 ;
      RECT 3580.425 189.04 3580.705 333.835 ;
      RECT 3579.865 189.04 3580.145 334.075 ;
      RECT 3579.305 189.04 3579.585 334.315 ;
      RECT 3578.745 189.04 3579.025 334.555 ;
      RECT 3578.185 189.04 3578.465 334.795 ;
      RECT 3577.625 189.04 3577.905 335.035 ;
      RECT 3577.065 189.04 3577.345 335.275 ;
      RECT 3576.505 189.04 3576.785 335.515 ;
      RECT 3575.945 189.04 3576.225 335.755 ;
      RECT 3575.385 189.04 3575.665 335.755 ;
      RECT 3574.825 187.94 3575.105 335.515 ;
      RECT 3574.265 189.04 3574.545 335.275 ;
      RECT 3573.705 187.94 3573.985 335.035 ;
      RECT 3573.145 189.04 3573.425 334.795 ;
      RECT 3572.585 189.04 3572.865 334.555 ;
      RECT 3572.025 189.04 3572.305 334.315 ;
      RECT 3571.465 187.94 3571.745 334.05 ;
      RECT 3570.905 189.04 3571.185 333.81 ;
      RECT 3570.345 187.94 3570.625 333.57 ;
      RECT 3569.785 189.04 3570.065 333.33 ;
      RECT 3560.825 187.94 3561.105 327.165 ;
      RECT 3560.265 189.04 3560.545 327.405 ;
      RECT 3559.705 189.04 3559.985 327.645 ;
      RECT 3559.145 189.04 3559.425 327.645 ;
      RECT 3558.585 189.04 3558.865 327.405 ;
      RECT 3558.025 189.04 3558.305 327.165 ;
      RECT 3557.465 189.04 3557.745 326.925 ;
      RECT 3556.905 189.04 3557.185 326.685 ;
      RECT 3556.345 189.04 3556.625 326.445 ;
      RECT 3555.785 189.04 3556.065 326.205 ;
      RECT 3555.225 189.04 3555.505 325.965 ;
      RECT 3554.665 189.04 3554.945 325.725 ;
      RECT 3554.105 189.04 3554.385 325.485 ;
      RECT 3553.545 187.94 3553.825 325.245 ;
      RECT 3551.025 189.04 3551.305 326.965 ;
      RECT 3550.465 187.94 3550.745 326.725 ;
      RECT 3549.905 189.04 3550.185 326.485 ;
      RECT 3549.345 187.94 3549.625 326.245 ;
      RECT 3548.785 189.04 3549.065 326.005 ;
      RECT 3548.225 189.04 3548.505 325.765 ;
      RECT 3547.665 189.04 3547.945 325.525 ;
      RECT 3521.625 189.04 3521.905 328.31 ;
      RECT 3521.065 189.04 3521.345 328.55 ;
      RECT 3520.505 189.04 3520.785 328.79 ;
      RECT 3519.945 189.04 3520.225 329.03 ;
      RECT 3519.385 189.04 3519.665 329.27 ;
      RECT 3518.825 187.94 3519.105 329.51 ;
      RECT 3518.265 189.04 3518.545 329.75 ;
      RECT 3517.705 187.94 3517.985 329.99 ;
      RECT 3517.145 189.04 3517.425 330.23 ;
      RECT 3516.585 189.04 3516.865 330.47 ;
      RECT 3516.025 189.04 3516.305 330.71 ;
      RECT 3515.465 189.04 3515.745 330.95 ;
      RECT 3514.905 189.04 3515.185 331.19 ;
      RECT 3514.345 189.04 3514.625 331.43 ;
      RECT 3513.785 189.04 3514.065 331.67 ;
      RECT 3513.225 189.04 3513.505 331.67 ;
      RECT 3512.665 189.04 3512.945 331.43 ;
      RECT 3512.105 189.04 3512.385 331.19 ;
      RECT 3511.545 189.04 3511.825 330.95 ;
      RECT 3510.985 189.04 3511.265 330.705 ;
      RECT 3510.425 189.04 3510.705 330.465 ;
      RECT 3509.865 189.04 3510.145 330.225 ;
      RECT 3509.305 187.94 3509.585 329.985 ;
      RECT 3508.745 189.04 3509.025 329.745 ;
      RECT 3495.305 187.94 3495.585 327.225 ;
      RECT 3494.745 189.04 3495.025 326.985 ;
      RECT 3494.185 189.04 3494.465 326.745 ;
      RECT 3493.625 189.04 3493.905 326.505 ;
      RECT 3493.065 187.94 3493.345 326.265 ;
      RECT 3492.505 189.04 3492.785 326.025 ;
      RECT 3491.945 187.94 3492.225 325.785 ;
      RECT 3491.385 189.04 3491.665 325.545 ;
      RECT 3490.825 187.94 3491.105 325.305 ;
      RECT 3490.265 189.04 3490.545 325.065 ;
      RECT 3489.705 189.04 3489.985 324.825 ;
      RECT 3489.145 189.04 3489.425 324.585 ;
      RECT 3488.585 189.04 3488.865 324.345 ;
      RECT 3488.025 189.04 3488.305 324.105 ;
      RECT 3487.465 189.04 3487.745 323.865 ;
      RECT 3486.905 189.04 3487.185 323.625 ;
      RECT 3486.345 189.04 3486.625 323.385 ;
      RECT 3485.785 189.04 3486.065 323.145 ;
      RECT 3485.225 189.04 3485.505 322.905 ;
      RECT 3484.665 189.04 3484.945 322.665 ;
      RECT 3484.105 189.04 3484.385 322.425 ;
      RECT 3483.545 187.94 3483.825 322.185 ;
      RECT 3482.985 189.04 3483.265 321.945 ;
      RECT 3482.425 187.94 3482.705 321.705 ;
      RECT 3442.665 189.04 3442.945 332.175 ;
      RECT 3442.105 187.94 3442.385 332.415 ;
      RECT 3441.545 189.04 3441.825 332.655 ;
      RECT 3440.985 189.04 3441.265 332.895 ;
      RECT 3440.425 189.04 3440.705 333.135 ;
      RECT 3439.865 189.04 3440.145 333.375 ;
      RECT 3439.305 189.04 3439.585 333.615 ;
      RECT 3438.745 189.04 3439.025 333.86 ;
      RECT 3438.185 189.04 3438.465 334.1 ;
      RECT 3437.625 189.04 3437.905 334.34 ;
      RECT 3437.065 187.94 3437.345 334.58 ;
      RECT 3436.505 189.04 3436.785 334.82 ;
      RECT 3435.945 187.94 3436.225 335.06 ;
      RECT 3435.385 189.04 3435.665 335.3 ;
      RECT 3434.825 189.04 3435.105 335.54 ;
      RECT 3434.265 189.04 3434.545 335.78 ;
      RECT 3433.705 189.04 3433.985 336.02 ;
      RECT 3433.145 189.04 3433.425 336.26 ;
      RECT 3432.585 189.04 3432.865 336.5 ;
      RECT 3432.025 189.04 3432.305 336.74 ;
      RECT 3431.465 189.04 3431.745 336.98 ;
      RECT 3430.905 189.04 3431.185 337.22 ;
      RECT 3430.345 189.04 3430.625 337.46 ;
      RECT 3429.785 189.04 3430.065 337.7 ;
      RECT 3420.825 189.04 3421.105 333.285 ;
      RECT 3420.265 189.04 3420.545 333.045 ;
      RECT 3419.705 189.04 3419.985 332.805 ;
      RECT 3419.145 187.94 3419.425 332.565 ;
      RECT 3418.585 189.04 3418.865 332.325 ;
      RECT 3418.025 187.94 3418.305 332.085 ;
      RECT 3417.465 189.04 3417.745 331.845 ;
      RECT 3416.905 189.04 3417.185 331.605 ;
      RECT 3416.345 189.04 3416.625 331.365 ;
      RECT 3415.785 187.94 3416.065 331.125 ;
      RECT 3415.225 189.04 3415.505 330.885 ;
      RECT 3414.665 187.94 3414.945 330.645 ;
      RECT 3414.105 189.04 3414.385 330.405 ;
      RECT 3413.545 187.94 3413.825 330.165 ;
      RECT 3411.025 189.04 3411.305 322.565 ;
      RECT 3410.465 189.04 3410.745 322.325 ;
      RECT 3409.905 189.04 3410.185 322.085 ;
      RECT 3409.345 189.04 3409.625 321.845 ;
      RECT 3408.785 189.04 3409.065 321.605 ;
      RECT 3408.225 189.04 3408.505 321.365 ;
      RECT 3407.665 189.04 3407.945 321.125 ;
      RECT 3381.625 189.04 3381.905 335 ;
      RECT 3381.065 189.04 3381.345 335.24 ;
      RECT 3380.505 189.04 3380.785 335.48 ;
      RECT 3379.945 189.04 3380.225 335.72 ;
      RECT 3379.385 189.04 3379.665 335.96 ;
      RECT 3378.825 187.94 3379.105 335.96 ;
      RECT 3378.265 189.04 3378.545 335.72 ;
      RECT 3377.705 187.94 3377.985 335.475 ;
      RECT 3377.145 189.04 3377.425 335.235 ;
      RECT 3376.585 187.94 3376.865 334.995 ;
      RECT 3376.025 189.04 3376.305 334.755 ;
      RECT 3375.465 189.04 3375.745 334.515 ;
      RECT 3374.905 189.04 3375.185 334.275 ;
      RECT 3374.345 189.04 3374.625 334.035 ;
      RECT 3373.785 189.04 3374.065 333.795 ;
      RECT 3373.225 189.04 3373.505 333.555 ;
      RECT 3372.665 189.04 3372.945 333.315 ;
      RECT 3372.105 189.04 3372.385 333.075 ;
      RECT 3371.545 187.94 3371.825 332.835 ;
      RECT 3370.985 189.04 3371.265 332.595 ;
      RECT 3370.425 187.94 3370.705 332.355 ;
      RECT 3369.865 189.04 3370.145 332.115 ;
      RECT 3369.305 189.04 3369.585 331.875 ;
      RECT 3368.745 189.04 3369.025 331.635 ;
      RECT 3355.305 189.04 3355.585 335.035 ;
      RECT 3354.745 189.04 3355.025 335.275 ;
      RECT 3354.185 189.04 3354.465 335.52 ;
      RECT 3353.625 189.04 3353.905 335.76 ;
      RECT 3353.065 189.04 3353.345 336 ;
      RECT 3352.505 189.04 3352.785 336 ;
      RECT 3351.945 189.04 3352.225 335.76 ;
      RECT 3351.385 189.04 3351.665 335.52 ;
      RECT 3350.825 189.04 3351.105 328.505 ;
      RECT 3350.265 189.04 3350.545 328.265 ;
      RECT 3349.705 189.04 3349.985 328.025 ;
      RECT 3349.145 187.94 3349.425 327.785 ;
      RECT 3348.585 189.04 3348.865 327.545 ;
      RECT 3348.025 187.94 3348.305 327.305 ;
      RECT 3347.465 189.04 3347.745 327.065 ;
      RECT 3346.905 189.04 3347.185 326.825 ;
      RECT 3346.345 189.04 3346.625 326.585 ;
      RECT 3345.785 187.94 3346.065 326.345 ;
      RECT 3345.225 189.04 3345.505 326.105 ;
      RECT 3344.665 187.94 3344.945 325.865 ;
      RECT 3344.105 189.04 3344.385 325.625 ;
      RECT 3343.545 187.94 3343.825 325.385 ;
      RECT 3342.985 189.04 3343.265 325.145 ;
      RECT 3342.425 189.04 3342.705 324.905 ;
      RECT 3302.105 189.04 3302.385 333.8 ;
      RECT 3301.545 189.04 3301.825 334.04 ;
      RECT 3300.985 189.04 3301.265 334.285 ;
      RECT 3300.425 189.04 3300.705 334.525 ;
      RECT 3299.865 189.04 3300.145 334.765 ;
      RECT 3299.305 189.04 3299.585 335.005 ;
      RECT 3298.745 189.04 3299.025 335.245 ;
      RECT 3298.185 189.04 3298.465 335.485 ;
      RECT 3297.625 189.04 3297.905 335.725 ;
      RECT 3297.065 189.04 3297.345 335.965 ;
      RECT 3296.505 187.94 3296.785 336.205 ;
      RECT 3295.945 189.04 3296.225 336.445 ;
      RECT 3295.385 187.94 3295.665 336.685 ;
      RECT 3294.825 189.04 3295.105 336.925 ;
      RECT 3294.265 187.94 3294.545 337.165 ;
      RECT 3293.705 189.04 3293.985 337.165 ;
      RECT 3293.145 189.04 3293.425 336.925 ;
      RECT 3292.585 189.04 3292.865 336.685 ;
      RECT 3292.025 189.04 3292.305 336.445 ;
      RECT 3291.465 189.04 3291.745 336.205 ;
      RECT 3290.905 189.04 3291.185 335.965 ;
      RECT 3290.345 189.04 3290.625 335.725 ;
      RECT 3289.785 189.04 3290.065 335.485 ;
      RECT 3280.825 187.94 3281.105 335.515 ;
      RECT 3280.265 189.04 3280.545 335.755 ;
      RECT 3279.705 187.94 3279.985 335.995 ;
      RECT 3279.145 189.04 3279.425 336.21 ;
      RECT 3278.585 189.04 3278.865 335.785 ;
      RECT 3278.025 189.04 3278.305 335.545 ;
      RECT 3277.465 189.04 3277.745 335.305 ;
      RECT 3276.905 189.04 3277.185 335.065 ;
      RECT 3276.345 189.04 3276.625 334.825 ;
      RECT 3275.785 189.04 3276.065 334.585 ;
      RECT 3275.225 189.04 3275.505 334.345 ;
      RECT 3274.665 189.04 3274.945 334.105 ;
      RECT 3274.105 189.04 3274.385 333.865 ;
      RECT 3273.545 189.04 3273.825 333.625 ;
      RECT 3271.025 189.04 3271.305 332.8 ;
      RECT 3270.465 189.04 3270.745 332.56 ;
      RECT 3269.905 189.04 3270.185 332.32 ;
      RECT 3269.345 187.94 3269.625 332.08 ;
      RECT 3268.785 189.04 3269.065 331.84 ;
      RECT 3268.225 187.94 3268.505 331.6 ;
      RECT 3267.665 189.04 3267.945 331.36 ;
      RECT 3267.105 189.04 3267.385 331.12 ;
      RECT 3240.505 189.04 3240.785 342.165 ;
      RECT 3239.945 187.94 3240.225 342.405 ;
      RECT 3239.385 189.04 3239.665 342.645 ;
      RECT 3238.825 187.94 3239.105 342.89 ;
      RECT 3238.265 189.04 3238.545 343.13 ;
      RECT 3237.705 187.94 3237.985 343.37 ;
      RECT 3237.145 189.04 3237.425 343.61 ;
      RECT 3236.585 189.04 3236.865 343.85 ;
      RECT 3236.025 189.04 3236.305 329.47 ;
      RECT 3235.465 189.04 3235.745 329.23 ;
      RECT 3234.905 189.04 3235.185 328.99 ;
      RECT 3234.345 189.04 3234.625 328.75 ;
      RECT 3233.785 189.04 3234.065 328.51 ;
      RECT 3233.225 189.04 3233.505 328.27 ;
      RECT 3232.665 189.04 3232.945 328.03 ;
      RECT 3232.105 189.04 3232.385 327.79 ;
      RECT 3231.545 189.04 3231.825 327.55 ;
      RECT 3230.985 189.04 3231.265 327.31 ;
      RECT 3230.425 187.94 3230.705 327.07 ;
      RECT 3229.865 189.04 3230.145 326.83 ;
      RECT 3229.305 187.94 3229.585 326.59 ;
      RECT 3228.745 189.04 3229.025 326.35 ;
      RECT 3214.745 187.94 3215.025 332.47 ;
      RECT 3214.185 189.04 3214.465 332.23 ;
      RECT 3213.625 189.04 3213.905 331.99 ;
      RECT 3213.065 189.04 3213.345 331.75 ;
      RECT 3212.505 189.04 3212.785 331.51 ;
      RECT 3211.945 189.04 3212.225 331.27 ;
      RECT 3211.385 189.04 3211.665 331.03 ;
      RECT 3210.825 189.04 3211.105 330.79 ;
      RECT 3210.265 189.04 3210.545 330.55 ;
      RECT 3209.705 187.94 3209.985 330.31 ;
      RECT 3209.145 189.04 3209.425 330.07 ;
      RECT 3208.585 187.94 3208.865 329.83 ;
      RECT 3208.025 189.04 3208.305 329.59 ;
      RECT 3207.465 189.04 3207.745 329.35 ;
      RECT 3206.905 189.04 3207.185 329.11 ;
      RECT 3206.345 189.04 3206.625 328.87 ;
      RECT 3205.785 189.04 3206.065 328.63 ;
      RECT 3205.225 189.04 3205.505 328.39 ;
      RECT 3204.665 189.04 3204.945 328.15 ;
      RECT 3204.105 189.04 3204.385 327.91 ;
      RECT 3203.545 189.04 3203.825 327.67 ;
      RECT 3202.985 189.04 3203.265 327.43 ;
      RECT 3202.425 189.04 3202.705 327.19 ;
      RECT 3163.225 189.04 3163.505 334.095 ;
      RECT 3162.665 189.04 3162.945 334.335 ;
      RECT 3162.105 189.04 3162.385 334.575 ;
      RECT 3161.545 187.94 3161.825 334.815 ;
      RECT 3160.985 189.04 3161.265 335.055 ;
      RECT 3160.425 187.94 3160.705 335.295 ;
      RECT 3159.865 189.04 3160.145 335.535 ;
      RECT 3159.305 189.04 3159.585 335.775 ;
      RECT 3158.745 189.04 3159.025 336.015 ;
      RECT 3158.185 187.94 3158.465 336.255 ;
      RECT 3157.625 189.04 3157.905 336.495 ;
      RECT 3157.065 187.94 3157.345 336.735 ;
      RECT 3156.505 189.04 3156.785 336.975 ;
      RECT 3155.945 187.94 3156.225 337.215 ;
      RECT 3155.385 189.04 3155.665 337.455 ;
      RECT 3154.825 189.04 3155.105 337.695 ;
      RECT 3154.265 189.04 3154.545 337.695 ;
      RECT 3153.705 189.04 3153.985 337.455 ;
      RECT 3153.145 189.04 3153.425 337.215 ;
      RECT 3152.585 189.04 3152.865 336.975 ;
      RECT 3152.025 189.04 3152.305 336.735 ;
      RECT 3151.465 189.04 3151.745 336.495 ;
      RECT 3150.905 189.04 3151.185 336.255 ;
      RECT 3150.345 189.04 3150.625 336.015 ;
      RECT 3149.785 189.04 3150.065 335.775 ;
      RECT 3140.825 189.04 3141.105 335.29 ;
      RECT 3140.265 187.94 3140.545 335.05 ;
      RECT 3139.705 189.04 3139.985 334.81 ;
      RECT 3139.145 187.94 3139.425 334.57 ;
      RECT 3138.585 189.04 3138.865 334.33 ;
      RECT 3138.025 187.94 3138.305 334.09 ;
      RECT 3137.465 189.04 3137.745 333.85 ;
      RECT 3136.905 189.04 3137.185 333.61 ;
      RECT 3136.345 189.04 3136.625 333.37 ;
      RECT 3135.785 189.04 3136.065 333.13 ;
      RECT 3135.225 189.04 3135.505 332.89 ;
      RECT 3134.665 189.04 3134.945 332.65 ;
      RECT 3134.105 189.04 3134.385 332.41 ;
      RECT 3133.545 189.04 3133.825 332.17 ;
      RECT 3131.025 187.94 3131.305 333.89 ;
      RECT 3130.465 189.04 3130.745 333.65 ;
      RECT 3129.905 187.94 3130.185 333.41 ;
      RECT 3129.345 189.04 3129.625 333.17 ;
      RECT 3128.785 189.04 3129.065 332.93 ;
      RECT 3128.225 189.04 3128.505 332.69 ;
      RECT 3127.665 189.04 3127.945 332.45 ;
      RECT 3127.105 189.04 3127.385 332.21 ;
      RECT 3101.065 189.04 3101.345 329.86 ;
      RECT 3100.505 189.04 3100.785 330.1 ;
      RECT 3099.945 189.04 3100.225 330.34 ;
      RECT 3099.385 189.04 3099.665 330.585 ;
      RECT 3098.825 189.04 3099.105 330.825 ;
      RECT 3098.265 189.04 3098.545 331.065 ;
      RECT 3097.705 189.04 3097.985 331.065 ;
      RECT 3097.145 189.04 3097.425 330.825 ;
      RECT 3096.585 189.04 3096.865 330.585 ;
      RECT 3096.025 187.94 3096.305 330.345 ;
      RECT 3095.465 189.04 3095.745 330.105 ;
      RECT 3094.905 187.94 3095.185 329.865 ;
      RECT 3094.345 189.04 3094.625 329.625 ;
      RECT 3093.785 189.04 3094.065 329.385 ;
      RECT 3093.225 189.04 3093.505 329.145 ;
      RECT 3092.665 187.94 3092.945 328.905 ;
      RECT 3092.105 189.04 3092.385 328.665 ;
      RECT 3091.545 187.94 3091.825 328.425 ;
      RECT 3090.985 189.04 3091.265 328.185 ;
      RECT 3090.425 187.94 3090.705 327.945 ;
      RECT 3089.865 189.04 3090.145 327.705 ;
      RECT 3089.305 189.04 3089.585 327.465 ;
      RECT 3088.745 189.04 3089.025 327.225 ;
      RECT 3088.185 189.04 3088.465 326.985 ;
      RECT 3074.745 189.04 3075.025 332.785 ;
      RECT 3074.185 189.04 3074.465 332.545 ;
      RECT 3073.625 189.04 3073.905 332.305 ;
      RECT 3073.065 189.04 3073.345 332.065 ;
      RECT 3072.505 189.04 3072.785 331.825 ;
      RECT 3071.945 189.04 3072.225 331.585 ;
      RECT 3071.385 189.04 3071.665 331.345 ;
      RECT 3070.825 189.04 3071.105 331.105 ;
      RECT 3070.265 187.94 3070.545 330.865 ;
      RECT 3069.705 189.04 3069.985 330.625 ;
      RECT 3069.145 187.94 3069.425 330.305 ;
      RECT 3068.585 189.04 3068.865 330.145 ;
      RECT 3068.025 187.94 3068.305 329.905 ;
      RECT 3067.465 189.04 3067.745 329.665 ;
      RECT 3066.905 189.04 3067.185 329.425 ;
      RECT 3066.345 189.04 3066.625 329.185 ;
      RECT 3065.785 189.04 3066.065 328.945 ;
      RECT 3065.225 189.04 3065.505 328.705 ;
      RECT 3064.665 189.04 3064.945 328.465 ;
      RECT 3064.105 189.04 3064.385 328.225 ;
      RECT 3063.545 189.04 3063.825 327.985 ;
      RECT 3062.985 187.94 3063.265 327.745 ;
      RECT 3062.425 189.04 3062.705 327.505 ;
      RECT 3061.865 187.94 3062.145 327.265 ;
      RECT 3022.665 189.04 3022.945 332.875 ;
      RECT 3022.105 189.04 3022.385 333.115 ;
      RECT 3021.545 189.04 3021.825 333.355 ;
      RECT 3020.985 189.04 3021.265 333.595 ;
      RECT 3020.425 189.04 3020.705 333.835 ;
      RECT 3019.865 189.04 3020.145 334.075 ;
      RECT 3019.305 189.04 3019.585 334.315 ;
      RECT 3018.745 189.04 3019.025 334.555 ;
      RECT 3018.185 189.04 3018.465 334.795 ;
      RECT 3017.625 189.04 3017.905 335.035 ;
      RECT 3017.065 189.04 3017.345 335.275 ;
      RECT 3016.505 189.04 3016.785 335.515 ;
      RECT 3015.945 189.04 3016.225 335.755 ;
      RECT 3015.385 189.04 3015.665 335.755 ;
      RECT 3014.825 187.94 3015.105 335.515 ;
      RECT 3014.265 189.04 3014.545 335.275 ;
      RECT 3013.705 187.94 3013.985 335.035 ;
      RECT 3013.145 189.04 3013.425 334.795 ;
      RECT 3012.585 189.04 3012.865 334.555 ;
      RECT 3012.025 189.04 3012.305 334.315 ;
      RECT 3011.465 187.94 3011.745 334.05 ;
      RECT 3010.905 189.04 3011.185 333.81 ;
      RECT 3010.345 187.94 3010.625 333.57 ;
      RECT 3009.785 189.04 3010.065 333.33 ;
      RECT 3000.825 187.94 3001.105 327.165 ;
      RECT 3000.265 189.04 3000.545 327.405 ;
      RECT 2999.705 189.04 2999.985 327.645 ;
      RECT 2999.145 189.04 2999.425 327.645 ;
      RECT 2998.585 189.04 2998.865 327.405 ;
      RECT 2998.025 189.04 2998.305 327.165 ;
      RECT 2997.465 189.04 2997.745 326.925 ;
      RECT 2996.905 189.04 2997.185 326.685 ;
      RECT 2996.345 189.04 2996.625 326.445 ;
      RECT 2995.785 189.04 2996.065 326.205 ;
      RECT 2995.225 189.04 2995.505 325.965 ;
      RECT 2994.665 189.04 2994.945 325.725 ;
      RECT 2994.105 189.04 2994.385 325.485 ;
      RECT 2993.545 187.94 2993.825 325.245 ;
      RECT 2991.025 189.04 2991.305 326.965 ;
      RECT 2990.465 187.94 2990.745 326.725 ;
      RECT 2989.905 189.04 2990.185 326.485 ;
      RECT 2989.345 187.94 2989.625 326.245 ;
      RECT 2988.785 189.04 2989.065 326.005 ;
      RECT 2988.225 189.04 2988.505 325.765 ;
      RECT 2987.665 189.04 2987.945 325.525 ;
      RECT 2961.625 189.04 2961.905 328.31 ;
      RECT 2961.065 189.04 2961.345 328.55 ;
      RECT 2960.505 189.04 2960.785 328.79 ;
      RECT 2959.945 189.04 2960.225 329.03 ;
      RECT 2959.385 189.04 2959.665 329.27 ;
      RECT 2958.825 187.94 2959.105 329.51 ;
      RECT 2958.265 189.04 2958.545 329.75 ;
      RECT 2957.705 187.94 2957.985 329.99 ;
      RECT 2957.145 189.04 2957.425 330.23 ;
      RECT 2956.585 189.04 2956.865 330.47 ;
      RECT 2956.025 189.04 2956.305 330.71 ;
      RECT 2955.465 189.04 2955.745 330.95 ;
      RECT 2954.905 189.04 2955.185 331.19 ;
      RECT 2954.345 189.04 2954.625 331.43 ;
      RECT 2953.785 189.04 2954.065 331.67 ;
      RECT 2953.225 189.04 2953.505 331.67 ;
      RECT 2952.665 189.04 2952.945 331.43 ;
      RECT 2952.105 189.04 2952.385 331.19 ;
      RECT 2951.545 189.04 2951.825 330.95 ;
      RECT 2950.985 189.04 2951.265 330.705 ;
      RECT 2950.425 189.04 2950.705 330.465 ;
      RECT 2949.865 189.04 2950.145 330.225 ;
      RECT 2949.305 187.94 2949.585 329.985 ;
      RECT 2948.745 189.04 2949.025 329.745 ;
      RECT 2935.305 187.94 2935.585 327.225 ;
      RECT 2934.745 189.04 2935.025 326.985 ;
      RECT 2934.185 189.04 2934.465 326.745 ;
      RECT 2933.625 189.04 2933.905 326.505 ;
      RECT 2933.065 187.94 2933.345 326.265 ;
      RECT 2932.505 189.04 2932.785 326.025 ;
      RECT 2931.945 187.94 2932.225 325.785 ;
      RECT 2931.385 189.04 2931.665 325.545 ;
      RECT 2930.825 187.94 2931.105 325.305 ;
      RECT 2930.265 189.04 2930.545 325.065 ;
      RECT 2929.705 189.04 2929.985 324.825 ;
      RECT 2929.145 189.04 2929.425 324.585 ;
      RECT 2928.585 189.04 2928.865 324.345 ;
      RECT 2928.025 189.04 2928.305 324.105 ;
      RECT 2927.465 189.04 2927.745 323.865 ;
      RECT 2926.905 189.04 2927.185 323.625 ;
      RECT 2926.345 189.04 2926.625 323.385 ;
      RECT 2925.785 189.04 2926.065 323.145 ;
      RECT 2925.225 189.04 2925.505 322.905 ;
      RECT 2924.665 189.04 2924.945 322.665 ;
      RECT 2924.105 189.04 2924.385 322.425 ;
      RECT 2923.545 187.94 2923.825 322.185 ;
      RECT 2922.985 189.04 2923.265 321.945 ;
      RECT 2922.425 187.94 2922.705 321.705 ;
      RECT 2882.665 189.04 2882.945 332.175 ;
      RECT 2882.105 187.94 2882.385 332.415 ;
      RECT 2881.545 189.04 2881.825 332.655 ;
      RECT 2880.985 189.04 2881.265 332.895 ;
      RECT 2880.425 189.04 2880.705 333.135 ;
      RECT 2879.865 189.04 2880.145 333.375 ;
      RECT 2879.305 189.04 2879.585 333.615 ;
      RECT 2878.745 189.04 2879.025 333.86 ;
      RECT 2878.185 189.04 2878.465 334.1 ;
      RECT 2877.625 189.04 2877.905 334.34 ;
      RECT 2877.065 187.94 2877.345 334.58 ;
      RECT 2876.505 189.04 2876.785 334.82 ;
      RECT 2875.945 187.94 2876.225 335.06 ;
      RECT 2875.385 189.04 2875.665 335.3 ;
      RECT 2874.825 189.04 2875.105 335.54 ;
      RECT 2874.265 189.04 2874.545 335.78 ;
      RECT 2873.705 189.04 2873.985 336.02 ;
      RECT 2873.145 189.04 2873.425 336.26 ;
      RECT 2872.585 189.04 2872.865 336.5 ;
      RECT 2872.025 189.04 2872.305 336.74 ;
      RECT 2871.465 189.04 2871.745 336.98 ;
      RECT 2870.905 189.04 2871.185 337.22 ;
      RECT 2870.345 189.04 2870.625 337.46 ;
      RECT 2869.785 189.04 2870.065 337.7 ;
      RECT 2860.825 189.04 2861.105 333.285 ;
      RECT 2860.265 189.04 2860.545 333.045 ;
      RECT 2859.705 189.04 2859.985 332.805 ;
      RECT 2859.145 187.94 2859.425 332.565 ;
      RECT 2858.585 189.04 2858.865 332.325 ;
      RECT 2858.025 187.94 2858.305 332.085 ;
      RECT 2857.465 189.04 2857.745 331.845 ;
      RECT 2856.905 189.04 2857.185 331.605 ;
      RECT 2856.345 189.04 2856.625 331.365 ;
      RECT 2855.785 187.94 2856.065 331.125 ;
      RECT 2855.225 189.04 2855.505 330.885 ;
      RECT 2854.665 187.94 2854.945 330.645 ;
      RECT 2854.105 189.04 2854.385 330.405 ;
      RECT 2853.545 187.94 2853.825 330.165 ;
      RECT 2851.025 189.04 2851.305 322.565 ;
      RECT 2850.465 189.04 2850.745 322.325 ;
      RECT 2849.905 189.04 2850.185 322.085 ;
      RECT 2849.345 189.04 2849.625 321.845 ;
      RECT 2848.785 189.04 2849.065 321.605 ;
      RECT 2848.225 189.04 2848.505 321.365 ;
      RECT 2847.665 189.04 2847.945 321.125 ;
      RECT 2821.625 189.04 2821.905 335 ;
      RECT 2821.065 189.04 2821.345 335.24 ;
      RECT 2820.505 189.04 2820.785 335.48 ;
      RECT 2819.945 189.04 2820.225 335.72 ;
      RECT 2819.385 189.04 2819.665 335.96 ;
      RECT 2818.825 187.94 2819.105 335.96 ;
      RECT 2818.265 189.04 2818.545 335.72 ;
      RECT 2817.705 187.94 2817.985 335.475 ;
      RECT 2817.145 189.04 2817.425 335.235 ;
      RECT 2816.585 187.94 2816.865 334.995 ;
      RECT 2816.025 189.04 2816.305 334.755 ;
      RECT 2815.465 189.04 2815.745 334.515 ;
      RECT 2814.905 189.04 2815.185 334.275 ;
      RECT 2814.345 189.04 2814.625 334.035 ;
      RECT 2813.785 189.04 2814.065 333.795 ;
      RECT 2813.225 189.04 2813.505 333.555 ;
      RECT 2812.665 189.04 2812.945 333.315 ;
      RECT 2812.105 189.04 2812.385 333.075 ;
      RECT 2811.545 187.94 2811.825 332.835 ;
      RECT 2810.985 189.04 2811.265 332.595 ;
      RECT 2810.425 187.94 2810.705 332.355 ;
      RECT 2809.865 189.04 2810.145 332.115 ;
      RECT 2809.305 189.04 2809.585 331.875 ;
      RECT 2808.745 189.04 2809.025 331.635 ;
      RECT 2795.305 189.04 2795.585 335.035 ;
      RECT 2794.745 189.04 2795.025 335.275 ;
      RECT 2794.185 189.04 2794.465 335.52 ;
      RECT 2793.625 189.04 2793.905 335.76 ;
      RECT 2793.065 189.04 2793.345 336 ;
      RECT 2792.505 189.04 2792.785 336 ;
      RECT 2791.945 189.04 2792.225 335.76 ;
      RECT 2791.385 189.04 2791.665 335.52 ;
      RECT 2790.825 189.04 2791.105 328.505 ;
      RECT 2790.265 189.04 2790.545 328.265 ;
      RECT 2789.705 189.04 2789.985 328.025 ;
      RECT 2789.145 187.94 2789.425 327.785 ;
      RECT 2788.585 189.04 2788.865 327.545 ;
      RECT 2788.025 187.94 2788.305 327.305 ;
      RECT 2787.465 189.04 2787.745 327.065 ;
      RECT 2786.905 189.04 2787.185 326.825 ;
      RECT 2786.345 189.04 2786.625 326.585 ;
      RECT 2785.785 187.94 2786.065 326.345 ;
      RECT 2785.225 189.04 2785.505 326.105 ;
      RECT 2784.665 187.94 2784.945 325.865 ;
      RECT 2784.105 189.04 2784.385 325.625 ;
      RECT 2783.545 187.94 2783.825 325.385 ;
      RECT 2782.985 189.04 2783.265 325.145 ;
      RECT 2782.425 189.04 2782.705 324.905 ;
      RECT 2742.105 189.04 2742.385 333.8 ;
      RECT 2741.545 189.04 2741.825 334.04 ;
      RECT 2740.985 189.04 2741.265 334.285 ;
      RECT 2740.425 189.04 2740.705 334.525 ;
      RECT 2739.865 189.04 2740.145 334.765 ;
      RECT 2739.305 189.04 2739.585 335.005 ;
      RECT 2738.745 189.04 2739.025 335.245 ;
      RECT 2738.185 189.04 2738.465 335.485 ;
      RECT 2737.625 189.04 2737.905 335.725 ;
      RECT 2737.065 189.04 2737.345 335.965 ;
      RECT 2736.505 187.94 2736.785 336.205 ;
      RECT 2735.945 189.04 2736.225 336.445 ;
      RECT 2735.385 187.94 2735.665 336.685 ;
      RECT 2734.825 189.04 2735.105 336.925 ;
      RECT 2734.265 187.94 2734.545 337.165 ;
      RECT 2733.705 189.04 2733.985 337.165 ;
      RECT 2733.145 189.04 2733.425 336.925 ;
      RECT 2732.585 189.04 2732.865 336.685 ;
      RECT 2732.025 189.04 2732.305 336.445 ;
      RECT 2731.465 189.04 2731.745 336.205 ;
      RECT 2730.905 189.04 2731.185 335.965 ;
      RECT 2730.345 189.04 2730.625 335.725 ;
      RECT 2729.785 189.04 2730.065 335.485 ;
      RECT 2720.825 187.94 2721.105 335.515 ;
      RECT 2720.265 189.04 2720.545 335.755 ;
      RECT 2719.705 187.94 2719.985 335.995 ;
      RECT 2719.145 189.04 2719.425 336.21 ;
      RECT 2718.585 189.04 2718.865 335.785 ;
      RECT 2718.025 189.04 2718.305 335.545 ;
      RECT 2717.465 189.04 2717.745 335.305 ;
      RECT 2716.905 189.04 2717.185 335.065 ;
      RECT 2716.345 189.04 2716.625 334.825 ;
      RECT 2715.785 189.04 2716.065 334.585 ;
      RECT 2715.225 189.04 2715.505 334.345 ;
      RECT 2714.665 189.04 2714.945 334.105 ;
      RECT 2714.105 189.04 2714.385 333.865 ;
      RECT 2713.545 189.04 2713.825 333.625 ;
      RECT 2711.025 189.04 2711.305 332.8 ;
      RECT 2710.465 189.04 2710.745 332.56 ;
      RECT 2709.905 189.04 2710.185 332.32 ;
      RECT 2709.345 187.94 2709.625 332.08 ;
      RECT 2708.785 189.04 2709.065 331.84 ;
      RECT 2708.225 187.94 2708.505 331.6 ;
      RECT 2707.665 189.04 2707.945 331.36 ;
      RECT 2707.105 189.04 2707.385 331.12 ;
      RECT 2680.505 189.04 2680.785 342.165 ;
      RECT 2679.945 187.94 2680.225 342.405 ;
      RECT 2679.385 189.04 2679.665 342.645 ;
      RECT 2678.825 187.94 2679.105 342.89 ;
      RECT 2678.265 189.04 2678.545 343.13 ;
      RECT 2677.705 187.94 2677.985 343.37 ;
      RECT 2677.145 189.04 2677.425 343.61 ;
      RECT 2676.585 189.04 2676.865 343.85 ;
      RECT 2676.025 189.04 2676.305 329.47 ;
      RECT 2675.465 189.04 2675.745 329.23 ;
      RECT 2674.905 189.04 2675.185 328.99 ;
      RECT 2674.345 189.04 2674.625 328.75 ;
      RECT 2673.785 189.04 2674.065 328.51 ;
      RECT 2673.225 189.04 2673.505 328.27 ;
      RECT 2672.665 189.04 2672.945 328.03 ;
      RECT 2672.105 189.04 2672.385 327.79 ;
      RECT 2671.545 189.04 2671.825 327.55 ;
      RECT 2670.985 189.04 2671.265 327.31 ;
      RECT 2670.425 187.94 2670.705 327.07 ;
      RECT 2669.865 189.04 2670.145 326.83 ;
      RECT 2669.305 187.94 2669.585 326.59 ;
      RECT 2668.745 189.04 2669.025 326.35 ;
      RECT 2654.745 187.94 2655.025 332.47 ;
      RECT 2654.185 189.04 2654.465 332.23 ;
      RECT 2653.625 189.04 2653.905 331.99 ;
      RECT 2653.065 189.04 2653.345 331.75 ;
      RECT 2652.505 189.04 2652.785 331.51 ;
      RECT 2651.945 189.04 2652.225 331.27 ;
      RECT 2651.385 189.04 2651.665 331.03 ;
      RECT 2650.825 189.04 2651.105 330.79 ;
      RECT 2650.265 189.04 2650.545 330.55 ;
      RECT 2649.705 187.94 2649.985 330.31 ;
      RECT 2649.145 189.04 2649.425 330.07 ;
      RECT 2648.585 187.94 2648.865 329.83 ;
      RECT 2648.025 189.04 2648.305 329.59 ;
      RECT 2647.465 189.04 2647.745 329.35 ;
      RECT 2646.905 189.04 2647.185 329.11 ;
      RECT 2646.345 189.04 2646.625 328.87 ;
      RECT 2645.785 189.04 2646.065 328.63 ;
      RECT 2645.225 189.04 2645.505 328.39 ;
      RECT 2644.665 189.04 2644.945 328.15 ;
      RECT 2644.105 189.04 2644.385 327.91 ;
      RECT 2643.545 189.04 2643.825 327.67 ;
      RECT 2642.985 189.04 2643.265 327.43 ;
      RECT 2642.425 189.04 2642.705 327.19 ;
      RECT 2603.225 189.04 2603.505 334.095 ;
      RECT 2602.665 189.04 2602.945 334.335 ;
      RECT 2602.105 189.04 2602.385 334.575 ;
      RECT 2601.545 187.94 2601.825 334.815 ;
      RECT 2600.985 189.04 2601.265 335.055 ;
      RECT 2600.425 187.94 2600.705 335.295 ;
      RECT 2599.865 189.04 2600.145 335.535 ;
      RECT 2599.305 189.04 2599.585 335.775 ;
      RECT 2598.745 189.04 2599.025 336.015 ;
      RECT 2598.185 187.94 2598.465 336.255 ;
      RECT 2597.625 189.04 2597.905 336.495 ;
      RECT 2597.065 187.94 2597.345 336.735 ;
      RECT 2596.505 189.04 2596.785 336.975 ;
      RECT 2595.945 187.94 2596.225 337.215 ;
      RECT 2595.385 189.04 2595.665 337.455 ;
      RECT 2594.825 189.04 2595.105 337.695 ;
      RECT 2594.265 189.04 2594.545 337.695 ;
      RECT 2593.705 189.04 2593.985 337.455 ;
      RECT 2593.145 189.04 2593.425 337.215 ;
      RECT 2592.585 189.04 2592.865 336.975 ;
      RECT 2592.025 189.04 2592.305 336.735 ;
      RECT 2591.465 189.04 2591.745 336.495 ;
      RECT 2590.905 189.04 2591.185 336.255 ;
      RECT 2590.345 189.04 2590.625 336.015 ;
      RECT 2589.785 189.04 2590.065 335.775 ;
      RECT 2580.825 189.04 2581.105 335.29 ;
      RECT 2580.265 187.94 2580.545 335.05 ;
      RECT 2579.705 189.04 2579.985 334.81 ;
      RECT 2579.145 187.94 2579.425 334.57 ;
      RECT 2578.585 189.04 2578.865 334.33 ;
      RECT 2578.025 187.94 2578.305 334.09 ;
      RECT 2577.465 189.04 2577.745 333.85 ;
      RECT 2576.905 189.04 2577.185 333.61 ;
      RECT 2576.345 189.04 2576.625 333.37 ;
      RECT 2575.785 189.04 2576.065 333.13 ;
      RECT 2575.225 189.04 2575.505 332.89 ;
      RECT 2574.665 189.04 2574.945 332.65 ;
      RECT 2574.105 189.04 2574.385 332.41 ;
      RECT 2573.545 189.04 2573.825 332.17 ;
      RECT 2571.025 187.94 2571.305 333.89 ;
      RECT 2570.465 189.04 2570.745 333.65 ;
      RECT 2569.905 187.94 2570.185 333.41 ;
      RECT 2569.345 189.04 2569.625 333.17 ;
      RECT 2568.785 189.04 2569.065 332.93 ;
      RECT 2568.225 189.04 2568.505 332.69 ;
      RECT 2567.665 189.04 2567.945 332.45 ;
      RECT 2567.105 189.04 2567.385 332.21 ;
      RECT 2541.065 189.04 2541.345 329.86 ;
      RECT 2540.505 189.04 2540.785 330.1 ;
      RECT 2539.945 189.04 2540.225 330.34 ;
      RECT 2539.385 189.04 2539.665 330.585 ;
      RECT 2538.825 189.04 2539.105 330.825 ;
      RECT 2538.265 189.04 2538.545 331.065 ;
      RECT 2537.705 189.04 2537.985 331.065 ;
      RECT 2537.145 189.04 2537.425 330.825 ;
      RECT 2536.585 189.04 2536.865 330.585 ;
      RECT 2536.025 187.94 2536.305 330.345 ;
      RECT 2535.465 189.04 2535.745 330.105 ;
      RECT 2534.905 187.94 2535.185 329.865 ;
      RECT 2534.345 189.04 2534.625 329.625 ;
      RECT 2533.785 189.04 2534.065 329.385 ;
      RECT 2533.225 189.04 2533.505 329.145 ;
      RECT 2532.665 187.94 2532.945 328.905 ;
      RECT 2532.105 189.04 2532.385 328.665 ;
      RECT 2531.545 187.94 2531.825 328.425 ;
      RECT 2530.985 189.04 2531.265 328.185 ;
      RECT 2530.425 187.94 2530.705 327.945 ;
      RECT 2529.865 189.04 2530.145 327.705 ;
      RECT 2529.305 189.04 2529.585 327.465 ;
      RECT 2528.745 189.04 2529.025 327.225 ;
      RECT 2528.185 189.04 2528.465 326.985 ;
      RECT 2514.745 189.04 2515.025 332.785 ;
      RECT 2514.185 189.04 2514.465 332.545 ;
      RECT 2513.625 189.04 2513.905 332.305 ;
      RECT 2513.065 189.04 2513.345 332.065 ;
      RECT 2512.505 189.04 2512.785 331.825 ;
      RECT 2511.945 189.04 2512.225 331.585 ;
      RECT 2511.385 189.04 2511.665 331.345 ;
      RECT 2510.825 189.04 2511.105 331.105 ;
      RECT 2510.265 187.94 2510.545 330.865 ;
      RECT 2509.705 189.04 2509.985 330.625 ;
      RECT 2509.145 187.94 2509.425 330.305 ;
      RECT 2508.585 189.04 2508.865 330.145 ;
      RECT 2508.025 187.94 2508.305 329.905 ;
      RECT 2507.465 189.04 2507.745 329.665 ;
      RECT 2506.905 189.04 2507.185 329.425 ;
      RECT 2506.345 189.04 2506.625 329.185 ;
      RECT 2505.785 189.04 2506.065 328.945 ;
      RECT 2505.225 189.04 2505.505 328.705 ;
      RECT 2504.665 189.04 2504.945 328.465 ;
      RECT 2504.105 189.04 2504.385 328.225 ;
      RECT 2503.545 189.04 2503.825 327.985 ;
      RECT 2502.985 187.94 2503.265 327.745 ;
      RECT 2502.425 189.04 2502.705 327.505 ;
      RECT 2501.865 187.94 2502.145 327.265 ;
      RECT 2462.665 189.04 2462.945 332.875 ;
      RECT 2462.105 189.04 2462.385 333.115 ;
      RECT 2461.545 189.04 2461.825 333.355 ;
      RECT 2460.985 189.04 2461.265 333.595 ;
      RECT 2460.425 189.04 2460.705 333.835 ;
      RECT 2459.865 189.04 2460.145 334.075 ;
      RECT 2459.305 189.04 2459.585 334.315 ;
      RECT 2458.745 189.04 2459.025 334.555 ;
      RECT 2458.185 189.04 2458.465 334.795 ;
      RECT 2457.625 189.04 2457.905 335.035 ;
      RECT 2457.065 189.04 2457.345 335.275 ;
      RECT 2456.505 189.04 2456.785 335.515 ;
      RECT 2455.945 189.04 2456.225 335.755 ;
      RECT 2455.385 189.04 2455.665 335.755 ;
      RECT 2454.825 187.94 2455.105 335.515 ;
      RECT 2454.265 189.04 2454.545 335.275 ;
      RECT 2453.705 187.94 2453.985 335.035 ;
      RECT 2453.145 189.04 2453.425 334.795 ;
      RECT 2452.585 189.04 2452.865 334.555 ;
      RECT 2452.025 189.04 2452.305 334.315 ;
      RECT 2451.465 187.94 2451.745 334.05 ;
      RECT 2450.905 189.04 2451.185 333.81 ;
      RECT 2450.345 187.94 2450.625 333.57 ;
      RECT 2449.785 189.04 2450.065 333.33 ;
      RECT 2440.825 187.94 2441.105 327.165 ;
      RECT 2440.265 189.04 2440.545 327.405 ;
      RECT 2439.705 189.04 2439.985 327.645 ;
      RECT 2439.145 189.04 2439.425 327.645 ;
      RECT 2438.585 189.04 2438.865 327.405 ;
      RECT 2438.025 189.04 2438.305 327.165 ;
      RECT 2437.465 189.04 2437.745 326.925 ;
      RECT 2436.905 189.04 2437.185 326.685 ;
      RECT 2436.345 189.04 2436.625 326.445 ;
      RECT 2435.785 189.04 2436.065 326.205 ;
      RECT 2435.225 189.04 2435.505 325.965 ;
      RECT 2434.665 189.04 2434.945 325.725 ;
      RECT 2434.105 189.04 2434.385 325.485 ;
      RECT 2433.545 187.94 2433.825 325.245 ;
      RECT 2431.025 189.04 2431.305 326.965 ;
      RECT 2430.465 187.94 2430.745 326.725 ;
      RECT 2429.905 189.04 2430.185 326.485 ;
      RECT 2429.345 187.94 2429.625 326.245 ;
      RECT 2428.785 189.04 2429.065 326.005 ;
      RECT 2428.225 189.04 2428.505 325.765 ;
      RECT 2427.665 189.04 2427.945 325.525 ;
      RECT 2401.625 189.04 2401.905 328.31 ;
      RECT 2401.065 189.04 2401.345 328.55 ;
      RECT 2400.505 189.04 2400.785 328.79 ;
      RECT 2399.945 189.04 2400.225 329.03 ;
      RECT 2399.385 189.04 2399.665 329.27 ;
      RECT 2398.825 187.94 2399.105 329.51 ;
      RECT 2398.265 189.04 2398.545 329.75 ;
      RECT 2397.705 187.94 2397.985 329.99 ;
      RECT 2397.145 189.04 2397.425 330.23 ;
      RECT 2396.585 189.04 2396.865 330.47 ;
      RECT 2396.025 189.04 2396.305 330.71 ;
      RECT 2395.465 189.04 2395.745 330.95 ;
      RECT 2394.905 189.04 2395.185 331.19 ;
      RECT 2394.345 189.04 2394.625 331.43 ;
      RECT 2393.785 189.04 2394.065 331.67 ;
      RECT 2393.225 189.04 2393.505 331.67 ;
      RECT 2392.665 189.04 2392.945 331.43 ;
      RECT 2392.105 189.04 2392.385 331.19 ;
      RECT 2391.545 189.04 2391.825 330.95 ;
      RECT 2390.985 189.04 2391.265 330.705 ;
      RECT 2390.425 189.04 2390.705 330.465 ;
      RECT 2389.865 189.04 2390.145 330.225 ;
      RECT 2389.305 187.94 2389.585 329.985 ;
      RECT 2388.745 189.04 2389.025 329.745 ;
      RECT 2375.305 187.94 2375.585 327.225 ;
      RECT 2374.745 189.04 2375.025 326.985 ;
      RECT 2374.185 189.04 2374.465 326.745 ;
      RECT 2373.625 189.04 2373.905 326.505 ;
      RECT 2373.065 187.94 2373.345 326.265 ;
      RECT 2372.505 189.04 2372.785 326.025 ;
      RECT 2371.945 187.94 2372.225 325.785 ;
      RECT 2371.385 189.04 2371.665 325.545 ;
      RECT 2370.825 187.94 2371.105 325.305 ;
      RECT 2370.265 189.04 2370.545 325.065 ;
      RECT 2369.705 189.04 2369.985 324.825 ;
      RECT 2369.145 189.04 2369.425 324.585 ;
      RECT 2368.585 189.04 2368.865 324.345 ;
      RECT 2368.025 189.04 2368.305 324.105 ;
      RECT 2367.465 189.04 2367.745 323.865 ;
      RECT 2366.905 189.04 2367.185 323.625 ;
      RECT 2366.345 189.04 2366.625 323.385 ;
      RECT 2365.785 189.04 2366.065 323.145 ;
      RECT 2365.225 189.04 2365.505 322.905 ;
      RECT 2364.665 189.04 2364.945 322.665 ;
      RECT 2364.105 189.04 2364.385 322.425 ;
      RECT 2363.545 187.94 2363.825 322.185 ;
      RECT 2362.985 189.04 2363.265 321.945 ;
      RECT 2362.425 187.94 2362.705 321.705 ;
      RECT 2322.665 189.04 2322.945 332.175 ;
      RECT 2322.105 187.94 2322.385 332.415 ;
      RECT 2321.545 189.04 2321.825 332.655 ;
      RECT 2320.985 189.04 2321.265 332.895 ;
      RECT 2320.425 189.04 2320.705 333.135 ;
      RECT 2319.865 189.04 2320.145 333.375 ;
      RECT 2319.305 189.04 2319.585 333.615 ;
      RECT 2318.745 189.04 2319.025 333.86 ;
      RECT 2318.185 189.04 2318.465 334.1 ;
      RECT 2317.625 189.04 2317.905 334.34 ;
      RECT 2317.065 187.94 2317.345 334.58 ;
      RECT 2316.505 189.04 2316.785 334.82 ;
      RECT 2315.945 187.94 2316.225 335.06 ;
      RECT 2315.385 189.04 2315.665 335.3 ;
      RECT 2314.825 189.04 2315.105 335.54 ;
      RECT 2314.265 189.04 2314.545 335.78 ;
      RECT 2313.705 189.04 2313.985 336.02 ;
      RECT 2313.145 189.04 2313.425 336.26 ;
      RECT 2312.585 189.04 2312.865 336.5 ;
      RECT 2312.025 189.04 2312.305 336.74 ;
      RECT 2311.465 189.04 2311.745 336.98 ;
      RECT 2310.905 189.04 2311.185 337.22 ;
      RECT 2310.345 189.04 2310.625 337.46 ;
      RECT 2309.785 189.04 2310.065 337.7 ;
      RECT 2300.825 189.04 2301.105 333.285 ;
      RECT 2300.265 189.04 2300.545 333.045 ;
      RECT 2299.705 189.04 2299.985 332.805 ;
      RECT 2299.145 187.94 2299.425 332.565 ;
      RECT 2298.585 189.04 2298.865 332.325 ;
      RECT 2298.025 187.94 2298.305 332.085 ;
      RECT 2297.465 189.04 2297.745 331.845 ;
      RECT 2296.905 189.04 2297.185 331.605 ;
      RECT 2296.345 189.04 2296.625 331.365 ;
      RECT 2295.785 187.94 2296.065 331.125 ;
      RECT 2295.225 189.04 2295.505 330.885 ;
      RECT 2294.665 187.94 2294.945 330.645 ;
      RECT 2294.105 189.04 2294.385 330.405 ;
      RECT 2293.545 187.94 2293.825 330.165 ;
      RECT 2291.025 189.04 2291.305 322.565 ;
      RECT 2290.465 189.04 2290.745 322.325 ;
      RECT 2289.905 189.04 2290.185 322.085 ;
      RECT 2289.345 189.04 2289.625 321.845 ;
      RECT 2288.785 189.04 2289.065 321.605 ;
      RECT 2288.225 189.04 2288.505 321.365 ;
      RECT 2287.665 189.04 2287.945 321.125 ;
      RECT 2261.625 189.04 2261.905 335 ;
      RECT 2261.065 189.04 2261.345 335.24 ;
      RECT 2260.505 189.04 2260.785 335.48 ;
      RECT 2259.945 189.04 2260.225 335.72 ;
      RECT 2259.385 189.04 2259.665 335.96 ;
      RECT 2258.825 187.94 2259.105 335.96 ;
      RECT 2258.265 189.04 2258.545 335.72 ;
      RECT 2257.705 187.94 2257.985 335.475 ;
      RECT 2257.145 189.04 2257.425 335.235 ;
      RECT 2256.585 187.94 2256.865 334.995 ;
      RECT 2256.025 189.04 2256.305 334.755 ;
      RECT 2255.465 189.04 2255.745 334.515 ;
      RECT 2254.905 189.04 2255.185 334.275 ;
      RECT 2254.345 189.04 2254.625 334.035 ;
      RECT 2253.785 189.04 2254.065 333.795 ;
      RECT 2253.225 189.04 2253.505 333.555 ;
      RECT 2252.665 189.04 2252.945 333.315 ;
      RECT 2252.105 189.04 2252.385 333.075 ;
      RECT 2251.545 187.94 2251.825 332.835 ;
      RECT 2250.985 189.04 2251.265 332.595 ;
      RECT 2250.425 187.94 2250.705 332.355 ;
      RECT 2249.865 189.04 2250.145 332.115 ;
      RECT 2249.305 189.04 2249.585 331.875 ;
      RECT 2248.745 189.04 2249.025 331.635 ;
      RECT 2235.305 189.04 2235.585 335.035 ;
      RECT 2234.745 189.04 2235.025 335.275 ;
      RECT 2234.185 189.04 2234.465 335.52 ;
      RECT 2233.625 189.04 2233.905 335.76 ;
      RECT 2233.065 189.04 2233.345 336 ;
      RECT 2232.505 189.04 2232.785 336 ;
      RECT 2231.945 189.04 2232.225 335.76 ;
      RECT 2231.385 189.04 2231.665 335.52 ;
      RECT 2230.825 189.04 2231.105 328.505 ;
      RECT 2230.265 189.04 2230.545 328.265 ;
      RECT 2229.705 189.04 2229.985 328.025 ;
      RECT 2229.145 187.94 2229.425 327.785 ;
      RECT 2228.585 189.04 2228.865 327.545 ;
      RECT 2228.025 187.94 2228.305 327.305 ;
      RECT 2227.465 189.04 2227.745 327.065 ;
      RECT 2226.905 189.04 2227.185 326.825 ;
      RECT 2226.345 189.04 2226.625 326.585 ;
      RECT 2225.785 187.94 2226.065 326.345 ;
      RECT 2225.225 189.04 2225.505 326.105 ;
      RECT 2224.665 187.94 2224.945 325.865 ;
      RECT 2224.105 189.04 2224.385 325.625 ;
      RECT 2223.545 187.94 2223.825 325.385 ;
      RECT 2222.985 189.04 2223.265 325.145 ;
      RECT 2222.425 189.04 2222.705 324.905 ;
      RECT 2182.105 189.04 2182.385 333.8 ;
      RECT 2181.545 189.04 2181.825 334.04 ;
      RECT 2180.985 189.04 2181.265 334.285 ;
      RECT 2180.425 189.04 2180.705 334.525 ;
      RECT 2179.865 189.04 2180.145 334.765 ;
      RECT 2179.305 189.04 2179.585 335.005 ;
      RECT 2178.745 189.04 2179.025 335.245 ;
      RECT 2178.185 189.04 2178.465 335.485 ;
      RECT 2177.625 189.04 2177.905 335.725 ;
      RECT 2177.065 189.04 2177.345 335.965 ;
      RECT 2176.505 187.94 2176.785 336.205 ;
      RECT 2175.945 189.04 2176.225 336.445 ;
      RECT 2175.385 187.94 2175.665 336.685 ;
      RECT 2174.825 189.04 2175.105 336.925 ;
      RECT 2174.265 187.94 2174.545 337.165 ;
      RECT 2173.705 189.04 2173.985 337.165 ;
      RECT 2173.145 189.04 2173.425 336.925 ;
      RECT 2172.585 189.04 2172.865 336.685 ;
      RECT 2172.025 189.04 2172.305 336.445 ;
      RECT 2171.465 189.04 2171.745 336.205 ;
      RECT 2170.905 189.04 2171.185 335.965 ;
      RECT 2170.345 189.04 2170.625 335.725 ;
      RECT 2169.785 189.04 2170.065 335.485 ;
      RECT 2160.825 187.94 2161.105 335.515 ;
      RECT 2160.265 189.04 2160.545 335.755 ;
      RECT 2159.705 187.94 2159.985 335.995 ;
      RECT 2159.145 189.04 2159.425 336.21 ;
      RECT 2158.585 189.04 2158.865 335.785 ;
      RECT 2158.025 189.04 2158.305 335.545 ;
      RECT 2157.465 189.04 2157.745 335.305 ;
      RECT 2156.905 189.04 2157.185 335.065 ;
      RECT 2156.345 189.04 2156.625 334.825 ;
      RECT 2155.785 189.04 2156.065 334.585 ;
      RECT 2155.225 189.04 2155.505 334.345 ;
      RECT 2154.665 189.04 2154.945 334.105 ;
      RECT 2154.105 189.04 2154.385 333.865 ;
      RECT 2153.545 189.04 2153.825 333.625 ;
      RECT 2151.025 189.04 2151.305 332.8 ;
      RECT 2150.465 189.04 2150.745 332.56 ;
      RECT 2149.905 189.04 2150.185 332.32 ;
      RECT 2149.345 187.94 2149.625 332.08 ;
      RECT 2148.785 189.04 2149.065 331.84 ;
      RECT 2148.225 187.94 2148.505 331.6 ;
      RECT 2147.665 189.04 2147.945 331.36 ;
      RECT 2147.105 189.04 2147.385 331.12 ;
      RECT 2120.505 189.04 2120.785 342.165 ;
      RECT 2119.945 187.94 2120.225 342.405 ;
      RECT 2119.385 189.04 2119.665 342.645 ;
      RECT 2118.825 187.94 2119.105 342.89 ;
      RECT 2118.265 189.04 2118.545 343.13 ;
      RECT 2117.705 187.94 2117.985 343.37 ;
      RECT 2117.145 189.04 2117.425 343.61 ;
      RECT 2116.585 189.04 2116.865 343.85 ;
      RECT 2116.025 189.04 2116.305 329.47 ;
      RECT 2115.465 189.04 2115.745 329.23 ;
      RECT 2114.905 189.04 2115.185 328.99 ;
      RECT 2114.345 189.04 2114.625 328.75 ;
      RECT 2113.785 189.04 2114.065 328.51 ;
      RECT 2113.225 189.04 2113.505 328.27 ;
      RECT 2112.665 189.04 2112.945 328.03 ;
      RECT 2112.105 189.04 2112.385 327.79 ;
      RECT 2111.545 189.04 2111.825 327.55 ;
      RECT 2110.985 189.04 2111.265 327.31 ;
      RECT 2110.425 187.94 2110.705 327.07 ;
      RECT 2109.865 189.04 2110.145 326.83 ;
      RECT 2109.305 187.94 2109.585 326.59 ;
      RECT 2108.745 189.04 2109.025 326.35 ;
      RECT 2094.745 187.94 2095.025 332.47 ;
      RECT 2094.185 189.04 2094.465 332.23 ;
      RECT 2093.625 189.04 2093.905 331.99 ;
      RECT 2093.065 189.04 2093.345 331.75 ;
      RECT 2092.505 189.04 2092.785 331.51 ;
      RECT 2091.945 189.04 2092.225 331.27 ;
      RECT 2091.385 189.04 2091.665 331.03 ;
      RECT 2090.825 189.04 2091.105 330.79 ;
      RECT 2090.265 189.04 2090.545 330.55 ;
      RECT 2089.705 187.94 2089.985 330.31 ;
      RECT 2089.145 189.04 2089.425 330.07 ;
      RECT 2088.585 187.94 2088.865 329.83 ;
      RECT 2088.025 189.04 2088.305 329.59 ;
      RECT 2087.465 189.04 2087.745 329.35 ;
      RECT 2086.905 189.04 2087.185 329.11 ;
      RECT 2086.345 189.04 2086.625 328.87 ;
      RECT 2085.785 189.04 2086.065 328.63 ;
      RECT 2085.225 189.04 2085.505 328.39 ;
      RECT 2084.665 189.04 2084.945 328.15 ;
      RECT 2084.105 189.04 2084.385 327.91 ;
      RECT 2083.545 189.04 2083.825 327.67 ;
      RECT 2082.985 189.04 2083.265 327.43 ;
      RECT 2082.425 189.04 2082.705 327.19 ;
      RECT 2043.225 189.04 2043.505 334.095 ;
      RECT 2042.665 189.04 2042.945 334.335 ;
      RECT 2042.105 189.04 2042.385 334.575 ;
      RECT 2041.545 187.94 2041.825 334.815 ;
      RECT 2040.985 189.04 2041.265 335.055 ;
      RECT 2040.425 187.94 2040.705 335.295 ;
      RECT 2039.865 189.04 2040.145 335.535 ;
      RECT 2039.305 189.04 2039.585 335.775 ;
      RECT 2038.745 189.04 2039.025 336.015 ;
      RECT 2038.185 187.94 2038.465 336.255 ;
      RECT 2037.625 189.04 2037.905 336.495 ;
      RECT 2037.065 187.94 2037.345 336.735 ;
      RECT 2036.505 189.04 2036.785 336.975 ;
      RECT 2035.945 187.94 2036.225 337.215 ;
      RECT 2035.385 189.04 2035.665 337.455 ;
      RECT 2034.825 189.04 2035.105 337.695 ;
      RECT 2034.265 189.04 2034.545 337.695 ;
      RECT 2033.705 189.04 2033.985 337.455 ;
      RECT 2033.145 189.04 2033.425 337.215 ;
      RECT 2032.585 189.04 2032.865 336.975 ;
      RECT 2032.025 189.04 2032.305 336.735 ;
      RECT 2031.465 189.04 2031.745 336.495 ;
      RECT 2030.905 189.04 2031.185 336.255 ;
      RECT 2030.345 189.04 2030.625 336.015 ;
      RECT 2029.785 189.04 2030.065 335.775 ;
      RECT 2020.825 189.04 2021.105 335.29 ;
      RECT 2020.265 187.94 2020.545 335.05 ;
      RECT 2019.705 189.04 2019.985 334.81 ;
      RECT 2019.145 187.94 2019.425 334.57 ;
      RECT 2018.585 189.04 2018.865 334.33 ;
      RECT 2018.025 187.94 2018.305 334.09 ;
      RECT 2017.465 189.04 2017.745 333.85 ;
      RECT 2016.905 189.04 2017.185 333.61 ;
      RECT 2016.345 189.04 2016.625 333.37 ;
      RECT 2015.785 189.04 2016.065 333.13 ;
      RECT 2015.225 189.04 2015.505 332.89 ;
      RECT 2014.665 189.04 2014.945 332.65 ;
      RECT 2014.105 189.04 2014.385 332.41 ;
      RECT 2013.545 189.04 2013.825 332.17 ;
      RECT 2011.025 187.94 2011.305 333.89 ;
      RECT 2010.465 189.04 2010.745 333.65 ;
      RECT 2009.905 187.94 2010.185 333.41 ;
      RECT 2009.345 189.04 2009.625 333.17 ;
      RECT 2008.785 189.04 2009.065 332.93 ;
      RECT 2008.225 189.04 2008.505 332.69 ;
      RECT 2007.665 189.04 2007.945 332.45 ;
      RECT 2007.105 189.04 2007.385 332.21 ;
      RECT 1981.065 189.04 1981.345 329.86 ;
      RECT 1980.505 189.04 1980.785 330.1 ;
      RECT 1979.945 189.04 1980.225 330.34 ;
      RECT 1979.385 189.04 1979.665 330.585 ;
      RECT 1978.825 189.04 1979.105 330.825 ;
      RECT 1978.265 189.04 1978.545 331.065 ;
      RECT 1977.705 189.04 1977.985 331.065 ;
      RECT 1977.145 189.04 1977.425 330.825 ;
      RECT 1976.585 189.04 1976.865 330.585 ;
      RECT 1976.025 187.94 1976.305 330.345 ;
      RECT 1975.465 189.04 1975.745 330.105 ;
      RECT 1974.905 187.94 1975.185 329.865 ;
      RECT 1974.345 189.04 1974.625 329.625 ;
      RECT 1973.785 189.04 1974.065 329.385 ;
      RECT 1973.225 189.04 1973.505 329.145 ;
      RECT 1972.665 187.94 1972.945 328.905 ;
      RECT 1972.105 189.04 1972.385 328.665 ;
      RECT 1971.545 187.94 1971.825 328.425 ;
      RECT 1970.985 189.04 1971.265 328.185 ;
      RECT 1970.425 187.94 1970.705 327.945 ;
      RECT 1969.865 189.04 1970.145 327.705 ;
      RECT 1969.305 189.04 1969.585 327.465 ;
      RECT 1968.745 189.04 1969.025 327.225 ;
      RECT 1968.185 189.04 1968.465 326.985 ;
      RECT 1954.745 189.04 1955.025 332.785 ;
      RECT 1954.185 189.04 1954.465 332.545 ;
      RECT 1953.625 189.04 1953.905 332.305 ;
      RECT 1953.065 189.04 1953.345 332.065 ;
      RECT 1952.505 189.04 1952.785 331.825 ;
      RECT 1951.945 189.04 1952.225 331.585 ;
      RECT 1951.385 189.04 1951.665 331.345 ;
      RECT 1950.825 189.04 1951.105 331.105 ;
      RECT 1950.265 187.94 1950.545 330.865 ;
      RECT 1949.705 189.04 1949.985 330.625 ;
      RECT 1949.145 187.94 1949.425 330.305 ;
      RECT 1948.585 189.04 1948.865 330.145 ;
      RECT 1948.025 187.94 1948.305 329.905 ;
      RECT 1947.465 189.04 1947.745 329.665 ;
      RECT 1946.905 189.04 1947.185 329.425 ;
      RECT 1946.345 189.04 1946.625 329.185 ;
      RECT 1945.785 189.04 1946.065 328.945 ;
      RECT 1945.225 189.04 1945.505 328.705 ;
      RECT 1944.665 189.04 1944.945 328.465 ;
      RECT 1944.105 189.04 1944.385 328.225 ;
      RECT 1943.545 189.04 1943.825 327.985 ;
      RECT 1942.985 187.94 1943.265 327.745 ;
      RECT 1942.425 189.04 1942.705 327.505 ;
      RECT 1941.865 187.94 1942.145 327.265 ;
      RECT 1902.665 189.04 1902.945 332.875 ;
      RECT 1902.105 189.04 1902.385 333.115 ;
      RECT 1901.545 189.04 1901.825 333.355 ;
      RECT 1900.985 189.04 1901.265 333.595 ;
      RECT 1900.425 189.04 1900.705 333.835 ;
      RECT 1899.865 189.04 1900.145 334.075 ;
      RECT 1899.305 189.04 1899.585 334.315 ;
      RECT 1898.745 189.04 1899.025 334.555 ;
      RECT 1898.185 189.04 1898.465 334.795 ;
      RECT 1897.625 189.04 1897.905 335.035 ;
      RECT 1897.065 189.04 1897.345 335.275 ;
      RECT 1896.505 189.04 1896.785 335.515 ;
      RECT 1895.945 189.04 1896.225 335.755 ;
      RECT 1895.385 189.04 1895.665 335.755 ;
      RECT 1894.825 187.94 1895.105 335.515 ;
      RECT 1894.265 189.04 1894.545 335.275 ;
      RECT 1893.705 187.94 1893.985 335.035 ;
      RECT 1893.145 189.04 1893.425 334.795 ;
      RECT 1892.585 189.04 1892.865 334.555 ;
      RECT 1892.025 189.04 1892.305 334.315 ;
      RECT 1891.465 187.94 1891.745 334.05 ;
      RECT 1890.905 189.04 1891.185 333.81 ;
      RECT 1890.345 187.94 1890.625 333.57 ;
      RECT 1889.785 189.04 1890.065 333.33 ;
      RECT 1880.825 187.94 1881.105 327.165 ;
      RECT 1880.265 189.04 1880.545 327.405 ;
      RECT 1879.705 189.04 1879.985 327.645 ;
      RECT 1879.145 189.04 1879.425 327.645 ;
      RECT 1878.585 189.04 1878.865 327.405 ;
      RECT 1878.025 189.04 1878.305 327.165 ;
      RECT 1877.465 189.04 1877.745 326.925 ;
      RECT 1876.905 189.04 1877.185 326.685 ;
      RECT 1876.345 189.04 1876.625 326.445 ;
      RECT 1875.785 189.04 1876.065 326.205 ;
      RECT 1875.225 189.04 1875.505 325.965 ;
      RECT 1874.665 189.04 1874.945 325.725 ;
      RECT 1874.105 189.04 1874.385 325.485 ;
      RECT 1873.545 187.94 1873.825 325.245 ;
      RECT 1871.025 189.04 1871.305 326.965 ;
      RECT 1870.465 187.94 1870.745 326.725 ;
      RECT 1869.905 189.04 1870.185 326.485 ;
      RECT 1869.345 187.94 1869.625 326.245 ;
      RECT 1868.785 189.04 1869.065 326.005 ;
      RECT 1868.225 189.04 1868.505 325.765 ;
      RECT 1867.665 189.04 1867.945 325.525 ;
      RECT 1841.625 189.04 1841.905 328.31 ;
      RECT 1841.065 189.04 1841.345 328.55 ;
      RECT 1840.505 189.04 1840.785 328.79 ;
      RECT 1839.945 189.04 1840.225 329.03 ;
      RECT 1839.385 189.04 1839.665 329.27 ;
      RECT 1838.825 187.94 1839.105 329.51 ;
      RECT 1838.265 189.04 1838.545 329.75 ;
      RECT 1837.705 187.94 1837.985 329.99 ;
      RECT 1837.145 189.04 1837.425 330.23 ;
      RECT 1836.585 189.04 1836.865 330.47 ;
      RECT 1836.025 189.04 1836.305 330.71 ;
      RECT 1835.465 189.04 1835.745 330.95 ;
      RECT 1834.905 189.04 1835.185 331.19 ;
      RECT 1834.345 189.04 1834.625 331.43 ;
      RECT 1833.785 189.04 1834.065 331.67 ;
      RECT 1833.225 189.04 1833.505 331.67 ;
      RECT 1832.665 189.04 1832.945 331.43 ;
      RECT 1832.105 189.04 1832.385 331.19 ;
      RECT 1831.545 189.04 1831.825 330.95 ;
      RECT 1830.985 189.04 1831.265 330.705 ;
      RECT 1830.425 189.04 1830.705 330.465 ;
      RECT 1829.865 189.04 1830.145 330.225 ;
      RECT 1829.305 187.94 1829.585 329.985 ;
      RECT 1828.745 189.04 1829.025 329.745 ;
      RECT 1815.305 187.94 1815.585 327.225 ;
      RECT 1814.745 189.04 1815.025 326.985 ;
      RECT 1814.185 189.04 1814.465 326.745 ;
      RECT 1813.625 189.04 1813.905 326.505 ;
      RECT 1813.065 187.94 1813.345 326.265 ;
      RECT 1812.505 189.04 1812.785 326.025 ;
      RECT 1811.945 187.94 1812.225 325.785 ;
      RECT 1811.385 189.04 1811.665 325.545 ;
      RECT 1810.825 187.94 1811.105 325.305 ;
      RECT 1810.265 189.04 1810.545 325.065 ;
      RECT 1809.705 189.04 1809.985 324.825 ;
      RECT 1809.145 189.04 1809.425 324.585 ;
      RECT 1808.585 189.04 1808.865 324.345 ;
      RECT 1808.025 189.04 1808.305 324.105 ;
      RECT 1807.465 189.04 1807.745 323.865 ;
      RECT 1806.905 189.04 1807.185 323.625 ;
      RECT 1806.345 189.04 1806.625 323.385 ;
      RECT 1805.785 189.04 1806.065 323.145 ;
      RECT 1805.225 189.04 1805.505 322.905 ;
      RECT 1804.665 189.04 1804.945 322.665 ;
      RECT 1804.105 189.04 1804.385 322.425 ;
      RECT 1803.545 187.94 1803.825 322.185 ;
      RECT 1802.985 189.04 1803.265 321.945 ;
      RECT 1802.425 187.94 1802.705 321.705 ;
      RECT 1762.665 189.04 1762.945 332.175 ;
      RECT 1762.105 187.94 1762.385 332.415 ;
      RECT 1761.545 189.04 1761.825 332.655 ;
      RECT 1760.985 189.04 1761.265 332.895 ;
      RECT 1760.425 189.04 1760.705 333.135 ;
      RECT 1759.865 189.04 1760.145 333.375 ;
      RECT 1759.305 189.04 1759.585 333.615 ;
      RECT 1758.745 189.04 1759.025 333.86 ;
      RECT 1758.185 189.04 1758.465 334.1 ;
      RECT 1757.625 189.04 1757.905 334.34 ;
      RECT 1757.065 187.94 1757.345 334.58 ;
      RECT 1756.505 189.04 1756.785 334.82 ;
      RECT 1755.945 187.94 1756.225 335.06 ;
      RECT 1755.385 189.04 1755.665 335.3 ;
      RECT 1754.825 189.04 1755.105 335.54 ;
      RECT 1754.265 189.04 1754.545 335.78 ;
      RECT 1753.705 189.04 1753.985 336.02 ;
      RECT 1753.145 189.04 1753.425 336.26 ;
      RECT 1752.585 189.04 1752.865 336.5 ;
      RECT 1752.025 189.04 1752.305 336.74 ;
      RECT 1751.465 189.04 1751.745 336.98 ;
      RECT 1750.905 189.04 1751.185 337.22 ;
      RECT 1750.345 189.04 1750.625 337.46 ;
      RECT 1749.785 189.04 1750.065 337.7 ;
      RECT 1740.825 189.04 1741.105 333.285 ;
      RECT 1740.265 189.04 1740.545 333.045 ;
      RECT 1739.705 189.04 1739.985 332.805 ;
      RECT 1739.145 187.94 1739.425 332.565 ;
      RECT 1738.585 189.04 1738.865 332.325 ;
      RECT 1738.025 187.94 1738.305 332.085 ;
      RECT 1737.465 189.04 1737.745 331.845 ;
      RECT 1736.905 189.04 1737.185 331.605 ;
      RECT 1736.345 189.04 1736.625 331.365 ;
      RECT 1735.785 187.94 1736.065 331.125 ;
      RECT 1735.225 189.04 1735.505 330.885 ;
      RECT 1734.665 187.94 1734.945 330.645 ;
      RECT 1734.105 189.04 1734.385 330.405 ;
      RECT 1733.545 187.94 1733.825 330.165 ;
      RECT 1731.025 189.04 1731.305 322.565 ;
      RECT 1730.465 189.04 1730.745 322.325 ;
      RECT 1729.905 189.04 1730.185 322.085 ;
      RECT 1729.345 189.04 1729.625 321.845 ;
      RECT 1728.785 189.04 1729.065 321.605 ;
      RECT 1728.225 189.04 1728.505 321.365 ;
      RECT 1727.665 189.04 1727.945 321.125 ;
      RECT 1701.625 189.04 1701.905 335 ;
      RECT 1701.065 189.04 1701.345 335.24 ;
      RECT 1700.505 189.04 1700.785 335.48 ;
      RECT 1699.945 189.04 1700.225 335.72 ;
      RECT 1699.385 189.04 1699.665 335.96 ;
      RECT 1698.825 187.94 1699.105 335.96 ;
      RECT 1698.265 189.04 1698.545 335.72 ;
      RECT 1697.705 187.94 1697.985 335.475 ;
      RECT 1697.145 189.04 1697.425 335.235 ;
      RECT 1696.585 187.94 1696.865 334.995 ;
      RECT 1696.025 189.04 1696.305 334.755 ;
      RECT 1695.465 189.04 1695.745 334.515 ;
      RECT 1694.905 189.04 1695.185 334.275 ;
      RECT 1694.345 189.04 1694.625 334.035 ;
      RECT 1693.785 189.04 1694.065 333.795 ;
      RECT 1693.225 189.04 1693.505 333.555 ;
      RECT 1692.665 189.04 1692.945 333.315 ;
      RECT 1692.105 189.04 1692.385 333.075 ;
      RECT 1691.545 187.94 1691.825 332.835 ;
      RECT 1690.985 189.04 1691.265 332.595 ;
      RECT 1690.425 187.94 1690.705 332.355 ;
      RECT 1689.865 189.04 1690.145 332.115 ;
      RECT 1689.305 189.04 1689.585 331.875 ;
      RECT 1688.745 189.04 1689.025 331.635 ;
      RECT 1675.305 189.04 1675.585 335.035 ;
      RECT 1674.745 189.04 1675.025 335.275 ;
      RECT 1674.185 189.04 1674.465 335.52 ;
      RECT 1673.625 189.04 1673.905 335.76 ;
      RECT 1673.065 189.04 1673.345 336 ;
      RECT 1672.505 189.04 1672.785 336 ;
      RECT 1671.945 189.04 1672.225 335.76 ;
      RECT 1671.385 189.04 1671.665 335.52 ;
      RECT 1670.825 189.04 1671.105 328.505 ;
      RECT 1670.265 189.04 1670.545 328.265 ;
      RECT 1669.705 189.04 1669.985 328.025 ;
      RECT 1669.145 187.94 1669.425 327.785 ;
      RECT 1668.585 189.04 1668.865 327.545 ;
      RECT 1668.025 187.94 1668.305 327.305 ;
      RECT 1667.465 189.04 1667.745 327.065 ;
      RECT 1666.905 189.04 1667.185 326.825 ;
      RECT 1666.345 189.04 1666.625 326.585 ;
      RECT 1665.785 187.94 1666.065 326.345 ;
      RECT 1665.225 189.04 1665.505 326.105 ;
      RECT 1664.665 187.94 1664.945 325.865 ;
      RECT 1664.105 189.04 1664.385 325.625 ;
      RECT 1663.545 187.94 1663.825 325.385 ;
      RECT 1662.985 189.04 1663.265 325.145 ;
      RECT 1662.425 189.04 1662.705 324.905 ;
      RECT 1622.105 189.04 1622.385 333.8 ;
      RECT 1621.545 189.04 1621.825 334.04 ;
      RECT 1620.985 189.04 1621.265 334.285 ;
      RECT 1620.425 189.04 1620.705 334.525 ;
      RECT 1619.865 189.04 1620.145 334.765 ;
      RECT 1619.305 189.04 1619.585 335.005 ;
      RECT 1618.745 189.04 1619.025 335.245 ;
      RECT 1618.185 189.04 1618.465 335.485 ;
      RECT 1617.625 189.04 1617.905 335.725 ;
      RECT 1617.065 189.04 1617.345 335.965 ;
      RECT 1616.505 187.94 1616.785 336.205 ;
      RECT 1615.945 189.04 1616.225 336.445 ;
      RECT 1615.385 187.94 1615.665 336.685 ;
      RECT 1614.825 189.04 1615.105 336.925 ;
      RECT 1614.265 187.94 1614.545 337.165 ;
      RECT 1613.705 189.04 1613.985 337.165 ;
      RECT 1613.145 189.04 1613.425 336.925 ;
      RECT 1612.585 189.04 1612.865 336.685 ;
      RECT 1612.025 189.04 1612.305 336.445 ;
      RECT 1611.465 189.04 1611.745 336.205 ;
      RECT 1610.905 189.04 1611.185 335.965 ;
      RECT 1610.345 189.04 1610.625 335.725 ;
      RECT 1609.785 189.04 1610.065 335.485 ;
      RECT 1600.825 187.94 1601.105 335.515 ;
      RECT 1600.265 189.04 1600.545 335.755 ;
      RECT 1599.705 187.94 1599.985 335.995 ;
      RECT 1599.145 189.04 1599.425 336.21 ;
      RECT 1598.585 189.04 1598.865 335.785 ;
      RECT 1598.025 189.04 1598.305 335.545 ;
      RECT 1597.465 189.04 1597.745 335.305 ;
      RECT 1596.905 189.04 1597.185 335.065 ;
      RECT 1596.345 189.04 1596.625 334.825 ;
      RECT 1595.785 189.04 1596.065 334.585 ;
      RECT 1595.225 189.04 1595.505 334.345 ;
      RECT 1594.665 189.04 1594.945 334.105 ;
      RECT 1594.105 189.04 1594.385 333.865 ;
      RECT 1593.545 189.04 1593.825 333.625 ;
      RECT 1591.025 189.04 1591.305 332.8 ;
      RECT 1590.465 189.04 1590.745 332.56 ;
      RECT 1589.905 189.04 1590.185 332.32 ;
      RECT 1589.345 187.94 1589.625 332.08 ;
      RECT 1588.785 189.04 1589.065 331.84 ;
      RECT 1588.225 187.94 1588.505 331.6 ;
      RECT 1587.665 189.04 1587.945 331.36 ;
      RECT 1587.105 189.04 1587.385 331.12 ;
      RECT 1560.505 189.04 1560.785 342.165 ;
      RECT 1559.945 187.94 1560.225 342.405 ;
      RECT 1559.385 189.04 1559.665 342.645 ;
      RECT 1558.825 187.94 1559.105 342.89 ;
      RECT 1558.265 189.04 1558.545 343.13 ;
      RECT 1557.705 187.94 1557.985 343.37 ;
      RECT 1557.145 189.04 1557.425 343.61 ;
      RECT 1556.585 189.04 1556.865 343.85 ;
      RECT 1556.025 189.04 1556.305 329.47 ;
      RECT 1555.465 189.04 1555.745 329.23 ;
      RECT 1554.905 189.04 1555.185 328.99 ;
      RECT 1554.345 189.04 1554.625 328.75 ;
      RECT 1553.785 189.04 1554.065 328.51 ;
      RECT 1553.225 189.04 1553.505 328.27 ;
      RECT 1552.665 189.04 1552.945 328.03 ;
      RECT 1552.105 189.04 1552.385 327.79 ;
      RECT 1551.545 189.04 1551.825 327.55 ;
      RECT 1550.985 189.04 1551.265 327.31 ;
      RECT 1550.425 187.94 1550.705 327.07 ;
      RECT 1549.865 189.04 1550.145 326.83 ;
      RECT 1549.305 187.94 1549.585 326.59 ;
      RECT 1548.745 189.04 1549.025 326.35 ;
      RECT 1534.745 187.94 1535.025 332.47 ;
      RECT 1534.185 189.04 1534.465 332.23 ;
      RECT 1533.625 189.04 1533.905 331.99 ;
      RECT 1533.065 189.04 1533.345 331.75 ;
      RECT 1532.505 189.04 1532.785 331.51 ;
      RECT 1531.945 189.04 1532.225 331.27 ;
      RECT 1531.385 189.04 1531.665 331.03 ;
      RECT 1530.825 189.04 1531.105 330.79 ;
      RECT 1530.265 189.04 1530.545 330.55 ;
      RECT 1529.705 187.94 1529.985 330.31 ;
      RECT 1529.145 189.04 1529.425 330.07 ;
      RECT 1528.585 187.94 1528.865 329.83 ;
      RECT 1528.025 189.04 1528.305 329.59 ;
      RECT 1527.465 189.04 1527.745 329.35 ;
      RECT 1526.905 189.04 1527.185 329.11 ;
      RECT 1526.345 189.04 1526.625 328.87 ;
      RECT 1525.785 189.04 1526.065 328.63 ;
      RECT 1525.225 189.04 1525.505 328.39 ;
      RECT 1524.665 189.04 1524.945 328.15 ;
      RECT 1524.105 189.04 1524.385 327.91 ;
      RECT 1523.545 189.04 1523.825 327.67 ;
      RECT 1522.985 189.04 1523.265 327.43 ;
      RECT 1522.425 189.04 1522.705 327.19 ;
      RECT 1483.225 189.04 1483.505 334.095 ;
      RECT 1482.665 189.04 1482.945 334.335 ;
      RECT 1482.105 189.04 1482.385 334.575 ;
      RECT 1481.545 187.94 1481.825 334.815 ;
      RECT 1480.985 189.04 1481.265 335.055 ;
      RECT 1480.425 187.94 1480.705 335.295 ;
      RECT 1479.865 189.04 1480.145 335.535 ;
      RECT 1479.305 189.04 1479.585 335.775 ;
      RECT 1478.745 189.04 1479.025 336.015 ;
      RECT 1478.185 187.94 1478.465 336.255 ;
      RECT 1477.625 189.04 1477.905 336.495 ;
      RECT 1477.065 187.94 1477.345 336.735 ;
      RECT 1476.505 189.04 1476.785 336.975 ;
      RECT 1475.945 187.94 1476.225 337.215 ;
      RECT 1475.385 189.04 1475.665 337.455 ;
      RECT 1474.825 189.04 1475.105 337.695 ;
      RECT 1474.265 189.04 1474.545 337.695 ;
      RECT 1473.705 189.04 1473.985 337.455 ;
      RECT 1473.145 189.04 1473.425 337.215 ;
      RECT 1472.585 189.04 1472.865 336.975 ;
      RECT 1472.025 189.04 1472.305 336.735 ;
      RECT 1471.465 189.04 1471.745 336.495 ;
      RECT 1470.905 189.04 1471.185 336.255 ;
      RECT 1470.345 189.04 1470.625 336.015 ;
      RECT 1469.785 189.04 1470.065 335.775 ;
      RECT 1460.825 189.04 1461.105 335.29 ;
      RECT 1460.265 187.94 1460.545 335.05 ;
      RECT 1459.705 189.04 1459.985 334.81 ;
      RECT 1459.145 187.94 1459.425 334.57 ;
      RECT 1458.585 189.04 1458.865 334.33 ;
      RECT 1458.025 187.94 1458.305 334.09 ;
      RECT 1457.465 189.04 1457.745 333.85 ;
      RECT 1456.905 189.04 1457.185 333.61 ;
      RECT 1456.345 189.04 1456.625 333.37 ;
      RECT 1455.785 189.04 1456.065 333.13 ;
      RECT 1455.225 189.04 1455.505 332.89 ;
      RECT 1454.665 189.04 1454.945 332.65 ;
      RECT 1454.105 189.04 1454.385 332.41 ;
      RECT 1453.545 189.04 1453.825 332.17 ;
      RECT 1451.025 187.94 1451.305 333.89 ;
      RECT 1450.465 189.04 1450.745 333.65 ;
      RECT 1449.905 187.94 1450.185 333.41 ;
      RECT 1449.345 189.04 1449.625 333.17 ;
      RECT 1448.785 189.04 1449.065 332.93 ;
      RECT 1448.225 189.04 1448.505 332.69 ;
      RECT 1447.665 189.04 1447.945 332.45 ;
      RECT 1447.105 189.04 1447.385 332.21 ;
      RECT 1421.065 189.04 1421.345 329.86 ;
      RECT 1420.505 189.04 1420.785 330.1 ;
      RECT 1419.945 189.04 1420.225 330.34 ;
      RECT 1419.385 189.04 1419.665 330.585 ;
      RECT 1418.825 189.04 1419.105 330.825 ;
      RECT 1418.265 189.04 1418.545 331.065 ;
      RECT 1417.705 189.04 1417.985 331.065 ;
      RECT 1417.145 189.04 1417.425 330.825 ;
      RECT 1416.585 189.04 1416.865 330.585 ;
      RECT 1416.025 187.94 1416.305 330.345 ;
      RECT 1415.465 189.04 1415.745 330.105 ;
      RECT 1414.905 187.94 1415.185 329.865 ;
      RECT 1414.345 189.04 1414.625 329.625 ;
      RECT 1413.785 189.04 1414.065 329.385 ;
      RECT 1413.225 189.04 1413.505 329.145 ;
      RECT 1412.665 187.94 1412.945 328.905 ;
      RECT 1412.105 189.04 1412.385 328.665 ;
      RECT 1411.545 187.94 1411.825 328.425 ;
      RECT 1410.985 189.04 1411.265 328.185 ;
      RECT 1410.425 187.94 1410.705 327.945 ;
      RECT 1409.865 189.04 1410.145 327.705 ;
      RECT 1409.305 189.04 1409.585 327.465 ;
      RECT 1408.745 189.04 1409.025 327.225 ;
      RECT 1408.185 189.04 1408.465 326.985 ;
      RECT 1394.745 189.04 1395.025 332.785 ;
      RECT 1394.185 189.04 1394.465 332.545 ;
      RECT 1393.625 189.04 1393.905 332.305 ;
      RECT 1393.065 189.04 1393.345 332.065 ;
      RECT 1392.505 189.04 1392.785 331.825 ;
      RECT 1391.945 189.04 1392.225 331.585 ;
      RECT 1391.385 189.04 1391.665 331.345 ;
      RECT 1390.825 189.04 1391.105 331.105 ;
      RECT 1390.265 187.94 1390.545 330.865 ;
      RECT 1389.705 189.04 1389.985 330.625 ;
      RECT 1389.145 187.94 1389.425 330.305 ;
      RECT 1388.585 189.04 1388.865 330.145 ;
      RECT 1388.025 187.94 1388.305 329.905 ;
      RECT 1387.465 189.04 1387.745 329.665 ;
      RECT 1386.905 189.04 1387.185 329.425 ;
      RECT 1386.345 189.04 1386.625 329.185 ;
      RECT 1385.785 189.04 1386.065 328.945 ;
      RECT 1385.225 189.04 1385.505 328.705 ;
      RECT 1384.665 189.04 1384.945 328.465 ;
      RECT 1384.105 189.04 1384.385 328.225 ;
      RECT 1383.545 189.04 1383.825 327.985 ;
      RECT 1382.985 187.94 1383.265 327.745 ;
      RECT 1382.425 189.04 1382.705 327.505 ;
      RECT 1381.865 187.94 1382.145 327.265 ;
      RECT 1342.665 189.04 1342.945 332.875 ;
      RECT 1342.105 189.04 1342.385 333.115 ;
      RECT 1341.545 189.04 1341.825 333.355 ;
      RECT 1340.985 189.04 1341.265 333.595 ;
      RECT 1340.425 189.04 1340.705 333.835 ;
      RECT 1339.865 189.04 1340.145 334.075 ;
      RECT 1339.305 189.04 1339.585 334.315 ;
      RECT 1338.745 189.04 1339.025 334.555 ;
      RECT 1338.185 189.04 1338.465 334.795 ;
      RECT 1337.625 189.04 1337.905 335.035 ;
      RECT 1337.065 189.04 1337.345 335.275 ;
      RECT 1336.505 189.04 1336.785 335.515 ;
      RECT 1335.945 189.04 1336.225 335.755 ;
      RECT 1335.385 189.04 1335.665 335.755 ;
      RECT 1334.825 187.94 1335.105 335.515 ;
      RECT 1334.265 189.04 1334.545 335.275 ;
      RECT 1333.705 187.94 1333.985 335.035 ;
      RECT 1333.145 189.04 1333.425 334.795 ;
      RECT 1332.585 189.04 1332.865 334.555 ;
      RECT 1332.025 189.04 1332.305 334.315 ;
      RECT 1331.465 187.94 1331.745 334.05 ;
      RECT 1330.905 189.04 1331.185 333.81 ;
      RECT 1330.345 187.94 1330.625 333.57 ;
      RECT 1329.785 189.04 1330.065 333.33 ;
      RECT 1320.825 187.94 1321.105 327.165 ;
      RECT 1320.265 189.04 1320.545 327.405 ;
      RECT 1319.705 189.04 1319.985 327.645 ;
      RECT 1319.145 189.04 1319.425 327.645 ;
      RECT 1318.585 189.04 1318.865 327.405 ;
      RECT 1318.025 189.04 1318.305 327.165 ;
      RECT 1317.465 189.04 1317.745 326.925 ;
      RECT 1316.905 189.04 1317.185 326.685 ;
      RECT 1316.345 189.04 1316.625 326.445 ;
      RECT 1315.785 189.04 1316.065 326.205 ;
      RECT 1315.225 189.04 1315.505 325.965 ;
      RECT 1314.665 189.04 1314.945 325.725 ;
      RECT 1314.105 189.04 1314.385 325.485 ;
      RECT 1313.545 187.94 1313.825 325.245 ;
      RECT 1311.025 189.04 1311.305 326.965 ;
      RECT 1310.465 187.94 1310.745 326.725 ;
      RECT 1309.905 189.04 1310.185 326.485 ;
      RECT 1309.345 187.94 1309.625 326.245 ;
      RECT 1308.785 189.04 1309.065 326.005 ;
      RECT 1308.225 189.04 1308.505 325.765 ;
      RECT 1307.665 189.04 1307.945 325.525 ;
      RECT 1281.625 189.04 1281.905 328.31 ;
      RECT 1281.065 189.04 1281.345 328.55 ;
      RECT 1280.505 189.04 1280.785 328.79 ;
      RECT 1279.945 189.04 1280.225 329.03 ;
      RECT 1279.385 189.04 1279.665 329.27 ;
      RECT 1278.825 187.94 1279.105 329.51 ;
      RECT 1278.265 189.04 1278.545 329.75 ;
      RECT 1277.705 187.94 1277.985 329.99 ;
      RECT 1277.145 189.04 1277.425 330.23 ;
      RECT 1276.585 189.04 1276.865 330.47 ;
      RECT 1276.025 189.04 1276.305 330.71 ;
      RECT 1275.465 189.04 1275.745 330.95 ;
      RECT 1274.905 189.04 1275.185 331.19 ;
      RECT 1274.345 189.04 1274.625 331.43 ;
      RECT 1273.785 189.04 1274.065 331.67 ;
      RECT 1273.225 189.04 1273.505 331.67 ;
      RECT 1272.665 189.04 1272.945 331.43 ;
      RECT 1272.105 189.04 1272.385 331.19 ;
      RECT 1271.545 189.04 1271.825 330.95 ;
      RECT 1270.985 189.04 1271.265 330.705 ;
      RECT 1270.425 189.04 1270.705 330.465 ;
      RECT 1269.865 189.04 1270.145 330.225 ;
      RECT 1269.305 187.94 1269.585 329.985 ;
      RECT 1268.745 189.04 1269.025 329.745 ;
      RECT 1255.305 187.94 1255.585 327.225 ;
      RECT 1254.745 189.04 1255.025 326.985 ;
      RECT 1254.185 189.04 1254.465 326.745 ;
      RECT 1253.625 189.04 1253.905 326.505 ;
      RECT 1253.065 187.94 1253.345 326.265 ;
      RECT 1252.505 189.04 1252.785 326.025 ;
      RECT 1251.945 187.94 1252.225 325.785 ;
      RECT 1251.385 189.04 1251.665 325.545 ;
      RECT 1250.825 187.94 1251.105 325.305 ;
      RECT 1250.265 189.04 1250.545 325.065 ;
      RECT 1249.705 189.04 1249.985 324.825 ;
      RECT 1249.145 189.04 1249.425 324.585 ;
      RECT 1248.585 189.04 1248.865 324.345 ;
      RECT 1248.025 189.04 1248.305 324.105 ;
      RECT 1247.465 189.04 1247.745 323.865 ;
      RECT 1246.905 189.04 1247.185 323.625 ;
      RECT 1246.345 189.04 1246.625 323.385 ;
      RECT 1245.785 189.04 1246.065 323.145 ;
      RECT 1245.225 189.04 1245.505 322.905 ;
      RECT 1244.665 189.04 1244.945 322.665 ;
      RECT 1244.105 189.04 1244.385 322.425 ;
      RECT 1243.545 187.94 1243.825 322.185 ;
      RECT 1242.985 189.04 1243.265 321.945 ;
      RECT 1242.425 187.94 1242.705 321.705 ;
      RECT 1202.665 189.04 1202.945 332.175 ;
      RECT 1202.105 187.94 1202.385 332.415 ;
      RECT 1201.545 189.04 1201.825 332.655 ;
      RECT 1200.985 189.04 1201.265 332.895 ;
      RECT 1200.425 189.04 1200.705 333.135 ;
      RECT 1199.865 189.04 1200.145 333.375 ;
      RECT 1199.305 189.04 1199.585 333.615 ;
      RECT 1198.745 189.04 1199.025 333.86 ;
      RECT 1198.185 189.04 1198.465 334.1 ;
      RECT 1197.625 189.04 1197.905 334.34 ;
      RECT 1197.065 187.94 1197.345 334.58 ;
      RECT 1196.505 189.04 1196.785 334.82 ;
      RECT 1195.945 187.94 1196.225 335.06 ;
      RECT 1195.385 189.04 1195.665 335.3 ;
      RECT 1194.825 189.04 1195.105 335.54 ;
      RECT 1194.265 189.04 1194.545 335.78 ;
      RECT 1193.705 189.04 1193.985 336.02 ;
      RECT 1193.145 189.04 1193.425 336.26 ;
      RECT 1192.585 189.04 1192.865 336.5 ;
      RECT 1192.025 189.04 1192.305 336.74 ;
      RECT 1191.465 189.04 1191.745 336.98 ;
      RECT 1190.905 189.04 1191.185 337.22 ;
      RECT 1190.345 189.04 1190.625 337.46 ;
      RECT 1189.785 189.04 1190.065 337.7 ;
      RECT 1180.825 189.04 1181.105 333.285 ;
      RECT 1180.265 189.04 1180.545 333.045 ;
      RECT 1179.705 189.04 1179.985 332.805 ;
      RECT 1179.145 187.94 1179.425 332.565 ;
      RECT 1178.585 189.04 1178.865 332.325 ;
      RECT 1178.025 187.94 1178.305 332.085 ;
      RECT 1177.465 189.04 1177.745 331.845 ;
      RECT 1176.905 189.04 1177.185 331.605 ;
      RECT 1176.345 189.04 1176.625 331.365 ;
      RECT 1175.785 187.94 1176.065 331.125 ;
      RECT 1175.225 189.04 1175.505 330.885 ;
      RECT 1174.665 187.94 1174.945 330.645 ;
      RECT 1174.105 189.04 1174.385 330.405 ;
      RECT 1173.545 187.94 1173.825 330.165 ;
      RECT 1171.025 189.04 1171.305 322.565 ;
      RECT 1170.465 189.04 1170.745 322.325 ;
      RECT 1169.905 189.04 1170.185 322.085 ;
      RECT 1169.345 189.04 1169.625 321.845 ;
      RECT 1168.785 189.04 1169.065 321.605 ;
      RECT 1168.225 189.04 1168.505 321.365 ;
      RECT 1167.665 189.04 1167.945 321.125 ;
      RECT 1141.625 189.04 1141.905 335 ;
      RECT 1141.065 189.04 1141.345 335.24 ;
      RECT 1140.505 189.04 1140.785 335.48 ;
      RECT 1139.945 189.04 1140.225 335.72 ;
      RECT 1139.385 189.04 1139.665 335.96 ;
      RECT 1138.825 187.94 1139.105 335.96 ;
      RECT 1138.265 189.04 1138.545 335.72 ;
      RECT 1137.705 187.94 1137.985 335.475 ;
      RECT 1137.145 189.04 1137.425 335.235 ;
      RECT 1136.585 187.94 1136.865 334.995 ;
      RECT 1136.025 189.04 1136.305 334.755 ;
      RECT 1135.465 189.04 1135.745 334.515 ;
      RECT 1134.905 189.04 1135.185 334.275 ;
      RECT 1134.345 189.04 1134.625 334.035 ;
      RECT 1133.785 189.04 1134.065 333.795 ;
      RECT 1133.225 189.04 1133.505 333.555 ;
      RECT 1132.665 189.04 1132.945 333.315 ;
      RECT 1132.105 189.04 1132.385 333.075 ;
      RECT 1131.545 187.94 1131.825 332.835 ;
      RECT 1130.985 189.04 1131.265 332.595 ;
      RECT 1130.425 187.94 1130.705 332.355 ;
      RECT 1129.865 189.04 1130.145 332.115 ;
      RECT 1129.305 189.04 1129.585 331.875 ;
      RECT 1128.745 189.04 1129.025 331.635 ;
      RECT 1115.305 189.04 1115.585 335.035 ;
      RECT 1114.745 189.04 1115.025 335.275 ;
      RECT 1114.185 189.04 1114.465 335.52 ;
      RECT 1113.625 189.04 1113.905 335.76 ;
      RECT 1113.065 189.04 1113.345 336 ;
      RECT 1112.505 189.04 1112.785 336 ;
      RECT 1111.945 189.04 1112.225 335.76 ;
      RECT 1111.385 189.04 1111.665 335.52 ;
      RECT 1110.825 189.04 1111.105 328.505 ;
      RECT 1110.265 189.04 1110.545 328.265 ;
      RECT 1109.705 189.04 1109.985 328.025 ;
      RECT 1109.145 187.94 1109.425 327.785 ;
      RECT 1108.585 189.04 1108.865 327.545 ;
      RECT 1108.025 187.94 1108.305 327.305 ;
      RECT 1107.465 189.04 1107.745 327.065 ;
      RECT 1106.905 189.04 1107.185 326.825 ;
      RECT 1106.345 189.04 1106.625 326.585 ;
      RECT 1105.785 187.94 1106.065 326.345 ;
      RECT 1105.225 189.04 1105.505 326.105 ;
      RECT 1104.665 187.94 1104.945 325.865 ;
      RECT 1104.105 189.04 1104.385 325.625 ;
      RECT 1103.545 187.94 1103.825 325.385 ;
      RECT 1102.985 189.04 1103.265 325.145 ;
      RECT 1102.425 189.04 1102.705 324.905 ;
      RECT 1062.105 189.04 1062.385 333.8 ;
      RECT 1061.545 189.04 1061.825 334.04 ;
      RECT 1060.985 189.04 1061.265 334.285 ;
      RECT 1060.425 189.04 1060.705 334.525 ;
      RECT 1059.865 189.04 1060.145 334.765 ;
      RECT 1059.305 189.04 1059.585 335.005 ;
      RECT 1058.745 189.04 1059.025 335.245 ;
      RECT 1058.185 189.04 1058.465 335.485 ;
      RECT 1057.625 189.04 1057.905 335.725 ;
      RECT 1057.065 189.04 1057.345 335.965 ;
      RECT 1056.505 187.94 1056.785 336.205 ;
      RECT 1055.945 189.04 1056.225 336.445 ;
      RECT 1055.385 187.94 1055.665 336.685 ;
      RECT 1054.825 189.04 1055.105 336.925 ;
      RECT 1054.265 187.94 1054.545 337.165 ;
      RECT 1053.705 189.04 1053.985 337.165 ;
      RECT 1053.145 189.04 1053.425 336.925 ;
      RECT 1052.585 189.04 1052.865 336.685 ;
      RECT 1052.025 189.04 1052.305 336.445 ;
      RECT 1051.465 189.04 1051.745 336.205 ;
      RECT 1050.905 189.04 1051.185 335.965 ;
      RECT 1050.345 189.04 1050.625 335.725 ;
      RECT 1049.785 189.04 1050.065 335.485 ;
      RECT 1040.825 187.94 1041.105 335.515 ;
      RECT 1040.265 189.04 1040.545 335.755 ;
      RECT 1039.705 187.94 1039.985 335.995 ;
      RECT 1039.145 189.04 1039.425 336.21 ;
      RECT 1038.585 189.04 1038.865 335.785 ;
      RECT 1038.025 189.04 1038.305 335.545 ;
      RECT 1037.465 189.04 1037.745 335.305 ;
      RECT 1036.905 189.04 1037.185 335.065 ;
      RECT 1036.345 189.04 1036.625 334.825 ;
      RECT 1035.785 189.04 1036.065 334.585 ;
      RECT 1035.225 189.04 1035.505 334.345 ;
      RECT 1034.665 189.04 1034.945 334.105 ;
      RECT 1034.105 189.04 1034.385 333.865 ;
      RECT 1033.545 189.04 1033.825 333.625 ;
      RECT 1031.025 189.04 1031.305 332.8 ;
      RECT 1030.465 189.04 1030.745 332.56 ;
      RECT 1029.905 189.04 1030.185 332.32 ;
      RECT 1029.345 187.94 1029.625 332.08 ;
      RECT 1028.785 189.04 1029.065 331.84 ;
      RECT 1028.225 187.94 1028.505 331.6 ;
      RECT 1027.665 189.04 1027.945 331.36 ;
      RECT 1027.105 189.04 1027.385 331.12 ;
      RECT 1000.505 189.04 1000.785 342.165 ;
      RECT 999.945 187.94 1000.225 342.405 ;
      RECT 999.385 189.04 999.665 342.645 ;
      RECT 998.825 187.94 999.105 342.89 ;
      RECT 998.265 189.04 998.545 343.13 ;
      RECT 997.705 187.94 997.985 343.37 ;
      RECT 997.145 189.04 997.425 343.61 ;
      RECT 996.585 189.04 996.865 343.85 ;
      RECT 996.025 189.04 996.305 329.47 ;
      RECT 995.465 189.04 995.745 329.23 ;
      RECT 994.905 189.04 995.185 328.99 ;
      RECT 994.345 189.04 994.625 328.75 ;
      RECT 993.785 189.04 994.065 328.51 ;
      RECT 993.225 189.04 993.505 328.27 ;
      RECT 992.665 189.04 992.945 328.03 ;
      RECT 992.105 189.04 992.385 327.79 ;
      RECT 991.545 189.04 991.825 327.55 ;
      RECT 990.985 189.04 991.265 327.31 ;
      RECT 990.425 187.94 990.705 327.07 ;
      RECT 989.865 189.04 990.145 326.83 ;
      RECT 989.305 187.94 989.585 326.59 ;
      RECT 988.745 189.04 989.025 326.35 ;
      RECT 974.745 187.94 975.025 332.47 ;
      RECT 974.185 189.04 974.465 332.23 ;
      RECT 973.625 189.04 973.905 331.99 ;
      RECT 973.065 189.04 973.345 331.75 ;
      RECT 972.505 189.04 972.785 331.51 ;
      RECT 971.945 189.04 972.225 331.27 ;
      RECT 971.385 189.04 971.665 331.03 ;
      RECT 970.825 189.04 971.105 330.79 ;
      RECT 970.265 189.04 970.545 330.55 ;
      RECT 969.705 187.94 969.985 330.31 ;
      RECT 969.145 189.04 969.425 330.07 ;
      RECT 968.585 187.94 968.865 329.83 ;
      RECT 968.025 189.04 968.305 329.59 ;
      RECT 967.465 189.04 967.745 329.35 ;
      RECT 966.905 189.04 967.185 329.11 ;
      RECT 966.345 189.04 966.625 328.87 ;
      RECT 965.785 189.04 966.065 328.63 ;
      RECT 965.225 189.04 965.505 328.39 ;
      RECT 964.665 189.04 964.945 328.15 ;
      RECT 964.105 189.04 964.385 327.91 ;
      RECT 963.545 189.04 963.825 327.67 ;
      RECT 962.985 189.04 963.265 327.43 ;
      RECT 962.425 189.04 962.705 327.19 ;
      RECT 923.225 189.04 923.505 334.095 ;
      RECT 922.665 189.04 922.945 334.335 ;
      RECT 922.105 189.04 922.385 334.575 ;
      RECT 921.545 187.94 921.825 334.815 ;
      RECT 920.985 189.04 921.265 335.055 ;
      RECT 920.425 187.94 920.705 335.295 ;
      RECT 919.865 189.04 920.145 335.535 ;
      RECT 919.305 189.04 919.585 335.775 ;
      RECT 918.745 189.04 919.025 336.015 ;
      RECT 918.185 187.94 918.465 336.255 ;
      RECT 917.625 189.04 917.905 336.495 ;
      RECT 917.065 187.94 917.345 336.735 ;
      RECT 916.505 189.04 916.785 336.975 ;
      RECT 915.945 187.94 916.225 337.215 ;
      RECT 915.385 189.04 915.665 337.455 ;
      RECT 914.825 189.04 915.105 337.695 ;
      RECT 914.265 189.04 914.545 337.695 ;
      RECT 913.705 189.04 913.985 337.455 ;
      RECT 913.145 189.04 913.425 337.215 ;
      RECT 912.585 189.04 912.865 336.975 ;
      RECT 912.025 189.04 912.305 336.735 ;
      RECT 911.465 189.04 911.745 336.495 ;
      RECT 910.905 189.04 911.185 336.255 ;
      RECT 910.345 189.04 910.625 336.015 ;
      RECT 909.785 189.04 910.065 335.775 ;
      RECT 900.825 189.04 901.105 335.29 ;
      RECT 900.265 187.94 900.545 335.05 ;
      RECT 899.705 189.04 899.985 334.81 ;
      RECT 899.145 187.94 899.425 334.57 ;
      RECT 898.585 189.04 898.865 334.33 ;
      RECT 898.025 187.94 898.305 334.09 ;
      RECT 897.465 189.04 897.745 333.85 ;
      RECT 896.905 189.04 897.185 333.61 ;
      RECT 896.345 189.04 896.625 333.37 ;
      RECT 895.785 189.04 896.065 333.13 ;
      RECT 895.225 189.04 895.505 332.89 ;
      RECT 894.665 189.04 894.945 332.65 ;
      RECT 894.105 189.04 894.385 332.41 ;
      RECT 893.545 189.04 893.825 332.17 ;
      RECT 891.025 187.94 891.305 333.89 ;
      RECT 890.465 189.04 890.745 333.65 ;
      RECT 889.905 187.94 890.185 333.41 ;
      RECT 889.345 189.04 889.625 333.17 ;
      RECT 888.785 189.04 889.065 332.93 ;
      RECT 888.225 189.04 888.505 332.69 ;
      RECT 887.665 189.04 887.945 332.45 ;
      RECT 887.105 189.04 887.385 332.21 ;
      RECT 861.065 189.04 861.345 329.86 ;
      RECT 860.505 189.04 860.785 330.1 ;
      RECT 859.945 189.04 860.225 330.34 ;
      RECT 859.385 189.04 859.665 330.585 ;
      RECT 858.825 189.04 859.105 330.825 ;
      RECT 858.265 189.04 858.545 331.065 ;
      RECT 857.705 189.04 857.985 331.065 ;
      RECT 857.145 189.04 857.425 330.825 ;
      RECT 856.585 189.04 856.865 330.585 ;
      RECT 856.025 187.94 856.305 330.345 ;
      RECT 855.465 189.04 855.745 330.105 ;
      RECT 854.905 187.94 855.185 329.865 ;
      RECT 854.345 189.04 854.625 329.625 ;
      RECT 853.785 189.04 854.065 329.385 ;
      RECT 853.225 189.04 853.505 329.145 ;
      RECT 852.665 187.94 852.945 328.905 ;
      RECT 852.105 189.04 852.385 328.665 ;
      RECT 851.545 187.94 851.825 328.425 ;
      RECT 850.985 189.04 851.265 328.185 ;
      RECT 850.425 187.94 850.705 327.945 ;
      RECT 849.865 189.04 850.145 327.705 ;
      RECT 849.305 189.04 849.585 327.465 ;
      RECT 848.745 189.04 849.025 327.225 ;
      RECT 848.185 189.04 848.465 326.985 ;
      RECT 834.745 189.04 835.025 332.785 ;
      RECT 834.185 189.04 834.465 332.545 ;
      RECT 833.625 189.04 833.905 332.305 ;
      RECT 833.065 189.04 833.345 332.065 ;
      RECT 832.505 189.04 832.785 331.825 ;
      RECT 831.945 189.04 832.225 331.585 ;
      RECT 831.385 189.04 831.665 331.345 ;
      RECT 830.825 189.04 831.105 331.105 ;
      RECT 830.265 187.94 830.545 330.865 ;
      RECT 829.705 189.04 829.985 330.625 ;
      RECT 829.145 187.94 829.425 330.305 ;
      RECT 828.585 189.04 828.865 330.145 ;
      RECT 828.025 187.94 828.305 329.905 ;
      RECT 827.465 189.04 827.745 329.665 ;
      RECT 826.905 189.04 827.185 329.425 ;
      RECT 826.345 189.04 826.625 329.185 ;
      RECT 825.785 189.04 826.065 328.945 ;
      RECT 825.225 189.04 825.505 328.705 ;
      RECT 824.665 189.04 824.945 328.465 ;
      RECT 824.105 189.04 824.385 328.225 ;
      RECT 823.545 189.04 823.825 327.985 ;
      RECT 822.985 187.94 823.265 327.745 ;
      RECT 822.425 189.04 822.705 327.505 ;
      RECT 821.865 187.94 822.145 327.265 ;
      RECT 782.665 189.04 782.945 332.875 ;
      RECT 782.105 189.04 782.385 333.115 ;
      RECT 781.545 189.04 781.825 333.355 ;
      RECT 780.985 189.04 781.265 333.595 ;
      RECT 780.425 189.04 780.705 333.835 ;
      RECT 779.865 189.04 780.145 334.075 ;
      RECT 779.305 189.04 779.585 334.315 ;
      RECT 778.745 189.04 779.025 334.555 ;
      RECT 778.185 189.04 778.465 334.795 ;
      RECT 777.625 189.04 777.905 335.035 ;
      RECT 777.065 189.04 777.345 335.275 ;
      RECT 776.505 189.04 776.785 335.515 ;
      RECT 775.945 189.04 776.225 335.755 ;
      RECT 775.385 189.04 775.665 335.755 ;
      RECT 774.825 187.94 775.105 335.515 ;
      RECT 774.265 189.04 774.545 335.275 ;
      RECT 773.705 187.94 773.985 335.035 ;
      RECT 773.145 189.04 773.425 334.795 ;
      RECT 772.585 189.04 772.865 334.555 ;
      RECT 772.025 189.04 772.305 334.315 ;
      RECT 771.465 187.94 771.745 334.05 ;
      RECT 770.905 189.04 771.185 333.81 ;
      RECT 770.345 187.94 770.625 333.57 ;
      RECT 769.785 189.04 770.065 333.33 ;
      RECT 760.825 187.94 761.105 327.165 ;
      RECT 760.265 189.04 760.545 327.405 ;
      RECT 759.705 189.04 759.985 327.645 ;
      RECT 759.145 189.04 759.425 327.645 ;
      RECT 758.585 189.04 758.865 327.405 ;
      RECT 758.025 189.04 758.305 327.165 ;
      RECT 757.465 189.04 757.745 326.925 ;
      RECT 756.905 189.04 757.185 326.685 ;
      RECT 756.345 189.04 756.625 326.445 ;
      RECT 755.785 189.04 756.065 326.205 ;
      RECT 755.225 189.04 755.505 325.965 ;
      RECT 754.665 189.04 754.945 325.725 ;
      RECT 754.105 189.04 754.385 325.485 ;
      RECT 753.545 187.94 753.825 325.245 ;
      RECT 751.025 189.04 751.305 326.965 ;
      RECT 750.465 187.94 750.745 326.725 ;
      RECT 749.905 189.04 750.185 326.485 ;
      RECT 749.345 187.94 749.625 326.245 ;
      RECT 748.785 189.04 749.065 326.005 ;
      RECT 748.225 189.04 748.505 325.765 ;
      RECT 747.665 189.04 747.945 325.525 ;
      RECT 721.625 189.04 721.905 328.31 ;
      RECT 721.065 189.04 721.345 328.55 ;
      RECT 720.505 189.04 720.785 328.79 ;
      RECT 719.945 189.04 720.225 329.03 ;
      RECT 719.385 189.04 719.665 329.27 ;
      RECT 718.825 187.94 719.105 329.51 ;
      RECT 718.265 189.04 718.545 329.75 ;
      RECT 717.705 187.94 717.985 329.99 ;
      RECT 717.145 189.04 717.425 330.23 ;
      RECT 716.585 189.04 716.865 330.47 ;
      RECT 716.025 189.04 716.305 330.71 ;
      RECT 715.465 189.04 715.745 330.95 ;
      RECT 714.905 189.04 715.185 331.19 ;
      RECT 714.345 189.04 714.625 331.43 ;
      RECT 713.785 189.04 714.065 331.67 ;
      RECT 713.225 189.04 713.505 331.67 ;
      RECT 712.665 189.04 712.945 331.43 ;
      RECT 712.105 189.04 712.385 331.19 ;
      RECT 711.545 189.04 711.825 330.95 ;
      RECT 710.985 189.04 711.265 330.705 ;
      RECT 710.425 189.04 710.705 330.465 ;
      RECT 709.865 189.04 710.145 330.225 ;
      RECT 709.305 187.94 709.585 329.985 ;
      RECT 708.745 189.04 709.025 329.745 ;
      RECT 695.305 187.94 695.585 327.225 ;
      RECT 694.745 189.04 695.025 326.985 ;
      RECT 694.185 189.04 694.465 326.745 ;
      RECT 693.625 189.04 693.905 326.505 ;
      RECT 693.065 187.94 693.345 326.265 ;
      RECT 692.505 189.04 692.785 326.025 ;
      RECT 691.945 187.94 692.225 325.785 ;
      RECT 691.385 189.04 691.665 325.545 ;
      RECT 690.825 187.94 691.105 325.305 ;
      RECT 690.265 189.04 690.545 325.065 ;
      RECT 689.705 189.04 689.985 324.825 ;
      RECT 689.145 189.04 689.425 324.585 ;
      RECT 688.585 189.04 688.865 324.345 ;
      RECT 688.025 189.04 688.305 324.105 ;
      RECT 687.465 189.04 687.745 323.865 ;
      RECT 686.905 189.04 687.185 323.625 ;
      RECT 686.345 189.04 686.625 323.385 ;
      RECT 685.785 189.04 686.065 323.145 ;
      RECT 685.225 189.04 685.505 322.905 ;
      RECT 684.665 189.04 684.945 322.665 ;
      RECT 684.105 189.04 684.385 322.425 ;
      RECT 683.545 187.94 683.825 322.185 ;
      RECT 682.985 189.04 683.265 321.945 ;
      RECT 682.425 187.94 682.705 321.705 ;
      RECT 642.665 189.04 642.945 332.175 ;
      RECT 642.105 187.94 642.385 332.415 ;
      RECT 641.545 189.04 641.825 332.655 ;
      RECT 640.985 189.04 641.265 332.895 ;
      RECT 640.425 189.04 640.705 333.135 ;
      RECT 639.865 189.04 640.145 333.375 ;
      RECT 639.305 189.04 639.585 333.615 ;
      RECT 638.745 189.04 639.025 333.86 ;
      RECT 638.185 189.04 638.465 334.1 ;
      RECT 637.625 189.04 637.905 334.34 ;
      RECT 637.065 187.94 637.345 334.58 ;
      RECT 636.505 189.04 636.785 334.82 ;
      RECT 635.945 187.94 636.225 335.06 ;
      RECT 635.385 189.04 635.665 335.3 ;
      RECT 634.825 189.04 635.105 335.54 ;
      RECT 634.265 189.04 634.545 335.78 ;
      RECT 633.705 189.04 633.985 336.02 ;
      RECT 633.145 189.04 633.425 336.26 ;
      RECT 632.585 189.04 632.865 336.5 ;
      RECT 632.025 189.04 632.305 336.74 ;
      RECT 631.465 189.04 631.745 336.98 ;
      RECT 630.905 189.04 631.185 337.22 ;
      RECT 630.345 189.04 630.625 337.46 ;
      RECT 629.785 189.04 630.065 337.7 ;
      RECT 620.825 189.04 621.105 333.285 ;
      RECT 620.265 189.04 620.545 333.045 ;
      RECT 619.705 189.04 619.985 332.805 ;
      RECT 619.145 187.94 619.425 332.565 ;
      RECT 618.585 189.04 618.865 332.325 ;
      RECT 618.025 187.94 618.305 332.085 ;
      RECT 617.465 189.04 617.745 331.845 ;
      RECT 616.905 189.04 617.185 331.605 ;
      RECT 616.345 189.04 616.625 331.365 ;
      RECT 615.785 187.94 616.065 331.125 ;
      RECT 615.225 189.04 615.505 330.885 ;
      RECT 614.665 187.94 614.945 330.645 ;
      RECT 614.105 189.04 614.385 330.405 ;
      RECT 613.545 187.94 613.825 330.165 ;
      RECT 611.025 189.04 611.305 322.565 ;
      RECT 610.465 189.04 610.745 322.325 ;
      RECT 609.905 189.04 610.185 322.085 ;
      RECT 609.345 189.04 609.625 321.845 ;
      RECT 608.785 189.04 609.065 321.605 ;
      RECT 608.225 189.04 608.505 321.365 ;
      RECT 607.665 189.04 607.945 321.125 ;
      RECT 581.625 189.04 581.905 335 ;
      RECT 581.065 189.04 581.345 335.24 ;
      RECT 580.505 189.04 580.785 335.48 ;
      RECT 579.945 189.04 580.225 335.72 ;
      RECT 579.385 189.04 579.665 335.96 ;
      RECT 578.825 187.94 579.105 335.96 ;
      RECT 578.265 189.04 578.545 335.72 ;
      RECT 577.705 187.94 577.985 335.475 ;
      RECT 577.145 189.04 577.425 335.235 ;
      RECT 576.585 187.94 576.865 334.995 ;
      RECT 576.025 189.04 576.305 334.755 ;
      RECT 575.465 189.04 575.745 334.515 ;
      RECT 574.905 189.04 575.185 334.275 ;
      RECT 574.345 189.04 574.625 334.035 ;
      RECT 573.785 189.04 574.065 333.795 ;
      RECT 573.225 189.04 573.505 333.555 ;
      RECT 572.665 189.04 572.945 333.315 ;
      RECT 572.105 189.04 572.385 333.075 ;
      RECT 571.545 187.94 571.825 332.835 ;
      RECT 570.985 189.04 571.265 332.595 ;
      RECT 570.425 187.94 570.705 332.355 ;
      RECT 569.865 189.04 570.145 332.115 ;
      RECT 569.305 189.04 569.585 331.875 ;
      RECT 568.745 189.04 569.025 331.635 ;
      RECT 555.305 189.04 555.585 335.035 ;
      RECT 554.745 189.04 555.025 335.275 ;
      RECT 554.185 189.04 554.465 335.52 ;
      RECT 553.625 189.04 553.905 335.76 ;
      RECT 553.065 189.04 553.345 336 ;
      RECT 552.505 189.04 552.785 336 ;
      RECT 551.945 189.04 552.225 335.76 ;
      RECT 551.385 189.04 551.665 335.52 ;
      RECT 550.825 189.04 551.105 328.505 ;
      RECT 550.265 189.04 550.545 328.265 ;
      RECT 549.705 189.04 549.985 328.025 ;
      RECT 549.145 187.94 549.425 327.785 ;
      RECT 548.585 189.04 548.865 327.545 ;
      RECT 548.025 187.94 548.305 327.305 ;
      RECT 547.465 189.04 547.745 327.065 ;
      RECT 546.905 189.04 547.185 326.825 ;
      RECT 546.345 189.04 546.625 326.585 ;
      RECT 545.785 187.94 546.065 326.345 ;
      RECT 545.225 189.04 545.505 326.105 ;
      RECT 544.665 187.94 544.945 325.865 ;
      RECT 544.105 189.04 544.385 325.625 ;
      RECT 543.545 187.94 543.825 325.385 ;
      RECT 542.985 189.04 543.265 325.145 ;
      RECT 542.425 189.04 542.705 324.905 ;
      RECT 502.105 189.04 502.385 333.8 ;
      RECT 501.545 189.04 501.825 334.04 ;
      RECT 500.985 189.04 501.265 334.285 ;
      RECT 500.425 189.04 500.705 334.525 ;
      RECT 499.865 189.04 500.145 334.765 ;
      RECT 499.305 189.04 499.585 335.005 ;
      RECT 498.745 189.04 499.025 335.245 ;
      RECT 498.185 189.04 498.465 335.485 ;
      RECT 497.625 189.04 497.905 335.725 ;
      RECT 497.065 189.04 497.345 335.965 ;
      RECT 496.505 187.94 496.785 336.205 ;
      RECT 495.945 189.04 496.225 336.445 ;
      RECT 495.385 187.94 495.665 336.685 ;
      RECT 494.825 189.04 495.105 336.925 ;
      RECT 494.265 187.94 494.545 337.165 ;
      RECT 493.705 189.04 493.985 337.165 ;
      RECT 493.145 189.04 493.425 336.925 ;
      RECT 492.585 189.04 492.865 336.685 ;
      RECT 492.025 189.04 492.305 336.445 ;
      RECT 491.465 189.04 491.745 336.205 ;
      RECT 490.905 189.04 491.185 335.965 ;
      RECT 490.345 189.04 490.625 335.725 ;
      RECT 489.785 189.04 490.065 335.485 ;
      RECT 480.825 187.94 481.105 335.515 ;
      RECT 480.265 189.04 480.545 335.755 ;
      RECT 479.705 187.94 479.985 335.995 ;
      RECT 479.145 189.04 479.425 336.21 ;
      RECT 478.585 189.04 478.865 335.785 ;
      RECT 478.025 189.04 478.305 335.545 ;
      RECT 477.465 189.04 477.745 335.305 ;
      RECT 476.905 189.04 477.185 335.065 ;
      RECT 476.345 189.04 476.625 334.825 ;
      RECT 475.785 189.04 476.065 334.585 ;
      RECT 475.225 189.04 475.505 334.345 ;
      RECT 474.665 189.04 474.945 334.105 ;
      RECT 474.105 189.04 474.385 333.865 ;
      RECT 473.545 189.04 473.825 333.625 ;
      RECT 471.025 189.04 471.305 332.8 ;
      RECT 470.465 189.04 470.745 332.56 ;
      RECT 469.905 189.04 470.185 332.32 ;
      RECT 469.345 187.94 469.625 332.08 ;
      RECT 468.785 189.04 469.065 331.84 ;
      RECT 468.225 187.94 468.505 331.6 ;
      RECT 467.665 189.04 467.945 331.36 ;
      RECT 467.105 189.04 467.385 331.12 ;
      RECT 466.545 189.04 466.825 295.135 ;
      RECT 328.26 8399.58 351.33 8401 ;
      RECT 328.26 8438.095 351.33 8439.515 ;
      RECT 328.26 8471.58 351.33 8473 ;
      RECT 328.26 8510.095 351.33 8511.515 ;
      RECT 328.26 8543.58 351.33 8545 ;
      RECT 328.26 8582.095 351.33 8583.515 ;
    LAYER M4 SPACING 0.28 ;
      RECT 13498.305 8583.935 18490.46 8613.565 ;
      RECT 13498.305 188.86 18489.04 8613.565 ;
      RECT 13498.305 8545.42 18490.46 8581.675 ;
      RECT 13498.305 8511.935 18490.46 8543.16 ;
      RECT 13498.305 8473.42 18490.46 8509.675 ;
      RECT 13498.305 8439.935 18490.46 8471.16 ;
      RECT 13498.305 8401.42 18490.46 8437.675 ;
      RECT 18361.765 187.44 18490.46 8399.16 ;
      RECT 18359.945 187.94 18360.225 8613.565 ;
      RECT 18358.825 187.94 18359.105 8613.565 ;
      RECT 18357.705 187.94 18357.985 8613.565 ;
      RECT 18350.425 187.94 18350.705 8613.565 ;
      RECT 18349.305 187.94 18349.585 8613.565 ;
      RECT 18334.745 187.94 18348.325 8613.565 ;
      RECT 18334.885 187.44 18348.325 8613.565 ;
      RECT 18329.705 187.94 18329.985 8613.565 ;
      RECT 18328.585 187.94 18328.865 8613.565 ;
      RECT 18283.925 187.44 18322.005 8613.565 ;
      RECT 18281.545 187.94 18281.825 8613.565 ;
      RECT 18280.425 187.94 18280.705 8613.565 ;
      RECT 18278.185 187.94 18278.465 8613.565 ;
      RECT 18277.065 187.94 18277.345 8613.565 ;
      RECT 18275.945 187.94 18276.225 8613.565 ;
      RECT 18261.525 187.44 18269.365 8613.565 ;
      RECT 18260.265 187.94 18260.545 8613.565 ;
      RECT 18259.145 187.94 18259.425 8613.565 ;
      RECT 18258.025 187.94 18258.305 8613.565 ;
      RECT 18251.025 187.94 18253.125 8613.565 ;
      RECT 18251.165 187.44 18253.125 8613.565 ;
      RECT 18249.905 187.94 18250.185 8613.565 ;
      RECT 18221.765 187.44 18246.685 8613.565 ;
      RECT 18216.025 187.94 18216.305 8613.565 ;
      RECT 18214.905 187.94 18215.185 8613.565 ;
      RECT 18212.665 187.94 18212.945 8613.565 ;
      RECT 18211.545 187.94 18211.825 8613.565 ;
      RECT 18210.425 187.94 18210.705 8613.565 ;
      RECT 18195.445 187.44 18207.765 8613.565 ;
      RECT 18190.265 187.94 18190.545 8613.565 ;
      RECT 18189.145 187.94 18189.425 8613.565 ;
      RECT 18188.025 187.94 18188.305 8613.565 ;
      RECT 18182.985 187.94 18183.265 8613.565 ;
      RECT 18143.365 187.94 18182.145 8613.565 ;
      RECT 18134.825 187.94 18135.105 8613.565 ;
      RECT 18133.705 187.94 18133.985 8613.565 ;
      RECT 18131.465 187.94 18131.745 8613.565 ;
      RECT 18130.345 187.94 18130.625 8613.565 ;
      RECT 18120.825 187.94 18129.365 8613.565 ;
      RECT 18120.965 187.44 18129.365 8613.565 ;
      RECT 18111.725 187.94 18113.825 8613.565 ;
      RECT 18110.465 187.94 18110.745 8613.565 ;
      RECT 18109.345 187.94 18109.625 8613.565 ;
      RECT 18082.325 187.44 18107.245 8613.565 ;
      RECT 18078.825 187.94 18079.105 8613.565 ;
      RECT 18077.705 187.94 18077.985 8613.565 ;
      RECT 18069.305 187.94 18069.585 8613.565 ;
      RECT 18055.305 187.94 18068.325 8613.565 ;
      RECT 18055.445 187.44 18068.325 8613.565 ;
      RECT 18053.065 187.94 18053.345 8613.565 ;
      RECT 18051.945 187.94 18052.225 8613.565 ;
      RECT 18050.825 187.94 18051.105 8613.565 ;
      RECT 18043.545 187.94 18043.825 8613.565 ;
      RECT 18003.365 187.94 18042.705 8613.565 ;
      RECT 18002.105 187.94 18002.385 8613.565 ;
      RECT 17997.065 187.94 17997.345 8613.565 ;
      RECT 17995.945 187.94 17996.225 8613.565 ;
      RECT 17981.525 187.44 17989.365 8613.565 ;
      RECT 17979.145 187.94 17979.425 8613.565 ;
      RECT 17978.025 187.94 17978.305 8613.565 ;
      RECT 17975.785 187.94 17976.065 8613.565 ;
      RECT 17974.665 187.94 17974.945 8613.565 ;
      RECT 17971.725 187.94 17973.825 8613.565 ;
      RECT 17942.325 187.44 17967.245 8613.565 ;
      RECT 17938.825 187.94 17939.105 8613.565 ;
      RECT 17937.705 187.94 17937.985 8613.565 ;
      RECT 17936.585 187.94 17936.865 8613.565 ;
      RECT 17931.545 187.94 17931.825 8613.565 ;
      RECT 17930.425 187.94 17930.705 8613.565 ;
      RECT 17916.005 187.44 17928.325 8613.565 ;
      RECT 17909.145 187.94 17909.425 8613.565 ;
      RECT 17908.025 187.94 17908.305 8613.565 ;
      RECT 17905.785 187.94 17906.065 8613.565 ;
      RECT 17904.665 187.94 17904.945 8613.565 ;
      RECT 17903.545 187.94 17903.825 8613.565 ;
      RECT 17862.805 187.44 17902.005 8613.565 ;
      RECT 17856.505 187.94 17856.785 8613.565 ;
      RECT 17855.385 187.94 17855.665 8613.565 ;
      RECT 17854.265 187.94 17854.545 8613.565 ;
      RECT 17840.825 187.94 17849.365 8613.565 ;
      RECT 17840.965 187.44 17849.365 8613.565 ;
      RECT 17839.705 187.94 17839.985 8613.565 ;
      RECT 17831.725 187.44 17833.125 8613.565 ;
      RECT 17829.345 187.94 17829.625 8613.565 ;
      RECT 17828.225 187.94 17828.505 8613.565 ;
      RECT 17801.205 187.44 17826.685 8613.565 ;
      RECT 17799.945 187.94 17800.225 8613.565 ;
      RECT 17798.825 187.94 17799.105 8613.565 ;
      RECT 17797.705 187.94 17797.985 8613.565 ;
      RECT 17790.425 187.94 17790.705 8613.565 ;
      RECT 17789.305 187.94 17789.585 8613.565 ;
      RECT 17774.745 187.94 17788.325 8613.565 ;
      RECT 17774.885 187.44 17788.325 8613.565 ;
      RECT 17769.705 187.94 17769.985 8613.565 ;
      RECT 17768.585 187.94 17768.865 8613.565 ;
      RECT 17723.925 187.44 17762.005 8613.565 ;
      RECT 17721.545 187.94 17721.825 8613.565 ;
      RECT 17720.425 187.94 17720.705 8613.565 ;
      RECT 17718.185 187.94 17718.465 8613.565 ;
      RECT 17717.065 187.94 17717.345 8613.565 ;
      RECT 17715.945 187.94 17716.225 8613.565 ;
      RECT 17701.525 187.44 17709.365 8613.565 ;
      RECT 17700.265 187.94 17700.545 8613.565 ;
      RECT 17699.145 187.94 17699.425 8613.565 ;
      RECT 17698.025 187.94 17698.305 8613.565 ;
      RECT 17691.025 187.94 17693.125 8613.565 ;
      RECT 17691.165 187.44 17693.125 8613.565 ;
      RECT 17689.905 187.94 17690.185 8613.565 ;
      RECT 17661.765 187.44 17686.685 8613.565 ;
      RECT 17656.025 187.94 17656.305 8613.565 ;
      RECT 17654.905 187.94 17655.185 8613.565 ;
      RECT 17652.665 187.94 17652.945 8613.565 ;
      RECT 17651.545 187.94 17651.825 8613.565 ;
      RECT 17650.425 187.94 17650.705 8613.565 ;
      RECT 17635.445 187.44 17647.765 8613.565 ;
      RECT 17630.265 187.94 17630.545 8613.565 ;
      RECT 17629.145 187.94 17629.425 8613.565 ;
      RECT 17628.025 187.94 17628.305 8613.565 ;
      RECT 17622.985 187.94 17623.265 8613.565 ;
      RECT 17583.365 187.94 17622.145 8613.565 ;
      RECT 17574.825 187.94 17575.105 8613.565 ;
      RECT 17573.705 187.94 17573.985 8613.565 ;
      RECT 17571.465 187.94 17571.745 8613.565 ;
      RECT 17570.345 187.94 17570.625 8613.565 ;
      RECT 17560.825 187.94 17569.365 8613.565 ;
      RECT 17560.965 187.44 17569.365 8613.565 ;
      RECT 17551.725 187.94 17553.825 8613.565 ;
      RECT 17550.465 187.94 17550.745 8613.565 ;
      RECT 17549.345 187.94 17549.625 8613.565 ;
      RECT 17522.325 187.44 17547.245 8613.565 ;
      RECT 17518.825 187.94 17519.105 8613.565 ;
      RECT 17517.705 187.94 17517.985 8613.565 ;
      RECT 17509.305 187.94 17509.585 8613.565 ;
      RECT 17495.305 187.94 17508.325 8613.565 ;
      RECT 17495.445 187.44 17508.325 8613.565 ;
      RECT 17493.065 187.94 17493.345 8613.565 ;
      RECT 17491.945 187.94 17492.225 8613.565 ;
      RECT 17490.825 187.94 17491.105 8613.565 ;
      RECT 17483.545 187.94 17483.825 8613.565 ;
      RECT 17443.365 187.94 17482.705 8613.565 ;
      RECT 17442.105 187.94 17442.385 8613.565 ;
      RECT 17437.065 187.94 17437.345 8613.565 ;
      RECT 17435.945 187.94 17436.225 8613.565 ;
      RECT 17421.525 187.44 17429.365 8613.565 ;
      RECT 17419.145 187.94 17419.425 8613.565 ;
      RECT 17418.025 187.94 17418.305 8613.565 ;
      RECT 17415.785 187.94 17416.065 8613.565 ;
      RECT 17414.665 187.94 17414.945 8613.565 ;
      RECT 17411.725 187.94 17413.825 8613.565 ;
      RECT 17382.325 187.44 17407.245 8613.565 ;
      RECT 17378.825 187.94 17379.105 8613.565 ;
      RECT 17377.705 187.94 17377.985 8613.565 ;
      RECT 17376.585 187.94 17376.865 8613.565 ;
      RECT 17371.545 187.94 17371.825 8613.565 ;
      RECT 17370.425 187.94 17370.705 8613.565 ;
      RECT 17356.005 187.44 17368.325 8613.565 ;
      RECT 17349.145 187.94 17349.425 8613.565 ;
      RECT 17348.025 187.94 17348.305 8613.565 ;
      RECT 17345.785 187.94 17346.065 8613.565 ;
      RECT 17344.665 187.94 17344.945 8613.565 ;
      RECT 17343.545 187.94 17343.825 8613.565 ;
      RECT 17302.805 187.44 17342.005 8613.565 ;
      RECT 17296.505 187.94 17296.785 8613.565 ;
      RECT 17295.385 187.94 17295.665 8613.565 ;
      RECT 17294.265 187.94 17294.545 8613.565 ;
      RECT 17280.825 187.94 17289.365 8613.565 ;
      RECT 17280.965 187.44 17289.365 8613.565 ;
      RECT 17279.705 187.94 17279.985 8613.565 ;
      RECT 17271.725 187.44 17273.125 8613.565 ;
      RECT 17269.345 187.94 17269.625 8613.565 ;
      RECT 17268.225 187.94 17268.505 8613.565 ;
      RECT 17241.205 187.44 17266.685 8613.565 ;
      RECT 17239.945 187.94 17240.225 8613.565 ;
      RECT 17238.825 187.94 17239.105 8613.565 ;
      RECT 17237.705 187.94 17237.985 8613.565 ;
      RECT 17230.425 187.94 17230.705 8613.565 ;
      RECT 17229.305 187.94 17229.585 8613.565 ;
      RECT 17214.745 187.94 17228.325 8613.565 ;
      RECT 17214.885 187.44 17228.325 8613.565 ;
      RECT 17209.705 187.94 17209.985 8613.565 ;
      RECT 17208.585 187.94 17208.865 8613.565 ;
      RECT 17163.925 187.44 17202.005 8613.565 ;
      RECT 17161.545 187.94 17161.825 8613.565 ;
      RECT 17160.425 187.94 17160.705 8613.565 ;
      RECT 17158.185 187.94 17158.465 8613.565 ;
      RECT 17157.065 187.94 17157.345 8613.565 ;
      RECT 17155.945 187.94 17156.225 8613.565 ;
      RECT 17141.525 187.44 17149.365 8613.565 ;
      RECT 17140.265 187.94 17140.545 8613.565 ;
      RECT 17139.145 187.94 17139.425 8613.565 ;
      RECT 17138.025 187.94 17138.305 8613.565 ;
      RECT 17131.025 187.94 17133.125 8613.565 ;
      RECT 17131.165 187.44 17133.125 8613.565 ;
      RECT 17129.905 187.94 17130.185 8613.565 ;
      RECT 17101.765 187.44 17126.685 8613.565 ;
      RECT 17096.025 187.94 17096.305 8613.565 ;
      RECT 17094.905 187.94 17095.185 8613.565 ;
      RECT 17092.665 187.94 17092.945 8613.565 ;
      RECT 17091.545 187.94 17091.825 8613.565 ;
      RECT 17090.425 187.94 17090.705 8613.565 ;
      RECT 17075.445 187.44 17087.765 8613.565 ;
      RECT 17070.265 187.94 17070.545 8613.565 ;
      RECT 17069.145 187.94 17069.425 8613.565 ;
      RECT 17068.025 187.94 17068.305 8613.565 ;
      RECT 17062.985 187.94 17063.265 8613.565 ;
      RECT 17023.365 187.94 17062.145 8613.565 ;
      RECT 17014.825 187.94 17015.105 8613.565 ;
      RECT 17013.705 187.94 17013.985 8613.565 ;
      RECT 17011.465 187.94 17011.745 8613.565 ;
      RECT 17010.345 187.94 17010.625 8613.565 ;
      RECT 17000.825 187.94 17009.365 8613.565 ;
      RECT 17000.965 187.44 17009.365 8613.565 ;
      RECT 16991.725 187.94 16993.825 8613.565 ;
      RECT 16990.465 187.94 16990.745 8613.565 ;
      RECT 16989.345 187.94 16989.625 8613.565 ;
      RECT 16962.325 187.44 16987.245 8613.565 ;
      RECT 16958.825 187.94 16959.105 8613.565 ;
      RECT 16957.705 187.94 16957.985 8613.565 ;
      RECT 16949.305 187.94 16949.585 8613.565 ;
      RECT 16935.305 187.94 16948.325 8613.565 ;
      RECT 16935.445 187.44 16948.325 8613.565 ;
      RECT 16933.065 187.94 16933.345 8613.565 ;
      RECT 16931.945 187.94 16932.225 8613.565 ;
      RECT 16930.825 187.94 16931.105 8613.565 ;
      RECT 16923.545 187.94 16923.825 8613.565 ;
      RECT 16883.365 187.94 16922.705 8613.565 ;
      RECT 16882.105 187.94 16882.385 8613.565 ;
      RECT 16877.065 187.94 16877.345 8613.565 ;
      RECT 16875.945 187.94 16876.225 8613.565 ;
      RECT 16861.525 187.44 16869.365 8613.565 ;
      RECT 16859.145 187.94 16859.425 8613.565 ;
      RECT 16858.025 187.94 16858.305 8613.565 ;
      RECT 16855.785 187.94 16856.065 8613.565 ;
      RECT 16854.665 187.94 16854.945 8613.565 ;
      RECT 16851.725 187.94 16853.825 8613.565 ;
      RECT 16822.325 187.44 16847.245 8613.565 ;
      RECT 16818.825 187.94 16819.105 8613.565 ;
      RECT 16817.705 187.94 16817.985 8613.565 ;
      RECT 16816.585 187.94 16816.865 8613.565 ;
      RECT 16811.545 187.94 16811.825 8613.565 ;
      RECT 16810.425 187.94 16810.705 8613.565 ;
      RECT 16796.005 187.44 16808.325 8613.565 ;
      RECT 16789.145 187.94 16789.425 8613.565 ;
      RECT 16788.025 187.94 16788.305 8613.565 ;
      RECT 16785.785 187.94 16786.065 8613.565 ;
      RECT 16784.665 187.94 16784.945 8613.565 ;
      RECT 16783.545 187.94 16783.825 8613.565 ;
      RECT 16742.805 187.44 16782.005 8613.565 ;
      RECT 16736.505 187.94 16736.785 8613.565 ;
      RECT 16735.385 187.94 16735.665 8613.565 ;
      RECT 16734.265 187.94 16734.545 8613.565 ;
      RECT 16720.825 187.94 16729.365 8613.565 ;
      RECT 16720.965 187.44 16729.365 8613.565 ;
      RECT 16719.705 187.94 16719.985 8613.565 ;
      RECT 16711.725 187.44 16713.125 8613.565 ;
      RECT 16709.345 187.94 16709.625 8613.565 ;
      RECT 16708.225 187.94 16708.505 8613.565 ;
      RECT 16681.205 187.44 16706.685 8613.565 ;
      RECT 16679.945 187.94 16680.225 8613.565 ;
      RECT 16678.825 187.94 16679.105 8613.565 ;
      RECT 16677.705 187.94 16677.985 8613.565 ;
      RECT 16670.425 187.94 16670.705 8613.565 ;
      RECT 16669.305 187.94 16669.585 8613.565 ;
      RECT 16654.745 187.94 16668.325 8613.565 ;
      RECT 16654.885 187.44 16668.325 8613.565 ;
      RECT 16649.705 187.94 16649.985 8613.565 ;
      RECT 16648.585 187.94 16648.865 8613.565 ;
      RECT 16603.925 187.44 16642.005 8613.565 ;
      RECT 16601.545 187.94 16601.825 8613.565 ;
      RECT 16600.425 187.94 16600.705 8613.565 ;
      RECT 16598.185 187.94 16598.465 8613.565 ;
      RECT 16597.065 187.94 16597.345 8613.565 ;
      RECT 16595.945 187.94 16596.225 8613.565 ;
      RECT 16581.525 187.44 16589.365 8613.565 ;
      RECT 16580.265 187.94 16580.545 8613.565 ;
      RECT 16579.145 187.94 16579.425 8613.565 ;
      RECT 16578.025 187.94 16578.305 8613.565 ;
      RECT 16571.025 187.94 16573.125 8613.565 ;
      RECT 16571.165 187.44 16573.125 8613.565 ;
      RECT 16569.905 187.94 16570.185 8613.565 ;
      RECT 16541.765 187.44 16566.685 8613.565 ;
      RECT 16536.025 187.94 16536.305 8613.565 ;
      RECT 16534.905 187.94 16535.185 8613.565 ;
      RECT 16532.665 187.94 16532.945 8613.565 ;
      RECT 16531.545 187.94 16531.825 8613.565 ;
      RECT 16530.425 187.94 16530.705 8613.565 ;
      RECT 16515.445 187.44 16527.765 8613.565 ;
      RECT 16510.265 187.94 16510.545 8613.565 ;
      RECT 16509.145 187.94 16509.425 8613.565 ;
      RECT 16508.025 187.94 16508.305 8613.565 ;
      RECT 16502.985 187.94 16503.265 8613.565 ;
      RECT 16463.365 187.94 16502.145 8613.565 ;
      RECT 16454.825 187.94 16455.105 8613.565 ;
      RECT 16453.705 187.94 16453.985 8613.565 ;
      RECT 16451.465 187.94 16451.745 8613.565 ;
      RECT 16450.345 187.94 16450.625 8613.565 ;
      RECT 16440.825 187.94 16449.365 8613.565 ;
      RECT 16440.965 187.44 16449.365 8613.565 ;
      RECT 16431.725 187.94 16433.825 8613.565 ;
      RECT 16430.465 187.94 16430.745 8613.565 ;
      RECT 16429.345 187.94 16429.625 8613.565 ;
      RECT 16402.325 187.44 16427.245 8613.565 ;
      RECT 16398.825 187.94 16399.105 8613.565 ;
      RECT 16397.705 187.94 16397.985 8613.565 ;
      RECT 16389.305 187.94 16389.585 8613.565 ;
      RECT 16375.305 187.94 16388.325 8613.565 ;
      RECT 16375.445 187.44 16388.325 8613.565 ;
      RECT 16373.065 187.94 16373.345 8613.565 ;
      RECT 16371.945 187.94 16372.225 8613.565 ;
      RECT 16370.825 187.94 16371.105 8613.565 ;
      RECT 16363.545 187.94 16363.825 8613.565 ;
      RECT 16323.365 187.94 16362.705 8613.565 ;
      RECT 16322.105 187.94 16322.385 8613.565 ;
      RECT 16317.065 187.94 16317.345 8613.565 ;
      RECT 16315.945 187.94 16316.225 8613.565 ;
      RECT 16301.525 187.44 16309.365 8613.565 ;
      RECT 16299.145 187.94 16299.425 8613.565 ;
      RECT 16298.025 187.94 16298.305 8613.565 ;
      RECT 16295.785 187.94 16296.065 8613.565 ;
      RECT 16294.665 187.94 16294.945 8613.565 ;
      RECT 16291.725 187.94 16293.825 8613.565 ;
      RECT 16262.325 187.44 16287.245 8613.565 ;
      RECT 16258.825 187.94 16259.105 8613.565 ;
      RECT 16257.705 187.94 16257.985 8613.565 ;
      RECT 16256.585 187.94 16256.865 8613.565 ;
      RECT 16251.545 187.94 16251.825 8613.565 ;
      RECT 16250.425 187.94 16250.705 8613.565 ;
      RECT 16236.005 187.44 16248.325 8613.565 ;
      RECT 16229.145 187.94 16229.425 8613.565 ;
      RECT 16228.025 187.94 16228.305 8613.565 ;
      RECT 16225.785 187.94 16226.065 8613.565 ;
      RECT 16224.665 187.94 16224.945 8613.565 ;
      RECT 16223.545 187.94 16223.825 8613.565 ;
      RECT 16182.805 187.44 16222.005 8613.565 ;
      RECT 16176.505 187.94 16176.785 8613.565 ;
      RECT 16175.385 187.94 16175.665 8613.565 ;
      RECT 16174.265 187.94 16174.545 8613.565 ;
      RECT 16160.825 187.94 16169.365 8613.565 ;
      RECT 16160.965 187.44 16169.365 8613.565 ;
      RECT 16159.705 187.94 16159.985 8613.565 ;
      RECT 16151.725 187.44 16153.125 8613.565 ;
      RECT 16149.345 187.94 16149.625 8613.565 ;
      RECT 16148.225 187.94 16148.505 8613.565 ;
      RECT 16121.205 187.44 16146.685 8613.565 ;
      RECT 16119.945 187.94 16120.225 8613.565 ;
      RECT 16118.825 187.94 16119.105 8613.565 ;
      RECT 16117.705 187.94 16117.985 8613.565 ;
      RECT 16110.425 187.94 16110.705 8613.565 ;
      RECT 16109.305 187.94 16109.585 8613.565 ;
      RECT 16094.745 187.94 16108.325 8613.565 ;
      RECT 16094.885 187.44 16108.325 8613.565 ;
      RECT 16089.705 187.94 16089.985 8613.565 ;
      RECT 16088.585 187.94 16088.865 8613.565 ;
      RECT 16043.925 187.44 16082.005 8613.565 ;
      RECT 16041.545 187.94 16041.825 8613.565 ;
      RECT 16040.425 187.94 16040.705 8613.565 ;
      RECT 16038.185 187.94 16038.465 8613.565 ;
      RECT 16037.065 187.94 16037.345 8613.565 ;
      RECT 16035.945 187.94 16036.225 8613.565 ;
      RECT 16021.525 187.44 16029.365 8613.565 ;
      RECT 16020.265 187.94 16020.545 8613.565 ;
      RECT 16019.145 187.94 16019.425 8613.565 ;
      RECT 16018.025 187.94 16018.305 8613.565 ;
      RECT 16011.025 187.94 16013.125 8613.565 ;
      RECT 16011.165 187.44 16013.125 8613.565 ;
      RECT 16009.905 187.94 16010.185 8613.565 ;
      RECT 15981.765 187.44 16006.685 8613.565 ;
      RECT 15976.025 187.94 15976.305 8613.565 ;
      RECT 15974.905 187.94 15975.185 8613.565 ;
      RECT 15972.665 187.94 15972.945 8613.565 ;
      RECT 15971.545 187.94 15971.825 8613.565 ;
      RECT 15970.425 187.94 15970.705 8613.565 ;
      RECT 15955.445 187.44 15967.765 8613.565 ;
      RECT 15950.265 187.94 15950.545 8613.565 ;
      RECT 15949.145 187.94 15949.425 8613.565 ;
      RECT 15948.025 187.94 15948.305 8613.565 ;
      RECT 15942.985 187.94 15943.265 8613.565 ;
      RECT 15903.365 187.94 15942.145 8613.565 ;
      RECT 15894.825 187.94 15895.105 8613.565 ;
      RECT 15893.705 187.94 15893.985 8613.565 ;
      RECT 15891.465 187.94 15891.745 8613.565 ;
      RECT 15890.345 187.94 15890.625 8613.565 ;
      RECT 15880.825 187.94 15889.365 8613.565 ;
      RECT 15880.965 187.44 15889.365 8613.565 ;
      RECT 15871.725 187.94 15873.825 8613.565 ;
      RECT 15870.465 187.94 15870.745 8613.565 ;
      RECT 15869.345 187.94 15869.625 8613.565 ;
      RECT 15842.325 187.44 15867.245 8613.565 ;
      RECT 15838.825 187.94 15839.105 8613.565 ;
      RECT 15837.705 187.94 15837.985 8613.565 ;
      RECT 15829.305 187.94 15829.585 8613.565 ;
      RECT 15815.305 187.94 15828.325 8613.565 ;
      RECT 15815.445 187.44 15828.325 8613.565 ;
      RECT 15813.065 187.94 15813.345 8613.565 ;
      RECT 15811.945 187.94 15812.225 8613.565 ;
      RECT 15810.825 187.94 15811.105 8613.565 ;
      RECT 15803.545 187.94 15803.825 8613.565 ;
      RECT 15763.365 187.94 15802.705 8613.565 ;
      RECT 15762.105 187.94 15762.385 8613.565 ;
      RECT 15757.065 187.94 15757.345 8613.565 ;
      RECT 15755.945 187.94 15756.225 8613.565 ;
      RECT 15741.525 187.44 15749.365 8613.565 ;
      RECT 15739.145 187.94 15739.425 8613.565 ;
      RECT 15738.025 187.94 15738.305 8613.565 ;
      RECT 15735.785 187.94 15736.065 8613.565 ;
      RECT 15734.665 187.94 15734.945 8613.565 ;
      RECT 15731.725 187.94 15733.825 8613.565 ;
      RECT 15702.325 187.44 15727.245 8613.565 ;
      RECT 15698.825 187.94 15699.105 8613.565 ;
      RECT 15697.705 187.94 15697.985 8613.565 ;
      RECT 15696.585 187.94 15696.865 8613.565 ;
      RECT 15691.545 187.94 15691.825 8613.565 ;
      RECT 15690.425 187.94 15690.705 8613.565 ;
      RECT 15676.005 187.44 15688.325 8613.565 ;
      RECT 15669.145 187.94 15669.425 8613.565 ;
      RECT 15668.025 187.94 15668.305 8613.565 ;
      RECT 15665.785 187.94 15666.065 8613.565 ;
      RECT 15664.665 187.94 15664.945 8613.565 ;
      RECT 15663.545 187.94 15663.825 8613.565 ;
      RECT 15622.805 187.44 15662.005 8613.565 ;
      RECT 15616.505 187.94 15616.785 8613.565 ;
      RECT 15615.385 187.94 15615.665 8613.565 ;
      RECT 15614.265 187.94 15614.545 8613.565 ;
      RECT 15600.825 187.94 15609.365 8613.565 ;
      RECT 15600.965 187.44 15609.365 8613.565 ;
      RECT 15599.705 187.94 15599.985 8613.565 ;
      RECT 15591.725 187.44 15593.125 8613.565 ;
      RECT 15589.345 187.94 15589.625 8613.565 ;
      RECT 15588.225 187.94 15588.505 8613.565 ;
      RECT 15561.205 187.44 15586.685 8613.565 ;
      RECT 15559.945 187.94 15560.225 8613.565 ;
      RECT 15558.825 187.94 15559.105 8613.565 ;
      RECT 15557.705 187.94 15557.985 8613.565 ;
      RECT 15550.425 187.94 15550.705 8613.565 ;
      RECT 15549.305 187.94 15549.585 8613.565 ;
      RECT 15534.745 187.94 15548.325 8613.565 ;
      RECT 15534.885 187.44 15548.325 8613.565 ;
      RECT 15529.705 187.94 15529.985 8613.565 ;
      RECT 15528.585 187.94 15528.865 8613.565 ;
      RECT 15483.925 187.44 15522.005 8613.565 ;
      RECT 15481.545 187.94 15481.825 8613.565 ;
      RECT 15480.425 187.94 15480.705 8613.565 ;
      RECT 15478.185 187.94 15478.465 8613.565 ;
      RECT 15477.065 187.94 15477.345 8613.565 ;
      RECT 15475.945 187.94 15476.225 8613.565 ;
      RECT 15461.525 187.44 15469.365 8613.565 ;
      RECT 15460.265 187.94 15460.545 8613.565 ;
      RECT 15459.145 187.94 15459.425 8613.565 ;
      RECT 15458.025 187.94 15458.305 8613.565 ;
      RECT 15451.025 187.94 15453.125 8613.565 ;
      RECT 15451.165 187.44 15453.125 8613.565 ;
      RECT 15449.905 187.94 15450.185 8613.565 ;
      RECT 15421.765 187.44 15446.685 8613.565 ;
      RECT 15416.025 187.94 15416.305 8613.565 ;
      RECT 15414.905 187.94 15415.185 8613.565 ;
      RECT 15412.665 187.94 15412.945 8613.565 ;
      RECT 15411.545 187.94 15411.825 8613.565 ;
      RECT 15410.425 187.94 15410.705 8613.565 ;
      RECT 15395.445 187.44 15407.765 8613.565 ;
      RECT 15390.265 187.94 15390.545 8613.565 ;
      RECT 15389.145 187.94 15389.425 8613.565 ;
      RECT 15388.025 187.94 15388.305 8613.565 ;
      RECT 15382.985 187.94 15383.265 8613.565 ;
      RECT 15343.365 187.94 15382.145 8613.565 ;
      RECT 15334.825 187.94 15335.105 8613.565 ;
      RECT 15333.705 187.94 15333.985 8613.565 ;
      RECT 15331.465 187.94 15331.745 8613.565 ;
      RECT 15330.345 187.94 15330.625 8613.565 ;
      RECT 15320.825 187.94 15329.365 8613.565 ;
      RECT 15320.965 187.44 15329.365 8613.565 ;
      RECT 15311.725 187.94 15313.825 8613.565 ;
      RECT 15310.465 187.94 15310.745 8613.565 ;
      RECT 15309.345 187.94 15309.625 8613.565 ;
      RECT 15282.325 187.44 15307.245 8613.565 ;
      RECT 15278.825 187.94 15279.105 8613.565 ;
      RECT 15277.705 187.94 15277.985 8613.565 ;
      RECT 15269.305 187.94 15269.585 8613.565 ;
      RECT 15255.305 187.94 15268.325 8613.565 ;
      RECT 15255.445 187.44 15268.325 8613.565 ;
      RECT 15253.065 187.94 15253.345 8613.565 ;
      RECT 15251.945 187.94 15252.225 8613.565 ;
      RECT 15250.825 187.94 15251.105 8613.565 ;
      RECT 15243.545 187.94 15243.825 8613.565 ;
      RECT 15203.365 187.94 15242.705 8613.565 ;
      RECT 15202.105 187.94 15202.385 8613.565 ;
      RECT 15197.065 187.94 15197.345 8613.565 ;
      RECT 15195.945 187.94 15196.225 8613.565 ;
      RECT 15181.525 187.44 15189.365 8613.565 ;
      RECT 15179.145 187.94 15179.425 8613.565 ;
      RECT 15178.025 187.94 15178.305 8613.565 ;
      RECT 15175.785 187.94 15176.065 8613.565 ;
      RECT 15174.665 187.94 15174.945 8613.565 ;
      RECT 15171.725 187.94 15173.825 8613.565 ;
      RECT 15142.325 187.44 15167.245 8613.565 ;
      RECT 15138.825 187.94 15139.105 8613.565 ;
      RECT 15137.705 187.94 15137.985 8613.565 ;
      RECT 15136.585 187.94 15136.865 8613.565 ;
      RECT 15131.545 187.94 15131.825 8613.565 ;
      RECT 15130.425 187.94 15130.705 8613.565 ;
      RECT 15116.005 187.44 15128.325 8613.565 ;
      RECT 15109.145 187.94 15109.425 8613.565 ;
      RECT 15108.025 187.94 15108.305 8613.565 ;
      RECT 15105.785 187.94 15106.065 8613.565 ;
      RECT 15104.665 187.94 15104.945 8613.565 ;
      RECT 15103.545 187.94 15103.825 8613.565 ;
      RECT 15062.805 187.44 15102.005 8613.565 ;
      RECT 15056.505 187.94 15056.785 8613.565 ;
      RECT 15055.385 187.94 15055.665 8613.565 ;
      RECT 15054.265 187.94 15054.545 8613.565 ;
      RECT 15040.825 187.94 15049.365 8613.565 ;
      RECT 15040.965 187.44 15049.365 8613.565 ;
      RECT 15039.705 187.94 15039.985 8613.565 ;
      RECT 15031.725 187.44 15033.125 8613.565 ;
      RECT 15029.345 187.94 15029.625 8613.565 ;
      RECT 15028.225 187.94 15028.505 8613.565 ;
      RECT 15001.205 187.44 15026.685 8613.565 ;
      RECT 14999.945 187.94 15000.225 8613.565 ;
      RECT 14998.825 187.94 14999.105 8613.565 ;
      RECT 14997.705 187.94 14997.985 8613.565 ;
      RECT 14990.425 187.94 14990.705 8613.565 ;
      RECT 14989.305 187.94 14989.585 8613.565 ;
      RECT 14974.745 187.94 14988.325 8613.565 ;
      RECT 14974.885 187.44 14988.325 8613.565 ;
      RECT 14969.705 187.94 14969.985 8613.565 ;
      RECT 14968.585 187.94 14968.865 8613.565 ;
      RECT 14923.925 187.44 14962.005 8613.565 ;
      RECT 14921.545 187.94 14921.825 8613.565 ;
      RECT 14920.425 187.94 14920.705 8613.565 ;
      RECT 14918.185 187.94 14918.465 8613.565 ;
      RECT 14917.065 187.94 14917.345 8613.565 ;
      RECT 14915.945 187.94 14916.225 8613.565 ;
      RECT 14901.525 187.44 14909.365 8613.565 ;
      RECT 14900.265 187.94 14900.545 8613.565 ;
      RECT 14899.145 187.94 14899.425 8613.565 ;
      RECT 14898.025 187.94 14898.305 8613.565 ;
      RECT 14891.025 187.94 14893.125 8613.565 ;
      RECT 14891.165 187.44 14893.125 8613.565 ;
      RECT 14889.905 187.94 14890.185 8613.565 ;
      RECT 14861.765 187.44 14886.685 8613.565 ;
      RECT 14856.025 187.94 14856.305 8613.565 ;
      RECT 14854.905 187.94 14855.185 8613.565 ;
      RECT 14852.665 187.94 14852.945 8613.565 ;
      RECT 14851.545 187.94 14851.825 8613.565 ;
      RECT 14850.425 187.94 14850.705 8613.565 ;
      RECT 14835.445 187.44 14847.765 8613.565 ;
      RECT 14830.265 187.94 14830.545 8613.565 ;
      RECT 14829.145 187.94 14829.425 8613.565 ;
      RECT 14828.025 187.94 14828.305 8613.565 ;
      RECT 14822.985 187.94 14823.265 8613.565 ;
      RECT 14783.365 187.94 14822.145 8613.565 ;
      RECT 14774.825 187.94 14775.105 8613.565 ;
      RECT 14773.705 187.94 14773.985 8613.565 ;
      RECT 14771.465 187.94 14771.745 8613.565 ;
      RECT 14770.345 187.94 14770.625 8613.565 ;
      RECT 14760.825 187.94 14769.365 8613.565 ;
      RECT 14760.965 187.44 14769.365 8613.565 ;
      RECT 14751.725 187.94 14753.825 8613.565 ;
      RECT 14750.465 187.94 14750.745 8613.565 ;
      RECT 14749.345 187.94 14749.625 8613.565 ;
      RECT 14722.325 187.44 14747.245 8613.565 ;
      RECT 14718.825 187.94 14719.105 8613.565 ;
      RECT 14717.705 187.94 14717.985 8613.565 ;
      RECT 14709.305 187.94 14709.585 8613.565 ;
      RECT 14695.305 187.94 14708.325 8613.565 ;
      RECT 14695.445 187.44 14708.325 8613.565 ;
      RECT 14693.065 187.94 14693.345 8613.565 ;
      RECT 14691.945 187.94 14692.225 8613.565 ;
      RECT 14690.825 187.94 14691.105 8613.565 ;
      RECT 14683.545 187.94 14683.825 8613.565 ;
      RECT 14643.365 187.94 14682.705 8613.565 ;
      RECT 14642.105 187.94 14642.385 8613.565 ;
      RECT 14637.065 187.94 14637.345 8613.565 ;
      RECT 14635.945 187.94 14636.225 8613.565 ;
      RECT 14621.525 187.44 14629.365 8613.565 ;
      RECT 14619.145 187.94 14619.425 8613.565 ;
      RECT 14618.025 187.94 14618.305 8613.565 ;
      RECT 14615.785 187.94 14616.065 8613.565 ;
      RECT 14614.665 187.94 14614.945 8613.565 ;
      RECT 14611.725 187.94 14613.825 8613.565 ;
      RECT 14582.325 187.44 14607.245 8613.565 ;
      RECT 14578.825 187.94 14579.105 8613.565 ;
      RECT 14577.705 187.94 14577.985 8613.565 ;
      RECT 14576.585 187.94 14576.865 8613.565 ;
      RECT 14571.545 187.94 14571.825 8613.565 ;
      RECT 14570.425 187.94 14570.705 8613.565 ;
      RECT 14556.005 187.44 14568.325 8613.565 ;
      RECT 14549.145 187.94 14549.425 8613.565 ;
      RECT 14548.025 187.94 14548.305 8613.565 ;
      RECT 14545.785 187.94 14546.065 8613.565 ;
      RECT 14544.665 187.94 14544.945 8613.565 ;
      RECT 14543.545 187.94 14543.825 8613.565 ;
      RECT 14502.805 187.44 14542.005 8613.565 ;
      RECT 14496.505 187.94 14496.785 8613.565 ;
      RECT 14495.385 187.94 14495.665 8613.565 ;
      RECT 14494.265 187.94 14494.545 8613.565 ;
      RECT 14480.825 187.94 14489.365 8613.565 ;
      RECT 14480.965 187.44 14489.365 8613.565 ;
      RECT 14479.705 187.94 14479.985 8613.565 ;
      RECT 14471.725 187.44 14473.125 8613.565 ;
      RECT 14469.345 187.94 14469.625 8613.565 ;
      RECT 14468.225 187.94 14468.505 8613.565 ;
      RECT 14441.205 187.44 14466.685 8613.565 ;
      RECT 14439.945 187.94 14440.225 8613.565 ;
      RECT 14438.825 187.94 14439.105 8613.565 ;
      RECT 14437.705 187.94 14437.985 8613.565 ;
      RECT 14430.425 187.94 14430.705 8613.565 ;
      RECT 14429.305 187.94 14429.585 8613.565 ;
      RECT 14414.745 187.94 14428.325 8613.565 ;
      RECT 14414.885 187.44 14428.325 8613.565 ;
      RECT 14409.705 187.94 14409.985 8613.565 ;
      RECT 14408.585 187.94 14408.865 8613.565 ;
      RECT 14363.925 187.44 14402.005 8613.565 ;
      RECT 14361.545 187.94 14361.825 8613.565 ;
      RECT 14360.425 187.94 14360.705 8613.565 ;
      RECT 14358.185 187.94 14358.465 8613.565 ;
      RECT 14357.065 187.94 14357.345 8613.565 ;
      RECT 14355.945 187.94 14356.225 8613.565 ;
      RECT 14341.525 187.44 14349.365 8613.565 ;
      RECT 14340.265 187.94 14340.545 8613.565 ;
      RECT 14339.145 187.94 14339.425 8613.565 ;
      RECT 14338.025 187.94 14338.305 8613.565 ;
      RECT 14331.025 187.94 14333.125 8613.565 ;
      RECT 14331.165 187.44 14333.125 8613.565 ;
      RECT 14329.905 187.94 14330.185 8613.565 ;
      RECT 14301.765 187.44 14326.685 8613.565 ;
      RECT 14296.025 187.94 14296.305 8613.565 ;
      RECT 14294.905 187.94 14295.185 8613.565 ;
      RECT 14292.665 187.94 14292.945 8613.565 ;
      RECT 14291.545 187.94 14291.825 8613.565 ;
      RECT 14290.425 187.94 14290.705 8613.565 ;
      RECT 14275.445 187.44 14287.765 8613.565 ;
      RECT 14270.265 187.94 14270.545 8613.565 ;
      RECT 14269.145 187.94 14269.425 8613.565 ;
      RECT 14268.025 187.94 14268.305 8613.565 ;
      RECT 14262.985 187.94 14263.265 8613.565 ;
      RECT 14223.365 187.94 14262.145 8613.565 ;
      RECT 14214.825 187.94 14215.105 8613.565 ;
      RECT 14213.705 187.94 14213.985 8613.565 ;
      RECT 14211.465 187.94 14211.745 8613.565 ;
      RECT 14210.345 187.94 14210.625 8613.565 ;
      RECT 14200.825 187.94 14209.365 8613.565 ;
      RECT 14200.965 187.44 14209.365 8613.565 ;
      RECT 14191.725 187.94 14193.825 8613.565 ;
      RECT 14190.465 187.94 14190.745 8613.565 ;
      RECT 14189.345 187.94 14189.625 8613.565 ;
      RECT 14162.325 187.44 14187.245 8613.565 ;
      RECT 14158.825 187.94 14159.105 8613.565 ;
      RECT 14157.705 187.94 14157.985 8613.565 ;
      RECT 14149.305 187.94 14149.585 8613.565 ;
      RECT 14135.305 187.94 14148.325 8613.565 ;
      RECT 14135.445 187.44 14148.325 8613.565 ;
      RECT 14133.065 187.94 14133.345 8613.565 ;
      RECT 14131.945 187.94 14132.225 8613.565 ;
      RECT 14130.825 187.94 14131.105 8613.565 ;
      RECT 14123.545 187.94 14123.825 8613.565 ;
      RECT 14083.365 187.94 14122.705 8613.565 ;
      RECT 14082.105 187.94 14082.385 8613.565 ;
      RECT 14077.065 187.94 14077.345 8613.565 ;
      RECT 14075.945 187.94 14076.225 8613.565 ;
      RECT 14061.525 187.44 14069.365 8613.565 ;
      RECT 14059.145 187.94 14059.425 8613.565 ;
      RECT 14058.025 187.94 14058.305 8613.565 ;
      RECT 14055.785 187.94 14056.065 8613.565 ;
      RECT 14054.665 187.94 14054.945 8613.565 ;
      RECT 14051.725 187.94 14053.825 8613.565 ;
      RECT 14022.325 187.44 14047.245 8613.565 ;
      RECT 14018.825 187.94 14019.105 8613.565 ;
      RECT 14017.705 187.94 14017.985 8613.565 ;
      RECT 14016.585 187.94 14016.865 8613.565 ;
      RECT 14011.545 187.94 14011.825 8613.565 ;
      RECT 14010.425 187.94 14010.705 8613.565 ;
      RECT 13996.005 187.44 14008.325 8613.565 ;
      RECT 13989.145 187.94 13989.425 8613.565 ;
      RECT 13988.025 187.94 13988.305 8613.565 ;
      RECT 13985.785 187.94 13986.065 8613.565 ;
      RECT 13984.665 187.94 13984.945 8613.565 ;
      RECT 13983.545 187.94 13983.825 8613.565 ;
      RECT 13942.805 187.44 13982.005 8613.565 ;
      RECT 13936.505 187.94 13936.785 8613.565 ;
      RECT 13935.385 187.94 13935.665 8613.565 ;
      RECT 13934.265 187.94 13934.545 8613.565 ;
      RECT 13920.825 187.94 13929.365 8613.565 ;
      RECT 13920.965 187.44 13929.365 8613.565 ;
      RECT 13919.705 187.94 13919.985 8613.565 ;
      RECT 13911.725 187.44 13913.125 8613.565 ;
      RECT 13909.345 187.94 13909.625 8613.565 ;
      RECT 13908.225 187.94 13908.505 8613.565 ;
      RECT 13881.205 187.44 13906.685 8613.565 ;
      RECT 13879.945 187.94 13880.225 8613.565 ;
      RECT 13878.825 187.94 13879.105 8613.565 ;
      RECT 13877.705 187.94 13877.985 8613.565 ;
      RECT 13870.425 187.94 13870.705 8613.565 ;
      RECT 13869.305 187.94 13869.585 8613.565 ;
      RECT 13854.745 187.94 13868.325 8613.565 ;
      RECT 13854.885 187.44 13868.325 8613.565 ;
      RECT 13849.705 187.94 13849.985 8613.565 ;
      RECT 13848.585 187.94 13848.865 8613.565 ;
      RECT 13803.925 187.44 13842.005 8613.565 ;
      RECT 13801.545 187.94 13801.825 8613.565 ;
      RECT 13800.425 187.94 13800.705 8613.565 ;
      RECT 13798.185 187.94 13798.465 8613.565 ;
      RECT 13797.065 187.94 13797.345 8613.565 ;
      RECT 13795.945 187.94 13796.225 8613.565 ;
      RECT 13781.525 187.44 13789.365 8613.565 ;
      RECT 13780.265 187.94 13780.545 8613.565 ;
      RECT 13779.145 187.94 13779.425 8613.565 ;
      RECT 13778.025 187.94 13778.305 8613.565 ;
      RECT 13771.025 187.94 13773.125 8613.565 ;
      RECT 13771.165 187.44 13773.125 8613.565 ;
      RECT 13769.905 187.94 13770.185 8613.565 ;
      RECT 13741.765 187.44 13766.685 8613.565 ;
      RECT 13736.025 187.94 13736.305 8613.565 ;
      RECT 13734.905 187.94 13735.185 8613.565 ;
      RECT 13732.665 187.94 13732.945 8613.565 ;
      RECT 13731.545 187.94 13731.825 8613.565 ;
      RECT 13730.425 187.94 13730.705 8613.565 ;
      RECT 13715.445 187.44 13727.765 8613.565 ;
      RECT 13710.265 187.94 13710.545 8613.565 ;
      RECT 13709.145 187.94 13709.425 8613.565 ;
      RECT 13708.025 187.94 13708.305 8613.565 ;
      RECT 13702.985 187.94 13703.265 8613.565 ;
      RECT 13663.365 187.94 13702.145 8613.565 ;
      RECT 13654.825 187.94 13655.105 8613.565 ;
      RECT 13653.705 187.94 13653.985 8613.565 ;
      RECT 13651.465 187.94 13651.745 8613.565 ;
      RECT 13650.345 187.94 13650.625 8613.565 ;
      RECT 13640.825 187.94 13649.365 8613.565 ;
      RECT 13640.965 187.44 13649.365 8613.565 ;
      RECT 13631.725 187.94 13633.825 8613.565 ;
      RECT 13630.465 187.94 13630.745 8613.565 ;
      RECT 13629.345 187.94 13629.625 8613.565 ;
      RECT 13602.325 187.44 13627.245 8613.565 ;
      RECT 13598.825 187.94 13599.105 8613.565 ;
      RECT 13597.705 187.94 13597.985 8613.565 ;
      RECT 13589.305 187.94 13589.585 8613.565 ;
      RECT 13575.305 187.94 13588.325 8613.565 ;
      RECT 13575.445 187.44 13588.325 8613.565 ;
      RECT 13573.065 187.94 13573.345 8613.565 ;
      RECT 13571.945 187.94 13572.225 8613.565 ;
      RECT 13570.825 187.94 13571.105 8613.565 ;
      RECT 13563.545 187.94 13563.825 8613.565 ;
      RECT 13523.365 187.94 13562.705 8613.565 ;
      RECT 13522.105 187.94 13522.385 8613.565 ;
      RECT 13517.065 187.94 13517.345 8613.565 ;
      RECT 13515.945 187.94 13516.225 8613.565 ;
      RECT 13501.525 187.44 13509.365 8613.565 ;
      RECT 13499.145 187.94 13499.425 8613.565 ;
      RECT 18143.365 187.44 18182.005 8613.565 ;
      RECT 18111.725 187.44 18113.685 8613.565 ;
      RECT 18003.365 187.44 18042.565 8613.565 ;
      RECT 17971.725 187.44 17973.685 8613.565 ;
      RECT 17583.365 187.44 17622.005 8613.565 ;
      RECT 17551.725 187.44 17553.685 8613.565 ;
      RECT 17443.365 187.44 17482.565 8613.565 ;
      RECT 17411.725 187.44 17413.685 8613.565 ;
      RECT 17023.365 187.44 17062.005 8613.565 ;
      RECT 16991.725 187.44 16993.685 8613.565 ;
      RECT 16883.365 187.44 16922.565 8613.565 ;
      RECT 16851.725 187.44 16853.685 8613.565 ;
      RECT 16463.365 187.44 16502.005 8613.565 ;
      RECT 16431.725 187.44 16433.685 8613.565 ;
      RECT 16323.365 187.44 16362.565 8613.565 ;
      RECT 16291.725 187.44 16293.685 8613.565 ;
      RECT 15903.365 187.44 15942.005 8613.565 ;
      RECT 15871.725 187.44 15873.685 8613.565 ;
      RECT 15763.365 187.44 15802.565 8613.565 ;
      RECT 15731.725 187.44 15733.685 8613.565 ;
      RECT 15343.365 187.44 15382.005 8613.565 ;
      RECT 15311.725 187.44 15313.685 8613.565 ;
      RECT 15203.365 187.44 15242.565 8613.565 ;
      RECT 15171.725 187.44 15173.685 8613.565 ;
      RECT 14783.365 187.44 14822.005 8613.565 ;
      RECT 14751.725 187.44 14753.685 8613.565 ;
      RECT 14643.365 187.44 14682.565 8613.565 ;
      RECT 14611.725 187.44 14613.685 8613.565 ;
      RECT 14223.365 187.44 14262.005 8613.565 ;
      RECT 14191.725 187.44 14193.685 8613.565 ;
      RECT 14083.365 187.44 14122.565 8613.565 ;
      RECT 14051.725 187.44 14053.685 8613.565 ;
      RECT 13663.365 187.44 13702.005 8613.565 ;
      RECT 13631.725 187.44 13633.685 8613.565 ;
      RECT 13523.365 187.44 13562.565 8613.565 ;
      RECT 6982.145 188.86 13498.305 8613.565 ;
      RECT 13498.025 187.94 13498.305 8613.565 ;
      RECT 13495.785 187.94 13496.065 8613.565 ;
      RECT 13494.665 187.94 13494.945 8613.565 ;
      RECT 13491.725 187.94 13493.825 8613.565 ;
      RECT 13462.325 187.44 13487.245 8613.565 ;
      RECT 13458.825 187.94 13459.105 8613.565 ;
      RECT 13457.705 187.94 13457.985 8613.565 ;
      RECT 13456.585 187.94 13456.865 8613.565 ;
      RECT 13451.545 187.94 13451.825 8613.565 ;
      RECT 13450.425 187.94 13450.705 8613.565 ;
      RECT 13436.005 187.44 13448.325 8613.565 ;
      RECT 13429.145 187.94 13429.425 8613.565 ;
      RECT 13428.025 187.94 13428.305 8613.565 ;
      RECT 13425.785 187.94 13426.065 8613.565 ;
      RECT 13424.665 187.94 13424.945 8613.565 ;
      RECT 13423.545 187.94 13423.825 8613.565 ;
      RECT 13382.805 187.44 13422.005 8613.565 ;
      RECT 13376.505 187.94 13376.785 8613.565 ;
      RECT 13375.385 187.94 13375.665 8613.565 ;
      RECT 13374.265 187.94 13374.545 8613.565 ;
      RECT 13360.825 187.94 13369.365 8613.565 ;
      RECT 13360.965 187.44 13369.365 8613.565 ;
      RECT 13359.705 187.94 13359.985 8613.565 ;
      RECT 13351.725 187.44 13353.125 8613.565 ;
      RECT 13349.345 187.94 13349.625 8613.565 ;
      RECT 13348.225 187.94 13348.505 8613.565 ;
      RECT 13321.205 187.44 13346.685 8613.565 ;
      RECT 13319.945 187.94 13320.225 8613.565 ;
      RECT 13318.825 187.94 13319.105 8613.565 ;
      RECT 13317.705 187.94 13317.985 8613.565 ;
      RECT 13310.425 187.94 13310.705 8613.565 ;
      RECT 13309.305 187.94 13309.585 8613.565 ;
      RECT 13294.745 187.94 13308.325 8613.565 ;
      RECT 13294.885 187.44 13308.325 8613.565 ;
      RECT 13289.705 187.94 13289.985 8613.565 ;
      RECT 13288.585 187.94 13288.865 8613.565 ;
      RECT 13243.925 187.44 13282.005 8613.565 ;
      RECT 13241.545 187.94 13241.825 8613.565 ;
      RECT 13240.425 187.94 13240.705 8613.565 ;
      RECT 13238.185 187.94 13238.465 8613.565 ;
      RECT 13237.065 187.94 13237.345 8613.565 ;
      RECT 13235.945 187.94 13236.225 8613.565 ;
      RECT 13221.525 187.44 13229.365 8613.565 ;
      RECT 13220.265 187.94 13220.545 8613.565 ;
      RECT 13219.145 187.94 13219.425 8613.565 ;
      RECT 13218.025 187.94 13218.305 8613.565 ;
      RECT 13211.025 187.94 13213.125 8613.565 ;
      RECT 13211.165 187.44 13213.125 8613.565 ;
      RECT 13209.905 187.94 13210.185 8613.565 ;
      RECT 13181.765 187.44 13206.685 8613.565 ;
      RECT 13176.025 187.94 13176.305 8613.565 ;
      RECT 13174.905 187.94 13175.185 8613.565 ;
      RECT 13172.665 187.94 13172.945 8613.565 ;
      RECT 13171.545 187.94 13171.825 8613.565 ;
      RECT 13170.425 187.94 13170.705 8613.565 ;
      RECT 13155.445 187.44 13167.765 8613.565 ;
      RECT 13150.265 187.94 13150.545 8613.565 ;
      RECT 13149.145 187.94 13149.425 8613.565 ;
      RECT 13148.025 187.94 13148.305 8613.565 ;
      RECT 13142.985 187.94 13143.265 8613.565 ;
      RECT 13103.365 187.94 13142.145 8613.565 ;
      RECT 13094.825 187.94 13095.105 8613.565 ;
      RECT 13093.705 187.94 13093.985 8613.565 ;
      RECT 13091.465 187.94 13091.745 8613.565 ;
      RECT 13090.345 187.94 13090.625 8613.565 ;
      RECT 13080.825 187.94 13089.365 8613.565 ;
      RECT 13080.965 187.44 13089.365 8613.565 ;
      RECT 13071.725 187.94 13073.825 8613.565 ;
      RECT 13070.465 187.94 13070.745 8613.565 ;
      RECT 13069.345 187.94 13069.625 8613.565 ;
      RECT 13042.325 187.44 13067.245 8613.565 ;
      RECT 13038.825 187.94 13039.105 8613.565 ;
      RECT 13037.705 187.94 13037.985 8613.565 ;
      RECT 13029.305 187.94 13029.585 8613.565 ;
      RECT 13015.305 187.94 13028.325 8613.565 ;
      RECT 13015.445 187.44 13028.325 8613.565 ;
      RECT 13013.065 187.94 13013.345 8613.565 ;
      RECT 13011.945 187.94 13012.225 8613.565 ;
      RECT 13010.825 187.94 13011.105 8613.565 ;
      RECT 13003.545 187.94 13003.825 8613.565 ;
      RECT 12963.365 187.94 13002.705 8613.565 ;
      RECT 12962.105 187.94 12962.385 8613.565 ;
      RECT 12957.065 187.94 12957.345 8613.565 ;
      RECT 12955.945 187.94 12956.225 8613.565 ;
      RECT 12941.525 187.44 12949.365 8613.565 ;
      RECT 12939.145 187.94 12939.425 8613.565 ;
      RECT 12938.025 187.94 12938.305 8613.565 ;
      RECT 12935.785 187.94 12936.065 8613.565 ;
      RECT 12934.665 187.94 12934.945 8613.565 ;
      RECT 12931.725 187.94 12933.825 8613.565 ;
      RECT 12902.325 187.44 12927.245 8613.565 ;
      RECT 12898.825 187.94 12899.105 8613.565 ;
      RECT 12897.705 187.94 12897.985 8613.565 ;
      RECT 12896.585 187.94 12896.865 8613.565 ;
      RECT 12891.545 187.94 12891.825 8613.565 ;
      RECT 12890.425 187.94 12890.705 8613.565 ;
      RECT 12876.005 187.44 12888.325 8613.565 ;
      RECT 12869.145 187.94 12869.425 8613.565 ;
      RECT 12868.025 187.94 12868.305 8613.565 ;
      RECT 12865.785 187.94 12866.065 8613.565 ;
      RECT 12864.665 187.94 12864.945 8613.565 ;
      RECT 12863.545 187.94 12863.825 8613.565 ;
      RECT 12822.805 187.44 12862.005 8613.565 ;
      RECT 12816.505 187.94 12816.785 8613.565 ;
      RECT 12815.385 187.94 12815.665 8613.565 ;
      RECT 12814.265 187.94 12814.545 8613.565 ;
      RECT 12800.825 187.94 12809.365 8613.565 ;
      RECT 12800.965 187.44 12809.365 8613.565 ;
      RECT 12799.705 187.94 12799.985 8613.565 ;
      RECT 12791.725 187.44 12793.125 8613.565 ;
      RECT 12789.345 187.94 12789.625 8613.565 ;
      RECT 12788.225 187.94 12788.505 8613.565 ;
      RECT 12761.205 187.44 12786.685 8613.565 ;
      RECT 12759.945 187.94 12760.225 8613.565 ;
      RECT 12758.825 187.94 12759.105 8613.565 ;
      RECT 12757.705 187.94 12757.985 8613.565 ;
      RECT 12750.425 187.94 12750.705 8613.565 ;
      RECT 12749.305 187.94 12749.585 8613.565 ;
      RECT 12734.745 187.94 12748.325 8613.565 ;
      RECT 12734.885 187.44 12748.325 8613.565 ;
      RECT 12729.705 187.94 12729.985 8613.565 ;
      RECT 12728.585 187.94 12728.865 8613.565 ;
      RECT 12683.925 187.44 12722.005 8613.565 ;
      RECT 12681.545 187.94 12681.825 8613.565 ;
      RECT 12680.425 187.94 12680.705 8613.565 ;
      RECT 12678.185 187.94 12678.465 8613.565 ;
      RECT 12677.065 187.94 12677.345 8613.565 ;
      RECT 12675.945 187.94 12676.225 8613.565 ;
      RECT 12661.525 187.44 12669.365 8613.565 ;
      RECT 12660.265 187.94 12660.545 8613.565 ;
      RECT 12659.145 187.94 12659.425 8613.565 ;
      RECT 12658.025 187.94 12658.305 8613.565 ;
      RECT 12651.025 187.94 12653.125 8613.565 ;
      RECT 12651.165 187.44 12653.125 8613.565 ;
      RECT 12649.905 187.94 12650.185 8613.565 ;
      RECT 12621.765 187.44 12646.685 8613.565 ;
      RECT 12616.025 187.94 12616.305 8613.565 ;
      RECT 12614.905 187.94 12615.185 8613.565 ;
      RECT 12612.665 187.94 12612.945 8613.565 ;
      RECT 12611.545 187.94 12611.825 8613.565 ;
      RECT 12610.425 187.94 12610.705 8613.565 ;
      RECT 12595.445 187.44 12607.765 8613.565 ;
      RECT 12590.265 187.94 12590.545 8613.565 ;
      RECT 12589.145 187.94 12589.425 8613.565 ;
      RECT 12588.025 187.94 12588.305 8613.565 ;
      RECT 12582.985 187.94 12583.265 8613.565 ;
      RECT 12543.365 187.94 12582.145 8613.565 ;
      RECT 12534.825 187.94 12535.105 8613.565 ;
      RECT 12533.705 187.94 12533.985 8613.565 ;
      RECT 12531.465 187.94 12531.745 8613.565 ;
      RECT 12530.345 187.94 12530.625 8613.565 ;
      RECT 12520.825 187.94 12529.365 8613.565 ;
      RECT 12520.965 187.44 12529.365 8613.565 ;
      RECT 12511.725 187.94 12513.825 8613.565 ;
      RECT 12510.465 187.94 12510.745 8613.565 ;
      RECT 12509.345 187.94 12509.625 8613.565 ;
      RECT 12482.325 187.44 12507.245 8613.565 ;
      RECT 12478.825 187.94 12479.105 8613.565 ;
      RECT 12477.705 187.94 12477.985 8613.565 ;
      RECT 12469.305 187.94 12469.585 8613.565 ;
      RECT 12455.305 187.94 12468.325 8613.565 ;
      RECT 12455.445 187.44 12468.325 8613.565 ;
      RECT 12453.065 187.94 12453.345 8613.565 ;
      RECT 12451.945 187.94 12452.225 8613.565 ;
      RECT 12450.825 187.94 12451.105 8613.565 ;
      RECT 12443.545 187.94 12443.825 8613.565 ;
      RECT 12403.365 187.94 12442.705 8613.565 ;
      RECT 12402.105 187.94 12402.385 8613.565 ;
      RECT 12397.065 187.94 12397.345 8613.565 ;
      RECT 12395.945 187.94 12396.225 8613.565 ;
      RECT 12381.525 187.44 12389.365 8613.565 ;
      RECT 12379.145 187.94 12379.425 8613.565 ;
      RECT 12378.025 187.94 12378.305 8613.565 ;
      RECT 12375.785 187.94 12376.065 8613.565 ;
      RECT 12374.665 187.94 12374.945 8613.565 ;
      RECT 12371.725 187.94 12373.825 8613.565 ;
      RECT 12342.325 187.44 12367.245 8613.565 ;
      RECT 12338.825 187.94 12339.105 8613.565 ;
      RECT 12337.705 187.94 12337.985 8613.565 ;
      RECT 12336.585 187.94 12336.865 8613.565 ;
      RECT 12331.545 187.94 12331.825 8613.565 ;
      RECT 12330.425 187.94 12330.705 8613.565 ;
      RECT 12316.005 187.44 12328.325 8613.565 ;
      RECT 12309.145 187.94 12309.425 8613.565 ;
      RECT 12308.025 187.94 12308.305 8613.565 ;
      RECT 12305.785 187.94 12306.065 8613.565 ;
      RECT 12304.665 187.94 12304.945 8613.565 ;
      RECT 12303.545 187.94 12303.825 8613.565 ;
      RECT 12262.805 187.44 12302.005 8613.565 ;
      RECT 12256.505 187.94 12256.785 8613.565 ;
      RECT 12255.385 187.94 12255.665 8613.565 ;
      RECT 12254.265 187.94 12254.545 8613.565 ;
      RECT 12240.825 187.94 12249.365 8613.565 ;
      RECT 12240.965 187.44 12249.365 8613.565 ;
      RECT 12239.705 187.94 12239.985 8613.565 ;
      RECT 12231.725 187.44 12233.125 8613.565 ;
      RECT 12229.345 187.94 12229.625 8613.565 ;
      RECT 12228.225 187.94 12228.505 8613.565 ;
      RECT 12201.205 187.44 12226.685 8613.565 ;
      RECT 12199.945 187.94 12200.225 8613.565 ;
      RECT 12198.825 187.94 12199.105 8613.565 ;
      RECT 12197.705 187.94 12197.985 8613.565 ;
      RECT 12190.425 187.94 12190.705 8613.565 ;
      RECT 12189.305 187.94 12189.585 8613.565 ;
      RECT 12174.745 187.94 12188.325 8613.565 ;
      RECT 12174.885 187.44 12188.325 8613.565 ;
      RECT 12169.705 187.94 12169.985 8613.565 ;
      RECT 12168.585 187.94 12168.865 8613.565 ;
      RECT 12123.925 187.44 12162.005 8613.565 ;
      RECT 12121.545 187.94 12121.825 8613.565 ;
      RECT 12120.425 187.94 12120.705 8613.565 ;
      RECT 12118.185 187.94 12118.465 8613.565 ;
      RECT 12117.065 187.94 12117.345 8613.565 ;
      RECT 12115.945 187.94 12116.225 8613.565 ;
      RECT 12101.525 187.44 12109.365 8613.565 ;
      RECT 12100.265 187.94 12100.545 8613.565 ;
      RECT 12099.145 187.94 12099.425 8613.565 ;
      RECT 12098.025 187.94 12098.305 8613.565 ;
      RECT 12091.025 187.94 12093.125 8613.565 ;
      RECT 12091.165 187.44 12093.125 8613.565 ;
      RECT 12089.905 187.94 12090.185 8613.565 ;
      RECT 12061.765 187.44 12086.685 8613.565 ;
      RECT 12056.025 187.94 12056.305 8613.565 ;
      RECT 12054.905 187.94 12055.185 8613.565 ;
      RECT 12052.665 187.94 12052.945 8613.565 ;
      RECT 12051.545 187.94 12051.825 8613.565 ;
      RECT 12050.425 187.94 12050.705 8613.565 ;
      RECT 12035.445 187.44 12047.765 8613.565 ;
      RECT 12030.265 187.94 12030.545 8613.565 ;
      RECT 12029.145 187.94 12029.425 8613.565 ;
      RECT 12028.025 187.94 12028.305 8613.565 ;
      RECT 12022.985 187.94 12023.265 8613.565 ;
      RECT 11983.365 187.94 12022.145 8613.565 ;
      RECT 11974.825 187.94 11975.105 8613.565 ;
      RECT 11973.705 187.94 11973.985 8613.565 ;
      RECT 11971.465 187.94 11971.745 8613.565 ;
      RECT 11970.345 187.94 11970.625 8613.565 ;
      RECT 11960.825 187.94 11969.365 8613.565 ;
      RECT 11960.965 187.44 11969.365 8613.565 ;
      RECT 11951.725 187.94 11953.825 8613.565 ;
      RECT 11950.465 187.94 11950.745 8613.565 ;
      RECT 11949.345 187.94 11949.625 8613.565 ;
      RECT 11922.325 187.44 11947.245 8613.565 ;
      RECT 11918.825 187.94 11919.105 8613.565 ;
      RECT 11917.705 187.94 11917.985 8613.565 ;
      RECT 11909.305 187.94 11909.585 8613.565 ;
      RECT 11895.305 187.94 11908.325 8613.565 ;
      RECT 11895.445 187.44 11908.325 8613.565 ;
      RECT 11893.065 187.94 11893.345 8613.565 ;
      RECT 11891.945 187.94 11892.225 8613.565 ;
      RECT 11890.825 187.94 11891.105 8613.565 ;
      RECT 11883.545 187.94 11883.825 8613.565 ;
      RECT 11843.365 187.94 11882.705 8613.565 ;
      RECT 11842.105 187.94 11842.385 8613.565 ;
      RECT 11837.065 187.94 11837.345 8613.565 ;
      RECT 11835.945 187.94 11836.225 8613.565 ;
      RECT 11821.525 187.44 11829.365 8613.565 ;
      RECT 11819.145 187.94 11819.425 8613.565 ;
      RECT 11818.025 187.94 11818.305 8613.565 ;
      RECT 11815.785 187.94 11816.065 8613.565 ;
      RECT 11814.665 187.94 11814.945 8613.565 ;
      RECT 11811.725 187.94 11813.825 8613.565 ;
      RECT 11782.325 187.44 11807.245 8613.565 ;
      RECT 11778.825 187.94 11779.105 8613.565 ;
      RECT 11777.705 187.94 11777.985 8613.565 ;
      RECT 11776.585 187.94 11776.865 8613.565 ;
      RECT 11771.545 187.94 11771.825 8613.565 ;
      RECT 11770.425 187.94 11770.705 8613.565 ;
      RECT 11756.005 187.44 11768.325 8613.565 ;
      RECT 11749.145 187.94 11749.425 8613.565 ;
      RECT 11748.025 187.94 11748.305 8613.565 ;
      RECT 11745.785 187.94 11746.065 8613.565 ;
      RECT 11744.665 187.94 11744.945 8613.565 ;
      RECT 11743.545 187.94 11743.825 8613.565 ;
      RECT 11702.805 187.44 11742.005 8613.565 ;
      RECT 11696.505 187.94 11696.785 8613.565 ;
      RECT 11695.385 187.94 11695.665 8613.565 ;
      RECT 11694.265 187.94 11694.545 8613.565 ;
      RECT 11680.825 187.94 11689.365 8613.565 ;
      RECT 11680.965 187.44 11689.365 8613.565 ;
      RECT 11679.705 187.94 11679.985 8613.565 ;
      RECT 11671.725 187.44 11673.125 8613.565 ;
      RECT 11669.345 187.94 11669.625 8613.565 ;
      RECT 11668.225 187.94 11668.505 8613.565 ;
      RECT 11641.205 187.44 11666.685 8613.565 ;
      RECT 11639.945 187.94 11640.225 8613.565 ;
      RECT 11638.825 187.94 11639.105 8613.565 ;
      RECT 11637.705 187.94 11637.985 8613.565 ;
      RECT 11630.425 187.94 11630.705 8613.565 ;
      RECT 11629.305 187.94 11629.585 8613.565 ;
      RECT 11614.745 187.94 11628.325 8613.565 ;
      RECT 11614.885 187.44 11628.325 8613.565 ;
      RECT 11609.705 187.94 11609.985 8613.565 ;
      RECT 11608.585 187.94 11608.865 8613.565 ;
      RECT 11563.925 187.44 11602.005 8613.565 ;
      RECT 11561.545 187.94 11561.825 8613.565 ;
      RECT 11560.425 187.94 11560.705 8613.565 ;
      RECT 11558.185 187.94 11558.465 8613.565 ;
      RECT 11557.065 187.94 11557.345 8613.565 ;
      RECT 11555.945 187.94 11556.225 8613.565 ;
      RECT 11541.525 187.44 11549.365 8613.565 ;
      RECT 11540.265 187.94 11540.545 8613.565 ;
      RECT 11539.145 187.94 11539.425 8613.565 ;
      RECT 11538.025 187.94 11538.305 8613.565 ;
      RECT 11531.025 187.94 11533.125 8613.565 ;
      RECT 11531.165 187.44 11533.125 8613.565 ;
      RECT 11529.905 187.94 11530.185 8613.565 ;
      RECT 11501.765 187.44 11526.685 8613.565 ;
      RECT 11496.025 187.94 11496.305 8613.565 ;
      RECT 11494.905 187.94 11495.185 8613.565 ;
      RECT 11492.665 187.94 11492.945 8613.565 ;
      RECT 11491.545 187.94 11491.825 8613.565 ;
      RECT 11490.425 187.94 11490.705 8613.565 ;
      RECT 11475.445 187.44 11487.765 8613.565 ;
      RECT 11470.265 187.94 11470.545 8613.565 ;
      RECT 11469.145 187.94 11469.425 8613.565 ;
      RECT 11468.025 187.94 11468.305 8613.565 ;
      RECT 11462.985 187.94 11463.265 8613.565 ;
      RECT 11423.365 187.94 11462.145 8613.565 ;
      RECT 11414.825 187.94 11415.105 8613.565 ;
      RECT 11413.705 187.94 11413.985 8613.565 ;
      RECT 11411.465 187.94 11411.745 8613.565 ;
      RECT 11410.345 187.94 11410.625 8613.565 ;
      RECT 11400.825 187.94 11409.365 8613.565 ;
      RECT 11400.965 187.44 11409.365 8613.565 ;
      RECT 11391.725 187.94 11393.825 8613.565 ;
      RECT 11390.465 187.94 11390.745 8613.565 ;
      RECT 11389.345 187.94 11389.625 8613.565 ;
      RECT 11362.325 187.44 11387.245 8613.565 ;
      RECT 11358.825 187.94 11359.105 8613.565 ;
      RECT 11357.705 187.94 11357.985 8613.565 ;
      RECT 11349.305 187.94 11349.585 8613.565 ;
      RECT 11335.305 187.94 11348.325 8613.565 ;
      RECT 11335.445 187.44 11348.325 8613.565 ;
      RECT 11333.065 187.94 11333.345 8613.565 ;
      RECT 11331.945 187.94 11332.225 8613.565 ;
      RECT 11330.825 187.94 11331.105 8613.565 ;
      RECT 11323.545 187.94 11323.825 8613.565 ;
      RECT 11283.365 187.94 11322.705 8613.565 ;
      RECT 11282.105 187.94 11282.385 8613.565 ;
      RECT 11277.065 187.94 11277.345 8613.565 ;
      RECT 11275.945 187.94 11276.225 8613.565 ;
      RECT 11261.525 187.44 11269.365 8613.565 ;
      RECT 11259.145 187.94 11259.425 8613.565 ;
      RECT 11258.025 187.94 11258.305 8613.565 ;
      RECT 11255.785 187.94 11256.065 8613.565 ;
      RECT 11254.665 187.94 11254.945 8613.565 ;
      RECT 11251.725 187.94 11253.825 8613.565 ;
      RECT 11222.325 187.44 11247.245 8613.565 ;
      RECT 11218.825 187.94 11219.105 8613.565 ;
      RECT 11217.705 187.94 11217.985 8613.565 ;
      RECT 11216.585 187.94 11216.865 8613.565 ;
      RECT 11211.545 187.94 11211.825 8613.565 ;
      RECT 11210.425 187.94 11210.705 8613.565 ;
      RECT 11196.005 187.44 11208.325 8613.565 ;
      RECT 11189.145 187.94 11189.425 8613.565 ;
      RECT 11188.025 187.94 11188.305 8613.565 ;
      RECT 11185.785 187.94 11186.065 8613.565 ;
      RECT 11184.665 187.94 11184.945 8613.565 ;
      RECT 11183.545 187.94 11183.825 8613.565 ;
      RECT 11142.805 187.44 11182.005 8613.565 ;
      RECT 11136.505 187.94 11136.785 8613.565 ;
      RECT 11135.385 187.94 11135.665 8613.565 ;
      RECT 11134.265 187.94 11134.545 8613.565 ;
      RECT 11120.825 187.94 11129.365 8613.565 ;
      RECT 11120.965 187.44 11129.365 8613.565 ;
      RECT 11119.705 187.94 11119.985 8613.565 ;
      RECT 11111.725 187.44 11113.125 8613.565 ;
      RECT 11109.345 187.94 11109.625 8613.565 ;
      RECT 11108.225 187.94 11108.505 8613.565 ;
      RECT 11081.205 187.44 11106.685 8613.565 ;
      RECT 11079.945 187.94 11080.225 8613.565 ;
      RECT 11078.825 187.94 11079.105 8613.565 ;
      RECT 11077.705 187.94 11077.985 8613.565 ;
      RECT 11070.425 187.94 11070.705 8613.565 ;
      RECT 11069.305 187.94 11069.585 8613.565 ;
      RECT 11054.745 187.94 11068.325 8613.565 ;
      RECT 11054.885 187.44 11068.325 8613.565 ;
      RECT 11049.705 187.94 11049.985 8613.565 ;
      RECT 11048.585 187.94 11048.865 8613.565 ;
      RECT 11003.925 187.44 11042.005 8613.565 ;
      RECT 11001.545 187.94 11001.825 8613.565 ;
      RECT 11000.425 187.94 11000.705 8613.565 ;
      RECT 10998.185 187.94 10998.465 8613.565 ;
      RECT 10997.065 187.94 10997.345 8613.565 ;
      RECT 10995.945 187.94 10996.225 8613.565 ;
      RECT 10981.525 187.44 10989.365 8613.565 ;
      RECT 10980.265 187.94 10980.545 8613.565 ;
      RECT 10979.145 187.94 10979.425 8613.565 ;
      RECT 10978.025 187.94 10978.305 8613.565 ;
      RECT 10971.025 187.94 10973.125 8613.565 ;
      RECT 10971.165 187.44 10973.125 8613.565 ;
      RECT 10969.905 187.94 10970.185 8613.565 ;
      RECT 10941.765 187.44 10966.685 8613.565 ;
      RECT 10936.025 187.94 10936.305 8613.565 ;
      RECT 10934.905 187.94 10935.185 8613.565 ;
      RECT 10932.665 187.94 10932.945 8613.565 ;
      RECT 10931.545 187.94 10931.825 8613.565 ;
      RECT 10930.425 187.94 10930.705 8613.565 ;
      RECT 10915.445 187.44 10927.765 8613.565 ;
      RECT 10910.265 187.94 10910.545 8613.565 ;
      RECT 10909.145 187.94 10909.425 8613.565 ;
      RECT 10908.025 187.94 10908.305 8613.565 ;
      RECT 10902.985 187.94 10903.265 8613.565 ;
      RECT 10863.365 187.94 10902.145 8613.565 ;
      RECT 10854.825 187.94 10855.105 8613.565 ;
      RECT 10853.705 187.94 10853.985 8613.565 ;
      RECT 10851.465 187.94 10851.745 8613.565 ;
      RECT 10850.345 187.94 10850.625 8613.565 ;
      RECT 10840.825 187.94 10849.365 8613.565 ;
      RECT 10840.965 187.44 10849.365 8613.565 ;
      RECT 10831.725 187.94 10833.825 8613.565 ;
      RECT 10830.465 187.94 10830.745 8613.565 ;
      RECT 10829.345 187.94 10829.625 8613.565 ;
      RECT 10802.325 187.44 10827.245 8613.565 ;
      RECT 10798.825 187.94 10799.105 8613.565 ;
      RECT 10797.705 187.94 10797.985 8613.565 ;
      RECT 10789.305 187.94 10789.585 8613.565 ;
      RECT 10775.305 187.94 10788.325 8613.565 ;
      RECT 10775.445 187.44 10788.325 8613.565 ;
      RECT 10773.065 187.94 10773.345 8613.565 ;
      RECT 10771.945 187.94 10772.225 8613.565 ;
      RECT 10770.825 187.94 10771.105 8613.565 ;
      RECT 10763.545 187.94 10763.825 8613.565 ;
      RECT 10723.365 187.94 10762.705 8613.565 ;
      RECT 10722.105 187.94 10722.385 8613.565 ;
      RECT 10717.065 187.94 10717.345 8613.565 ;
      RECT 10715.945 187.94 10716.225 8613.565 ;
      RECT 10701.525 187.44 10709.365 8613.565 ;
      RECT 10699.145 187.94 10699.425 8613.565 ;
      RECT 10698.025 187.94 10698.305 8613.565 ;
      RECT 10695.785 187.94 10696.065 8613.565 ;
      RECT 10694.665 187.94 10694.945 8613.565 ;
      RECT 10691.725 187.94 10693.825 8613.565 ;
      RECT 10662.325 187.44 10687.245 8613.565 ;
      RECT 10658.825 187.94 10659.105 8613.565 ;
      RECT 10657.705 187.94 10657.985 8613.565 ;
      RECT 10656.585 187.94 10656.865 8613.565 ;
      RECT 10651.545 187.94 10651.825 8613.565 ;
      RECT 10650.425 187.94 10650.705 8613.565 ;
      RECT 10636.005 187.44 10648.325 8613.565 ;
      RECT 10629.145 187.94 10629.425 8613.565 ;
      RECT 10628.025 187.94 10628.305 8613.565 ;
      RECT 10625.785 187.94 10626.065 8613.565 ;
      RECT 10624.665 187.94 10624.945 8613.565 ;
      RECT 10623.545 187.94 10623.825 8613.565 ;
      RECT 10582.805 187.44 10622.005 8613.565 ;
      RECT 10576.505 187.94 10576.785 8613.565 ;
      RECT 10575.385 187.94 10575.665 8613.565 ;
      RECT 10574.265 187.94 10574.545 8613.565 ;
      RECT 10560.825 187.94 10569.365 8613.565 ;
      RECT 10560.965 187.44 10569.365 8613.565 ;
      RECT 10559.705 187.94 10559.985 8613.565 ;
      RECT 10551.725 187.44 10553.125 8613.565 ;
      RECT 10549.345 187.94 10549.625 8613.565 ;
      RECT 10548.225 187.94 10548.505 8613.565 ;
      RECT 10521.205 187.44 10546.685 8613.565 ;
      RECT 10519.945 187.94 10520.225 8613.565 ;
      RECT 10518.825 187.94 10519.105 8613.565 ;
      RECT 10517.705 187.94 10517.985 8613.565 ;
      RECT 10510.425 187.94 10510.705 8613.565 ;
      RECT 10509.305 187.94 10509.585 8613.565 ;
      RECT 10494.745 187.94 10508.325 8613.565 ;
      RECT 10494.885 187.44 10508.325 8613.565 ;
      RECT 10489.705 187.94 10489.985 8613.565 ;
      RECT 10488.585 187.94 10488.865 8613.565 ;
      RECT 10443.925 187.44 10482.005 8613.565 ;
      RECT 10441.545 187.94 10441.825 8613.565 ;
      RECT 10440.425 187.94 10440.705 8613.565 ;
      RECT 10438.185 187.94 10438.465 8613.565 ;
      RECT 10437.065 187.94 10437.345 8613.565 ;
      RECT 10435.945 187.94 10436.225 8613.565 ;
      RECT 10421.525 187.44 10429.365 8613.565 ;
      RECT 10420.265 187.94 10420.545 8613.565 ;
      RECT 10419.145 187.94 10419.425 8613.565 ;
      RECT 10418.025 187.94 10418.305 8613.565 ;
      RECT 10411.025 187.94 10413.125 8613.565 ;
      RECT 10411.165 187.44 10413.125 8613.565 ;
      RECT 10409.905 187.94 10410.185 8613.565 ;
      RECT 10381.765 187.44 10406.685 8613.565 ;
      RECT 10376.025 187.94 10376.305 8613.565 ;
      RECT 10374.905 187.94 10375.185 8613.565 ;
      RECT 10372.665 187.94 10372.945 8613.565 ;
      RECT 10371.545 187.94 10371.825 8613.565 ;
      RECT 10370.425 187.94 10370.705 8613.565 ;
      RECT 10355.445 187.44 10367.765 8613.565 ;
      RECT 10350.265 187.94 10350.545 8613.565 ;
      RECT 10349.145 187.94 10349.425 8613.565 ;
      RECT 10348.025 187.94 10348.305 8613.565 ;
      RECT 10342.985 187.94 10343.265 8613.565 ;
      RECT 10303.365 187.94 10342.145 8613.565 ;
      RECT 10294.825 187.94 10295.105 8613.565 ;
      RECT 10293.705 187.94 10293.985 8613.565 ;
      RECT 10291.465 187.94 10291.745 8613.565 ;
      RECT 10290.345 187.94 10290.625 8613.565 ;
      RECT 10280.825 187.94 10289.365 8613.565 ;
      RECT 10280.965 187.44 10289.365 8613.565 ;
      RECT 10271.725 187.94 10273.825 8613.565 ;
      RECT 10270.465 187.94 10270.745 8613.565 ;
      RECT 10269.345 187.94 10269.625 8613.565 ;
      RECT 10242.325 187.44 10267.245 8613.565 ;
      RECT 10238.825 187.94 10239.105 8613.565 ;
      RECT 10237.705 187.94 10237.985 8613.565 ;
      RECT 10229.305 187.94 10229.585 8613.565 ;
      RECT 10215.305 187.94 10228.325 8613.565 ;
      RECT 10215.445 187.44 10228.325 8613.565 ;
      RECT 10213.065 187.94 10213.345 8613.565 ;
      RECT 10211.945 187.94 10212.225 8613.565 ;
      RECT 10210.825 187.94 10211.105 8613.565 ;
      RECT 10203.545 187.94 10203.825 8613.565 ;
      RECT 10163.365 187.94 10202.705 8613.565 ;
      RECT 10162.105 187.94 10162.385 8613.565 ;
      RECT 10157.065 187.94 10157.345 8613.565 ;
      RECT 10155.945 187.94 10156.225 8613.565 ;
      RECT 10141.525 187.44 10149.365 8613.565 ;
      RECT 10139.145 187.94 10139.425 8613.565 ;
      RECT 10138.025 187.94 10138.305 8613.565 ;
      RECT 10135.785 187.94 10136.065 8613.565 ;
      RECT 10134.665 187.94 10134.945 8613.565 ;
      RECT 10131.725 187.94 10133.825 8613.565 ;
      RECT 10102.325 187.44 10127.245 8613.565 ;
      RECT 10098.825 187.94 10099.105 8613.565 ;
      RECT 10097.705 187.94 10097.985 8613.565 ;
      RECT 10096.585 187.94 10096.865 8613.565 ;
      RECT 10091.545 187.94 10091.825 8613.565 ;
      RECT 10090.425 187.94 10090.705 8613.565 ;
      RECT 10076.005 187.44 10088.325 8613.565 ;
      RECT 10069.145 187.94 10069.425 8613.565 ;
      RECT 10068.025 187.94 10068.305 8613.565 ;
      RECT 10065.785 187.94 10066.065 8613.565 ;
      RECT 10064.665 187.94 10064.945 8613.565 ;
      RECT 10063.545 187.94 10063.825 8613.565 ;
      RECT 10022.805 187.44 10062.005 8613.565 ;
      RECT 10016.505 187.94 10016.785 8613.565 ;
      RECT 10015.385 187.94 10015.665 8613.565 ;
      RECT 10014.265 187.94 10014.545 8613.565 ;
      RECT 10000.825 187.94 10009.365 8613.565 ;
      RECT 10000.965 187.44 10009.365 8613.565 ;
      RECT 9999.705 187.94 9999.985 8613.565 ;
      RECT 9991.725 187.44 9993.125 8613.565 ;
      RECT 9989.345 187.94 9989.625 8613.565 ;
      RECT 9988.225 187.94 9988.505 8613.565 ;
      RECT 9961.205 187.44 9986.685 8613.565 ;
      RECT 9959.945 187.94 9960.225 8613.565 ;
      RECT 9958.825 187.94 9959.105 8613.565 ;
      RECT 9957.705 187.94 9957.985 8613.565 ;
      RECT 9950.425 187.94 9950.705 8613.565 ;
      RECT 9949.305 187.94 9949.585 8613.565 ;
      RECT 9934.745 187.94 9948.325 8613.565 ;
      RECT 9934.885 187.44 9948.325 8613.565 ;
      RECT 9929.705 187.94 9929.985 8613.565 ;
      RECT 9928.585 187.94 9928.865 8613.565 ;
      RECT 9883.925 187.44 9922.005 8613.565 ;
      RECT 9881.545 187.94 9881.825 8613.565 ;
      RECT 9880.425 187.94 9880.705 8613.565 ;
      RECT 9878.185 187.94 9878.465 8613.565 ;
      RECT 9877.065 187.94 9877.345 8613.565 ;
      RECT 9875.945 187.94 9876.225 8613.565 ;
      RECT 9861.525 187.44 9869.365 8613.565 ;
      RECT 9860.265 187.94 9860.545 8613.565 ;
      RECT 9859.145 187.94 9859.425 8613.565 ;
      RECT 9858.025 187.94 9858.305 8613.565 ;
      RECT 9851.025 187.94 9853.125 8613.565 ;
      RECT 9851.165 187.44 9853.125 8613.565 ;
      RECT 9849.905 187.94 9850.185 8613.565 ;
      RECT 9821.765 187.44 9846.685 8613.565 ;
      RECT 9816.025 187.94 9816.305 8613.565 ;
      RECT 9814.905 187.94 9815.185 8613.565 ;
      RECT 9812.665 187.94 9812.945 8613.565 ;
      RECT 9811.545 187.94 9811.825 8613.565 ;
      RECT 9810.425 187.94 9810.705 8613.565 ;
      RECT 9795.445 187.44 9807.765 8613.565 ;
      RECT 9790.265 187.94 9790.545 8613.565 ;
      RECT 9789.145 187.94 9789.425 8613.565 ;
      RECT 9788.025 187.94 9788.305 8613.565 ;
      RECT 9782.985 187.94 9783.265 8613.565 ;
      RECT 9743.365 187.94 9782.145 8613.565 ;
      RECT 9734.825 187.94 9735.105 8613.565 ;
      RECT 9733.705 187.94 9733.985 8613.565 ;
      RECT 9731.465 187.94 9731.745 8613.565 ;
      RECT 9730.345 187.94 9730.625 8613.565 ;
      RECT 9720.825 187.94 9729.365 8613.565 ;
      RECT 9720.965 187.44 9729.365 8613.565 ;
      RECT 9711.725 187.94 9713.825 8613.565 ;
      RECT 9710.465 187.94 9710.745 8613.565 ;
      RECT 9709.345 187.94 9709.625 8613.565 ;
      RECT 9682.325 187.44 9707.245 8613.565 ;
      RECT 9678.825 187.94 9679.105 8613.565 ;
      RECT 9677.705 187.94 9677.985 8613.565 ;
      RECT 9669.305 187.94 9669.585 8613.565 ;
      RECT 9655.305 187.94 9668.325 8613.565 ;
      RECT 9655.445 187.44 9668.325 8613.565 ;
      RECT 9653.065 187.94 9653.345 8613.565 ;
      RECT 9651.945 187.94 9652.225 8613.565 ;
      RECT 9650.825 187.94 9651.105 8613.565 ;
      RECT 9643.545 187.94 9643.825 8613.565 ;
      RECT 9603.365 187.94 9642.705 8613.565 ;
      RECT 9602.105 187.94 9602.385 8613.565 ;
      RECT 9597.065 187.94 9597.345 8613.565 ;
      RECT 9595.945 187.94 9596.225 8613.565 ;
      RECT 9581.525 187.44 9589.365 8613.565 ;
      RECT 9579.145 187.94 9579.425 8613.565 ;
      RECT 9578.025 187.94 9578.305 8613.565 ;
      RECT 9575.785 187.94 9576.065 8613.565 ;
      RECT 9574.665 187.94 9574.945 8613.565 ;
      RECT 9571.725 187.94 9573.825 8613.565 ;
      RECT 9542.325 187.44 9567.245 8613.565 ;
      RECT 9538.825 187.94 9539.105 8613.565 ;
      RECT 9537.705 187.94 9537.985 8613.565 ;
      RECT 9536.585 187.94 9536.865 8613.565 ;
      RECT 9531.545 187.94 9531.825 8613.565 ;
      RECT 9530.425 187.94 9530.705 8613.565 ;
      RECT 9516.005 187.44 9528.325 8613.565 ;
      RECT 9509.145 187.94 9509.425 8613.565 ;
      RECT 9508.025 187.94 9508.305 8613.565 ;
      RECT 9505.785 187.94 9506.065 8613.565 ;
      RECT 9504.665 187.94 9504.945 8613.565 ;
      RECT 9503.545 187.94 9503.825 8613.565 ;
      RECT 9462.805 187.44 9502.005 8613.565 ;
      RECT 9456.505 187.94 9456.785 8613.565 ;
      RECT 9455.385 187.94 9455.665 8613.565 ;
      RECT 9454.265 187.94 9454.545 8613.565 ;
      RECT 9440.825 187.94 9449.365 8613.565 ;
      RECT 9440.965 187.44 9449.365 8613.565 ;
      RECT 9439.705 187.94 9439.985 8613.565 ;
      RECT 9431.725 187.44 9433.125 8613.565 ;
      RECT 9429.345 187.94 9429.625 8613.565 ;
      RECT 9428.225 187.94 9428.505 8613.565 ;
      RECT 9401.205 187.44 9426.685 8613.565 ;
      RECT 9399.945 187.94 9400.225 8613.565 ;
      RECT 9398.825 187.94 9399.105 8613.565 ;
      RECT 9397.705 187.94 9397.985 8613.565 ;
      RECT 9390.425 187.94 9390.705 8613.565 ;
      RECT 9389.305 187.94 9389.585 8613.565 ;
      RECT 9374.745 187.94 9388.325 8613.565 ;
      RECT 9374.885 187.44 9388.325 8613.565 ;
      RECT 9369.705 187.94 9369.985 8613.565 ;
      RECT 9368.585 187.94 9368.865 8613.565 ;
      RECT 9323.925 187.44 9362.005 8613.565 ;
      RECT 9321.545 187.94 9321.825 8613.565 ;
      RECT 9320.425 187.94 9320.705 8613.565 ;
      RECT 9318.185 187.94 9318.465 8613.565 ;
      RECT 9317.065 187.94 9317.345 8613.565 ;
      RECT 9315.945 187.94 9316.225 8613.565 ;
      RECT 9301.525 187.44 9309.365 8613.565 ;
      RECT 9300.265 187.94 9300.545 8613.565 ;
      RECT 9299.145 187.94 9299.425 8613.565 ;
      RECT 9298.025 187.94 9298.305 8613.565 ;
      RECT 9291.025 187.94 9293.125 8613.565 ;
      RECT 9291.165 187.44 9293.125 8613.565 ;
      RECT 9289.905 187.94 9290.185 8613.565 ;
      RECT 9261.765 187.44 9286.685 8613.565 ;
      RECT 9256.025 187.94 9256.305 8613.565 ;
      RECT 9254.905 187.94 9255.185 8613.565 ;
      RECT 9252.665 187.94 9252.945 8613.565 ;
      RECT 9251.545 187.94 9251.825 8613.565 ;
      RECT 9250.425 187.94 9250.705 8613.565 ;
      RECT 9235.445 187.44 9247.765 8613.565 ;
      RECT 9230.265 187.94 9230.545 8613.565 ;
      RECT 9229.145 187.94 9229.425 8613.565 ;
      RECT 9228.025 187.94 9228.305 8613.565 ;
      RECT 9222.985 187.94 9223.265 8613.565 ;
      RECT 9183.365 187.94 9222.145 8613.565 ;
      RECT 9174.825 187.94 9175.105 8613.565 ;
      RECT 9173.705 187.94 9173.985 8613.565 ;
      RECT 9171.465 187.94 9171.745 8613.565 ;
      RECT 9170.345 187.94 9170.625 8613.565 ;
      RECT 9160.825 187.94 9169.365 8613.565 ;
      RECT 9160.965 187.44 9169.365 8613.565 ;
      RECT 9151.725 187.94 9153.825 8613.565 ;
      RECT 9150.465 187.94 9150.745 8613.565 ;
      RECT 9149.345 187.94 9149.625 8613.565 ;
      RECT 9122.325 187.44 9147.245 8613.565 ;
      RECT 9118.825 187.94 9119.105 8613.565 ;
      RECT 9117.705 187.94 9117.985 8613.565 ;
      RECT 9109.305 187.94 9109.585 8613.565 ;
      RECT 9095.305 187.94 9108.325 8613.565 ;
      RECT 9095.445 187.44 9108.325 8613.565 ;
      RECT 9093.065 187.94 9093.345 8613.565 ;
      RECT 9091.945 187.94 9092.225 8613.565 ;
      RECT 9090.825 187.94 9091.105 8613.565 ;
      RECT 9083.545 187.94 9083.825 8613.565 ;
      RECT 9043.365 187.94 9082.705 8613.565 ;
      RECT 9042.105 187.94 9042.385 8613.565 ;
      RECT 9037.065 187.94 9037.345 8613.565 ;
      RECT 9035.945 187.94 9036.225 8613.565 ;
      RECT 9021.525 187.44 9029.365 8613.565 ;
      RECT 9019.145 187.94 9019.425 8613.565 ;
      RECT 9018.025 187.94 9018.305 8613.565 ;
      RECT 9015.785 187.94 9016.065 8613.565 ;
      RECT 9014.665 187.94 9014.945 8613.565 ;
      RECT 9011.725 187.94 9013.825 8613.565 ;
      RECT 8982.325 187.44 9007.245 8613.565 ;
      RECT 8978.825 187.94 8979.105 8613.565 ;
      RECT 8977.705 187.94 8977.985 8613.565 ;
      RECT 8976.585 187.94 8976.865 8613.565 ;
      RECT 8971.545 187.94 8971.825 8613.565 ;
      RECT 8970.425 187.94 8970.705 8613.565 ;
      RECT 8956.005 187.44 8968.325 8613.565 ;
      RECT 8949.145 187.94 8949.425 8613.565 ;
      RECT 8948.025 187.94 8948.305 8613.565 ;
      RECT 8945.785 187.94 8946.065 8613.565 ;
      RECT 8944.665 187.94 8944.945 8613.565 ;
      RECT 8943.545 187.94 8943.825 8613.565 ;
      RECT 8902.805 187.44 8942.005 8613.565 ;
      RECT 8896.505 187.94 8896.785 8613.565 ;
      RECT 8895.385 187.94 8895.665 8613.565 ;
      RECT 8894.265 187.94 8894.545 8613.565 ;
      RECT 8880.825 187.94 8889.365 8613.565 ;
      RECT 8880.965 187.44 8889.365 8613.565 ;
      RECT 8879.705 187.94 8879.985 8613.565 ;
      RECT 8871.725 187.44 8873.125 8613.565 ;
      RECT 8869.345 187.94 8869.625 8613.565 ;
      RECT 8868.225 187.94 8868.505 8613.565 ;
      RECT 8841.205 187.44 8866.685 8613.565 ;
      RECT 8839.945 187.94 8840.225 8613.565 ;
      RECT 8838.825 187.94 8839.105 8613.565 ;
      RECT 8837.705 187.94 8837.985 8613.565 ;
      RECT 8830.425 187.94 8830.705 8613.565 ;
      RECT 8829.305 187.94 8829.585 8613.565 ;
      RECT 8814.745 187.94 8828.325 8613.565 ;
      RECT 8814.885 187.44 8828.325 8613.565 ;
      RECT 8809.705 187.94 8809.985 8613.565 ;
      RECT 8808.585 187.94 8808.865 8613.565 ;
      RECT 8763.925 187.44 8802.005 8613.565 ;
      RECT 8761.545 187.94 8761.825 8613.565 ;
      RECT 8760.425 187.94 8760.705 8613.565 ;
      RECT 8758.185 187.94 8758.465 8613.565 ;
      RECT 8757.065 187.94 8757.345 8613.565 ;
      RECT 8755.945 187.94 8756.225 8613.565 ;
      RECT 8741.525 187.44 8749.365 8613.565 ;
      RECT 8740.265 187.94 8740.545 8613.565 ;
      RECT 8739.145 187.94 8739.425 8613.565 ;
      RECT 8738.025 187.94 8738.305 8613.565 ;
      RECT 8731.025 187.94 8733.125 8613.565 ;
      RECT 8731.165 187.44 8733.125 8613.565 ;
      RECT 8729.905 187.94 8730.185 8613.565 ;
      RECT 8701.765 187.44 8726.685 8613.565 ;
      RECT 8696.025 187.94 8696.305 8613.565 ;
      RECT 8694.905 187.94 8695.185 8613.565 ;
      RECT 8692.665 187.94 8692.945 8613.565 ;
      RECT 8691.545 187.94 8691.825 8613.565 ;
      RECT 8690.425 187.94 8690.705 8613.565 ;
      RECT 8675.445 187.44 8687.765 8613.565 ;
      RECT 8670.265 187.94 8670.545 8613.565 ;
      RECT 8669.145 187.94 8669.425 8613.565 ;
      RECT 8668.025 187.94 8668.305 8613.565 ;
      RECT 8662.985 187.94 8663.265 8613.565 ;
      RECT 8623.365 187.94 8662.145 8613.565 ;
      RECT 8614.825 187.94 8615.105 8613.565 ;
      RECT 8613.705 187.94 8613.985 8613.565 ;
      RECT 8611.465 187.94 8611.745 8613.565 ;
      RECT 8610.345 187.94 8610.625 8613.565 ;
      RECT 8600.825 187.94 8609.365 8613.565 ;
      RECT 8600.965 187.44 8609.365 8613.565 ;
      RECT 8591.725 187.94 8593.825 8613.565 ;
      RECT 8590.465 187.94 8590.745 8613.565 ;
      RECT 8589.345 187.94 8589.625 8613.565 ;
      RECT 8562.325 187.44 8587.245 8613.565 ;
      RECT 8558.825 187.94 8559.105 8613.565 ;
      RECT 8557.705 187.94 8557.985 8613.565 ;
      RECT 8549.305 187.94 8549.585 8613.565 ;
      RECT 8535.305 187.94 8548.325 8613.565 ;
      RECT 8535.445 187.44 8548.325 8613.565 ;
      RECT 8533.065 187.94 8533.345 8613.565 ;
      RECT 8531.945 187.94 8532.225 8613.565 ;
      RECT 8530.825 187.94 8531.105 8613.565 ;
      RECT 8523.545 187.94 8523.825 8613.565 ;
      RECT 8483.365 187.94 8522.705 8613.565 ;
      RECT 8482.105 187.94 8482.385 8613.565 ;
      RECT 8477.065 187.94 8477.345 8613.565 ;
      RECT 8475.945 187.94 8476.225 8613.565 ;
      RECT 8461.525 187.44 8469.365 8613.565 ;
      RECT 8459.145 187.94 8459.425 8613.565 ;
      RECT 8458.025 187.94 8458.305 8613.565 ;
      RECT 8455.785 187.94 8456.065 8613.565 ;
      RECT 8454.665 187.94 8454.945 8613.565 ;
      RECT 8451.725 187.94 8453.825 8613.565 ;
      RECT 8422.325 187.44 8447.245 8613.565 ;
      RECT 8418.825 187.94 8419.105 8613.565 ;
      RECT 8417.705 187.94 8417.985 8613.565 ;
      RECT 8416.585 187.94 8416.865 8613.565 ;
      RECT 8411.545 187.94 8411.825 8613.565 ;
      RECT 8410.425 187.94 8410.705 8613.565 ;
      RECT 8396.005 187.44 8408.325 8613.565 ;
      RECT 8389.145 187.94 8389.425 8613.565 ;
      RECT 8388.025 187.94 8388.305 8613.565 ;
      RECT 8385.785 187.94 8386.065 8613.565 ;
      RECT 8384.665 187.94 8384.945 8613.565 ;
      RECT 8383.545 187.94 8383.825 8613.565 ;
      RECT 8342.805 187.44 8382.005 8613.565 ;
      RECT 8336.505 187.94 8336.785 8613.565 ;
      RECT 8335.385 187.94 8335.665 8613.565 ;
      RECT 8334.265 187.94 8334.545 8613.565 ;
      RECT 8320.825 187.94 8329.365 8613.565 ;
      RECT 8320.965 187.44 8329.365 8613.565 ;
      RECT 8319.705 187.94 8319.985 8613.565 ;
      RECT 8311.725 187.44 8313.125 8613.565 ;
      RECT 8309.345 187.94 8309.625 8613.565 ;
      RECT 8308.225 187.94 8308.505 8613.565 ;
      RECT 8281.205 187.44 8306.685 8613.565 ;
      RECT 8279.945 187.94 8280.225 8613.565 ;
      RECT 8278.825 187.94 8279.105 8613.565 ;
      RECT 8277.705 187.94 8277.985 8613.565 ;
      RECT 8270.425 187.94 8270.705 8613.565 ;
      RECT 8269.305 187.94 8269.585 8613.565 ;
      RECT 8254.745 187.94 8268.325 8613.565 ;
      RECT 8254.885 187.44 8268.325 8613.565 ;
      RECT 8249.705 187.94 8249.985 8613.565 ;
      RECT 8248.585 187.94 8248.865 8613.565 ;
      RECT 8203.925 187.44 8242.005 8613.565 ;
      RECT 8201.545 187.94 8201.825 8613.565 ;
      RECT 8200.425 187.94 8200.705 8613.565 ;
      RECT 8198.185 187.94 8198.465 8613.565 ;
      RECT 8197.065 187.94 8197.345 8613.565 ;
      RECT 8195.945 187.94 8196.225 8613.565 ;
      RECT 8181.525 187.44 8189.365 8613.565 ;
      RECT 8180.265 187.94 8180.545 8613.565 ;
      RECT 8179.145 187.94 8179.425 8613.565 ;
      RECT 8178.025 187.94 8178.305 8613.565 ;
      RECT 8171.025 187.94 8173.125 8613.565 ;
      RECT 8171.165 187.44 8173.125 8613.565 ;
      RECT 8169.905 187.94 8170.185 8613.565 ;
      RECT 8141.765 187.44 8166.685 8613.565 ;
      RECT 8136.025 187.94 8136.305 8613.565 ;
      RECT 8134.905 187.94 8135.185 8613.565 ;
      RECT 8132.665 187.94 8132.945 8613.565 ;
      RECT 8131.545 187.94 8131.825 8613.565 ;
      RECT 8130.425 187.94 8130.705 8613.565 ;
      RECT 8115.445 187.44 8127.765 8613.565 ;
      RECT 8110.265 187.94 8110.545 8613.565 ;
      RECT 8109.145 187.94 8109.425 8613.565 ;
      RECT 8108.025 187.94 8108.305 8613.565 ;
      RECT 8102.985 187.94 8103.265 8613.565 ;
      RECT 8063.365 187.94 8102.145 8613.565 ;
      RECT 8054.825 187.94 8055.105 8613.565 ;
      RECT 8053.705 187.94 8053.985 8613.565 ;
      RECT 8051.465 187.94 8051.745 8613.565 ;
      RECT 8050.345 187.94 8050.625 8613.565 ;
      RECT 8040.825 187.94 8049.365 8613.565 ;
      RECT 8040.965 187.44 8049.365 8613.565 ;
      RECT 8031.725 187.94 8033.825 8613.565 ;
      RECT 8030.465 187.94 8030.745 8613.565 ;
      RECT 8029.345 187.94 8029.625 8613.565 ;
      RECT 8002.325 187.44 8027.245 8613.565 ;
      RECT 7998.825 187.94 7999.105 8613.565 ;
      RECT 7997.705 187.94 7997.985 8613.565 ;
      RECT 7989.305 187.94 7989.585 8613.565 ;
      RECT 7975.305 187.94 7988.325 8613.565 ;
      RECT 7975.445 187.44 7988.325 8613.565 ;
      RECT 7973.065 187.94 7973.345 8613.565 ;
      RECT 7971.945 187.94 7972.225 8613.565 ;
      RECT 7970.825 187.94 7971.105 8613.565 ;
      RECT 7963.545 187.94 7963.825 8613.565 ;
      RECT 7923.365 187.94 7962.705 8613.565 ;
      RECT 7922.105 187.94 7922.385 8613.565 ;
      RECT 7917.065 187.94 7917.345 8613.565 ;
      RECT 7915.945 187.94 7916.225 8613.565 ;
      RECT 7901.525 187.44 7909.365 8613.565 ;
      RECT 7899.145 187.94 7899.425 8613.565 ;
      RECT 7898.025 187.94 7898.305 8613.565 ;
      RECT 7895.785 187.94 7896.065 8613.565 ;
      RECT 7894.665 187.94 7894.945 8613.565 ;
      RECT 7891.725 187.94 7893.825 8613.565 ;
      RECT 7862.325 187.44 7887.245 8613.565 ;
      RECT 7858.825 187.94 7859.105 8613.565 ;
      RECT 7857.705 187.94 7857.985 8613.565 ;
      RECT 7856.585 187.94 7856.865 8613.565 ;
      RECT 7851.545 187.94 7851.825 8613.565 ;
      RECT 7850.425 187.94 7850.705 8613.565 ;
      RECT 7836.005 187.44 7848.325 8613.565 ;
      RECT 7829.145 187.94 7829.425 8613.565 ;
      RECT 7828.025 187.94 7828.305 8613.565 ;
      RECT 7825.785 187.94 7826.065 8613.565 ;
      RECT 7824.665 187.94 7824.945 8613.565 ;
      RECT 7823.545 187.94 7823.825 8613.565 ;
      RECT 7782.805 187.44 7822.005 8613.565 ;
      RECT 7776.505 187.94 7776.785 8613.565 ;
      RECT 7775.385 187.94 7775.665 8613.565 ;
      RECT 7774.265 187.94 7774.545 8613.565 ;
      RECT 7760.825 187.94 7769.365 8613.565 ;
      RECT 7760.965 187.44 7769.365 8613.565 ;
      RECT 7759.705 187.94 7759.985 8613.565 ;
      RECT 7751.725 187.44 7753.125 8613.565 ;
      RECT 7749.345 187.94 7749.625 8613.565 ;
      RECT 7748.225 187.94 7748.505 8613.565 ;
      RECT 7721.205 187.44 7746.685 8613.565 ;
      RECT 7719.945 187.94 7720.225 8613.565 ;
      RECT 7718.825 187.94 7719.105 8613.565 ;
      RECT 7717.705 187.94 7717.985 8613.565 ;
      RECT 7710.425 187.94 7710.705 8613.565 ;
      RECT 7709.305 187.94 7709.585 8613.565 ;
      RECT 7694.745 187.94 7708.325 8613.565 ;
      RECT 7694.885 187.44 7708.325 8613.565 ;
      RECT 7689.705 187.94 7689.985 8613.565 ;
      RECT 7688.585 187.94 7688.865 8613.565 ;
      RECT 7643.925 187.44 7682.005 8613.565 ;
      RECT 7641.545 187.94 7641.825 8613.565 ;
      RECT 7640.425 187.94 7640.705 8613.565 ;
      RECT 7638.185 187.94 7638.465 8613.565 ;
      RECT 7637.065 187.94 7637.345 8613.565 ;
      RECT 7635.945 187.94 7636.225 8613.565 ;
      RECT 7621.525 187.44 7629.365 8613.565 ;
      RECT 7620.265 187.94 7620.545 8613.565 ;
      RECT 7619.145 187.94 7619.425 8613.565 ;
      RECT 7618.025 187.94 7618.305 8613.565 ;
      RECT 7611.025 187.94 7613.125 8613.565 ;
      RECT 7611.165 187.44 7613.125 8613.565 ;
      RECT 7609.905 187.94 7610.185 8613.565 ;
      RECT 7581.765 187.44 7606.685 8613.565 ;
      RECT 7576.025 187.94 7576.305 8613.565 ;
      RECT 7574.905 187.94 7575.185 8613.565 ;
      RECT 7572.665 187.94 7572.945 8613.565 ;
      RECT 7571.545 187.94 7571.825 8613.565 ;
      RECT 7570.425 187.94 7570.705 8613.565 ;
      RECT 7555.445 187.44 7567.765 8613.565 ;
      RECT 7550.265 187.94 7550.545 8613.565 ;
      RECT 7549.145 187.94 7549.425 8613.565 ;
      RECT 7548.025 187.94 7548.305 8613.565 ;
      RECT 7542.985 187.94 7543.265 8613.565 ;
      RECT 7503.365 187.94 7542.145 8613.565 ;
      RECT 7494.825 187.94 7495.105 8613.565 ;
      RECT 7493.705 187.94 7493.985 8613.565 ;
      RECT 7491.465 187.94 7491.745 8613.565 ;
      RECT 7490.345 187.94 7490.625 8613.565 ;
      RECT 7480.825 187.94 7489.365 8613.565 ;
      RECT 7480.965 187.44 7489.365 8613.565 ;
      RECT 7471.725 187.94 7473.825 8613.565 ;
      RECT 7470.465 187.94 7470.745 8613.565 ;
      RECT 7469.345 187.94 7469.625 8613.565 ;
      RECT 7442.325 187.44 7467.245 8613.565 ;
      RECT 7438.825 187.94 7439.105 8613.565 ;
      RECT 7437.705 187.94 7437.985 8613.565 ;
      RECT 7429.305 187.94 7429.585 8613.565 ;
      RECT 7415.305 187.94 7428.325 8613.565 ;
      RECT 7415.445 187.44 7428.325 8613.565 ;
      RECT 7413.065 187.94 7413.345 8613.565 ;
      RECT 7411.945 187.94 7412.225 8613.565 ;
      RECT 7410.825 187.94 7411.105 8613.565 ;
      RECT 7403.545 187.94 7403.825 8613.565 ;
      RECT 7363.365 187.94 7402.705 8613.565 ;
      RECT 7362.105 187.94 7362.385 8613.565 ;
      RECT 7357.065 187.94 7357.345 8613.565 ;
      RECT 7355.945 187.94 7356.225 8613.565 ;
      RECT 7341.525 187.44 7349.365 8613.565 ;
      RECT 7339.145 187.94 7339.425 8613.565 ;
      RECT 7338.025 187.94 7338.305 8613.565 ;
      RECT 7335.785 187.94 7336.065 8613.565 ;
      RECT 7334.665 187.94 7334.945 8613.565 ;
      RECT 7331.725 187.94 7333.825 8613.565 ;
      RECT 7302.325 187.44 7327.245 8613.565 ;
      RECT 7298.825 187.94 7299.105 8613.565 ;
      RECT 7297.705 187.94 7297.985 8613.565 ;
      RECT 7296.585 187.94 7296.865 8613.565 ;
      RECT 7291.545 187.94 7291.825 8613.565 ;
      RECT 7290.425 187.94 7290.705 8613.565 ;
      RECT 7276.005 187.44 7288.325 8613.565 ;
      RECT 7269.145 187.94 7269.425 8613.565 ;
      RECT 7268.025 187.94 7268.305 8613.565 ;
      RECT 7265.785 187.94 7266.065 8613.565 ;
      RECT 7264.665 187.94 7264.945 8613.565 ;
      RECT 7263.545 187.94 7263.825 8613.565 ;
      RECT 7222.805 187.44 7262.005 8613.565 ;
      RECT 7216.505 187.94 7216.785 8613.565 ;
      RECT 7215.385 187.94 7215.665 8613.565 ;
      RECT 7214.265 187.94 7214.545 8613.565 ;
      RECT 7200.825 187.94 7209.365 8613.565 ;
      RECT 7200.965 187.44 7209.365 8613.565 ;
      RECT 7199.705 187.94 7199.985 8613.565 ;
      RECT 7191.725 187.44 7193.125 8613.565 ;
      RECT 7189.345 187.94 7189.625 8613.565 ;
      RECT 7188.225 187.94 7188.505 8613.565 ;
      RECT 7161.205 187.44 7186.685 8613.565 ;
      RECT 7159.945 187.94 7160.225 8613.565 ;
      RECT 7158.825 187.94 7159.105 8613.565 ;
      RECT 7157.705 187.94 7157.985 8613.565 ;
      RECT 7150.425 187.94 7150.705 8613.565 ;
      RECT 7149.305 187.94 7149.585 8613.565 ;
      RECT 7134.745 187.94 7148.325 8613.565 ;
      RECT 7134.885 187.44 7148.325 8613.565 ;
      RECT 7129.705 187.94 7129.985 8613.565 ;
      RECT 7128.585 187.94 7128.865 8613.565 ;
      RECT 7083.925 187.44 7122.005 8613.565 ;
      RECT 7081.545 187.94 7081.825 8613.565 ;
      RECT 7080.425 187.94 7080.705 8613.565 ;
      RECT 7078.185 187.94 7078.465 8613.565 ;
      RECT 7077.065 187.94 7077.345 8613.565 ;
      RECT 7075.945 187.94 7076.225 8613.565 ;
      RECT 7061.525 187.44 7069.365 8613.565 ;
      RECT 7060.265 187.94 7060.545 8613.565 ;
      RECT 7059.145 187.94 7059.425 8613.565 ;
      RECT 7058.025 187.94 7058.305 8613.565 ;
      RECT 7051.025 187.94 7053.125 8613.565 ;
      RECT 7051.165 187.44 7053.125 8613.565 ;
      RECT 7049.905 187.94 7050.185 8613.565 ;
      RECT 7021.765 187.44 7046.685 8613.565 ;
      RECT 7016.025 187.94 7016.305 8613.565 ;
      RECT 7014.905 187.94 7015.185 8613.565 ;
      RECT 7012.665 187.94 7012.945 8613.565 ;
      RECT 7011.545 187.94 7011.825 8613.565 ;
      RECT 7010.425 187.94 7010.705 8613.565 ;
      RECT 6995.445 187.44 7007.765 8613.565 ;
      RECT 6990.265 187.94 6990.545 8613.565 ;
      RECT 6989.145 187.94 6989.425 8613.565 ;
      RECT 6988.025 187.94 6988.305 8613.565 ;
      RECT 6982.985 187.94 6983.265 8613.565 ;
      RECT 13491.725 187.44 13493.685 8613.565 ;
      RECT 13103.365 187.44 13142.005 8613.565 ;
      RECT 13071.725 187.44 13073.685 8613.565 ;
      RECT 12963.365 187.44 13002.565 8613.565 ;
      RECT 12931.725 187.44 12933.685 8613.565 ;
      RECT 12543.365 187.44 12582.005 8613.565 ;
      RECT 12511.725 187.44 12513.685 8613.565 ;
      RECT 12403.365 187.44 12442.565 8613.565 ;
      RECT 12371.725 187.44 12373.685 8613.565 ;
      RECT 11983.365 187.44 12022.005 8613.565 ;
      RECT 11951.725 187.44 11953.685 8613.565 ;
      RECT 11843.365 187.44 11882.565 8613.565 ;
      RECT 11811.725 187.44 11813.685 8613.565 ;
      RECT 11423.365 187.44 11462.005 8613.565 ;
      RECT 11391.725 187.44 11393.685 8613.565 ;
      RECT 11283.365 187.44 11322.565 8613.565 ;
      RECT 11251.725 187.44 11253.685 8613.565 ;
      RECT 10863.365 187.44 10902.005 8613.565 ;
      RECT 10831.725 187.44 10833.685 8613.565 ;
      RECT 10723.365 187.44 10762.565 8613.565 ;
      RECT 10691.725 187.44 10693.685 8613.565 ;
      RECT 10303.365 187.44 10342.005 8613.565 ;
      RECT 10271.725 187.44 10273.685 8613.565 ;
      RECT 10163.365 187.44 10202.565 8613.565 ;
      RECT 10131.725 187.44 10133.685 8613.565 ;
      RECT 9743.365 187.44 9782.005 8613.565 ;
      RECT 9711.725 187.44 9713.685 8613.565 ;
      RECT 9603.365 187.44 9642.565 8613.565 ;
      RECT 9571.725 187.44 9573.685 8613.565 ;
      RECT 9183.365 187.44 9222.005 8613.565 ;
      RECT 9151.725 187.44 9153.685 8613.565 ;
      RECT 9043.365 187.44 9082.565 8613.565 ;
      RECT 9011.725 187.44 9013.685 8613.565 ;
      RECT 8623.365 187.44 8662.005 8613.565 ;
      RECT 8591.725 187.44 8593.685 8613.565 ;
      RECT 8483.365 187.44 8522.565 8613.565 ;
      RECT 8451.725 187.44 8453.685 8613.565 ;
      RECT 8063.365 187.44 8102.005 8613.565 ;
      RECT 8031.725 187.44 8033.685 8613.565 ;
      RECT 7923.365 187.44 7962.565 8613.565 ;
      RECT 7891.725 187.44 7893.685 8613.565 ;
      RECT 7503.365 187.44 7542.005 8613.565 ;
      RECT 7471.725 187.44 7473.685 8613.565 ;
      RECT 7363.365 187.44 7402.565 8613.565 ;
      RECT 7331.725 187.44 7333.685 8613.565 ;
      RECT 326.66 8583.935 6982.145 8613.565 ;
      RECT 6943.365 187.94 6982.145 8613.565 ;
      RECT 328.08 188.86 6982.145 8613.565 ;
      RECT 326.66 8545.42 6982.145 8581.675 ;
      RECT 326.66 8511.935 6982.145 8543.16 ;
      RECT 326.66 8473.42 6982.145 8509.675 ;
      RECT 326.66 8439.935 6982.145 8471.16 ;
      RECT 326.66 8401.42 6982.145 8437.675 ;
      RECT 326.66 187.44 466.125 8399.16 ;
      RECT 6934.825 187.94 6935.105 8613.565 ;
      RECT 6933.705 187.94 6933.985 8613.565 ;
      RECT 6931.465 187.94 6931.745 8613.565 ;
      RECT 6930.345 187.94 6930.625 8613.565 ;
      RECT 6920.825 187.94 6929.365 8613.565 ;
      RECT 6920.965 187.44 6929.365 8613.565 ;
      RECT 6911.725 187.94 6913.825 8613.565 ;
      RECT 6910.465 187.94 6910.745 8613.565 ;
      RECT 6909.345 187.94 6909.625 8613.565 ;
      RECT 6882.325 187.44 6907.245 8613.565 ;
      RECT 6878.825 187.94 6879.105 8613.565 ;
      RECT 6877.705 187.94 6877.985 8613.565 ;
      RECT 6869.305 187.94 6869.585 8613.565 ;
      RECT 6855.305 187.94 6868.325 8613.565 ;
      RECT 6855.445 187.44 6868.325 8613.565 ;
      RECT 6853.065 187.94 6853.345 8613.565 ;
      RECT 6851.945 187.94 6852.225 8613.565 ;
      RECT 6850.825 187.94 6851.105 8613.565 ;
      RECT 6843.545 187.94 6843.825 8613.565 ;
      RECT 6803.365 187.94 6842.705 8613.565 ;
      RECT 6802.105 187.94 6802.385 8613.565 ;
      RECT 6797.065 187.94 6797.345 8613.565 ;
      RECT 6795.945 187.94 6796.225 8613.565 ;
      RECT 6781.525 187.44 6789.365 8613.565 ;
      RECT 6779.145 187.94 6779.425 8613.565 ;
      RECT 6778.025 187.94 6778.305 8613.565 ;
      RECT 6775.785 187.94 6776.065 8613.565 ;
      RECT 6774.665 187.94 6774.945 8613.565 ;
      RECT 6771.725 187.94 6773.825 8613.565 ;
      RECT 6742.325 187.44 6767.245 8613.565 ;
      RECT 6738.825 187.94 6739.105 8613.565 ;
      RECT 6737.705 187.94 6737.985 8613.565 ;
      RECT 6736.585 187.94 6736.865 8613.565 ;
      RECT 6731.545 187.94 6731.825 8613.565 ;
      RECT 6730.425 187.94 6730.705 8613.565 ;
      RECT 6716.005 187.44 6728.325 8613.565 ;
      RECT 6709.145 187.94 6709.425 8613.565 ;
      RECT 6708.025 187.94 6708.305 8613.565 ;
      RECT 6705.785 187.94 6706.065 8613.565 ;
      RECT 6704.665 187.94 6704.945 8613.565 ;
      RECT 6703.545 187.94 6703.825 8613.565 ;
      RECT 6662.805 187.44 6702.005 8613.565 ;
      RECT 6656.505 187.94 6656.785 8613.565 ;
      RECT 6655.385 187.94 6655.665 8613.565 ;
      RECT 6654.265 187.94 6654.545 8613.565 ;
      RECT 6640.825 187.94 6649.365 8613.565 ;
      RECT 6640.965 187.44 6649.365 8613.565 ;
      RECT 6639.705 187.94 6639.985 8613.565 ;
      RECT 6631.725 187.44 6633.125 8613.565 ;
      RECT 6629.345 187.94 6629.625 8613.565 ;
      RECT 6628.225 187.94 6628.505 8613.565 ;
      RECT 6601.205 187.44 6626.685 8613.565 ;
      RECT 6599.945 187.94 6600.225 8613.565 ;
      RECT 6598.825 187.94 6599.105 8613.565 ;
      RECT 6597.705 187.94 6597.985 8613.565 ;
      RECT 6590.425 187.94 6590.705 8613.565 ;
      RECT 6589.305 187.94 6589.585 8613.565 ;
      RECT 6574.745 187.94 6588.325 8613.565 ;
      RECT 6574.885 187.44 6588.325 8613.565 ;
      RECT 6569.705 187.94 6569.985 8613.565 ;
      RECT 6568.585 187.94 6568.865 8613.565 ;
      RECT 6523.925 187.44 6562.005 8613.565 ;
      RECT 6521.545 187.94 6521.825 8613.565 ;
      RECT 6520.425 187.94 6520.705 8613.565 ;
      RECT 6518.185 187.94 6518.465 8613.565 ;
      RECT 6517.065 187.94 6517.345 8613.565 ;
      RECT 6515.945 187.94 6516.225 8613.565 ;
      RECT 6501.525 187.44 6509.365 8613.565 ;
      RECT 6500.265 187.94 6500.545 8613.565 ;
      RECT 6499.145 187.94 6499.425 8613.565 ;
      RECT 6498.025 187.94 6498.305 8613.565 ;
      RECT 6491.025 187.94 6493.125 8613.565 ;
      RECT 6491.165 187.44 6493.125 8613.565 ;
      RECT 6489.905 187.94 6490.185 8613.565 ;
      RECT 6461.765 187.44 6486.685 8613.565 ;
      RECT 6456.025 187.94 6456.305 8613.565 ;
      RECT 6454.905 187.94 6455.185 8613.565 ;
      RECT 6452.665 187.94 6452.945 8613.565 ;
      RECT 6451.545 187.94 6451.825 8613.565 ;
      RECT 6450.425 187.94 6450.705 8613.565 ;
      RECT 6435.445 187.44 6447.765 8613.565 ;
      RECT 6430.265 187.94 6430.545 8613.565 ;
      RECT 6429.145 187.94 6429.425 8613.565 ;
      RECT 6428.025 187.94 6428.305 8613.565 ;
      RECT 6422.985 187.94 6423.265 8613.565 ;
      RECT 6383.365 187.94 6422.145 8613.565 ;
      RECT 6374.825 187.94 6375.105 8613.565 ;
      RECT 6373.705 187.94 6373.985 8613.565 ;
      RECT 6371.465 187.94 6371.745 8613.565 ;
      RECT 6370.345 187.94 6370.625 8613.565 ;
      RECT 6360.825 187.94 6369.365 8613.565 ;
      RECT 6360.965 187.44 6369.365 8613.565 ;
      RECT 6351.725 187.94 6353.825 8613.565 ;
      RECT 6350.465 187.94 6350.745 8613.565 ;
      RECT 6349.345 187.94 6349.625 8613.565 ;
      RECT 6322.325 187.44 6347.245 8613.565 ;
      RECT 6318.825 187.94 6319.105 8613.565 ;
      RECT 6317.705 187.94 6317.985 8613.565 ;
      RECT 6309.305 187.94 6309.585 8613.565 ;
      RECT 6295.305 187.94 6308.325 8613.565 ;
      RECT 6295.445 187.44 6308.325 8613.565 ;
      RECT 6293.065 187.94 6293.345 8613.565 ;
      RECT 6291.945 187.94 6292.225 8613.565 ;
      RECT 6290.825 187.94 6291.105 8613.565 ;
      RECT 6283.545 187.94 6283.825 8613.565 ;
      RECT 6243.365 187.94 6282.705 8613.565 ;
      RECT 6242.105 187.94 6242.385 8613.565 ;
      RECT 6237.065 187.94 6237.345 8613.565 ;
      RECT 6235.945 187.94 6236.225 8613.565 ;
      RECT 6221.525 187.44 6229.365 8613.565 ;
      RECT 6219.145 187.94 6219.425 8613.565 ;
      RECT 6218.025 187.94 6218.305 8613.565 ;
      RECT 6215.785 187.94 6216.065 8613.565 ;
      RECT 6214.665 187.94 6214.945 8613.565 ;
      RECT 6211.725 187.94 6213.825 8613.565 ;
      RECT 6182.325 187.44 6207.245 8613.565 ;
      RECT 6178.825 187.94 6179.105 8613.565 ;
      RECT 6177.705 187.94 6177.985 8613.565 ;
      RECT 6176.585 187.94 6176.865 8613.565 ;
      RECT 6171.545 187.94 6171.825 8613.565 ;
      RECT 6170.425 187.94 6170.705 8613.565 ;
      RECT 6156.005 187.44 6168.325 8613.565 ;
      RECT 6149.145 187.94 6149.425 8613.565 ;
      RECT 6148.025 187.94 6148.305 8613.565 ;
      RECT 6145.785 187.94 6146.065 8613.565 ;
      RECT 6144.665 187.94 6144.945 8613.565 ;
      RECT 6143.545 187.94 6143.825 8613.565 ;
      RECT 6102.805 187.44 6142.005 8613.565 ;
      RECT 6096.505 187.94 6096.785 8613.565 ;
      RECT 6095.385 187.94 6095.665 8613.565 ;
      RECT 6094.265 187.94 6094.545 8613.565 ;
      RECT 6080.825 187.94 6089.365 8613.565 ;
      RECT 6080.965 187.44 6089.365 8613.565 ;
      RECT 6079.705 187.94 6079.985 8613.565 ;
      RECT 6071.725 187.44 6073.125 8613.565 ;
      RECT 6069.345 187.94 6069.625 8613.565 ;
      RECT 6068.225 187.94 6068.505 8613.565 ;
      RECT 6041.205 187.44 6066.685 8613.565 ;
      RECT 6039.945 187.94 6040.225 8613.565 ;
      RECT 6038.825 187.94 6039.105 8613.565 ;
      RECT 6037.705 187.94 6037.985 8613.565 ;
      RECT 6030.425 187.94 6030.705 8613.565 ;
      RECT 6029.305 187.94 6029.585 8613.565 ;
      RECT 6014.745 187.94 6028.325 8613.565 ;
      RECT 6014.885 187.44 6028.325 8613.565 ;
      RECT 6009.705 187.94 6009.985 8613.565 ;
      RECT 6008.585 187.94 6008.865 8613.565 ;
      RECT 5963.925 187.44 6002.005 8613.565 ;
      RECT 5961.545 187.94 5961.825 8613.565 ;
      RECT 5960.425 187.94 5960.705 8613.565 ;
      RECT 5958.185 187.94 5958.465 8613.565 ;
      RECT 5957.065 187.94 5957.345 8613.565 ;
      RECT 5955.945 187.94 5956.225 8613.565 ;
      RECT 5941.525 187.44 5949.365 8613.565 ;
      RECT 5940.265 187.94 5940.545 8613.565 ;
      RECT 5939.145 187.94 5939.425 8613.565 ;
      RECT 5938.025 187.94 5938.305 8613.565 ;
      RECT 5931.025 187.94 5933.125 8613.565 ;
      RECT 5931.165 187.44 5933.125 8613.565 ;
      RECT 5929.905 187.94 5930.185 8613.565 ;
      RECT 5901.765 187.44 5926.685 8613.565 ;
      RECT 5896.025 187.94 5896.305 8613.565 ;
      RECT 5894.905 187.94 5895.185 8613.565 ;
      RECT 5892.665 187.94 5892.945 8613.565 ;
      RECT 5891.545 187.94 5891.825 8613.565 ;
      RECT 5890.425 187.94 5890.705 8613.565 ;
      RECT 5875.445 187.44 5887.765 8613.565 ;
      RECT 5870.265 187.94 5870.545 8613.565 ;
      RECT 5869.145 187.94 5869.425 8613.565 ;
      RECT 5868.025 187.94 5868.305 8613.565 ;
      RECT 5862.985 187.94 5863.265 8613.565 ;
      RECT 5823.365 187.94 5862.145 8613.565 ;
      RECT 5814.825 187.94 5815.105 8613.565 ;
      RECT 5813.705 187.94 5813.985 8613.565 ;
      RECT 5811.465 187.94 5811.745 8613.565 ;
      RECT 5810.345 187.94 5810.625 8613.565 ;
      RECT 5800.825 187.94 5809.365 8613.565 ;
      RECT 5800.965 187.44 5809.365 8613.565 ;
      RECT 5791.725 187.94 5793.825 8613.565 ;
      RECT 5790.465 187.94 5790.745 8613.565 ;
      RECT 5789.345 187.94 5789.625 8613.565 ;
      RECT 5762.325 187.44 5787.245 8613.565 ;
      RECT 5758.825 187.94 5759.105 8613.565 ;
      RECT 5757.705 187.94 5757.985 8613.565 ;
      RECT 5749.305 187.94 5749.585 8613.565 ;
      RECT 5735.305 187.94 5748.325 8613.565 ;
      RECT 5735.445 187.44 5748.325 8613.565 ;
      RECT 5733.065 187.94 5733.345 8613.565 ;
      RECT 5731.945 187.94 5732.225 8613.565 ;
      RECT 5730.825 187.94 5731.105 8613.565 ;
      RECT 5723.545 187.94 5723.825 8613.565 ;
      RECT 5683.365 187.94 5722.705 8613.565 ;
      RECT 5682.105 187.94 5682.385 8613.565 ;
      RECT 5677.065 187.94 5677.345 8613.565 ;
      RECT 5675.945 187.94 5676.225 8613.565 ;
      RECT 5661.525 187.44 5669.365 8613.565 ;
      RECT 5659.145 187.94 5659.425 8613.565 ;
      RECT 5658.025 187.94 5658.305 8613.565 ;
      RECT 5655.785 187.94 5656.065 8613.565 ;
      RECT 5654.665 187.94 5654.945 8613.565 ;
      RECT 5651.725 187.94 5653.825 8613.565 ;
      RECT 5622.325 187.44 5647.245 8613.565 ;
      RECT 5618.825 187.94 5619.105 8613.565 ;
      RECT 5617.705 187.94 5617.985 8613.565 ;
      RECT 5616.585 187.94 5616.865 8613.565 ;
      RECT 5611.545 187.94 5611.825 8613.565 ;
      RECT 5610.425 187.94 5610.705 8613.565 ;
      RECT 5596.005 187.44 5608.325 8613.565 ;
      RECT 5589.145 187.94 5589.425 8613.565 ;
      RECT 5588.025 187.94 5588.305 8613.565 ;
      RECT 5585.785 187.94 5586.065 8613.565 ;
      RECT 5584.665 187.94 5584.945 8613.565 ;
      RECT 5583.545 187.94 5583.825 8613.565 ;
      RECT 5542.805 187.44 5582.005 8613.565 ;
      RECT 5536.505 187.94 5536.785 8613.565 ;
      RECT 5535.385 187.94 5535.665 8613.565 ;
      RECT 5534.265 187.94 5534.545 8613.565 ;
      RECT 5520.825 187.94 5529.365 8613.565 ;
      RECT 5520.965 187.44 5529.365 8613.565 ;
      RECT 5519.705 187.94 5519.985 8613.565 ;
      RECT 5511.725 187.44 5513.125 8613.565 ;
      RECT 5509.345 187.94 5509.625 8613.565 ;
      RECT 5508.225 187.94 5508.505 8613.565 ;
      RECT 5481.205 187.44 5506.685 8613.565 ;
      RECT 5479.945 187.94 5480.225 8613.565 ;
      RECT 5478.825 187.94 5479.105 8613.565 ;
      RECT 5477.705 187.94 5477.985 8613.565 ;
      RECT 5470.425 187.94 5470.705 8613.565 ;
      RECT 5469.305 187.94 5469.585 8613.565 ;
      RECT 5454.745 187.94 5468.325 8613.565 ;
      RECT 5454.885 187.44 5468.325 8613.565 ;
      RECT 5449.705 187.94 5449.985 8613.565 ;
      RECT 5448.585 187.94 5448.865 8613.565 ;
      RECT 5403.925 187.44 5442.005 8613.565 ;
      RECT 5401.545 187.94 5401.825 8613.565 ;
      RECT 5400.425 187.94 5400.705 8613.565 ;
      RECT 5398.185 187.94 5398.465 8613.565 ;
      RECT 5397.065 187.94 5397.345 8613.565 ;
      RECT 5395.945 187.94 5396.225 8613.565 ;
      RECT 5381.525 187.44 5389.365 8613.565 ;
      RECT 5380.265 187.94 5380.545 8613.565 ;
      RECT 5379.145 187.94 5379.425 8613.565 ;
      RECT 5378.025 187.94 5378.305 8613.565 ;
      RECT 5371.025 187.94 5373.125 8613.565 ;
      RECT 5371.165 187.44 5373.125 8613.565 ;
      RECT 5369.905 187.94 5370.185 8613.565 ;
      RECT 5341.765 187.44 5366.685 8613.565 ;
      RECT 5336.025 187.94 5336.305 8613.565 ;
      RECT 5334.905 187.94 5335.185 8613.565 ;
      RECT 5332.665 187.94 5332.945 8613.565 ;
      RECT 5331.545 187.94 5331.825 8613.565 ;
      RECT 5330.425 187.94 5330.705 8613.565 ;
      RECT 5315.445 187.44 5327.765 8613.565 ;
      RECT 5310.265 187.94 5310.545 8613.565 ;
      RECT 5309.145 187.94 5309.425 8613.565 ;
      RECT 5308.025 187.94 5308.305 8613.565 ;
      RECT 5302.985 187.94 5303.265 8613.565 ;
      RECT 5263.365 187.94 5302.145 8613.565 ;
      RECT 5254.825 187.94 5255.105 8613.565 ;
      RECT 5253.705 187.94 5253.985 8613.565 ;
      RECT 5251.465 187.94 5251.745 8613.565 ;
      RECT 5250.345 187.94 5250.625 8613.565 ;
      RECT 5240.825 187.94 5249.365 8613.565 ;
      RECT 5240.965 187.44 5249.365 8613.565 ;
      RECT 5231.725 187.94 5233.825 8613.565 ;
      RECT 5230.465 187.94 5230.745 8613.565 ;
      RECT 5229.345 187.94 5229.625 8613.565 ;
      RECT 5202.325 187.44 5227.245 8613.565 ;
      RECT 5198.825 187.94 5199.105 8613.565 ;
      RECT 5197.705 187.94 5197.985 8613.565 ;
      RECT 5189.305 187.94 5189.585 8613.565 ;
      RECT 5175.305 187.94 5188.325 8613.565 ;
      RECT 5175.445 187.44 5188.325 8613.565 ;
      RECT 5173.065 187.94 5173.345 8613.565 ;
      RECT 5171.945 187.94 5172.225 8613.565 ;
      RECT 5170.825 187.94 5171.105 8613.565 ;
      RECT 5163.545 187.94 5163.825 8613.565 ;
      RECT 5123.365 187.94 5162.705 8613.565 ;
      RECT 5122.105 187.94 5122.385 8613.565 ;
      RECT 5117.065 187.94 5117.345 8613.565 ;
      RECT 5115.945 187.94 5116.225 8613.565 ;
      RECT 5101.525 187.44 5109.365 8613.565 ;
      RECT 5099.145 187.94 5099.425 8613.565 ;
      RECT 5098.025 187.94 5098.305 8613.565 ;
      RECT 5095.785 187.94 5096.065 8613.565 ;
      RECT 5094.665 187.94 5094.945 8613.565 ;
      RECT 5091.725 187.94 5093.825 8613.565 ;
      RECT 5062.325 187.44 5087.245 8613.565 ;
      RECT 5058.825 187.94 5059.105 8613.565 ;
      RECT 5057.705 187.94 5057.985 8613.565 ;
      RECT 5056.585 187.94 5056.865 8613.565 ;
      RECT 5051.545 187.94 5051.825 8613.565 ;
      RECT 5050.425 187.94 5050.705 8613.565 ;
      RECT 5036.005 187.44 5048.325 8613.565 ;
      RECT 5029.145 187.94 5029.425 8613.565 ;
      RECT 5028.025 187.94 5028.305 8613.565 ;
      RECT 5025.785 187.94 5026.065 8613.565 ;
      RECT 5024.665 187.94 5024.945 8613.565 ;
      RECT 5023.545 187.94 5023.825 8613.565 ;
      RECT 4982.805 187.44 5022.005 8613.565 ;
      RECT 4976.505 187.94 4976.785 8613.565 ;
      RECT 4975.385 187.94 4975.665 8613.565 ;
      RECT 4974.265 187.94 4974.545 8613.565 ;
      RECT 4960.825 187.94 4969.365 8613.565 ;
      RECT 4960.965 187.44 4969.365 8613.565 ;
      RECT 4959.705 187.94 4959.985 8613.565 ;
      RECT 4951.725 187.44 4953.125 8613.565 ;
      RECT 4949.345 187.94 4949.625 8613.565 ;
      RECT 4948.225 187.94 4948.505 8613.565 ;
      RECT 4921.205 187.44 4946.685 8613.565 ;
      RECT 4919.945 187.94 4920.225 8613.565 ;
      RECT 4918.825 187.94 4919.105 8613.565 ;
      RECT 4917.705 187.94 4917.985 8613.565 ;
      RECT 4910.425 187.94 4910.705 8613.565 ;
      RECT 4909.305 187.94 4909.585 8613.565 ;
      RECT 4894.745 187.94 4908.325 8613.565 ;
      RECT 4894.885 187.44 4908.325 8613.565 ;
      RECT 4889.705 187.94 4889.985 8613.565 ;
      RECT 4888.585 187.94 4888.865 8613.565 ;
      RECT 4843.925 187.44 4882.005 8613.565 ;
      RECT 4841.545 187.94 4841.825 8613.565 ;
      RECT 4840.425 187.94 4840.705 8613.565 ;
      RECT 4838.185 187.94 4838.465 8613.565 ;
      RECT 4837.065 187.94 4837.345 8613.565 ;
      RECT 4835.945 187.94 4836.225 8613.565 ;
      RECT 4821.525 187.44 4829.365 8613.565 ;
      RECT 4820.265 187.94 4820.545 8613.565 ;
      RECT 4819.145 187.94 4819.425 8613.565 ;
      RECT 4818.025 187.94 4818.305 8613.565 ;
      RECT 4811.025 187.94 4813.125 8613.565 ;
      RECT 4811.165 187.44 4813.125 8613.565 ;
      RECT 4809.905 187.94 4810.185 8613.565 ;
      RECT 4781.765 187.44 4806.685 8613.565 ;
      RECT 4776.025 187.94 4776.305 8613.565 ;
      RECT 4774.905 187.94 4775.185 8613.565 ;
      RECT 4772.665 187.94 4772.945 8613.565 ;
      RECT 4771.545 187.94 4771.825 8613.565 ;
      RECT 4770.425 187.94 4770.705 8613.565 ;
      RECT 4755.445 187.44 4767.765 8613.565 ;
      RECT 4750.265 187.94 4750.545 8613.565 ;
      RECT 4749.145 187.94 4749.425 8613.565 ;
      RECT 4748.025 187.94 4748.305 8613.565 ;
      RECT 4742.985 187.94 4743.265 8613.565 ;
      RECT 4703.365 187.94 4742.145 8613.565 ;
      RECT 4694.825 187.94 4695.105 8613.565 ;
      RECT 4693.705 187.94 4693.985 8613.565 ;
      RECT 4691.465 187.94 4691.745 8613.565 ;
      RECT 4690.345 187.94 4690.625 8613.565 ;
      RECT 4680.825 187.94 4689.365 8613.565 ;
      RECT 4680.965 187.44 4689.365 8613.565 ;
      RECT 4671.725 187.94 4673.825 8613.565 ;
      RECT 4670.465 187.94 4670.745 8613.565 ;
      RECT 4669.345 187.94 4669.625 8613.565 ;
      RECT 4642.325 187.44 4667.245 8613.565 ;
      RECT 4638.825 187.94 4639.105 8613.565 ;
      RECT 4637.705 187.94 4637.985 8613.565 ;
      RECT 4629.305 187.94 4629.585 8613.565 ;
      RECT 4615.305 187.94 4628.325 8613.565 ;
      RECT 4615.445 187.44 4628.325 8613.565 ;
      RECT 4613.065 187.94 4613.345 8613.565 ;
      RECT 4611.945 187.94 4612.225 8613.565 ;
      RECT 4610.825 187.94 4611.105 8613.565 ;
      RECT 4603.545 187.94 4603.825 8613.565 ;
      RECT 4563.365 187.94 4602.705 8613.565 ;
      RECT 4562.105 187.94 4562.385 8613.565 ;
      RECT 4557.065 187.94 4557.345 8613.565 ;
      RECT 4555.945 187.94 4556.225 8613.565 ;
      RECT 4541.525 187.44 4549.365 8613.565 ;
      RECT 4539.145 187.94 4539.425 8613.565 ;
      RECT 4538.025 187.94 4538.305 8613.565 ;
      RECT 4535.785 187.94 4536.065 8613.565 ;
      RECT 4534.665 187.94 4534.945 8613.565 ;
      RECT 4531.725 187.94 4533.825 8613.565 ;
      RECT 4502.325 187.44 4527.245 8613.565 ;
      RECT 4498.825 187.94 4499.105 8613.565 ;
      RECT 4497.705 187.94 4497.985 8613.565 ;
      RECT 4496.585 187.94 4496.865 8613.565 ;
      RECT 4491.545 187.94 4491.825 8613.565 ;
      RECT 4490.425 187.94 4490.705 8613.565 ;
      RECT 4476.005 187.44 4488.325 8613.565 ;
      RECT 4469.145 187.94 4469.425 8613.565 ;
      RECT 4468.025 187.94 4468.305 8613.565 ;
      RECT 4465.785 187.94 4466.065 8613.565 ;
      RECT 4464.665 187.94 4464.945 8613.565 ;
      RECT 4463.545 187.94 4463.825 8613.565 ;
      RECT 4422.805 187.44 4462.005 8613.565 ;
      RECT 4416.505 187.94 4416.785 8613.565 ;
      RECT 4415.385 187.94 4415.665 8613.565 ;
      RECT 4414.265 187.94 4414.545 8613.565 ;
      RECT 4400.825 187.94 4409.365 8613.565 ;
      RECT 4400.965 187.44 4409.365 8613.565 ;
      RECT 4399.705 187.94 4399.985 8613.565 ;
      RECT 4391.725 187.44 4393.125 8613.565 ;
      RECT 4389.345 187.94 4389.625 8613.565 ;
      RECT 4388.225 187.94 4388.505 8613.565 ;
      RECT 4361.205 187.44 4386.685 8613.565 ;
      RECT 4359.945 187.94 4360.225 8613.565 ;
      RECT 4358.825 187.94 4359.105 8613.565 ;
      RECT 4357.705 187.94 4357.985 8613.565 ;
      RECT 4350.425 187.94 4350.705 8613.565 ;
      RECT 4349.305 187.94 4349.585 8613.565 ;
      RECT 4334.745 187.94 4348.325 8613.565 ;
      RECT 4334.885 187.44 4348.325 8613.565 ;
      RECT 4329.705 187.94 4329.985 8613.565 ;
      RECT 4328.585 187.94 4328.865 8613.565 ;
      RECT 4283.925 187.44 4322.005 8613.565 ;
      RECT 4281.545 187.94 4281.825 8613.565 ;
      RECT 4280.425 187.94 4280.705 8613.565 ;
      RECT 4278.185 187.94 4278.465 8613.565 ;
      RECT 4277.065 187.94 4277.345 8613.565 ;
      RECT 4275.945 187.94 4276.225 8613.565 ;
      RECT 4261.525 187.44 4269.365 8613.565 ;
      RECT 4260.265 187.94 4260.545 8613.565 ;
      RECT 4259.145 187.94 4259.425 8613.565 ;
      RECT 4258.025 187.94 4258.305 8613.565 ;
      RECT 4251.025 187.94 4253.125 8613.565 ;
      RECT 4251.165 187.44 4253.125 8613.565 ;
      RECT 4249.905 187.94 4250.185 8613.565 ;
      RECT 4221.765 187.44 4246.685 8613.565 ;
      RECT 4216.025 187.94 4216.305 8613.565 ;
      RECT 4214.905 187.94 4215.185 8613.565 ;
      RECT 4212.665 187.94 4212.945 8613.565 ;
      RECT 4211.545 187.94 4211.825 8613.565 ;
      RECT 4210.425 187.94 4210.705 8613.565 ;
      RECT 4195.445 187.44 4207.765 8613.565 ;
      RECT 4190.265 187.94 4190.545 8613.565 ;
      RECT 4189.145 187.94 4189.425 8613.565 ;
      RECT 4188.025 187.94 4188.305 8613.565 ;
      RECT 4182.985 187.94 4183.265 8613.565 ;
      RECT 4143.365 187.94 4182.145 8613.565 ;
      RECT 4134.825 187.94 4135.105 8613.565 ;
      RECT 4133.705 187.94 4133.985 8613.565 ;
      RECT 4131.465 187.94 4131.745 8613.565 ;
      RECT 4130.345 187.94 4130.625 8613.565 ;
      RECT 4120.825 187.94 4129.365 8613.565 ;
      RECT 4120.965 187.44 4129.365 8613.565 ;
      RECT 4111.725 187.94 4113.825 8613.565 ;
      RECT 4110.465 187.94 4110.745 8613.565 ;
      RECT 4109.345 187.94 4109.625 8613.565 ;
      RECT 4082.325 187.44 4107.245 8613.565 ;
      RECT 4078.825 187.94 4079.105 8613.565 ;
      RECT 4077.705 187.94 4077.985 8613.565 ;
      RECT 4069.305 187.94 4069.585 8613.565 ;
      RECT 4055.305 187.94 4068.325 8613.565 ;
      RECT 4055.445 187.44 4068.325 8613.565 ;
      RECT 4053.065 187.94 4053.345 8613.565 ;
      RECT 4051.945 187.94 4052.225 8613.565 ;
      RECT 4050.825 187.94 4051.105 8613.565 ;
      RECT 4043.545 187.94 4043.825 8613.565 ;
      RECT 4003.365 187.94 4042.705 8613.565 ;
      RECT 4002.105 187.94 4002.385 8613.565 ;
      RECT 3997.065 187.94 3997.345 8613.565 ;
      RECT 3995.945 187.94 3996.225 8613.565 ;
      RECT 3981.525 187.44 3989.365 8613.565 ;
      RECT 3979.145 187.94 3979.425 8613.565 ;
      RECT 3978.025 187.94 3978.305 8613.565 ;
      RECT 3975.785 187.94 3976.065 8613.565 ;
      RECT 3974.665 187.94 3974.945 8613.565 ;
      RECT 3971.725 187.94 3973.825 8613.565 ;
      RECT 3942.325 187.44 3967.245 8613.565 ;
      RECT 3938.825 187.94 3939.105 8613.565 ;
      RECT 3937.705 187.94 3937.985 8613.565 ;
      RECT 3936.585 187.94 3936.865 8613.565 ;
      RECT 3931.545 187.94 3931.825 8613.565 ;
      RECT 3930.425 187.94 3930.705 8613.565 ;
      RECT 3916.005 187.44 3928.325 8613.565 ;
      RECT 3909.145 187.94 3909.425 8613.565 ;
      RECT 3908.025 187.94 3908.305 8613.565 ;
      RECT 3905.785 187.94 3906.065 8613.565 ;
      RECT 3904.665 187.94 3904.945 8613.565 ;
      RECT 3903.545 187.94 3903.825 8613.565 ;
      RECT 3862.805 187.44 3902.005 8613.565 ;
      RECT 3856.505 187.94 3856.785 8613.565 ;
      RECT 3855.385 187.94 3855.665 8613.565 ;
      RECT 3854.265 187.94 3854.545 8613.565 ;
      RECT 3840.825 187.94 3849.365 8613.565 ;
      RECT 3840.965 187.44 3849.365 8613.565 ;
      RECT 3839.705 187.94 3839.985 8613.565 ;
      RECT 3831.725 187.44 3833.125 8613.565 ;
      RECT 3829.345 187.94 3829.625 8613.565 ;
      RECT 3828.225 187.94 3828.505 8613.565 ;
      RECT 3801.205 187.44 3826.685 8613.565 ;
      RECT 3799.945 187.94 3800.225 8613.565 ;
      RECT 3798.825 187.94 3799.105 8613.565 ;
      RECT 3797.705 187.94 3797.985 8613.565 ;
      RECT 3790.425 187.94 3790.705 8613.565 ;
      RECT 3789.305 187.94 3789.585 8613.565 ;
      RECT 3774.745 187.94 3788.325 8613.565 ;
      RECT 3774.885 187.44 3788.325 8613.565 ;
      RECT 3769.705 187.94 3769.985 8613.565 ;
      RECT 3768.585 187.94 3768.865 8613.565 ;
      RECT 3723.925 187.44 3762.005 8613.565 ;
      RECT 3721.545 187.94 3721.825 8613.565 ;
      RECT 3720.425 187.94 3720.705 8613.565 ;
      RECT 3718.185 187.94 3718.465 8613.565 ;
      RECT 3717.065 187.94 3717.345 8613.565 ;
      RECT 3715.945 187.94 3716.225 8613.565 ;
      RECT 3701.525 187.44 3709.365 8613.565 ;
      RECT 3700.265 187.94 3700.545 8613.565 ;
      RECT 3699.145 187.94 3699.425 8613.565 ;
      RECT 3698.025 187.94 3698.305 8613.565 ;
      RECT 3691.025 187.94 3693.125 8613.565 ;
      RECT 3691.165 187.44 3693.125 8613.565 ;
      RECT 3689.905 187.94 3690.185 8613.565 ;
      RECT 3661.765 187.44 3686.685 8613.565 ;
      RECT 3656.025 187.94 3656.305 8613.565 ;
      RECT 3654.905 187.94 3655.185 8613.565 ;
      RECT 3652.665 187.94 3652.945 8613.565 ;
      RECT 3651.545 187.94 3651.825 8613.565 ;
      RECT 3650.425 187.94 3650.705 8613.565 ;
      RECT 3635.445 187.44 3647.765 8613.565 ;
      RECT 3630.265 187.94 3630.545 8613.565 ;
      RECT 3629.145 187.94 3629.425 8613.565 ;
      RECT 3628.025 187.94 3628.305 8613.565 ;
      RECT 3622.985 187.94 3623.265 8613.565 ;
      RECT 3583.365 187.94 3622.145 8613.565 ;
      RECT 3574.825 187.94 3575.105 8613.565 ;
      RECT 3573.705 187.94 3573.985 8613.565 ;
      RECT 3571.465 187.94 3571.745 8613.565 ;
      RECT 3570.345 187.94 3570.625 8613.565 ;
      RECT 3560.825 187.94 3569.365 8613.565 ;
      RECT 3560.965 187.44 3569.365 8613.565 ;
      RECT 3551.725 187.94 3553.825 8613.565 ;
      RECT 3550.465 187.94 3550.745 8613.565 ;
      RECT 3549.345 187.94 3549.625 8613.565 ;
      RECT 3522.325 187.44 3547.245 8613.565 ;
      RECT 3518.825 187.94 3519.105 8613.565 ;
      RECT 3517.705 187.94 3517.985 8613.565 ;
      RECT 3509.305 187.94 3509.585 8613.565 ;
      RECT 3495.305 187.94 3508.325 8613.565 ;
      RECT 3495.445 187.44 3508.325 8613.565 ;
      RECT 3493.065 187.94 3493.345 8613.565 ;
      RECT 3491.945 187.94 3492.225 8613.565 ;
      RECT 3490.825 187.94 3491.105 8613.565 ;
      RECT 3483.545 187.94 3483.825 8613.565 ;
      RECT 3443.365 187.94 3482.705 8613.565 ;
      RECT 3442.105 187.94 3442.385 8613.565 ;
      RECT 3437.065 187.94 3437.345 8613.565 ;
      RECT 3435.945 187.94 3436.225 8613.565 ;
      RECT 3421.525 187.44 3429.365 8613.565 ;
      RECT 3419.145 187.94 3419.425 8613.565 ;
      RECT 3418.025 187.94 3418.305 8613.565 ;
      RECT 3415.785 187.94 3416.065 8613.565 ;
      RECT 3414.665 187.94 3414.945 8613.565 ;
      RECT 3411.725 187.94 3413.825 8613.565 ;
      RECT 3382.325 187.44 3407.245 8613.565 ;
      RECT 3378.825 187.94 3379.105 8613.565 ;
      RECT 3377.705 187.94 3377.985 8613.565 ;
      RECT 3376.585 187.94 3376.865 8613.565 ;
      RECT 3371.545 187.94 3371.825 8613.565 ;
      RECT 3370.425 187.94 3370.705 8613.565 ;
      RECT 3356.005 187.44 3368.325 8613.565 ;
      RECT 3349.145 187.94 3349.425 8613.565 ;
      RECT 3348.025 187.94 3348.305 8613.565 ;
      RECT 3345.785 187.94 3346.065 8613.565 ;
      RECT 3344.665 187.94 3344.945 8613.565 ;
      RECT 3343.545 187.94 3343.825 8613.565 ;
      RECT 3302.805 187.44 3342.005 8613.565 ;
      RECT 3296.505 187.94 3296.785 8613.565 ;
      RECT 3295.385 187.94 3295.665 8613.565 ;
      RECT 3294.265 187.94 3294.545 8613.565 ;
      RECT 3280.825 187.94 3289.365 8613.565 ;
      RECT 3280.965 187.44 3289.365 8613.565 ;
      RECT 3279.705 187.94 3279.985 8613.565 ;
      RECT 3271.725 187.44 3273.125 8613.565 ;
      RECT 3269.345 187.94 3269.625 8613.565 ;
      RECT 3268.225 187.94 3268.505 8613.565 ;
      RECT 3241.205 187.44 3266.685 8613.565 ;
      RECT 3239.945 187.94 3240.225 8613.565 ;
      RECT 3238.825 187.94 3239.105 8613.565 ;
      RECT 3237.705 187.94 3237.985 8613.565 ;
      RECT 3230.425 187.94 3230.705 8613.565 ;
      RECT 3229.305 187.94 3229.585 8613.565 ;
      RECT 3214.745 187.94 3228.325 8613.565 ;
      RECT 3214.885 187.44 3228.325 8613.565 ;
      RECT 3209.705 187.94 3209.985 8613.565 ;
      RECT 3208.585 187.94 3208.865 8613.565 ;
      RECT 3163.925 187.44 3202.005 8613.565 ;
      RECT 3161.545 187.94 3161.825 8613.565 ;
      RECT 3160.425 187.94 3160.705 8613.565 ;
      RECT 3158.185 187.94 3158.465 8613.565 ;
      RECT 3157.065 187.94 3157.345 8613.565 ;
      RECT 3155.945 187.94 3156.225 8613.565 ;
      RECT 3141.525 187.44 3149.365 8613.565 ;
      RECT 3140.265 187.94 3140.545 8613.565 ;
      RECT 3139.145 187.94 3139.425 8613.565 ;
      RECT 3138.025 187.94 3138.305 8613.565 ;
      RECT 3131.025 187.94 3133.125 8613.565 ;
      RECT 3131.165 187.44 3133.125 8613.565 ;
      RECT 3129.905 187.94 3130.185 8613.565 ;
      RECT 3101.765 187.44 3126.685 8613.565 ;
      RECT 3096.025 187.94 3096.305 8613.565 ;
      RECT 3094.905 187.94 3095.185 8613.565 ;
      RECT 3092.665 187.94 3092.945 8613.565 ;
      RECT 3091.545 187.94 3091.825 8613.565 ;
      RECT 3090.425 187.94 3090.705 8613.565 ;
      RECT 3075.445 187.44 3087.765 8613.565 ;
      RECT 3070.265 187.94 3070.545 8613.565 ;
      RECT 3069.145 187.94 3069.425 8613.565 ;
      RECT 3068.025 187.94 3068.305 8613.565 ;
      RECT 3062.985 187.94 3063.265 8613.565 ;
      RECT 3023.365 187.94 3062.145 8613.565 ;
      RECT 3014.825 187.94 3015.105 8613.565 ;
      RECT 3013.705 187.94 3013.985 8613.565 ;
      RECT 3011.465 187.94 3011.745 8613.565 ;
      RECT 3010.345 187.94 3010.625 8613.565 ;
      RECT 3000.825 187.94 3009.365 8613.565 ;
      RECT 3000.965 187.44 3009.365 8613.565 ;
      RECT 2991.725 187.94 2993.825 8613.565 ;
      RECT 2990.465 187.94 2990.745 8613.565 ;
      RECT 2989.345 187.94 2989.625 8613.565 ;
      RECT 2962.325 187.44 2987.245 8613.565 ;
      RECT 2958.825 187.94 2959.105 8613.565 ;
      RECT 2957.705 187.94 2957.985 8613.565 ;
      RECT 2949.305 187.94 2949.585 8613.565 ;
      RECT 2935.305 187.94 2948.325 8613.565 ;
      RECT 2935.445 187.44 2948.325 8613.565 ;
      RECT 2933.065 187.94 2933.345 8613.565 ;
      RECT 2931.945 187.94 2932.225 8613.565 ;
      RECT 2930.825 187.94 2931.105 8613.565 ;
      RECT 2923.545 187.94 2923.825 8613.565 ;
      RECT 2883.365 187.94 2922.705 8613.565 ;
      RECT 2882.105 187.94 2882.385 8613.565 ;
      RECT 2877.065 187.94 2877.345 8613.565 ;
      RECT 2875.945 187.94 2876.225 8613.565 ;
      RECT 2861.525 187.44 2869.365 8613.565 ;
      RECT 2859.145 187.94 2859.425 8613.565 ;
      RECT 2858.025 187.94 2858.305 8613.565 ;
      RECT 2855.785 187.94 2856.065 8613.565 ;
      RECT 2854.665 187.94 2854.945 8613.565 ;
      RECT 2851.725 187.94 2853.825 8613.565 ;
      RECT 2822.325 187.44 2847.245 8613.565 ;
      RECT 2818.825 187.94 2819.105 8613.565 ;
      RECT 2817.705 187.94 2817.985 8613.565 ;
      RECT 2816.585 187.94 2816.865 8613.565 ;
      RECT 2811.545 187.94 2811.825 8613.565 ;
      RECT 2810.425 187.94 2810.705 8613.565 ;
      RECT 2796.005 187.44 2808.325 8613.565 ;
      RECT 2789.145 187.94 2789.425 8613.565 ;
      RECT 2788.025 187.94 2788.305 8613.565 ;
      RECT 2785.785 187.94 2786.065 8613.565 ;
      RECT 2784.665 187.94 2784.945 8613.565 ;
      RECT 2783.545 187.94 2783.825 8613.565 ;
      RECT 2742.805 187.44 2782.005 8613.565 ;
      RECT 2736.505 187.94 2736.785 8613.565 ;
      RECT 2735.385 187.94 2735.665 8613.565 ;
      RECT 2734.265 187.94 2734.545 8613.565 ;
      RECT 2720.825 187.94 2729.365 8613.565 ;
      RECT 2720.965 187.44 2729.365 8613.565 ;
      RECT 2719.705 187.94 2719.985 8613.565 ;
      RECT 2711.725 187.44 2713.125 8613.565 ;
      RECT 2709.345 187.94 2709.625 8613.565 ;
      RECT 2708.225 187.94 2708.505 8613.565 ;
      RECT 2681.205 187.44 2706.685 8613.565 ;
      RECT 2679.945 187.94 2680.225 8613.565 ;
      RECT 2678.825 187.94 2679.105 8613.565 ;
      RECT 2677.705 187.94 2677.985 8613.565 ;
      RECT 2670.425 187.94 2670.705 8613.565 ;
      RECT 2669.305 187.94 2669.585 8613.565 ;
      RECT 2654.745 187.94 2668.325 8613.565 ;
      RECT 2654.885 187.44 2668.325 8613.565 ;
      RECT 2649.705 187.94 2649.985 8613.565 ;
      RECT 2648.585 187.94 2648.865 8613.565 ;
      RECT 2603.925 187.44 2642.005 8613.565 ;
      RECT 2601.545 187.94 2601.825 8613.565 ;
      RECT 2600.425 187.94 2600.705 8613.565 ;
      RECT 2598.185 187.94 2598.465 8613.565 ;
      RECT 2597.065 187.94 2597.345 8613.565 ;
      RECT 2595.945 187.94 2596.225 8613.565 ;
      RECT 2581.525 187.44 2589.365 8613.565 ;
      RECT 2580.265 187.94 2580.545 8613.565 ;
      RECT 2579.145 187.94 2579.425 8613.565 ;
      RECT 2578.025 187.94 2578.305 8613.565 ;
      RECT 2571.025 187.94 2573.125 8613.565 ;
      RECT 2571.165 187.44 2573.125 8613.565 ;
      RECT 2569.905 187.94 2570.185 8613.565 ;
      RECT 2541.765 187.44 2566.685 8613.565 ;
      RECT 2536.025 187.94 2536.305 8613.565 ;
      RECT 2534.905 187.94 2535.185 8613.565 ;
      RECT 2532.665 187.94 2532.945 8613.565 ;
      RECT 2531.545 187.94 2531.825 8613.565 ;
      RECT 2530.425 187.94 2530.705 8613.565 ;
      RECT 2515.445 187.44 2527.765 8613.565 ;
      RECT 2510.265 187.94 2510.545 8613.565 ;
      RECT 2509.145 187.94 2509.425 8613.565 ;
      RECT 2508.025 187.94 2508.305 8613.565 ;
      RECT 2502.985 187.94 2503.265 8613.565 ;
      RECT 2463.365 187.94 2502.145 8613.565 ;
      RECT 2454.825 187.94 2455.105 8613.565 ;
      RECT 2453.705 187.94 2453.985 8613.565 ;
      RECT 2451.465 187.94 2451.745 8613.565 ;
      RECT 2450.345 187.94 2450.625 8613.565 ;
      RECT 2440.825 187.94 2449.365 8613.565 ;
      RECT 2440.965 187.44 2449.365 8613.565 ;
      RECT 2431.725 187.94 2433.825 8613.565 ;
      RECT 2430.465 187.94 2430.745 8613.565 ;
      RECT 2429.345 187.94 2429.625 8613.565 ;
      RECT 2402.325 187.44 2427.245 8613.565 ;
      RECT 2398.825 187.94 2399.105 8613.565 ;
      RECT 2397.705 187.94 2397.985 8613.565 ;
      RECT 2389.305 187.94 2389.585 8613.565 ;
      RECT 2375.305 187.94 2388.325 8613.565 ;
      RECT 2375.445 187.44 2388.325 8613.565 ;
      RECT 2373.065 187.94 2373.345 8613.565 ;
      RECT 2371.945 187.94 2372.225 8613.565 ;
      RECT 2370.825 187.94 2371.105 8613.565 ;
      RECT 2363.545 187.94 2363.825 8613.565 ;
      RECT 2323.365 187.94 2362.705 8613.565 ;
      RECT 2322.105 187.94 2322.385 8613.565 ;
      RECT 2317.065 187.94 2317.345 8613.565 ;
      RECT 2315.945 187.94 2316.225 8613.565 ;
      RECT 2301.525 187.44 2309.365 8613.565 ;
      RECT 2299.145 187.94 2299.425 8613.565 ;
      RECT 2298.025 187.94 2298.305 8613.565 ;
      RECT 2295.785 187.94 2296.065 8613.565 ;
      RECT 2294.665 187.94 2294.945 8613.565 ;
      RECT 2291.725 187.94 2293.825 8613.565 ;
      RECT 2262.325 187.44 2287.245 8613.565 ;
      RECT 2258.825 187.94 2259.105 8613.565 ;
      RECT 2257.705 187.94 2257.985 8613.565 ;
      RECT 2256.585 187.94 2256.865 8613.565 ;
      RECT 2251.545 187.94 2251.825 8613.565 ;
      RECT 2250.425 187.94 2250.705 8613.565 ;
      RECT 2236.005 187.44 2248.325 8613.565 ;
      RECT 2229.145 187.94 2229.425 8613.565 ;
      RECT 2228.025 187.94 2228.305 8613.565 ;
      RECT 2225.785 187.94 2226.065 8613.565 ;
      RECT 2224.665 187.94 2224.945 8613.565 ;
      RECT 2223.545 187.94 2223.825 8613.565 ;
      RECT 2182.805 187.44 2222.005 8613.565 ;
      RECT 2176.505 187.94 2176.785 8613.565 ;
      RECT 2175.385 187.94 2175.665 8613.565 ;
      RECT 2174.265 187.94 2174.545 8613.565 ;
      RECT 2160.825 187.94 2169.365 8613.565 ;
      RECT 2160.965 187.44 2169.365 8613.565 ;
      RECT 2159.705 187.94 2159.985 8613.565 ;
      RECT 2151.725 187.44 2153.125 8613.565 ;
      RECT 2149.345 187.94 2149.625 8613.565 ;
      RECT 2148.225 187.94 2148.505 8613.565 ;
      RECT 2121.205 187.44 2146.685 8613.565 ;
      RECT 2119.945 187.94 2120.225 8613.565 ;
      RECT 2118.825 187.94 2119.105 8613.565 ;
      RECT 2117.705 187.94 2117.985 8613.565 ;
      RECT 2110.425 187.94 2110.705 8613.565 ;
      RECT 2109.305 187.94 2109.585 8613.565 ;
      RECT 2094.745 187.94 2108.325 8613.565 ;
      RECT 2094.885 187.44 2108.325 8613.565 ;
      RECT 2089.705 187.94 2089.985 8613.565 ;
      RECT 2088.585 187.94 2088.865 8613.565 ;
      RECT 2043.925 187.44 2082.005 8613.565 ;
      RECT 2041.545 187.94 2041.825 8613.565 ;
      RECT 2040.425 187.94 2040.705 8613.565 ;
      RECT 2038.185 187.94 2038.465 8613.565 ;
      RECT 2037.065 187.94 2037.345 8613.565 ;
      RECT 2035.945 187.94 2036.225 8613.565 ;
      RECT 2021.525 187.44 2029.365 8613.565 ;
      RECT 2020.265 187.94 2020.545 8613.565 ;
      RECT 2019.145 187.94 2019.425 8613.565 ;
      RECT 2018.025 187.94 2018.305 8613.565 ;
      RECT 2011.025 187.94 2013.125 8613.565 ;
      RECT 2011.165 187.44 2013.125 8613.565 ;
      RECT 2009.905 187.94 2010.185 8613.565 ;
      RECT 1981.765 187.44 2006.685 8613.565 ;
      RECT 1976.025 187.94 1976.305 8613.565 ;
      RECT 1974.905 187.94 1975.185 8613.565 ;
      RECT 1972.665 187.94 1972.945 8613.565 ;
      RECT 1971.545 187.94 1971.825 8613.565 ;
      RECT 1970.425 187.94 1970.705 8613.565 ;
      RECT 1955.445 187.44 1967.765 8613.565 ;
      RECT 1950.265 187.94 1950.545 8613.565 ;
      RECT 1949.145 187.94 1949.425 8613.565 ;
      RECT 1948.025 187.94 1948.305 8613.565 ;
      RECT 1942.985 187.94 1943.265 8613.565 ;
      RECT 1903.365 187.94 1942.145 8613.565 ;
      RECT 1894.825 187.94 1895.105 8613.565 ;
      RECT 1893.705 187.94 1893.985 8613.565 ;
      RECT 1891.465 187.94 1891.745 8613.565 ;
      RECT 1890.345 187.94 1890.625 8613.565 ;
      RECT 1880.825 187.94 1889.365 8613.565 ;
      RECT 1880.965 187.44 1889.365 8613.565 ;
      RECT 1871.725 187.94 1873.825 8613.565 ;
      RECT 1870.465 187.94 1870.745 8613.565 ;
      RECT 1869.345 187.94 1869.625 8613.565 ;
      RECT 1842.325 187.44 1867.245 8613.565 ;
      RECT 1838.825 187.94 1839.105 8613.565 ;
      RECT 1837.705 187.94 1837.985 8613.565 ;
      RECT 1829.305 187.94 1829.585 8613.565 ;
      RECT 1815.305 187.94 1828.325 8613.565 ;
      RECT 1815.445 187.44 1828.325 8613.565 ;
      RECT 1813.065 187.94 1813.345 8613.565 ;
      RECT 1811.945 187.94 1812.225 8613.565 ;
      RECT 1810.825 187.94 1811.105 8613.565 ;
      RECT 1803.545 187.94 1803.825 8613.565 ;
      RECT 1763.365 187.94 1802.705 8613.565 ;
      RECT 1762.105 187.94 1762.385 8613.565 ;
      RECT 1757.065 187.94 1757.345 8613.565 ;
      RECT 1755.945 187.94 1756.225 8613.565 ;
      RECT 1741.525 187.44 1749.365 8613.565 ;
      RECT 1739.145 187.94 1739.425 8613.565 ;
      RECT 1738.025 187.94 1738.305 8613.565 ;
      RECT 1735.785 187.94 1736.065 8613.565 ;
      RECT 1734.665 187.94 1734.945 8613.565 ;
      RECT 1731.725 187.94 1733.825 8613.565 ;
      RECT 1702.325 187.44 1727.245 8613.565 ;
      RECT 1698.825 187.94 1699.105 8613.565 ;
      RECT 1697.705 187.94 1697.985 8613.565 ;
      RECT 1696.585 187.94 1696.865 8613.565 ;
      RECT 1691.545 187.94 1691.825 8613.565 ;
      RECT 1690.425 187.94 1690.705 8613.565 ;
      RECT 1676.005 187.44 1688.325 8613.565 ;
      RECT 1669.145 187.94 1669.425 8613.565 ;
      RECT 1668.025 187.94 1668.305 8613.565 ;
      RECT 1665.785 187.94 1666.065 8613.565 ;
      RECT 1664.665 187.94 1664.945 8613.565 ;
      RECT 1663.545 187.94 1663.825 8613.565 ;
      RECT 1622.805 187.44 1662.005 8613.565 ;
      RECT 1616.505 187.94 1616.785 8613.565 ;
      RECT 1615.385 187.94 1615.665 8613.565 ;
      RECT 1614.265 187.94 1614.545 8613.565 ;
      RECT 1600.825 187.94 1609.365 8613.565 ;
      RECT 1600.965 187.44 1609.365 8613.565 ;
      RECT 1599.705 187.94 1599.985 8613.565 ;
      RECT 1591.725 187.44 1593.125 8613.565 ;
      RECT 1589.345 187.94 1589.625 8613.565 ;
      RECT 1588.225 187.94 1588.505 8613.565 ;
      RECT 1561.205 187.44 1586.685 8613.565 ;
      RECT 1559.945 187.94 1560.225 8613.565 ;
      RECT 1558.825 187.94 1559.105 8613.565 ;
      RECT 1557.705 187.94 1557.985 8613.565 ;
      RECT 1550.425 187.94 1550.705 8613.565 ;
      RECT 1549.305 187.94 1549.585 8613.565 ;
      RECT 1534.745 187.94 1548.325 8613.565 ;
      RECT 1534.885 187.44 1548.325 8613.565 ;
      RECT 1529.705 187.94 1529.985 8613.565 ;
      RECT 1528.585 187.94 1528.865 8613.565 ;
      RECT 1483.925 187.44 1522.005 8613.565 ;
      RECT 1481.545 187.94 1481.825 8613.565 ;
      RECT 1480.425 187.94 1480.705 8613.565 ;
      RECT 1478.185 187.94 1478.465 8613.565 ;
      RECT 1477.065 187.94 1477.345 8613.565 ;
      RECT 1475.945 187.94 1476.225 8613.565 ;
      RECT 1461.525 187.44 1469.365 8613.565 ;
      RECT 1460.265 187.94 1460.545 8613.565 ;
      RECT 1459.145 187.94 1459.425 8613.565 ;
      RECT 1458.025 187.94 1458.305 8613.565 ;
      RECT 1451.025 187.94 1453.125 8613.565 ;
      RECT 1451.165 187.44 1453.125 8613.565 ;
      RECT 1449.905 187.94 1450.185 8613.565 ;
      RECT 1421.765 187.44 1446.685 8613.565 ;
      RECT 1416.025 187.94 1416.305 8613.565 ;
      RECT 1414.905 187.94 1415.185 8613.565 ;
      RECT 1412.665 187.94 1412.945 8613.565 ;
      RECT 1411.545 187.94 1411.825 8613.565 ;
      RECT 1410.425 187.94 1410.705 8613.565 ;
      RECT 1395.445 187.44 1407.765 8613.565 ;
      RECT 1390.265 187.94 1390.545 8613.565 ;
      RECT 1389.145 187.94 1389.425 8613.565 ;
      RECT 1388.025 187.94 1388.305 8613.565 ;
      RECT 1382.985 187.94 1383.265 8613.565 ;
      RECT 1343.365 187.94 1382.145 8613.565 ;
      RECT 1334.825 187.94 1335.105 8613.565 ;
      RECT 1333.705 187.94 1333.985 8613.565 ;
      RECT 1331.465 187.94 1331.745 8613.565 ;
      RECT 1330.345 187.94 1330.625 8613.565 ;
      RECT 1320.825 187.94 1329.365 8613.565 ;
      RECT 1320.965 187.44 1329.365 8613.565 ;
      RECT 1311.725 187.94 1313.825 8613.565 ;
      RECT 1310.465 187.94 1310.745 8613.565 ;
      RECT 1309.345 187.94 1309.625 8613.565 ;
      RECT 1282.325 187.44 1307.245 8613.565 ;
      RECT 1278.825 187.94 1279.105 8613.565 ;
      RECT 1277.705 187.94 1277.985 8613.565 ;
      RECT 1269.305 187.94 1269.585 8613.565 ;
      RECT 1255.305 187.94 1268.325 8613.565 ;
      RECT 1255.445 187.44 1268.325 8613.565 ;
      RECT 1253.065 187.94 1253.345 8613.565 ;
      RECT 1251.945 187.94 1252.225 8613.565 ;
      RECT 1250.825 187.94 1251.105 8613.565 ;
      RECT 1243.545 187.94 1243.825 8613.565 ;
      RECT 1203.365 187.94 1242.705 8613.565 ;
      RECT 1202.105 187.94 1202.385 8613.565 ;
      RECT 1197.065 187.94 1197.345 8613.565 ;
      RECT 1195.945 187.94 1196.225 8613.565 ;
      RECT 1181.525 187.44 1189.365 8613.565 ;
      RECT 1179.145 187.94 1179.425 8613.565 ;
      RECT 1178.025 187.94 1178.305 8613.565 ;
      RECT 1175.785 187.94 1176.065 8613.565 ;
      RECT 1174.665 187.94 1174.945 8613.565 ;
      RECT 1171.725 187.94 1173.825 8613.565 ;
      RECT 1142.325 187.44 1167.245 8613.565 ;
      RECT 1138.825 187.94 1139.105 8613.565 ;
      RECT 1137.705 187.94 1137.985 8613.565 ;
      RECT 1136.585 187.94 1136.865 8613.565 ;
      RECT 1131.545 187.94 1131.825 8613.565 ;
      RECT 1130.425 187.94 1130.705 8613.565 ;
      RECT 1116.005 187.44 1128.325 8613.565 ;
      RECT 1109.145 187.94 1109.425 8613.565 ;
      RECT 1108.025 187.94 1108.305 8613.565 ;
      RECT 1105.785 187.94 1106.065 8613.565 ;
      RECT 1104.665 187.94 1104.945 8613.565 ;
      RECT 1103.545 187.94 1103.825 8613.565 ;
      RECT 1062.805 187.44 1102.005 8613.565 ;
      RECT 1056.505 187.94 1056.785 8613.565 ;
      RECT 1055.385 187.94 1055.665 8613.565 ;
      RECT 1054.265 187.94 1054.545 8613.565 ;
      RECT 1040.825 187.94 1049.365 8613.565 ;
      RECT 1040.965 187.44 1049.365 8613.565 ;
      RECT 1039.705 187.94 1039.985 8613.565 ;
      RECT 1031.725 187.44 1033.125 8613.565 ;
      RECT 1029.345 187.94 1029.625 8613.565 ;
      RECT 1028.225 187.94 1028.505 8613.565 ;
      RECT 1001.205 187.44 1026.685 8613.565 ;
      RECT 999.945 187.94 1000.225 8613.565 ;
      RECT 998.825 187.94 999.105 8613.565 ;
      RECT 997.705 187.94 997.985 8613.565 ;
      RECT 990.425 187.94 990.705 8613.565 ;
      RECT 989.305 187.94 989.585 8613.565 ;
      RECT 974.745 187.94 988.325 8613.565 ;
      RECT 974.885 187.44 988.325 8613.565 ;
      RECT 969.705 187.94 969.985 8613.565 ;
      RECT 968.585 187.94 968.865 8613.565 ;
      RECT 923.925 187.44 962.005 8613.565 ;
      RECT 921.545 187.94 921.825 8613.565 ;
      RECT 920.425 187.94 920.705 8613.565 ;
      RECT 918.185 187.94 918.465 8613.565 ;
      RECT 917.065 187.94 917.345 8613.565 ;
      RECT 915.945 187.94 916.225 8613.565 ;
      RECT 901.525 187.44 909.365 8613.565 ;
      RECT 900.265 187.94 900.545 8613.565 ;
      RECT 899.145 187.94 899.425 8613.565 ;
      RECT 898.025 187.94 898.305 8613.565 ;
      RECT 891.025 187.94 893.125 8613.565 ;
      RECT 891.165 187.44 893.125 8613.565 ;
      RECT 889.905 187.94 890.185 8613.565 ;
      RECT 861.765 187.44 886.685 8613.565 ;
      RECT 856.025 187.94 856.305 8613.565 ;
      RECT 854.905 187.94 855.185 8613.565 ;
      RECT 852.665 187.94 852.945 8613.565 ;
      RECT 851.545 187.94 851.825 8613.565 ;
      RECT 850.425 187.94 850.705 8613.565 ;
      RECT 835.445 187.44 847.765 8613.565 ;
      RECT 830.265 187.94 830.545 8613.565 ;
      RECT 829.145 187.94 829.425 8613.565 ;
      RECT 828.025 187.94 828.305 8613.565 ;
      RECT 822.985 187.94 823.265 8613.565 ;
      RECT 783.365 187.94 822.145 8613.565 ;
      RECT 774.825 187.94 775.105 8613.565 ;
      RECT 773.705 187.94 773.985 8613.565 ;
      RECT 771.465 187.94 771.745 8613.565 ;
      RECT 770.345 187.94 770.625 8613.565 ;
      RECT 760.825 187.94 769.365 8613.565 ;
      RECT 760.965 187.44 769.365 8613.565 ;
      RECT 751.725 187.94 753.825 8613.565 ;
      RECT 750.465 187.94 750.745 8613.565 ;
      RECT 749.345 187.94 749.625 8613.565 ;
      RECT 722.325 187.44 747.245 8613.565 ;
      RECT 718.825 187.94 719.105 8613.565 ;
      RECT 717.705 187.94 717.985 8613.565 ;
      RECT 709.305 187.94 709.585 8613.565 ;
      RECT 695.305 187.94 708.325 8613.565 ;
      RECT 695.445 187.44 708.325 8613.565 ;
      RECT 693.065 187.94 693.345 8613.565 ;
      RECT 691.945 187.94 692.225 8613.565 ;
      RECT 690.825 187.94 691.105 8613.565 ;
      RECT 683.545 187.94 683.825 8613.565 ;
      RECT 643.365 187.94 682.705 8613.565 ;
      RECT 642.105 187.94 642.385 8613.565 ;
      RECT 637.065 187.94 637.345 8613.565 ;
      RECT 635.945 187.94 636.225 8613.565 ;
      RECT 621.525 187.44 629.365 8613.565 ;
      RECT 619.145 187.94 619.425 8613.565 ;
      RECT 618.025 187.94 618.305 8613.565 ;
      RECT 615.785 187.94 616.065 8613.565 ;
      RECT 614.665 187.94 614.945 8613.565 ;
      RECT 611.725 187.94 613.825 8613.565 ;
      RECT 582.325 187.44 607.245 8613.565 ;
      RECT 578.825 187.94 579.105 8613.565 ;
      RECT 577.705 187.94 577.985 8613.565 ;
      RECT 576.585 187.94 576.865 8613.565 ;
      RECT 571.545 187.94 571.825 8613.565 ;
      RECT 570.425 187.94 570.705 8613.565 ;
      RECT 556.005 187.44 568.325 8613.565 ;
      RECT 549.145 187.94 549.425 8613.565 ;
      RECT 548.025 187.94 548.305 8613.565 ;
      RECT 545.785 187.94 546.065 8613.565 ;
      RECT 544.665 187.94 544.945 8613.565 ;
      RECT 543.545 187.94 543.825 8613.565 ;
      RECT 502.805 187.44 542.005 8613.565 ;
      RECT 496.505 187.94 496.785 8613.565 ;
      RECT 495.385 187.94 495.665 8613.565 ;
      RECT 494.265 187.94 494.545 8613.565 ;
      RECT 480.825 187.94 489.365 8613.565 ;
      RECT 480.965 187.44 489.365 8613.565 ;
      RECT 479.705 187.94 479.985 8613.565 ;
      RECT 471.725 187.44 473.125 8613.565 ;
      RECT 469.345 187.94 469.625 8613.565 ;
      RECT 468.225 187.94 468.505 8613.565 ;
      RECT 6943.365 187.44 6982.005 8613.565 ;
      RECT 6911.725 187.44 6913.685 8613.565 ;
      RECT 6803.365 187.44 6842.565 8613.565 ;
      RECT 6771.725 187.44 6773.685 8613.565 ;
      RECT 6383.365 187.44 6422.005 8613.565 ;
      RECT 6351.725 187.44 6353.685 8613.565 ;
      RECT 6243.365 187.44 6282.565 8613.565 ;
      RECT 6211.725 187.44 6213.685 8613.565 ;
      RECT 5823.365 187.44 5862.005 8613.565 ;
      RECT 5791.725 187.44 5793.685 8613.565 ;
      RECT 5683.365 187.44 5722.565 8613.565 ;
      RECT 5651.725 187.44 5653.685 8613.565 ;
      RECT 5263.365 187.44 5302.005 8613.565 ;
      RECT 5231.725 187.44 5233.685 8613.565 ;
      RECT 5123.365 187.44 5162.565 8613.565 ;
      RECT 5091.725 187.44 5093.685 8613.565 ;
      RECT 4703.365 187.44 4742.005 8613.565 ;
      RECT 4671.725 187.44 4673.685 8613.565 ;
      RECT 4563.365 187.44 4602.565 8613.565 ;
      RECT 4531.725 187.44 4533.685 8613.565 ;
      RECT 4143.365 187.44 4182.005 8613.565 ;
      RECT 4111.725 187.44 4113.685 8613.565 ;
      RECT 4003.365 187.44 4042.565 8613.565 ;
      RECT 3971.725 187.44 3973.685 8613.565 ;
      RECT 3583.365 187.44 3622.005 8613.565 ;
      RECT 3551.725 187.44 3553.685 8613.565 ;
      RECT 3443.365 187.44 3482.565 8613.565 ;
      RECT 3411.725 187.44 3413.685 8613.565 ;
      RECT 3023.365 187.44 3062.005 8613.565 ;
      RECT 2991.725 187.44 2993.685 8613.565 ;
      RECT 2883.365 187.44 2922.565 8613.565 ;
      RECT 2851.725 187.44 2853.685 8613.565 ;
      RECT 2463.365 187.44 2502.005 8613.565 ;
      RECT 2431.725 187.44 2433.685 8613.565 ;
      RECT 2323.365 187.44 2362.565 8613.565 ;
      RECT 2291.725 187.44 2293.685 8613.565 ;
      RECT 1903.365 187.44 1942.005 8613.565 ;
      RECT 1871.725 187.44 1873.685 8613.565 ;
      RECT 1763.365 187.44 1802.565 8613.565 ;
      RECT 1731.725 187.44 1733.685 8613.565 ;
      RECT 1343.365 187.44 1382.005 8613.565 ;
      RECT 1311.725 187.44 1313.685 8613.565 ;
      RECT 1203.365 187.44 1242.565 8613.565 ;
      RECT 1171.725 187.44 1173.685 8613.565 ;
      RECT 783.365 187.44 822.005 8613.565 ;
      RECT 751.725 187.44 753.685 8613.565 ;
      RECT 643.365 187.44 682.565 8613.565 ;
      RECT 611.725 187.44 613.685 8613.565 ;
    LAYER M5 ;
      RECT 18362.06 307.445 18369.035 329.445 ;
      RECT 18369.035 268.27 18375.06 321.445 ;
      RECT 18362.06 189.04 18364.125 329.445 ;
      RECT 18362.06 268.27 18375.06 291.075 ;
      RECT 18362.06 228.445 18368.425 291.075 ;
      RECT 18362.06 228.445 18375.06 235.785 ;
      RECT 18371.12 189.04 18375.06 235.785 ;
      RECT 18369.035 194.415 18375.06 235.785 ;
      RECT 18362.06 194.415 18375.06 212.075 ;
      RECT 18362.06 189.04 18367.63 212.075 ;
      RECT 18362.06 189.04 18375.06 190.115 ;
      RECT 18345.08 307.445 18358.08 350.165 ;
      RECT 18346.705 189.04 18358.08 350.165 ;
      RECT 18345.08 228.445 18358.08 291.075 ;
      RECT 18345.08 189.04 18358.08 212.075 ;
      RECT 18314.56 324.445 18342.56 350.165 ;
      RECT 18320.705 189.04 18337.125 350.165 ;
      RECT 18314.56 211.445 18315.795 350.165 ;
      RECT 18314.56 211.445 18341.795 308.075 ;
      RECT 18314.56 228.445 18342.56 291.075 ;
      RECT 18316.925 189.04 18337.125 308.075 ;
      RECT 18314.56 189.04 18342.56 195.075 ;
      RECT 18299.04 228.445 18312.04 350.165 ;
      RECT 18299.04 189.04 18305.395 350.165 ;
      RECT 18299.04 189.04 18312.04 212.075 ;
      RECT 18282.06 290.445 18295.06 330.165 ;
      RECT 18293.19 189.04 18295.06 330.165 ;
      RECT 18291.425 194.425 18295.06 330.165 ;
      RECT 18282.06 189.04 18283.675 330.165 ;
      RECT 18282.06 194.425 18295.06 259.875 ;
      RECT 18282.06 189.04 18290.41 259.875 ;
      RECT 18282.06 189.04 18295.06 190.125 ;
      RECT 18265.08 211.445 18278.08 350.165 ;
      RECT 18265.425 189.04 18278.08 350.165 ;
      RECT 18265.08 189.04 18278.08 195.075 ;
      RECT 18234.56 259.445 18262.56 350.165 ;
      RECT 18246.935 211.445 18262.56 350.165 ;
      RECT 18234.56 189.04 18239.185 350.165 ;
      RECT 18234.56 189.04 18260.515 228.875 ;
      RECT 18234.56 189.04 18262.56 195.075 ;
      RECT 18219.04 307.445 18232.04 350.165 ;
      RECT 18229.035 194.37 18232.04 350.165 ;
      RECT 18219.04 189.04 18224.125 350.165 ;
      RECT 18219.04 228.445 18232.04 291.075 ;
      RECT 18219.04 194.37 18232.04 212.075 ;
      RECT 18219.04 189.04 18227.37 212.075 ;
      RECT 18219.04 189.04 18232.04 190.17 ;
      RECT 18202.06 307.445 18215.06 330.165 ;
      RECT 18206.705 189.04 18215.06 330.165 ;
      RECT 18206.54 228.445 18215.06 330.165 ;
      RECT 18202.06 228.445 18215.06 291.075 ;
      RECT 18202.06 189.04 18215.06 212.075 ;
      RECT 18185.08 324.445 18198.08 350.165 ;
      RECT 18185.08 189.04 18197.125 350.165 ;
      RECT 18185.08 211.445 18198.08 308.075 ;
      RECT 18185.08 189.04 18198.08 195.075 ;
      RECT 18154.56 324.445 18182.56 350.165 ;
      RECT 18180.705 189.04 18182.56 350.165 ;
      RECT 18154.56 228.445 18175.795 350.165 ;
      RECT 18178.115 189.04 18182.56 308.075 ;
      RECT 18161.11 211.445 18182.56 308.075 ;
      RECT 18154.56 189.04 18173.205 212.075 ;
      RECT 18154.56 189.04 18182.56 195.075 ;
      RECT 18139.04 290.445 18152.04 350.165 ;
      RECT 18151.425 194.42 18152.04 350.165 ;
      RECT 18139.04 189.04 18143.675 350.165 ;
      RECT 18139.04 194.42 18152.04 259.875 ;
      RECT 18139.04 189.04 18150.41 259.875 ;
      RECT 18139.04 189.04 18152.04 190.125 ;
      RECT 18122.06 211.445 18135.06 330.165 ;
      RECT 18125.425 189.04 18135.06 330.165 ;
      RECT 18122.06 189.04 18135.06 195.075 ;
      RECT 18105.08 259.445 18118.08 350.165 ;
      RECT 18106.935 189.04 18118.08 350.165 ;
      RECT 18105.08 189.04 18118.08 228.875 ;
      RECT 18074.56 307.445 18102.56 350.165 ;
      RECT 18089.035 259.445 18102.56 350.165 ;
      RECT 18074.56 189.04 18084.125 350.165 ;
      RECT 18074.56 228.445 18099.185 291.075 ;
      RECT 18093.09 189.04 18102.56 228.875 ;
      RECT 18089.035 194.37 18102.56 228.875 ;
      RECT 18074.56 194.37 18102.56 212.075 ;
      RECT 18074.56 189.04 18087.37 212.075 ;
      RECT 18074.56 189.04 18102.56 190.17 ;
      RECT 18059.04 324.445 18072.04 350.165 ;
      RECT 18066.705 189.04 18072.04 350.165 ;
      RECT 18062.035 307.445 18072.04 350.165 ;
      RECT 18059.04 307.445 18072.04 308.075 ;
      RECT 18059.04 211.445 18061.795 308.075 ;
      RECT 18059.04 228.445 18072.04 291.075 ;
      RECT 18059.04 211.445 18072.04 212.075 ;
      RECT 18062.035 189.04 18072.04 212.075 ;
      RECT 18059.04 189.04 18072.04 195.075 ;
      RECT 18025.08 324.445 18038.08 350.165 ;
      RECT 18025.08 228.445 18035.795 350.165 ;
      RECT 18030.31 211.445 18038.08 308.075 ;
      RECT 18025.08 189.04 18033.125 212.075 ;
      RECT 18025.08 189.04 18038.08 195.075 ;
      RECT 17994.56 290.445 18022.56 350.165 ;
      RECT 18013.19 189.04 18022.56 350.165 ;
      RECT 18011.425 194.425 18022.56 350.165 ;
      RECT 17994.56 189.04 18003.675 350.165 ;
      RECT 17994.56 194.425 18022.56 259.875 ;
      RECT 17994.56 189.04 18010.41 259.875 ;
      RECT 17994.56 189.04 18022.56 190.125 ;
      RECT 17979.04 211.445 17992.04 350.165 ;
      RECT 17985.425 189.04 17992.04 350.165 ;
      RECT 17979.04 189.04 17980.515 350.165 ;
      RECT 17979.04 189.04 17992.04 195.075 ;
      RECT 17962.06 259.445 17975.06 330.165 ;
      RECT 17966.935 189.04 17975.06 330.165 ;
      RECT 17962.06 189.04 17975.06 228.875 ;
      RECT 17945.08 307.445 17958.08 350.165 ;
      RECT 17953.09 189.04 17958.08 350.165 ;
      RECT 17949.035 194.37 17958.08 350.165 ;
      RECT 17945.08 228.445 17958.08 291.075 ;
      RECT 17945.08 194.37 17958.08 212.075 ;
      RECT 17945.08 189.04 17947.37 212.075 ;
      RECT 17945.08 189.04 17958.08 190.38 ;
      RECT 17914.56 324.445 17942.56 350.165 ;
      RECT 17926.705 189.04 17942.56 350.165 ;
      RECT 17922.035 307.445 17942.56 350.165 ;
      RECT 17914.56 189.04 17917.125 350.165 ;
      RECT 17914.56 307.445 17942.56 308.075 ;
      RECT 17914.56 211.445 17921.795 308.075 ;
      RECT 17914.56 228.445 17942.56 291.075 ;
      RECT 17914.56 211.445 17942.56 212.075 ;
      RECT 17922.035 189.04 17942.56 212.075 ;
      RECT 17914.56 189.04 17942.56 195.075 ;
      RECT 17899.04 324.445 17912.04 350.165 ;
      RECT 17900.705 189.04 17912.04 350.165 ;
      RECT 17899.04 189.04 17912.04 308.075 ;
      RECT 17882.06 228.445 17895.06 330.165 ;
      RECT 17888.69 211.445 17895.06 330.165 ;
      RECT 17882.06 189.04 17892.015 212.075 ;
      RECT 17882.06 189.04 17895.06 195.075 ;
      RECT 17865.08 290.445 17878.08 350.165 ;
      RECT 17873.19 189.04 17878.08 350.165 ;
      RECT 17871.425 194.425 17878.08 350.165 ;
      RECT 17865.08 194.425 17878.08 259.875 ;
      RECT 17865.08 189.04 17870.41 259.875 ;
      RECT 17865.08 189.04 17878.08 190.125 ;
      RECT 17834.56 211.445 17862.56 350.165 ;
      RECT 17845.425 189.04 17862.56 350.165 ;
      RECT 17834.56 189.04 17840.515 350.165 ;
      RECT 17834.56 189.04 17862.56 195.075 ;
      RECT 17819.04 259.445 17832.04 350.165 ;
      RECT 17826.935 189.04 17832.04 350.165 ;
      RECT 17819.04 189.04 17832.04 228.875 ;
      RECT 17802.06 307.445 17815.06 330.165 ;
      RECT 17812.99 189.04 17815.06 330.165 ;
      RECT 17809.035 194.37 17815.06 330.165 ;
      RECT 17802.06 189.04 17804.125 330.165 ;
      RECT 17802.06 228.445 17815.06 291.075 ;
      RECT 17802.06 194.37 17815.06 212.075 ;
      RECT 17802.06 189.04 17807.37 212.075 ;
      RECT 17802.06 189.04 17815.06 190.17 ;
      RECT 17785.08 307.445 17798.08 350.165 ;
      RECT 17786.705 189.04 17798.08 350.165 ;
      RECT 17785.08 228.445 17798.08 291.075 ;
      RECT 17785.08 189.04 17798.08 212.075 ;
      RECT 17754.56 324.445 17782.56 350.165 ;
      RECT 17760.705 189.04 17777.125 350.165 ;
      RECT 17754.56 211.445 17755.795 350.165 ;
      RECT 17754.56 211.445 17781.795 308.075 ;
      RECT 17754.56 228.445 17782.56 291.075 ;
      RECT 17756.925 189.04 17777.125 308.075 ;
      RECT 17754.56 189.04 17782.56 195.075 ;
      RECT 17739.04 228.445 17752.04 350.165 ;
      RECT 17739.04 189.04 17745.395 350.165 ;
      RECT 17739.04 189.04 17752.04 212.075 ;
      RECT 17722.06 290.445 17735.06 330.165 ;
      RECT 17733.19 189.04 17735.06 330.165 ;
      RECT 17731.425 194.425 17735.06 330.165 ;
      RECT 17722.06 189.04 17723.675 330.165 ;
      RECT 17722.06 194.425 17735.06 259.875 ;
      RECT 17722.06 189.04 17730.41 259.875 ;
      RECT 17722.06 189.04 17735.06 190.125 ;
      RECT 17705.08 211.445 17718.08 350.165 ;
      RECT 17705.425 189.04 17718.08 350.165 ;
      RECT 17705.08 189.04 17718.08 195.075 ;
      RECT 17674.56 259.445 17702.56 350.165 ;
      RECT 17686.935 211.445 17702.56 350.165 ;
      RECT 17674.56 189.04 17679.185 350.165 ;
      RECT 17674.56 189.04 17700.515 228.875 ;
      RECT 17674.56 189.04 17702.56 195.075 ;
      RECT 17659.04 307.445 17672.04 350.165 ;
      RECT 17669.035 194.37 17672.04 350.165 ;
      RECT 17659.04 189.04 17664.125 350.165 ;
      RECT 17659.04 228.445 17672.04 291.075 ;
      RECT 17659.04 194.37 17672.04 212.075 ;
      RECT 17659.04 189.04 17667.37 212.075 ;
      RECT 17659.04 189.04 17672.04 190.17 ;
      RECT 17642.06 307.445 17655.06 330.165 ;
      RECT 17646.705 189.04 17655.06 330.165 ;
      RECT 17646.54 228.445 17655.06 330.165 ;
      RECT 17642.06 228.445 17655.06 291.075 ;
      RECT 17642.06 189.04 17655.06 212.075 ;
      RECT 17625.08 324.445 17638.08 350.165 ;
      RECT 17625.08 189.04 17637.125 350.165 ;
      RECT 17625.08 211.445 17638.08 308.075 ;
      RECT 17625.08 189.04 17638.08 195.075 ;
      RECT 17594.56 324.445 17622.56 350.165 ;
      RECT 17620.705 189.04 17622.56 350.165 ;
      RECT 17594.56 228.445 17615.795 350.165 ;
      RECT 17618.115 189.04 17622.56 308.075 ;
      RECT 17601.11 211.445 17622.56 308.075 ;
      RECT 17594.56 189.04 17613.205 212.075 ;
      RECT 17594.56 189.04 17622.56 195.075 ;
      RECT 17579.04 290.445 17592.04 350.165 ;
      RECT 17591.425 194.42 17592.04 350.165 ;
      RECT 17579.04 189.04 17583.675 350.165 ;
      RECT 17579.04 194.42 17592.04 259.875 ;
      RECT 17579.04 189.04 17590.41 259.875 ;
      RECT 17579.04 189.04 17592.04 190.125 ;
      RECT 17562.06 211.445 17575.06 330.165 ;
      RECT 17565.425 189.04 17575.06 330.165 ;
      RECT 17562.06 189.04 17575.06 195.075 ;
      RECT 17545.08 259.445 17558.08 350.165 ;
      RECT 17546.935 189.04 17558.08 350.165 ;
      RECT 17545.08 189.04 17558.08 228.875 ;
      RECT 17514.56 307.445 17542.56 350.165 ;
      RECT 17529.035 259.445 17542.56 350.165 ;
      RECT 17514.56 189.04 17524.125 350.165 ;
      RECT 17514.56 228.445 17539.185 291.075 ;
      RECT 17533.09 189.04 17542.56 228.875 ;
      RECT 17529.035 194.37 17542.56 228.875 ;
      RECT 17514.56 194.37 17542.56 212.075 ;
      RECT 17514.56 189.04 17527.37 212.075 ;
      RECT 17514.56 189.04 17542.56 190.17 ;
      RECT 17499.04 324.445 17512.04 350.165 ;
      RECT 17506.705 189.04 17512.04 350.165 ;
      RECT 17502.035 307.445 17512.04 350.165 ;
      RECT 17499.04 307.445 17512.04 308.075 ;
      RECT 17499.04 211.445 17501.795 308.075 ;
      RECT 17499.04 228.445 17512.04 291.075 ;
      RECT 17499.04 211.445 17512.04 212.075 ;
      RECT 17502.035 189.04 17512.04 212.075 ;
      RECT 17499.04 189.04 17512.04 195.075 ;
      RECT 17465.08 324.445 17478.08 350.165 ;
      RECT 17465.08 228.445 17475.795 350.165 ;
      RECT 17470.31 211.445 17478.08 308.075 ;
      RECT 17465.08 189.04 17473.125 212.075 ;
      RECT 17465.08 189.04 17478.08 195.075 ;
      RECT 17434.56 290.445 17462.56 350.165 ;
      RECT 17453.19 189.04 17462.56 350.165 ;
      RECT 17451.425 194.425 17462.56 350.165 ;
      RECT 17434.56 189.04 17443.675 350.165 ;
      RECT 17434.56 194.425 17462.56 259.875 ;
      RECT 17434.56 189.04 17450.41 259.875 ;
      RECT 17434.56 189.04 17462.56 190.125 ;
      RECT 17419.04 211.445 17432.04 350.165 ;
      RECT 17425.425 189.04 17432.04 350.165 ;
      RECT 17419.04 189.04 17420.515 350.165 ;
      RECT 17419.04 189.04 17432.04 195.075 ;
      RECT 17402.06 259.445 17415.06 330.165 ;
      RECT 17406.935 189.04 17415.06 330.165 ;
      RECT 17402.06 189.04 17415.06 228.875 ;
      RECT 17385.08 307.445 17398.08 350.165 ;
      RECT 17393.09 189.04 17398.08 350.165 ;
      RECT 17389.035 194.37 17398.08 350.165 ;
      RECT 17385.08 228.445 17398.08 291.075 ;
      RECT 17385.08 194.37 17398.08 212.075 ;
      RECT 17385.08 189.04 17387.37 212.075 ;
      RECT 17385.08 189.04 17398.08 190.38 ;
      RECT 17354.56 324.445 17382.56 350.165 ;
      RECT 17366.705 189.04 17382.56 350.165 ;
      RECT 17362.035 307.445 17382.56 350.165 ;
      RECT 17354.56 189.04 17357.125 350.165 ;
      RECT 17354.56 307.445 17382.56 308.075 ;
      RECT 17354.56 211.445 17361.795 308.075 ;
      RECT 17354.56 228.445 17382.56 291.075 ;
      RECT 17354.56 211.445 17382.56 212.075 ;
      RECT 17362.035 189.04 17382.56 212.075 ;
      RECT 17354.56 189.04 17382.56 195.075 ;
      RECT 17339.04 324.445 17352.04 350.165 ;
      RECT 17340.705 189.04 17352.04 350.165 ;
      RECT 17339.04 189.04 17352.04 308.075 ;
      RECT 17322.06 228.445 17335.06 330.165 ;
      RECT 17328.69 211.445 17335.06 330.165 ;
      RECT 17322.06 189.04 17332.015 212.075 ;
      RECT 17322.06 189.04 17335.06 195.075 ;
      RECT 17305.08 290.445 17318.08 350.165 ;
      RECT 17313.19 189.04 17318.08 350.165 ;
      RECT 17311.425 194.425 17318.08 350.165 ;
      RECT 17305.08 194.425 17318.08 259.875 ;
      RECT 17305.08 189.04 17310.41 259.875 ;
      RECT 17305.08 189.04 17318.08 190.125 ;
      RECT 17274.56 211.445 17302.56 350.165 ;
      RECT 17285.425 189.04 17302.56 350.165 ;
      RECT 17274.56 189.04 17280.515 350.165 ;
      RECT 17274.56 189.04 17302.56 195.075 ;
      RECT 17259.04 259.445 17272.04 350.165 ;
      RECT 17266.935 189.04 17272.04 350.165 ;
      RECT 17259.04 189.04 17272.04 228.875 ;
      RECT 17242.06 307.445 17255.06 330.165 ;
      RECT 17252.99 189.04 17255.06 330.165 ;
      RECT 17249.035 194.37 17255.06 330.165 ;
      RECT 17242.06 189.04 17244.125 330.165 ;
      RECT 17242.06 228.445 17255.06 291.075 ;
      RECT 17242.06 194.37 17255.06 212.075 ;
      RECT 17242.06 189.04 17247.37 212.075 ;
      RECT 17242.06 189.04 17255.06 190.17 ;
      RECT 17225.08 307.445 17238.08 350.165 ;
      RECT 17226.705 189.04 17238.08 350.165 ;
      RECT 17225.08 228.445 17238.08 291.075 ;
      RECT 17225.08 189.04 17238.08 212.075 ;
      RECT 17194.56 324.445 17222.56 350.165 ;
      RECT 17200.705 189.04 17217.125 350.165 ;
      RECT 17194.56 211.445 17195.795 350.165 ;
      RECT 17194.56 211.445 17221.795 308.075 ;
      RECT 17194.56 228.445 17222.56 291.075 ;
      RECT 17196.925 189.04 17217.125 308.075 ;
      RECT 17194.56 189.04 17222.56 195.075 ;
      RECT 17179.04 228.445 17192.04 350.165 ;
      RECT 17179.04 189.04 17185.395 350.165 ;
      RECT 17179.04 189.04 17192.04 212.075 ;
      RECT 17162.06 290.445 17175.06 330.165 ;
      RECT 17173.19 189.04 17175.06 330.165 ;
      RECT 17171.425 194.425 17175.06 330.165 ;
      RECT 17162.06 189.04 17163.675 330.165 ;
      RECT 17162.06 194.425 17175.06 259.875 ;
      RECT 17162.06 189.04 17170.41 259.875 ;
      RECT 17162.06 189.04 17175.06 190.125 ;
      RECT 17145.08 211.445 17158.08 350.165 ;
      RECT 17145.425 189.04 17158.08 350.165 ;
      RECT 17145.08 189.04 17158.08 195.075 ;
      RECT 17114.56 259.445 17142.56 350.165 ;
      RECT 17126.935 211.445 17142.56 350.165 ;
      RECT 17114.56 189.04 17119.185 350.165 ;
      RECT 17114.56 189.04 17140.515 228.875 ;
      RECT 17114.56 189.04 17142.56 195.075 ;
      RECT 17099.04 307.445 17112.04 350.165 ;
      RECT 17109.035 194.37 17112.04 350.165 ;
      RECT 17099.04 189.04 17104.125 350.165 ;
      RECT 17099.04 228.445 17112.04 291.075 ;
      RECT 17099.04 194.37 17112.04 212.075 ;
      RECT 17099.04 189.04 17107.37 212.075 ;
      RECT 17099.04 189.04 17112.04 190.17 ;
      RECT 17082.06 307.445 17095.06 330.165 ;
      RECT 17086.705 189.04 17095.06 330.165 ;
      RECT 17086.54 228.445 17095.06 330.165 ;
      RECT 17082.06 228.445 17095.06 291.075 ;
      RECT 17082.06 189.04 17095.06 212.075 ;
      RECT 17065.08 324.445 17078.08 350.165 ;
      RECT 17065.08 189.04 17077.125 350.165 ;
      RECT 17065.08 211.445 17078.08 308.075 ;
      RECT 17065.08 189.04 17078.08 195.075 ;
      RECT 17034.56 324.445 17062.56 350.165 ;
      RECT 17060.705 189.04 17062.56 350.165 ;
      RECT 17034.56 228.445 17055.795 350.165 ;
      RECT 17058.115 189.04 17062.56 308.075 ;
      RECT 17041.11 211.445 17062.56 308.075 ;
      RECT 17034.56 189.04 17053.205 212.075 ;
      RECT 17034.56 189.04 17062.56 195.075 ;
      RECT 17019.04 290.445 17032.04 350.165 ;
      RECT 17031.425 194.42 17032.04 350.165 ;
      RECT 17019.04 189.04 17023.675 350.165 ;
      RECT 17019.04 194.42 17032.04 259.875 ;
      RECT 17019.04 189.04 17030.41 259.875 ;
      RECT 17019.04 189.04 17032.04 190.125 ;
      RECT 17002.06 211.445 17015.06 330.165 ;
      RECT 17005.425 189.04 17015.06 330.165 ;
      RECT 17002.06 189.04 17015.06 195.075 ;
      RECT 16985.08 259.445 16998.08 350.165 ;
      RECT 16986.935 189.04 16998.08 350.165 ;
      RECT 16985.08 189.04 16998.08 228.875 ;
      RECT 16954.56 307.445 16982.56 350.165 ;
      RECT 16969.035 259.445 16982.56 350.165 ;
      RECT 16954.56 189.04 16964.125 350.165 ;
      RECT 16954.56 228.445 16979.185 291.075 ;
      RECT 16973.09 189.04 16982.56 228.875 ;
      RECT 16969.035 194.37 16982.56 228.875 ;
      RECT 16954.56 194.37 16982.56 212.075 ;
      RECT 16954.56 189.04 16967.37 212.075 ;
      RECT 16954.56 189.04 16982.56 190.17 ;
      RECT 16939.04 324.445 16952.04 350.165 ;
      RECT 16946.705 189.04 16952.04 350.165 ;
      RECT 16942.035 307.445 16952.04 350.165 ;
      RECT 16939.04 307.445 16952.04 308.075 ;
      RECT 16939.04 211.445 16941.795 308.075 ;
      RECT 16939.04 228.445 16952.04 291.075 ;
      RECT 16939.04 211.445 16952.04 212.075 ;
      RECT 16942.035 189.04 16952.04 212.075 ;
      RECT 16939.04 189.04 16952.04 195.075 ;
      RECT 16905.08 324.445 16918.08 350.165 ;
      RECT 16905.08 228.445 16915.795 350.165 ;
      RECT 16910.31 211.445 16918.08 308.075 ;
      RECT 16905.08 189.04 16913.125 212.075 ;
      RECT 16905.08 189.04 16918.08 195.075 ;
      RECT 16874.56 290.445 16902.56 350.165 ;
      RECT 16893.19 189.04 16902.56 350.165 ;
      RECT 16891.425 194.425 16902.56 350.165 ;
      RECT 16874.56 189.04 16883.675 350.165 ;
      RECT 16874.56 194.425 16902.56 259.875 ;
      RECT 16874.56 189.04 16890.41 259.875 ;
      RECT 16874.56 189.04 16902.56 190.125 ;
      RECT 16859.04 211.445 16872.04 350.165 ;
      RECT 16865.425 189.04 16872.04 350.165 ;
      RECT 16859.04 189.04 16860.515 350.165 ;
      RECT 16859.04 189.04 16872.04 195.075 ;
      RECT 16842.06 259.445 16855.06 330.165 ;
      RECT 16846.935 189.04 16855.06 330.165 ;
      RECT 16842.06 189.04 16855.06 228.875 ;
      RECT 16825.08 307.445 16838.08 350.165 ;
      RECT 16833.09 189.04 16838.08 350.165 ;
      RECT 16829.035 194.37 16838.08 350.165 ;
      RECT 16825.08 228.445 16838.08 291.075 ;
      RECT 16825.08 194.37 16838.08 212.075 ;
      RECT 16825.08 189.04 16827.37 212.075 ;
      RECT 16825.08 189.04 16838.08 190.38 ;
      RECT 16794.56 324.445 16822.56 350.165 ;
      RECT 16806.705 189.04 16822.56 350.165 ;
      RECT 16802.035 307.445 16822.56 350.165 ;
      RECT 16794.56 189.04 16797.125 350.165 ;
      RECT 16794.56 307.445 16822.56 308.075 ;
      RECT 16794.56 211.445 16801.795 308.075 ;
      RECT 16794.56 228.445 16822.56 291.075 ;
      RECT 16794.56 211.445 16822.56 212.075 ;
      RECT 16802.035 189.04 16822.56 212.075 ;
      RECT 16794.56 189.04 16822.56 195.075 ;
      RECT 16779.04 324.445 16792.04 350.165 ;
      RECT 16780.705 189.04 16792.04 350.165 ;
      RECT 16779.04 189.04 16792.04 308.075 ;
      RECT 16762.06 228.445 16775.06 330.165 ;
      RECT 16768.69 211.445 16775.06 330.165 ;
      RECT 16762.06 189.04 16772.015 212.075 ;
      RECT 16762.06 189.04 16775.06 195.075 ;
      RECT 16745.08 290.445 16758.08 350.165 ;
      RECT 16753.19 189.04 16758.08 350.165 ;
      RECT 16751.425 194.425 16758.08 350.165 ;
      RECT 16745.08 194.425 16758.08 259.875 ;
      RECT 16745.08 189.04 16750.41 259.875 ;
      RECT 16745.08 189.04 16758.08 190.125 ;
      RECT 16714.56 211.445 16742.56 350.165 ;
      RECT 16725.425 189.04 16742.56 350.165 ;
      RECT 16714.56 189.04 16720.515 350.165 ;
      RECT 16714.56 189.04 16742.56 195.075 ;
      RECT 16699.04 259.445 16712.04 350.165 ;
      RECT 16706.935 189.04 16712.04 350.165 ;
      RECT 16699.04 189.04 16712.04 228.875 ;
      RECT 16682.06 307.445 16695.06 330.165 ;
      RECT 16692.99 189.04 16695.06 330.165 ;
      RECT 16689.035 194.37 16695.06 330.165 ;
      RECT 16682.06 189.04 16684.125 330.165 ;
      RECT 16682.06 228.445 16695.06 291.075 ;
      RECT 16682.06 194.37 16695.06 212.075 ;
      RECT 16682.06 189.04 16687.37 212.075 ;
      RECT 16682.06 189.04 16695.06 190.17 ;
      RECT 16665.08 307.445 16678.08 350.165 ;
      RECT 16666.705 189.04 16678.08 350.165 ;
      RECT 16665.08 228.445 16678.08 291.075 ;
      RECT 16665.08 189.04 16678.08 212.075 ;
      RECT 16634.56 324.445 16662.56 350.165 ;
      RECT 16640.705 189.04 16657.125 350.165 ;
      RECT 16634.56 211.445 16635.795 350.165 ;
      RECT 16634.56 211.445 16661.795 308.075 ;
      RECT 16634.56 228.445 16662.56 291.075 ;
      RECT 16636.925 189.04 16657.125 308.075 ;
      RECT 16634.56 189.04 16662.56 195.075 ;
      RECT 16619.04 228.445 16632.04 350.165 ;
      RECT 16619.04 189.04 16625.395 350.165 ;
      RECT 16619.04 189.04 16632.04 212.075 ;
      RECT 16602.06 290.445 16615.06 330.165 ;
      RECT 16613.19 189.04 16615.06 330.165 ;
      RECT 16611.425 194.425 16615.06 330.165 ;
      RECT 16602.06 189.04 16603.675 330.165 ;
      RECT 16602.06 194.425 16615.06 259.875 ;
      RECT 16602.06 189.04 16610.41 259.875 ;
      RECT 16602.06 189.04 16615.06 190.125 ;
      RECT 16585.08 211.445 16598.08 350.165 ;
      RECT 16585.425 189.04 16598.08 350.165 ;
      RECT 16585.08 189.04 16598.08 195.075 ;
      RECT 16554.56 259.445 16582.56 350.165 ;
      RECT 16566.935 211.445 16582.56 350.165 ;
      RECT 16554.56 189.04 16559.185 350.165 ;
      RECT 16554.56 189.04 16580.515 228.875 ;
      RECT 16554.56 189.04 16582.56 195.075 ;
      RECT 16539.04 307.445 16552.04 350.165 ;
      RECT 16549.035 194.37 16552.04 350.165 ;
      RECT 16539.04 189.04 16544.125 350.165 ;
      RECT 16539.04 228.445 16552.04 291.075 ;
      RECT 16539.04 194.37 16552.04 212.075 ;
      RECT 16539.04 189.04 16547.37 212.075 ;
      RECT 16539.04 189.04 16552.04 190.17 ;
      RECT 16522.06 307.445 16535.06 330.165 ;
      RECT 16526.705 189.04 16535.06 330.165 ;
      RECT 16526.54 228.445 16535.06 330.165 ;
      RECT 16522.06 228.445 16535.06 291.075 ;
      RECT 16522.06 189.04 16535.06 212.075 ;
      RECT 16505.08 324.445 16518.08 350.165 ;
      RECT 16505.08 189.04 16517.125 350.165 ;
      RECT 16505.08 211.445 16518.08 308.075 ;
      RECT 16505.08 189.04 16518.08 195.075 ;
      RECT 16474.56 324.445 16502.56 350.165 ;
      RECT 16500.705 189.04 16502.56 350.165 ;
      RECT 16474.56 228.445 16495.795 350.165 ;
      RECT 16498.115 189.04 16502.56 308.075 ;
      RECT 16481.11 211.445 16502.56 308.075 ;
      RECT 16474.56 189.04 16493.205 212.075 ;
      RECT 16474.56 189.04 16502.56 195.075 ;
      RECT 16459.04 290.445 16472.04 350.165 ;
      RECT 16471.425 194.42 16472.04 350.165 ;
      RECT 16459.04 189.04 16463.675 350.165 ;
      RECT 16459.04 194.42 16472.04 259.875 ;
      RECT 16459.04 189.04 16470.41 259.875 ;
      RECT 16459.04 189.04 16472.04 190.125 ;
      RECT 16442.06 211.445 16455.06 330.165 ;
      RECT 16445.425 189.04 16455.06 330.165 ;
      RECT 16442.06 189.04 16455.06 195.075 ;
      RECT 16425.08 259.445 16438.08 350.165 ;
      RECT 16426.935 189.04 16438.08 350.165 ;
      RECT 16425.08 189.04 16438.08 228.875 ;
      RECT 16394.56 307.445 16422.56 350.165 ;
      RECT 16409.035 259.445 16422.56 350.165 ;
      RECT 16394.56 189.04 16404.125 350.165 ;
      RECT 16394.56 228.445 16419.185 291.075 ;
      RECT 16413.09 189.04 16422.56 228.875 ;
      RECT 16409.035 194.37 16422.56 228.875 ;
      RECT 16394.56 194.37 16422.56 212.075 ;
      RECT 16394.56 189.04 16407.37 212.075 ;
      RECT 16394.56 189.04 16422.56 190.17 ;
      RECT 16379.04 324.445 16392.04 350.165 ;
      RECT 16386.705 189.04 16392.04 350.165 ;
      RECT 16382.035 307.445 16392.04 350.165 ;
      RECT 16379.04 307.445 16392.04 308.075 ;
      RECT 16379.04 211.445 16381.795 308.075 ;
      RECT 16379.04 228.445 16392.04 291.075 ;
      RECT 16379.04 211.445 16392.04 212.075 ;
      RECT 16382.035 189.04 16392.04 212.075 ;
      RECT 16379.04 189.04 16392.04 195.075 ;
      RECT 16345.08 324.445 16358.08 350.165 ;
      RECT 16345.08 228.445 16355.795 350.165 ;
      RECT 16350.31 211.445 16358.08 308.075 ;
      RECT 16345.08 189.04 16353.125 212.075 ;
      RECT 16345.08 189.04 16358.08 195.075 ;
      RECT 16314.56 290.445 16342.56 350.165 ;
      RECT 16333.19 189.04 16342.56 350.165 ;
      RECT 16331.425 194.425 16342.56 350.165 ;
      RECT 16314.56 189.04 16323.675 350.165 ;
      RECT 16314.56 194.425 16342.56 259.875 ;
      RECT 16314.56 189.04 16330.41 259.875 ;
      RECT 16314.56 189.04 16342.56 190.125 ;
      RECT 16299.04 211.445 16312.04 350.165 ;
      RECT 16305.425 189.04 16312.04 350.165 ;
      RECT 16299.04 189.04 16300.515 350.165 ;
      RECT 16299.04 189.04 16312.04 195.075 ;
      RECT 16282.06 259.445 16295.06 330.165 ;
      RECT 16286.935 189.04 16295.06 330.165 ;
      RECT 16282.06 189.04 16295.06 228.875 ;
      RECT 16265.08 307.445 16278.08 350.165 ;
      RECT 16273.09 189.04 16278.08 350.165 ;
      RECT 16269.035 194.37 16278.08 350.165 ;
      RECT 16265.08 228.445 16278.08 291.075 ;
      RECT 16265.08 194.37 16278.08 212.075 ;
      RECT 16265.08 189.04 16267.37 212.075 ;
      RECT 16265.08 189.04 16278.08 190.38 ;
      RECT 16234.56 324.445 16262.56 350.165 ;
      RECT 16246.705 189.04 16262.56 350.165 ;
      RECT 16242.035 307.445 16262.56 350.165 ;
      RECT 16234.56 189.04 16237.125 350.165 ;
      RECT 16234.56 307.445 16262.56 308.075 ;
      RECT 16234.56 211.445 16241.795 308.075 ;
      RECT 16234.56 228.445 16262.56 291.075 ;
      RECT 16234.56 211.445 16262.56 212.075 ;
      RECT 16242.035 189.04 16262.56 212.075 ;
      RECT 16234.56 189.04 16262.56 195.075 ;
      RECT 16219.04 324.445 16232.04 350.165 ;
      RECT 16220.705 189.04 16232.04 350.165 ;
      RECT 16219.04 189.04 16232.04 308.075 ;
      RECT 16202.06 228.445 16215.06 330.165 ;
      RECT 16208.69 211.445 16215.06 330.165 ;
      RECT 16202.06 189.04 16212.015 212.075 ;
      RECT 16202.06 189.04 16215.06 195.075 ;
      RECT 16185.08 290.445 16198.08 350.165 ;
      RECT 16193.19 189.04 16198.08 350.165 ;
      RECT 16191.425 194.425 16198.08 350.165 ;
      RECT 16185.08 194.425 16198.08 259.875 ;
      RECT 16185.08 189.04 16190.41 259.875 ;
      RECT 16185.08 189.04 16198.08 190.125 ;
      RECT 16154.56 211.445 16182.56 350.165 ;
      RECT 16165.425 189.04 16182.56 350.165 ;
      RECT 16154.56 189.04 16160.515 350.165 ;
      RECT 16154.56 189.04 16182.56 195.075 ;
      RECT 16139.04 259.445 16152.04 350.165 ;
      RECT 16146.935 189.04 16152.04 350.165 ;
      RECT 16139.04 189.04 16152.04 228.875 ;
      RECT 16122.06 307.445 16135.06 330.165 ;
      RECT 16132.99 189.04 16135.06 330.165 ;
      RECT 16129.035 194.37 16135.06 330.165 ;
      RECT 16122.06 189.04 16124.125 330.165 ;
      RECT 16122.06 228.445 16135.06 291.075 ;
      RECT 16122.06 194.37 16135.06 212.075 ;
      RECT 16122.06 189.04 16127.37 212.075 ;
      RECT 16122.06 189.04 16135.06 190.17 ;
      RECT 16105.08 307.445 16118.08 350.165 ;
      RECT 16106.705 189.04 16118.08 350.165 ;
      RECT 16105.08 228.445 16118.08 291.075 ;
      RECT 16105.08 189.04 16118.08 212.075 ;
      RECT 16074.56 324.445 16102.56 350.165 ;
      RECT 16080.705 189.04 16097.125 350.165 ;
      RECT 16074.56 211.445 16075.795 350.165 ;
      RECT 16074.56 211.445 16101.795 308.075 ;
      RECT 16074.56 228.445 16102.56 291.075 ;
      RECT 16076.925 189.04 16097.125 308.075 ;
      RECT 16074.56 189.04 16102.56 195.075 ;
      RECT 16059.04 228.445 16072.04 350.165 ;
      RECT 16059.04 189.04 16065.395 350.165 ;
      RECT 16059.04 189.04 16072.04 212.075 ;
      RECT 16042.06 290.445 16055.06 330.165 ;
      RECT 16053.19 189.04 16055.06 330.165 ;
      RECT 16051.425 194.425 16055.06 330.165 ;
      RECT 16042.06 189.04 16043.675 330.165 ;
      RECT 16042.06 194.425 16055.06 259.875 ;
      RECT 16042.06 189.04 16050.41 259.875 ;
      RECT 16042.06 189.04 16055.06 190.125 ;
      RECT 16025.08 211.445 16038.08 350.165 ;
      RECT 16025.425 189.04 16038.08 350.165 ;
      RECT 16025.08 189.04 16038.08 195.075 ;
      RECT 15994.56 259.445 16022.56 350.165 ;
      RECT 16006.935 211.445 16022.56 350.165 ;
      RECT 15994.56 189.04 15999.185 350.165 ;
      RECT 15994.56 189.04 16020.515 228.875 ;
      RECT 15994.56 189.04 16022.56 195.075 ;
      RECT 15979.04 307.445 15992.04 350.165 ;
      RECT 15989.035 194.37 15992.04 350.165 ;
      RECT 15979.04 189.04 15984.125 350.165 ;
      RECT 15979.04 228.445 15992.04 291.075 ;
      RECT 15979.04 194.37 15992.04 212.075 ;
      RECT 15979.04 189.04 15987.37 212.075 ;
      RECT 15979.04 189.04 15992.04 190.17 ;
      RECT 15962.06 307.445 15975.06 330.165 ;
      RECT 15966.705 189.04 15975.06 330.165 ;
      RECT 15966.54 228.445 15975.06 330.165 ;
      RECT 15962.06 228.445 15975.06 291.075 ;
      RECT 15962.06 189.04 15975.06 212.075 ;
      RECT 15945.08 324.445 15958.08 350.165 ;
      RECT 15945.08 189.04 15957.125 350.165 ;
      RECT 15945.08 211.445 15958.08 308.075 ;
      RECT 15945.08 189.04 15958.08 195.075 ;
      RECT 15914.56 324.445 15942.56 350.165 ;
      RECT 15940.705 189.04 15942.56 350.165 ;
      RECT 15914.56 228.445 15935.795 350.165 ;
      RECT 15938.115 189.04 15942.56 308.075 ;
      RECT 15921.11 211.445 15942.56 308.075 ;
      RECT 15914.56 189.04 15933.205 212.075 ;
      RECT 15914.56 189.04 15942.56 195.075 ;
      RECT 15899.04 290.445 15912.04 350.165 ;
      RECT 15911.425 194.42 15912.04 350.165 ;
      RECT 15899.04 189.04 15903.675 350.165 ;
      RECT 15899.04 194.42 15912.04 259.875 ;
      RECT 15899.04 189.04 15910.41 259.875 ;
      RECT 15899.04 189.04 15912.04 190.125 ;
      RECT 15882.06 211.445 15895.06 330.165 ;
      RECT 15885.425 189.04 15895.06 330.165 ;
      RECT 15882.06 189.04 15895.06 195.075 ;
      RECT 15865.08 259.445 15878.08 350.165 ;
      RECT 15866.935 189.04 15878.08 350.165 ;
      RECT 15865.08 189.04 15878.08 228.875 ;
      RECT 15834.56 307.445 15862.56 350.165 ;
      RECT 15849.035 259.445 15862.56 350.165 ;
      RECT 15834.56 189.04 15844.125 350.165 ;
      RECT 15834.56 228.445 15859.185 291.075 ;
      RECT 15853.09 189.04 15862.56 228.875 ;
      RECT 15849.035 194.37 15862.56 228.875 ;
      RECT 15834.56 194.37 15862.56 212.075 ;
      RECT 15834.56 189.04 15847.37 212.075 ;
      RECT 15834.56 189.04 15862.56 190.17 ;
      RECT 15819.04 324.445 15832.04 350.165 ;
      RECT 15826.705 189.04 15832.04 350.165 ;
      RECT 15822.035 307.445 15832.04 350.165 ;
      RECT 15819.04 307.445 15832.04 308.075 ;
      RECT 15819.04 211.445 15821.795 308.075 ;
      RECT 15819.04 228.445 15832.04 291.075 ;
      RECT 15819.04 211.445 15832.04 212.075 ;
      RECT 15822.035 189.04 15832.04 212.075 ;
      RECT 15819.04 189.04 15832.04 195.075 ;
      RECT 15785.08 324.445 15798.08 350.165 ;
      RECT 15785.08 228.445 15795.795 350.165 ;
      RECT 15790.31 211.445 15798.08 308.075 ;
      RECT 15785.08 189.04 15793.125 212.075 ;
      RECT 15785.08 189.04 15798.08 195.075 ;
      RECT 15754.56 290.445 15782.56 350.165 ;
      RECT 15773.19 189.04 15782.56 350.165 ;
      RECT 15771.425 194.425 15782.56 350.165 ;
      RECT 15754.56 189.04 15763.675 350.165 ;
      RECT 15754.56 194.425 15782.56 259.875 ;
      RECT 15754.56 189.04 15770.41 259.875 ;
      RECT 15754.56 189.04 15782.56 190.125 ;
      RECT 15739.04 211.445 15752.04 350.165 ;
      RECT 15745.425 189.04 15752.04 350.165 ;
      RECT 15739.04 189.04 15740.515 350.165 ;
      RECT 15739.04 189.04 15752.04 195.075 ;
      RECT 15722.06 259.445 15735.06 330.165 ;
      RECT 15726.935 189.04 15735.06 330.165 ;
      RECT 15722.06 189.04 15735.06 228.875 ;
      RECT 15705.08 307.445 15718.08 350.165 ;
      RECT 15713.09 189.04 15718.08 350.165 ;
      RECT 15709.035 194.37 15718.08 350.165 ;
      RECT 15705.08 228.445 15718.08 291.075 ;
      RECT 15705.08 194.37 15718.08 212.075 ;
      RECT 15705.08 189.04 15707.37 212.075 ;
      RECT 15705.08 189.04 15718.08 190.38 ;
      RECT 15674.56 324.445 15702.56 350.165 ;
      RECT 15686.705 189.04 15702.56 350.165 ;
      RECT 15682.035 307.445 15702.56 350.165 ;
      RECT 15674.56 189.04 15677.125 350.165 ;
      RECT 15674.56 307.445 15702.56 308.075 ;
      RECT 15674.56 211.445 15681.795 308.075 ;
      RECT 15674.56 228.445 15702.56 291.075 ;
      RECT 15674.56 211.445 15702.56 212.075 ;
      RECT 15682.035 189.04 15702.56 212.075 ;
      RECT 15674.56 189.04 15702.56 195.075 ;
      RECT 15659.04 324.445 15672.04 350.165 ;
      RECT 15660.705 189.04 15672.04 350.165 ;
      RECT 15659.04 189.04 15672.04 308.075 ;
      RECT 15642.06 228.445 15655.06 330.165 ;
      RECT 15648.69 211.445 15655.06 330.165 ;
      RECT 15642.06 189.04 15652.015 212.075 ;
      RECT 15642.06 189.04 15655.06 195.075 ;
      RECT 15625.08 290.445 15638.08 350.165 ;
      RECT 15633.19 189.04 15638.08 350.165 ;
      RECT 15631.425 194.425 15638.08 350.165 ;
      RECT 15625.08 194.425 15638.08 259.875 ;
      RECT 15625.08 189.04 15630.41 259.875 ;
      RECT 15625.08 189.04 15638.08 190.125 ;
      RECT 15594.56 211.445 15622.56 350.165 ;
      RECT 15605.425 189.04 15622.56 350.165 ;
      RECT 15594.56 189.04 15600.515 350.165 ;
      RECT 15594.56 189.04 15622.56 195.075 ;
      RECT 15579.04 259.445 15592.04 350.165 ;
      RECT 15586.935 189.04 15592.04 350.165 ;
      RECT 15579.04 189.04 15592.04 228.875 ;
      RECT 15562.06 307.445 15575.06 330.165 ;
      RECT 15572.99 189.04 15575.06 330.165 ;
      RECT 15569.035 194.37 15575.06 330.165 ;
      RECT 15562.06 189.04 15564.125 330.165 ;
      RECT 15562.06 228.445 15575.06 291.075 ;
      RECT 15562.06 194.37 15575.06 212.075 ;
      RECT 15562.06 189.04 15567.37 212.075 ;
      RECT 15562.06 189.04 15575.06 190.17 ;
      RECT 15545.08 307.445 15558.08 350.165 ;
      RECT 15546.705 189.04 15558.08 350.165 ;
      RECT 15545.08 228.445 15558.08 291.075 ;
      RECT 15545.08 189.04 15558.08 212.075 ;
      RECT 15514.56 324.445 15542.56 350.165 ;
      RECT 15520.705 189.04 15537.125 350.165 ;
      RECT 15514.56 211.445 15515.795 350.165 ;
      RECT 15514.56 211.445 15541.795 308.075 ;
      RECT 15514.56 228.445 15542.56 291.075 ;
      RECT 15516.925 189.04 15537.125 308.075 ;
      RECT 15514.56 189.04 15542.56 195.075 ;
      RECT 15499.04 228.445 15512.04 350.165 ;
      RECT 15499.04 189.04 15505.395 350.165 ;
      RECT 15499.04 189.04 15512.04 212.075 ;
      RECT 15482.06 290.445 15495.06 330.165 ;
      RECT 15493.19 189.04 15495.06 330.165 ;
      RECT 15491.425 194.425 15495.06 330.165 ;
      RECT 15482.06 189.04 15483.675 330.165 ;
      RECT 15482.06 194.425 15495.06 259.875 ;
      RECT 15482.06 189.04 15490.41 259.875 ;
      RECT 15482.06 189.04 15495.06 190.125 ;
      RECT 15465.08 211.445 15478.08 350.165 ;
      RECT 15465.425 189.04 15478.08 350.165 ;
      RECT 15465.08 189.04 15478.08 195.075 ;
      RECT 15434.56 259.445 15462.56 350.165 ;
      RECT 15446.935 211.445 15462.56 350.165 ;
      RECT 15434.56 189.04 15439.185 350.165 ;
      RECT 15434.56 189.04 15460.515 228.875 ;
      RECT 15434.56 189.04 15462.56 195.075 ;
      RECT 15419.04 307.445 15432.04 350.165 ;
      RECT 15429.035 194.37 15432.04 350.165 ;
      RECT 15419.04 189.04 15424.125 350.165 ;
      RECT 15419.04 228.445 15432.04 291.075 ;
      RECT 15419.04 194.37 15432.04 212.075 ;
      RECT 15419.04 189.04 15427.37 212.075 ;
      RECT 15419.04 189.04 15432.04 190.17 ;
      RECT 15402.06 307.445 15415.06 330.165 ;
      RECT 15406.705 189.04 15415.06 330.165 ;
      RECT 15406.54 228.445 15415.06 330.165 ;
      RECT 15402.06 228.445 15415.06 291.075 ;
      RECT 15402.06 189.04 15415.06 212.075 ;
      RECT 15385.08 324.445 15398.08 350.165 ;
      RECT 15385.08 189.04 15397.125 350.165 ;
      RECT 15385.08 211.445 15398.08 308.075 ;
      RECT 15385.08 189.04 15398.08 195.075 ;
      RECT 15354.56 324.445 15382.56 350.165 ;
      RECT 15380.705 189.04 15382.56 350.165 ;
      RECT 15354.56 228.445 15375.795 350.165 ;
      RECT 15378.115 189.04 15382.56 308.075 ;
      RECT 15361.11 211.445 15382.56 308.075 ;
      RECT 15354.56 189.04 15373.205 212.075 ;
      RECT 15354.56 189.04 15382.56 195.075 ;
      RECT 15339.04 290.445 15352.04 350.165 ;
      RECT 15351.425 194.42 15352.04 350.165 ;
      RECT 15339.04 189.04 15343.675 350.165 ;
      RECT 15339.04 194.42 15352.04 259.875 ;
      RECT 15339.04 189.04 15350.41 259.875 ;
      RECT 15339.04 189.04 15352.04 190.125 ;
      RECT 15322.06 211.445 15335.06 330.165 ;
      RECT 15325.425 189.04 15335.06 330.165 ;
      RECT 15322.06 189.04 15335.06 195.075 ;
      RECT 15305.08 259.445 15318.08 350.165 ;
      RECT 15306.935 189.04 15318.08 350.165 ;
      RECT 15305.08 189.04 15318.08 228.875 ;
      RECT 15274.56 307.445 15302.56 350.165 ;
      RECT 15289.035 259.445 15302.56 350.165 ;
      RECT 15274.56 189.04 15284.125 350.165 ;
      RECT 15274.56 228.445 15299.185 291.075 ;
      RECT 15293.09 189.04 15302.56 228.875 ;
      RECT 15289.035 194.37 15302.56 228.875 ;
      RECT 15274.56 194.37 15302.56 212.075 ;
      RECT 15274.56 189.04 15287.37 212.075 ;
      RECT 15274.56 189.04 15302.56 190.17 ;
      RECT 15259.04 324.445 15272.04 350.165 ;
      RECT 15266.705 189.04 15272.04 350.165 ;
      RECT 15262.035 307.445 15272.04 350.165 ;
      RECT 15259.04 307.445 15272.04 308.075 ;
      RECT 15259.04 211.445 15261.795 308.075 ;
      RECT 15259.04 228.445 15272.04 291.075 ;
      RECT 15259.04 211.445 15272.04 212.075 ;
      RECT 15262.035 189.04 15272.04 212.075 ;
      RECT 15259.04 189.04 15272.04 195.075 ;
      RECT 15225.08 324.445 15238.08 350.165 ;
      RECT 15225.08 228.445 15235.795 350.165 ;
      RECT 15230.31 211.445 15238.08 308.075 ;
      RECT 15225.08 189.04 15233.125 212.075 ;
      RECT 15225.08 189.04 15238.08 195.075 ;
      RECT 15194.56 290.445 15222.56 350.165 ;
      RECT 15213.19 189.04 15222.56 350.165 ;
      RECT 15211.425 194.425 15222.56 350.165 ;
      RECT 15194.56 189.04 15203.675 350.165 ;
      RECT 15194.56 194.425 15222.56 259.875 ;
      RECT 15194.56 189.04 15210.41 259.875 ;
      RECT 15194.56 189.04 15222.56 190.125 ;
      RECT 15179.04 211.445 15192.04 350.165 ;
      RECT 15185.425 189.04 15192.04 350.165 ;
      RECT 15179.04 189.04 15180.515 350.165 ;
      RECT 15179.04 189.04 15192.04 195.075 ;
      RECT 15162.06 259.445 15175.06 330.165 ;
      RECT 15166.935 189.04 15175.06 330.165 ;
      RECT 15162.06 189.04 15175.06 228.875 ;
      RECT 15145.08 307.445 15158.08 350.165 ;
      RECT 15153.09 189.04 15158.08 350.165 ;
      RECT 15149.035 194.37 15158.08 350.165 ;
      RECT 15145.08 228.445 15158.08 291.075 ;
      RECT 15145.08 194.37 15158.08 212.075 ;
      RECT 15145.08 189.04 15147.37 212.075 ;
      RECT 15145.08 189.04 15158.08 190.38 ;
      RECT 15114.56 324.445 15142.56 350.165 ;
      RECT 15126.705 189.04 15142.56 350.165 ;
      RECT 15122.035 307.445 15142.56 350.165 ;
      RECT 15114.56 189.04 15117.125 350.165 ;
      RECT 15114.56 307.445 15142.56 308.075 ;
      RECT 15114.56 211.445 15121.795 308.075 ;
      RECT 15114.56 228.445 15142.56 291.075 ;
      RECT 15114.56 211.445 15142.56 212.075 ;
      RECT 15122.035 189.04 15142.56 212.075 ;
      RECT 15114.56 189.04 15142.56 195.075 ;
      RECT 15099.04 324.445 15112.04 350.165 ;
      RECT 15100.705 189.04 15112.04 350.165 ;
      RECT 15099.04 189.04 15112.04 308.075 ;
      RECT 15082.06 228.445 15095.06 330.165 ;
      RECT 15088.69 211.445 15095.06 330.165 ;
      RECT 15082.06 189.04 15092.015 212.075 ;
      RECT 15082.06 189.04 15095.06 195.075 ;
      RECT 15065.08 290.445 15078.08 350.165 ;
      RECT 15073.19 189.04 15078.08 350.165 ;
      RECT 15071.425 194.425 15078.08 350.165 ;
      RECT 15065.08 194.425 15078.08 259.875 ;
      RECT 15065.08 189.04 15070.41 259.875 ;
      RECT 15065.08 189.04 15078.08 190.125 ;
      RECT 15034.56 211.445 15062.56 350.165 ;
      RECT 15045.425 189.04 15062.56 350.165 ;
      RECT 15034.56 189.04 15040.515 350.165 ;
      RECT 15034.56 189.04 15062.56 195.075 ;
      RECT 15019.04 259.445 15032.04 350.165 ;
      RECT 15026.935 189.04 15032.04 350.165 ;
      RECT 15019.04 189.04 15032.04 228.875 ;
      RECT 15002.06 307.445 15015.06 330.165 ;
      RECT 15012.99 189.04 15015.06 330.165 ;
      RECT 15009.035 194.37 15015.06 330.165 ;
      RECT 15002.06 189.04 15004.125 330.165 ;
      RECT 15002.06 228.445 15015.06 291.075 ;
      RECT 15002.06 194.37 15015.06 212.075 ;
      RECT 15002.06 189.04 15007.37 212.075 ;
      RECT 15002.06 189.04 15015.06 190.17 ;
      RECT 14985.08 307.445 14998.08 350.165 ;
      RECT 14986.705 189.04 14998.08 350.165 ;
      RECT 14985.08 228.445 14998.08 291.075 ;
      RECT 14985.08 189.04 14998.08 212.075 ;
      RECT 14954.56 324.445 14982.56 350.165 ;
      RECT 14960.705 189.04 14977.125 350.165 ;
      RECT 14954.56 211.445 14955.795 350.165 ;
      RECT 14954.56 211.445 14981.795 308.075 ;
      RECT 14954.56 228.445 14982.56 291.075 ;
      RECT 14956.925 189.04 14977.125 308.075 ;
      RECT 14954.56 189.04 14982.56 195.075 ;
      RECT 14939.04 228.445 14952.04 350.165 ;
      RECT 14939.04 189.04 14945.395 350.165 ;
      RECT 14939.04 189.04 14952.04 212.075 ;
      RECT 14922.06 290.445 14935.06 330.165 ;
      RECT 14933.19 189.04 14935.06 330.165 ;
      RECT 14931.425 194.425 14935.06 330.165 ;
      RECT 14922.06 189.04 14923.675 330.165 ;
      RECT 14922.06 194.425 14935.06 259.875 ;
      RECT 14922.06 189.04 14930.41 259.875 ;
      RECT 14922.06 189.04 14935.06 190.125 ;
      RECT 14905.08 211.445 14918.08 350.165 ;
      RECT 14905.425 189.04 14918.08 350.165 ;
      RECT 14905.08 189.04 14918.08 195.075 ;
      RECT 14874.56 259.445 14902.56 350.165 ;
      RECT 14886.935 211.445 14902.56 350.165 ;
      RECT 14874.56 189.04 14879.185 350.165 ;
      RECT 14874.56 189.04 14900.515 228.875 ;
      RECT 14874.56 189.04 14902.56 195.075 ;
      RECT 14859.04 307.445 14872.04 350.165 ;
      RECT 14869.035 194.37 14872.04 350.165 ;
      RECT 14859.04 189.04 14864.125 350.165 ;
      RECT 14859.04 228.445 14872.04 291.075 ;
      RECT 14859.04 194.37 14872.04 212.075 ;
      RECT 14859.04 189.04 14867.37 212.075 ;
      RECT 14859.04 189.04 14872.04 190.17 ;
      RECT 14842.06 307.445 14855.06 330.165 ;
      RECT 14846.705 189.04 14855.06 330.165 ;
      RECT 14846.54 228.445 14855.06 330.165 ;
      RECT 14842.06 228.445 14855.06 291.075 ;
      RECT 14842.06 189.04 14855.06 212.075 ;
      RECT 14825.08 324.445 14838.08 350.165 ;
      RECT 14825.08 189.04 14837.125 350.165 ;
      RECT 14825.08 211.445 14838.08 308.075 ;
      RECT 14825.08 189.04 14838.08 195.075 ;
      RECT 14794.56 324.445 14822.56 350.165 ;
      RECT 14820.705 189.04 14822.56 350.165 ;
      RECT 14794.56 228.445 14815.795 350.165 ;
      RECT 14818.115 189.04 14822.56 308.075 ;
      RECT 14801.11 211.445 14822.56 308.075 ;
      RECT 14794.56 189.04 14813.205 212.075 ;
      RECT 14794.56 189.04 14822.56 195.075 ;
      RECT 14779.04 290.445 14792.04 350.165 ;
      RECT 14791.425 194.42 14792.04 350.165 ;
      RECT 14779.04 189.04 14783.675 350.165 ;
      RECT 14779.04 194.42 14792.04 259.875 ;
      RECT 14779.04 189.04 14790.41 259.875 ;
      RECT 14779.04 189.04 14792.04 190.125 ;
      RECT 14762.06 211.445 14775.06 330.165 ;
      RECT 14765.425 189.04 14775.06 330.165 ;
      RECT 14762.06 189.04 14775.06 195.075 ;
      RECT 14745.08 259.445 14758.08 350.165 ;
      RECT 14746.935 189.04 14758.08 350.165 ;
      RECT 14745.08 189.04 14758.08 228.875 ;
      RECT 14714.56 307.445 14742.56 350.165 ;
      RECT 14729.035 259.445 14742.56 350.165 ;
      RECT 14714.56 189.04 14724.125 350.165 ;
      RECT 14714.56 228.445 14739.185 291.075 ;
      RECT 14733.09 189.04 14742.56 228.875 ;
      RECT 14729.035 194.37 14742.56 228.875 ;
      RECT 14714.56 194.37 14742.56 212.075 ;
      RECT 14714.56 189.04 14727.37 212.075 ;
      RECT 14714.56 189.04 14742.56 190.17 ;
      RECT 14699.04 324.445 14712.04 350.165 ;
      RECT 14706.705 189.04 14712.04 350.165 ;
      RECT 14702.035 307.445 14712.04 350.165 ;
      RECT 14699.04 307.445 14712.04 308.075 ;
      RECT 14699.04 211.445 14701.795 308.075 ;
      RECT 14699.04 228.445 14712.04 291.075 ;
      RECT 14699.04 211.445 14712.04 212.075 ;
      RECT 14702.035 189.04 14712.04 212.075 ;
      RECT 14699.04 189.04 14712.04 195.075 ;
      RECT 14665.08 324.445 14678.08 350.165 ;
      RECT 14665.08 228.445 14675.795 350.165 ;
      RECT 14670.31 211.445 14678.08 308.075 ;
      RECT 14665.08 189.04 14673.125 212.075 ;
      RECT 14665.08 189.04 14678.08 195.075 ;
      RECT 14634.56 290.445 14662.56 350.165 ;
      RECT 14653.19 189.04 14662.56 350.165 ;
      RECT 14651.425 194.425 14662.56 350.165 ;
      RECT 14634.56 189.04 14643.675 350.165 ;
      RECT 14634.56 194.425 14662.56 259.875 ;
      RECT 14634.56 189.04 14650.41 259.875 ;
      RECT 14634.56 189.04 14662.56 190.125 ;
      RECT 14619.04 211.445 14632.04 350.165 ;
      RECT 14625.425 189.04 14632.04 350.165 ;
      RECT 14619.04 189.04 14620.515 350.165 ;
      RECT 14619.04 189.04 14632.04 195.075 ;
      RECT 14602.06 259.445 14615.06 330.165 ;
      RECT 14606.935 189.04 14615.06 330.165 ;
      RECT 14602.06 189.04 14615.06 228.875 ;
      RECT 14585.08 307.445 14598.08 350.165 ;
      RECT 14593.09 189.04 14598.08 350.165 ;
      RECT 14589.035 194.37 14598.08 350.165 ;
      RECT 14585.08 228.445 14598.08 291.075 ;
      RECT 14585.08 194.37 14598.08 212.075 ;
      RECT 14585.08 189.04 14587.37 212.075 ;
      RECT 14585.08 189.04 14598.08 190.38 ;
      RECT 14554.56 324.445 14582.56 350.165 ;
      RECT 14566.705 189.04 14582.56 350.165 ;
      RECT 14562.035 307.445 14582.56 350.165 ;
      RECT 14554.56 189.04 14557.125 350.165 ;
      RECT 14554.56 307.445 14582.56 308.075 ;
      RECT 14554.56 211.445 14561.795 308.075 ;
      RECT 14554.56 228.445 14582.56 291.075 ;
      RECT 14554.56 211.445 14582.56 212.075 ;
      RECT 14562.035 189.04 14582.56 212.075 ;
      RECT 14554.56 189.04 14582.56 195.075 ;
      RECT 14539.04 324.445 14552.04 350.165 ;
      RECT 14540.705 189.04 14552.04 350.165 ;
      RECT 14539.04 189.04 14552.04 308.075 ;
      RECT 14522.06 228.445 14535.06 330.165 ;
      RECT 14528.69 211.445 14535.06 330.165 ;
      RECT 14522.06 189.04 14532.015 212.075 ;
      RECT 14522.06 189.04 14535.06 195.075 ;
      RECT 14505.08 290.445 14518.08 350.165 ;
      RECT 14513.19 189.04 14518.08 350.165 ;
      RECT 14511.425 194.425 14518.08 350.165 ;
      RECT 14505.08 194.425 14518.08 259.875 ;
      RECT 14505.08 189.04 14510.41 259.875 ;
      RECT 14505.08 189.04 14518.08 190.125 ;
      RECT 14474.56 211.445 14502.56 350.165 ;
      RECT 14485.425 189.04 14502.56 350.165 ;
      RECT 14474.56 189.04 14480.515 350.165 ;
      RECT 14474.56 189.04 14502.56 195.075 ;
      RECT 14459.04 259.445 14472.04 350.165 ;
      RECT 14466.935 189.04 14472.04 350.165 ;
      RECT 14459.04 189.04 14472.04 228.875 ;
      RECT 14442.06 307.445 14455.06 330.165 ;
      RECT 14452.99 189.04 14455.06 330.165 ;
      RECT 14449.035 194.37 14455.06 330.165 ;
      RECT 14442.06 189.04 14444.125 330.165 ;
      RECT 14442.06 228.445 14455.06 291.075 ;
      RECT 14442.06 194.37 14455.06 212.075 ;
      RECT 14442.06 189.04 14447.37 212.075 ;
      RECT 14442.06 189.04 14455.06 190.17 ;
      RECT 14425.08 307.445 14438.08 350.165 ;
      RECT 14426.705 189.04 14438.08 350.165 ;
      RECT 14425.08 228.445 14438.08 291.075 ;
      RECT 14425.08 189.04 14438.08 212.075 ;
      RECT 14394.56 324.445 14422.56 350.165 ;
      RECT 14400.705 189.04 14417.125 350.165 ;
      RECT 14394.56 211.445 14395.795 350.165 ;
      RECT 14394.56 211.445 14421.795 308.075 ;
      RECT 14394.56 228.445 14422.56 291.075 ;
      RECT 14396.925 189.04 14417.125 308.075 ;
      RECT 14394.56 189.04 14422.56 195.075 ;
      RECT 14379.04 228.445 14392.04 350.165 ;
      RECT 14379.04 189.04 14385.395 350.165 ;
      RECT 14379.04 189.04 14392.04 212.075 ;
      RECT 14362.06 290.445 14375.06 330.165 ;
      RECT 14373.19 189.04 14375.06 330.165 ;
      RECT 14371.425 194.425 14375.06 330.165 ;
      RECT 14362.06 189.04 14363.675 330.165 ;
      RECT 14362.06 194.425 14375.06 259.875 ;
      RECT 14362.06 189.04 14370.41 259.875 ;
      RECT 14362.06 189.04 14375.06 190.125 ;
      RECT 14345.08 211.445 14358.08 350.165 ;
      RECT 14345.425 189.04 14358.08 350.165 ;
      RECT 14345.08 189.04 14358.08 195.075 ;
      RECT 14314.56 259.445 14342.56 350.165 ;
      RECT 14326.935 211.445 14342.56 350.165 ;
      RECT 14314.56 189.04 14319.185 350.165 ;
      RECT 14314.56 189.04 14340.515 228.875 ;
      RECT 14314.56 189.04 14342.56 195.075 ;
      RECT 14299.04 307.445 14312.04 350.165 ;
      RECT 14309.035 194.37 14312.04 350.165 ;
      RECT 14299.04 189.04 14304.125 350.165 ;
      RECT 14299.04 228.445 14312.04 291.075 ;
      RECT 14299.04 194.37 14312.04 212.075 ;
      RECT 14299.04 189.04 14307.37 212.075 ;
      RECT 14299.04 189.04 14312.04 190.17 ;
      RECT 14282.06 307.445 14295.06 330.165 ;
      RECT 14286.705 189.04 14295.06 330.165 ;
      RECT 14286.54 228.445 14295.06 330.165 ;
      RECT 14282.06 228.445 14295.06 291.075 ;
      RECT 14282.06 189.04 14295.06 212.075 ;
      RECT 14265.08 324.445 14278.08 350.165 ;
      RECT 14265.08 189.04 14277.125 350.165 ;
      RECT 14265.08 211.445 14278.08 308.075 ;
      RECT 14265.08 189.04 14278.08 195.075 ;
      RECT 14234.56 324.445 14262.56 350.165 ;
      RECT 14260.705 189.04 14262.56 350.165 ;
      RECT 14234.56 228.445 14255.795 350.165 ;
      RECT 14258.115 189.04 14262.56 308.075 ;
      RECT 14241.11 211.445 14262.56 308.075 ;
      RECT 14234.56 189.04 14253.205 212.075 ;
      RECT 14234.56 189.04 14262.56 195.075 ;
      RECT 14219.04 290.445 14232.04 350.165 ;
      RECT 14231.425 194.42 14232.04 350.165 ;
      RECT 14219.04 189.04 14223.675 350.165 ;
      RECT 14219.04 194.42 14232.04 259.875 ;
      RECT 14219.04 189.04 14230.41 259.875 ;
      RECT 14219.04 189.04 14232.04 190.125 ;
      RECT 14202.06 211.445 14215.06 330.165 ;
      RECT 14205.425 189.04 14215.06 330.165 ;
      RECT 14202.06 189.04 14215.06 195.075 ;
      RECT 14185.08 259.445 14198.08 350.165 ;
      RECT 14186.935 189.04 14198.08 350.165 ;
      RECT 14185.08 189.04 14198.08 228.875 ;
      RECT 14154.56 307.445 14182.56 350.165 ;
      RECT 14169.035 259.445 14182.56 350.165 ;
      RECT 14154.56 189.04 14164.125 350.165 ;
      RECT 14154.56 228.445 14179.185 291.075 ;
      RECT 14173.09 189.04 14182.56 228.875 ;
      RECT 14169.035 194.37 14182.56 228.875 ;
      RECT 14154.56 194.37 14182.56 212.075 ;
      RECT 14154.56 189.04 14167.37 212.075 ;
      RECT 14154.56 189.04 14182.56 190.17 ;
      RECT 14139.04 324.445 14152.04 350.165 ;
      RECT 14146.705 189.04 14152.04 350.165 ;
      RECT 14142.035 307.445 14152.04 350.165 ;
      RECT 14139.04 307.445 14152.04 308.075 ;
      RECT 14139.04 211.445 14141.795 308.075 ;
      RECT 14139.04 228.445 14152.04 291.075 ;
      RECT 14139.04 211.445 14152.04 212.075 ;
      RECT 14142.035 189.04 14152.04 212.075 ;
      RECT 14139.04 189.04 14152.04 195.075 ;
      RECT 14105.08 324.445 14118.08 350.165 ;
      RECT 14105.08 228.445 14115.795 350.165 ;
      RECT 14110.31 211.445 14118.08 308.075 ;
      RECT 14105.08 189.04 14113.125 212.075 ;
      RECT 14105.08 189.04 14118.08 195.075 ;
      RECT 14074.56 290.445 14102.56 350.165 ;
      RECT 14093.19 189.04 14102.56 350.165 ;
      RECT 14091.425 194.425 14102.56 350.165 ;
      RECT 14074.56 189.04 14083.675 350.165 ;
      RECT 14074.56 194.425 14102.56 259.875 ;
      RECT 14074.56 189.04 14090.41 259.875 ;
      RECT 14074.56 189.04 14102.56 190.125 ;
      RECT 14059.04 211.445 14072.04 350.165 ;
      RECT 14065.425 189.04 14072.04 350.165 ;
      RECT 14059.04 189.04 14060.515 350.165 ;
      RECT 14059.04 189.04 14072.04 195.075 ;
      RECT 14042.06 259.445 14055.06 330.165 ;
      RECT 14046.935 189.04 14055.06 330.165 ;
      RECT 14042.06 189.04 14055.06 228.875 ;
      RECT 14025.08 307.445 14038.08 350.165 ;
      RECT 14033.09 189.04 14038.08 350.165 ;
      RECT 14029.035 194.37 14038.08 350.165 ;
      RECT 14025.08 228.445 14038.08 291.075 ;
      RECT 14025.08 194.37 14038.08 212.075 ;
      RECT 14025.08 189.04 14027.37 212.075 ;
      RECT 14025.08 189.04 14038.08 190.38 ;
      RECT 13994.56 324.445 14022.56 350.165 ;
      RECT 14006.705 189.04 14022.56 350.165 ;
      RECT 14002.035 307.445 14022.56 350.165 ;
      RECT 13994.56 189.04 13997.125 350.165 ;
      RECT 13994.56 307.445 14022.56 308.075 ;
      RECT 13994.56 211.445 14001.795 308.075 ;
      RECT 13994.56 228.445 14022.56 291.075 ;
      RECT 13994.56 211.445 14022.56 212.075 ;
      RECT 14002.035 189.04 14022.56 212.075 ;
      RECT 13994.56 189.04 14022.56 195.075 ;
      RECT 13979.04 324.445 13992.04 350.165 ;
      RECT 13980.705 189.04 13992.04 350.165 ;
      RECT 13979.04 189.04 13992.04 308.075 ;
      RECT 13962.06 228.445 13975.06 330.165 ;
      RECT 13968.69 211.445 13975.06 330.165 ;
      RECT 13962.06 189.04 13972.015 212.075 ;
      RECT 13962.06 189.04 13975.06 195.075 ;
      RECT 13945.08 290.445 13958.08 350.165 ;
      RECT 13953.19 189.04 13958.08 350.165 ;
      RECT 13951.425 194.425 13958.08 350.165 ;
      RECT 13945.08 194.425 13958.08 259.875 ;
      RECT 13945.08 189.04 13950.41 259.875 ;
      RECT 13945.08 189.04 13958.08 190.125 ;
      RECT 13914.56 211.445 13942.56 350.165 ;
      RECT 13925.425 189.04 13942.56 350.165 ;
      RECT 13914.56 189.04 13920.515 350.165 ;
      RECT 13914.56 189.04 13942.56 195.075 ;
      RECT 13899.04 259.445 13912.04 350.165 ;
      RECT 13906.935 189.04 13912.04 350.165 ;
      RECT 13899.04 189.04 13912.04 228.875 ;
      RECT 13882.06 307.445 13895.06 330.165 ;
      RECT 13892.99 189.04 13895.06 330.165 ;
      RECT 13889.035 194.37 13895.06 330.165 ;
      RECT 13882.06 189.04 13884.125 330.165 ;
      RECT 13882.06 228.445 13895.06 291.075 ;
      RECT 13882.06 194.37 13895.06 212.075 ;
      RECT 13882.06 189.04 13887.37 212.075 ;
      RECT 13882.06 189.04 13895.06 190.17 ;
      RECT 13865.08 307.445 13878.08 350.165 ;
      RECT 13866.705 189.04 13878.08 350.165 ;
      RECT 13865.08 228.445 13878.08 291.075 ;
      RECT 13865.08 189.04 13878.08 212.075 ;
      RECT 13834.56 324.445 13862.56 350.165 ;
      RECT 13840.705 189.04 13857.125 350.165 ;
      RECT 13834.56 211.445 13835.795 350.165 ;
      RECT 13834.56 211.445 13861.795 308.075 ;
      RECT 13834.56 228.445 13862.56 291.075 ;
      RECT 13836.925 189.04 13857.125 308.075 ;
      RECT 13834.56 189.04 13862.56 195.075 ;
      RECT 13819.04 228.445 13832.04 350.165 ;
      RECT 13819.04 189.04 13825.395 350.165 ;
      RECT 13819.04 189.04 13832.04 212.075 ;
      RECT 13802.06 290.445 13815.06 330.165 ;
      RECT 13813.19 189.04 13815.06 330.165 ;
      RECT 13811.425 194.425 13815.06 330.165 ;
      RECT 13802.06 189.04 13803.675 330.165 ;
      RECT 13802.06 194.425 13815.06 259.875 ;
      RECT 13802.06 189.04 13810.41 259.875 ;
      RECT 13802.06 189.04 13815.06 190.125 ;
      RECT 13785.08 211.445 13798.08 350.165 ;
      RECT 13785.425 189.04 13798.08 350.165 ;
      RECT 13785.08 189.04 13798.08 195.075 ;
      RECT 13754.56 259.445 13782.56 350.165 ;
      RECT 13766.935 211.445 13782.56 350.165 ;
      RECT 13754.56 189.04 13759.185 350.165 ;
      RECT 13754.56 189.04 13780.515 228.875 ;
      RECT 13754.56 189.04 13782.56 195.075 ;
      RECT 13739.04 307.445 13752.04 350.165 ;
      RECT 13749.035 194.37 13752.04 350.165 ;
      RECT 13739.04 189.04 13744.125 350.165 ;
      RECT 13739.04 228.445 13752.04 291.075 ;
      RECT 13739.04 194.37 13752.04 212.075 ;
      RECT 13739.04 189.04 13747.37 212.075 ;
      RECT 13739.04 189.04 13752.04 190.17 ;
      RECT 13722.06 307.445 13735.06 330.165 ;
      RECT 13726.705 189.04 13735.06 330.165 ;
      RECT 13726.54 228.445 13735.06 330.165 ;
      RECT 13722.06 228.445 13735.06 291.075 ;
      RECT 13722.06 189.04 13735.06 212.075 ;
      RECT 13705.08 324.445 13718.08 350.165 ;
      RECT 13705.08 189.04 13717.125 350.165 ;
      RECT 13705.08 211.445 13718.08 308.075 ;
      RECT 13705.08 189.04 13718.08 195.075 ;
      RECT 13674.56 324.445 13702.56 350.165 ;
      RECT 13700.705 189.04 13702.56 350.165 ;
      RECT 13674.56 228.445 13695.795 350.165 ;
      RECT 13698.115 189.04 13702.56 308.075 ;
      RECT 13681.11 211.445 13702.56 308.075 ;
      RECT 13674.56 189.04 13693.205 212.075 ;
      RECT 13674.56 189.04 13702.56 195.075 ;
      RECT 13659.04 290.445 13672.04 350.165 ;
      RECT 13671.425 194.42 13672.04 350.165 ;
      RECT 13659.04 189.04 13663.675 350.165 ;
      RECT 13659.04 194.42 13672.04 259.875 ;
      RECT 13659.04 189.04 13670.41 259.875 ;
      RECT 13659.04 189.04 13672.04 190.125 ;
      RECT 13642.06 211.445 13655.06 330.165 ;
      RECT 13645.425 189.04 13655.06 330.165 ;
      RECT 13642.06 189.04 13655.06 195.075 ;
      RECT 13625.08 259.445 13638.08 350.165 ;
      RECT 13626.935 189.04 13638.08 350.165 ;
      RECT 13625.08 189.04 13638.08 228.875 ;
      RECT 13594.56 307.445 13622.56 350.165 ;
      RECT 13609.035 259.445 13622.56 350.165 ;
      RECT 13594.56 189.04 13604.125 350.165 ;
      RECT 13594.56 228.445 13619.185 291.075 ;
      RECT 13613.09 189.04 13622.56 228.875 ;
      RECT 13609.035 194.37 13622.56 228.875 ;
      RECT 13594.56 194.37 13622.56 212.075 ;
      RECT 13594.56 189.04 13607.37 212.075 ;
      RECT 13594.56 189.04 13622.56 190.17 ;
      RECT 13579.04 324.445 13592.04 350.165 ;
      RECT 13586.705 189.04 13592.04 350.165 ;
      RECT 13582.035 307.445 13592.04 350.165 ;
      RECT 13579.04 307.445 13592.04 308.075 ;
      RECT 13579.04 211.445 13581.795 308.075 ;
      RECT 13579.04 228.445 13592.04 291.075 ;
      RECT 13579.04 211.445 13592.04 212.075 ;
      RECT 13582.035 189.04 13592.04 212.075 ;
      RECT 13579.04 189.04 13592.04 195.075 ;
      RECT 13545.08 324.445 13558.08 350.165 ;
      RECT 13545.08 228.445 13555.795 350.165 ;
      RECT 13550.31 211.445 13558.08 308.075 ;
      RECT 13545.08 189.04 13553.125 212.075 ;
      RECT 13545.08 189.04 13558.08 195.075 ;
      RECT 13514.56 290.445 13542.56 350.165 ;
      RECT 13533.19 189.04 13542.56 350.165 ;
      RECT 13531.425 194.425 13542.56 350.165 ;
      RECT 13514.56 189.04 13523.675 350.165 ;
      RECT 13514.56 194.425 13542.56 259.875 ;
      RECT 13514.56 189.04 13530.41 259.875 ;
      RECT 13514.56 189.04 13542.56 190.125 ;
      RECT 13499.04 211.445 13512.04 350.165 ;
      RECT 13505.425 189.04 13512.04 350.165 ;
      RECT 13499.04 189.04 13500.515 350.165 ;
      RECT 13499.04 189.04 13512.04 195.075 ;
      RECT 13482.06 259.445 13495.06 330.165 ;
      RECT 13486.935 189.04 13495.06 330.165 ;
      RECT 13482.06 189.04 13495.06 228.875 ;
      RECT 13465.08 307.445 13478.08 350.165 ;
      RECT 13473.09 189.04 13478.08 350.165 ;
      RECT 13469.035 194.37 13478.08 350.165 ;
      RECT 13465.08 228.445 13478.08 291.075 ;
      RECT 13465.08 194.37 13478.08 212.075 ;
      RECT 13465.08 189.04 13467.37 212.075 ;
      RECT 13465.08 189.04 13478.08 190.38 ;
      RECT 13434.56 324.445 13462.56 350.165 ;
      RECT 13446.705 189.04 13462.56 350.165 ;
      RECT 13442.035 307.445 13462.56 350.165 ;
      RECT 13434.56 189.04 13437.125 350.165 ;
      RECT 13434.56 307.445 13462.56 308.075 ;
      RECT 13434.56 211.445 13441.795 308.075 ;
      RECT 13434.56 228.445 13462.56 291.075 ;
      RECT 13434.56 211.445 13462.56 212.075 ;
      RECT 13442.035 189.04 13462.56 212.075 ;
      RECT 13434.56 189.04 13462.56 195.075 ;
      RECT 13419.04 324.445 13432.04 350.165 ;
      RECT 13420.705 189.04 13432.04 350.165 ;
      RECT 13419.04 189.04 13432.04 308.075 ;
      RECT 13402.06 228.445 13415.06 330.165 ;
      RECT 13408.69 211.445 13415.06 330.165 ;
      RECT 13402.06 189.04 13412.015 212.075 ;
      RECT 13402.06 189.04 13415.06 195.075 ;
      RECT 13385.08 290.445 13398.08 350.165 ;
      RECT 13393.19 189.04 13398.08 350.165 ;
      RECT 13391.425 194.425 13398.08 350.165 ;
      RECT 13385.08 194.425 13398.08 259.875 ;
      RECT 13385.08 189.04 13390.41 259.875 ;
      RECT 13385.08 189.04 13398.08 190.125 ;
      RECT 13354.56 211.445 13382.56 350.165 ;
      RECT 13365.425 189.04 13382.56 350.165 ;
      RECT 13354.56 189.04 13360.515 350.165 ;
      RECT 13354.56 189.04 13382.56 195.075 ;
      RECT 13339.04 259.445 13352.04 350.165 ;
      RECT 13346.935 189.04 13352.04 350.165 ;
      RECT 13339.04 189.04 13352.04 228.875 ;
      RECT 13322.06 307.445 13335.06 330.165 ;
      RECT 13332.99 189.04 13335.06 330.165 ;
      RECT 13329.035 194.37 13335.06 330.165 ;
      RECT 13322.06 189.04 13324.125 330.165 ;
      RECT 13322.06 228.445 13335.06 291.075 ;
      RECT 13322.06 194.37 13335.06 212.075 ;
      RECT 13322.06 189.04 13327.37 212.075 ;
      RECT 13322.06 189.04 13335.06 190.17 ;
      RECT 13305.08 307.445 13318.08 350.165 ;
      RECT 13306.705 189.04 13318.08 350.165 ;
      RECT 13305.08 228.445 13318.08 291.075 ;
      RECT 13305.08 189.04 13318.08 212.075 ;
      RECT 13274.56 324.445 13302.56 350.165 ;
      RECT 13280.705 189.04 13297.125 350.165 ;
      RECT 13274.56 211.445 13275.795 350.165 ;
      RECT 13274.56 211.445 13301.795 308.075 ;
      RECT 13274.56 228.445 13302.56 291.075 ;
      RECT 13276.925 189.04 13297.125 308.075 ;
      RECT 13274.56 189.04 13302.56 195.075 ;
      RECT 13259.04 228.445 13272.04 350.165 ;
      RECT 13259.04 189.04 13265.395 350.165 ;
      RECT 13259.04 189.04 13272.04 212.075 ;
      RECT 13242.06 290.445 13255.06 330.165 ;
      RECT 13253.19 189.04 13255.06 330.165 ;
      RECT 13251.425 194.425 13255.06 330.165 ;
      RECT 13242.06 189.04 13243.675 330.165 ;
      RECT 13242.06 194.425 13255.06 259.875 ;
      RECT 13242.06 189.04 13250.41 259.875 ;
      RECT 13242.06 189.04 13255.06 190.125 ;
      RECT 13225.08 211.445 13238.08 350.165 ;
      RECT 13225.425 189.04 13238.08 350.165 ;
      RECT 13225.08 189.04 13238.08 195.075 ;
      RECT 13194.56 259.445 13222.56 350.165 ;
      RECT 13206.935 211.445 13222.56 350.165 ;
      RECT 13194.56 189.04 13199.185 350.165 ;
      RECT 13194.56 189.04 13220.515 228.875 ;
      RECT 13194.56 189.04 13222.56 195.075 ;
      RECT 13179.04 307.445 13192.04 350.165 ;
      RECT 13189.035 194.37 13192.04 350.165 ;
      RECT 13179.04 189.04 13184.125 350.165 ;
      RECT 13179.04 228.445 13192.04 291.075 ;
      RECT 13179.04 194.37 13192.04 212.075 ;
      RECT 13179.04 189.04 13187.37 212.075 ;
      RECT 13179.04 189.04 13192.04 190.17 ;
      RECT 13162.06 307.445 13175.06 330.165 ;
      RECT 13166.705 189.04 13175.06 330.165 ;
      RECT 13166.54 228.445 13175.06 330.165 ;
      RECT 13162.06 228.445 13175.06 291.075 ;
      RECT 13162.06 189.04 13175.06 212.075 ;
      RECT 13145.08 324.445 13158.08 350.165 ;
      RECT 13145.08 189.04 13157.125 350.165 ;
      RECT 13145.08 211.445 13158.08 308.075 ;
      RECT 13145.08 189.04 13158.08 195.075 ;
      RECT 13114.56 324.445 13142.56 350.165 ;
      RECT 13140.705 189.04 13142.56 350.165 ;
      RECT 13114.56 228.445 13135.795 350.165 ;
      RECT 13138.115 189.04 13142.56 308.075 ;
      RECT 13121.11 211.445 13142.56 308.075 ;
      RECT 13114.56 189.04 13133.205 212.075 ;
      RECT 13114.56 189.04 13142.56 195.075 ;
      RECT 13099.04 290.445 13112.04 350.165 ;
      RECT 13111.425 194.42 13112.04 350.165 ;
      RECT 13099.04 189.04 13103.675 350.165 ;
      RECT 13099.04 194.42 13112.04 259.875 ;
      RECT 13099.04 189.04 13110.41 259.875 ;
      RECT 13099.04 189.04 13112.04 190.125 ;
      RECT 13082.06 211.445 13095.06 330.165 ;
      RECT 13085.425 189.04 13095.06 330.165 ;
      RECT 13082.06 189.04 13095.06 195.075 ;
      RECT 13065.08 259.445 13078.08 350.165 ;
      RECT 13066.935 189.04 13078.08 350.165 ;
      RECT 13065.08 189.04 13078.08 228.875 ;
      RECT 13034.56 307.445 13062.56 350.165 ;
      RECT 13049.035 259.445 13062.56 350.165 ;
      RECT 13034.56 189.04 13044.125 350.165 ;
      RECT 13034.56 228.445 13059.185 291.075 ;
      RECT 13053.09 189.04 13062.56 228.875 ;
      RECT 13049.035 194.37 13062.56 228.875 ;
      RECT 13034.56 194.37 13062.56 212.075 ;
      RECT 13034.56 189.04 13047.37 212.075 ;
      RECT 13034.56 189.04 13062.56 190.17 ;
      RECT 13019.04 324.445 13032.04 350.165 ;
      RECT 13026.705 189.04 13032.04 350.165 ;
      RECT 13022.035 307.445 13032.04 350.165 ;
      RECT 13019.04 307.445 13032.04 308.075 ;
      RECT 13019.04 211.445 13021.795 308.075 ;
      RECT 13019.04 228.445 13032.04 291.075 ;
      RECT 13019.04 211.445 13032.04 212.075 ;
      RECT 13022.035 189.04 13032.04 212.075 ;
      RECT 13019.04 189.04 13032.04 195.075 ;
      RECT 12985.08 324.445 12998.08 350.165 ;
      RECT 12985.08 228.445 12995.795 350.165 ;
      RECT 12990.31 211.445 12998.08 308.075 ;
      RECT 12985.08 189.04 12993.125 212.075 ;
      RECT 12985.08 189.04 12998.08 195.075 ;
      RECT 12954.56 290.445 12982.56 350.165 ;
      RECT 12973.19 189.04 12982.56 350.165 ;
      RECT 12971.425 194.425 12982.56 350.165 ;
      RECT 12954.56 189.04 12963.675 350.165 ;
      RECT 12954.56 194.425 12982.56 259.875 ;
      RECT 12954.56 189.04 12970.41 259.875 ;
      RECT 12954.56 189.04 12982.56 190.125 ;
      RECT 12939.04 211.445 12952.04 350.165 ;
      RECT 12945.425 189.04 12952.04 350.165 ;
      RECT 12939.04 189.04 12940.515 350.165 ;
      RECT 12939.04 189.04 12952.04 195.075 ;
      RECT 12922.06 259.445 12935.06 330.165 ;
      RECT 12926.935 189.04 12935.06 330.165 ;
      RECT 12922.06 189.04 12935.06 228.875 ;
      RECT 12905.08 307.445 12918.08 350.165 ;
      RECT 12913.09 189.04 12918.08 350.165 ;
      RECT 12909.035 194.37 12918.08 350.165 ;
      RECT 12905.08 228.445 12918.08 291.075 ;
      RECT 12905.08 194.37 12918.08 212.075 ;
      RECT 12905.08 189.04 12907.37 212.075 ;
      RECT 12905.08 189.04 12918.08 190.38 ;
      RECT 12874.56 324.445 12902.56 350.165 ;
      RECT 12886.705 189.04 12902.56 350.165 ;
      RECT 12882.035 307.445 12902.56 350.165 ;
      RECT 12874.56 189.04 12877.125 350.165 ;
      RECT 12874.56 307.445 12902.56 308.075 ;
      RECT 12874.56 211.445 12881.795 308.075 ;
      RECT 12874.56 228.445 12902.56 291.075 ;
      RECT 12874.56 211.445 12902.56 212.075 ;
      RECT 12882.035 189.04 12902.56 212.075 ;
      RECT 12874.56 189.04 12902.56 195.075 ;
      RECT 12859.04 324.445 12872.04 350.165 ;
      RECT 12860.705 189.04 12872.04 350.165 ;
      RECT 12859.04 189.04 12872.04 308.075 ;
      RECT 12842.06 228.445 12855.06 330.165 ;
      RECT 12848.69 211.445 12855.06 330.165 ;
      RECT 12842.06 189.04 12852.015 212.075 ;
      RECT 12842.06 189.04 12855.06 195.075 ;
      RECT 12825.08 290.445 12838.08 350.165 ;
      RECT 12833.19 189.04 12838.08 350.165 ;
      RECT 12831.425 194.425 12838.08 350.165 ;
      RECT 12825.08 194.425 12838.08 259.875 ;
      RECT 12825.08 189.04 12830.41 259.875 ;
      RECT 12825.08 189.04 12838.08 190.125 ;
      RECT 12794.56 211.445 12822.56 350.165 ;
      RECT 12805.425 189.04 12822.56 350.165 ;
      RECT 12794.56 189.04 12800.515 350.165 ;
      RECT 12794.56 189.04 12822.56 195.075 ;
      RECT 12779.04 259.445 12792.04 350.165 ;
      RECT 12786.935 189.04 12792.04 350.165 ;
      RECT 12779.04 189.04 12792.04 228.875 ;
      RECT 12762.06 307.445 12775.06 330.165 ;
      RECT 12772.99 189.04 12775.06 330.165 ;
      RECT 12769.035 194.37 12775.06 330.165 ;
      RECT 12762.06 189.04 12764.125 330.165 ;
      RECT 12762.06 228.445 12775.06 291.075 ;
      RECT 12762.06 194.37 12775.06 212.075 ;
      RECT 12762.06 189.04 12767.37 212.075 ;
      RECT 12762.06 189.04 12775.06 190.17 ;
      RECT 12745.08 307.445 12758.08 350.165 ;
      RECT 12746.705 189.04 12758.08 350.165 ;
      RECT 12745.08 228.445 12758.08 291.075 ;
      RECT 12745.08 189.04 12758.08 212.075 ;
      RECT 12714.56 324.445 12742.56 350.165 ;
      RECT 12720.705 189.04 12737.125 350.165 ;
      RECT 12714.56 211.445 12715.795 350.165 ;
      RECT 12714.56 211.445 12741.795 308.075 ;
      RECT 12714.56 228.445 12742.56 291.075 ;
      RECT 12716.925 189.04 12737.125 308.075 ;
      RECT 12714.56 189.04 12742.56 195.075 ;
      RECT 12699.04 228.445 12712.04 350.165 ;
      RECT 12699.04 189.04 12705.395 350.165 ;
      RECT 12699.04 189.04 12712.04 212.075 ;
      RECT 12682.06 290.445 12695.06 330.165 ;
      RECT 12693.19 189.04 12695.06 330.165 ;
      RECT 12691.425 194.425 12695.06 330.165 ;
      RECT 12682.06 189.04 12683.675 330.165 ;
      RECT 12682.06 194.425 12695.06 259.875 ;
      RECT 12682.06 189.04 12690.41 259.875 ;
      RECT 12682.06 189.04 12695.06 190.125 ;
      RECT 12665.08 211.445 12678.08 350.165 ;
      RECT 12665.425 189.04 12678.08 350.165 ;
      RECT 12665.08 189.04 12678.08 195.075 ;
      RECT 12634.56 259.445 12662.56 350.165 ;
      RECT 12646.935 211.445 12662.56 350.165 ;
      RECT 12634.56 189.04 12639.185 350.165 ;
      RECT 12634.56 189.04 12660.515 228.875 ;
      RECT 12634.56 189.04 12662.56 195.075 ;
      RECT 12619.04 307.445 12632.04 350.165 ;
      RECT 12629.035 194.37 12632.04 350.165 ;
      RECT 12619.04 189.04 12624.125 350.165 ;
      RECT 12619.04 228.445 12632.04 291.075 ;
      RECT 12619.04 194.37 12632.04 212.075 ;
      RECT 12619.04 189.04 12627.37 212.075 ;
      RECT 12619.04 189.04 12632.04 190.17 ;
      RECT 12602.06 307.445 12615.06 330.165 ;
      RECT 12606.705 189.04 12615.06 330.165 ;
      RECT 12606.54 228.445 12615.06 330.165 ;
      RECT 12602.06 228.445 12615.06 291.075 ;
      RECT 12602.06 189.04 12615.06 212.075 ;
      RECT 12585.08 324.445 12598.08 350.165 ;
      RECT 12585.08 189.04 12597.125 350.165 ;
      RECT 12585.08 211.445 12598.08 308.075 ;
      RECT 12585.08 189.04 12598.08 195.075 ;
      RECT 12554.56 324.445 12582.56 350.165 ;
      RECT 12580.705 189.04 12582.56 350.165 ;
      RECT 12554.56 228.445 12575.795 350.165 ;
      RECT 12578.115 189.04 12582.56 308.075 ;
      RECT 12561.11 211.445 12582.56 308.075 ;
      RECT 12554.56 189.04 12573.205 212.075 ;
      RECT 12554.56 189.04 12582.56 195.075 ;
      RECT 12539.04 290.445 12552.04 350.165 ;
      RECT 12551.425 194.42 12552.04 350.165 ;
      RECT 12539.04 189.04 12543.675 350.165 ;
      RECT 12539.04 194.42 12552.04 259.875 ;
      RECT 12539.04 189.04 12550.41 259.875 ;
      RECT 12539.04 189.04 12552.04 190.125 ;
      RECT 12522.06 211.445 12535.06 330.165 ;
      RECT 12525.425 189.04 12535.06 330.165 ;
      RECT 12522.06 189.04 12535.06 195.075 ;
      RECT 12505.08 259.445 12518.08 350.165 ;
      RECT 12506.935 189.04 12518.08 350.165 ;
      RECT 12505.08 189.04 12518.08 228.875 ;
      RECT 12474.56 307.445 12502.56 350.165 ;
      RECT 12489.035 259.445 12502.56 350.165 ;
      RECT 12474.56 189.04 12484.125 350.165 ;
      RECT 12474.56 228.445 12499.185 291.075 ;
      RECT 12493.09 189.04 12502.56 228.875 ;
      RECT 12489.035 194.37 12502.56 228.875 ;
      RECT 12474.56 194.37 12502.56 212.075 ;
      RECT 12474.56 189.04 12487.37 212.075 ;
      RECT 12474.56 189.04 12502.56 190.17 ;
      RECT 12459.04 324.445 12472.04 350.165 ;
      RECT 12466.705 189.04 12472.04 350.165 ;
      RECT 12462.035 307.445 12472.04 350.165 ;
      RECT 12459.04 307.445 12472.04 308.075 ;
      RECT 12459.04 211.445 12461.795 308.075 ;
      RECT 12459.04 228.445 12472.04 291.075 ;
      RECT 12459.04 211.445 12472.04 212.075 ;
      RECT 12462.035 189.04 12472.04 212.075 ;
      RECT 12459.04 189.04 12472.04 195.075 ;
      RECT 12425.08 324.445 12438.08 350.165 ;
      RECT 12425.08 228.445 12435.795 350.165 ;
      RECT 12430.31 211.445 12438.08 308.075 ;
      RECT 12425.08 189.04 12433.125 212.075 ;
      RECT 12425.08 189.04 12438.08 195.075 ;
      RECT 12394.56 290.445 12422.56 350.165 ;
      RECT 12413.19 189.04 12422.56 350.165 ;
      RECT 12411.425 194.425 12422.56 350.165 ;
      RECT 12394.56 189.04 12403.675 350.165 ;
      RECT 12394.56 194.425 12422.56 259.875 ;
      RECT 12394.56 189.04 12410.41 259.875 ;
      RECT 12394.56 189.04 12422.56 190.125 ;
      RECT 12379.04 211.445 12392.04 350.165 ;
      RECT 12385.425 189.04 12392.04 350.165 ;
      RECT 12379.04 189.04 12380.515 350.165 ;
      RECT 12379.04 189.04 12392.04 195.075 ;
      RECT 12362.06 259.445 12375.06 330.165 ;
      RECT 12366.935 189.04 12375.06 330.165 ;
      RECT 12362.06 189.04 12375.06 228.875 ;
      RECT 12345.08 307.445 12358.08 350.165 ;
      RECT 12353.09 189.04 12358.08 350.165 ;
      RECT 12349.035 194.37 12358.08 350.165 ;
      RECT 12345.08 228.445 12358.08 291.075 ;
      RECT 12345.08 194.37 12358.08 212.075 ;
      RECT 12345.08 189.04 12347.37 212.075 ;
      RECT 12345.08 189.04 12358.08 190.38 ;
      RECT 12314.56 324.445 12342.56 350.165 ;
      RECT 12326.705 189.04 12342.56 350.165 ;
      RECT 12322.035 307.445 12342.56 350.165 ;
      RECT 12314.56 189.04 12317.125 350.165 ;
      RECT 12314.56 307.445 12342.56 308.075 ;
      RECT 12314.56 211.445 12321.795 308.075 ;
      RECT 12314.56 228.445 12342.56 291.075 ;
      RECT 12314.56 211.445 12342.56 212.075 ;
      RECT 12322.035 189.04 12342.56 212.075 ;
      RECT 12314.56 189.04 12342.56 195.075 ;
      RECT 12299.04 324.445 12312.04 350.165 ;
      RECT 12300.705 189.04 12312.04 350.165 ;
      RECT 12299.04 189.04 12312.04 308.075 ;
      RECT 12282.06 228.445 12295.06 330.165 ;
      RECT 12288.69 211.445 12295.06 330.165 ;
      RECT 12282.06 189.04 12292.015 212.075 ;
      RECT 12282.06 189.04 12295.06 195.075 ;
      RECT 12265.08 290.445 12278.08 350.165 ;
      RECT 12273.19 189.04 12278.08 350.165 ;
      RECT 12271.425 194.425 12278.08 350.165 ;
      RECT 12265.08 194.425 12278.08 259.875 ;
      RECT 12265.08 189.04 12270.41 259.875 ;
      RECT 12265.08 189.04 12278.08 190.125 ;
      RECT 12234.56 211.445 12262.56 350.165 ;
      RECT 12245.425 189.04 12262.56 350.165 ;
      RECT 12234.56 189.04 12240.515 350.165 ;
      RECT 12234.56 189.04 12262.56 195.075 ;
      RECT 12219.04 259.445 12232.04 350.165 ;
      RECT 12226.935 189.04 12232.04 350.165 ;
      RECT 12219.04 189.04 12232.04 228.875 ;
      RECT 12202.06 307.445 12215.06 330.165 ;
      RECT 12212.99 189.04 12215.06 330.165 ;
      RECT 12209.035 194.37 12215.06 330.165 ;
      RECT 12202.06 189.04 12204.125 330.165 ;
      RECT 12202.06 228.445 12215.06 291.075 ;
      RECT 12202.06 194.37 12215.06 212.075 ;
      RECT 12202.06 189.04 12207.37 212.075 ;
      RECT 12202.06 189.04 12215.06 190.17 ;
      RECT 12185.08 307.445 12198.08 350.165 ;
      RECT 12186.705 189.04 12198.08 350.165 ;
      RECT 12185.08 228.445 12198.08 291.075 ;
      RECT 12185.08 189.04 12198.08 212.075 ;
      RECT 12154.56 324.445 12182.56 350.165 ;
      RECT 12160.705 189.04 12177.125 350.165 ;
      RECT 12154.56 211.445 12155.795 350.165 ;
      RECT 12154.56 211.445 12181.795 308.075 ;
      RECT 12154.56 228.445 12182.56 291.075 ;
      RECT 12156.925 189.04 12177.125 308.075 ;
      RECT 12154.56 189.04 12182.56 195.075 ;
      RECT 12139.04 228.445 12152.04 350.165 ;
      RECT 12139.04 189.04 12145.395 350.165 ;
      RECT 12139.04 189.04 12152.04 212.075 ;
      RECT 12122.06 290.445 12135.06 330.165 ;
      RECT 12133.19 189.04 12135.06 330.165 ;
      RECT 12131.425 194.425 12135.06 330.165 ;
      RECT 12122.06 189.04 12123.675 330.165 ;
      RECT 12122.06 194.425 12135.06 259.875 ;
      RECT 12122.06 189.04 12130.41 259.875 ;
      RECT 12122.06 189.04 12135.06 190.125 ;
      RECT 12105.08 211.445 12118.08 350.165 ;
      RECT 12105.425 189.04 12118.08 350.165 ;
      RECT 12105.08 189.04 12118.08 195.075 ;
      RECT 12074.56 259.445 12102.56 350.165 ;
      RECT 12086.935 211.445 12102.56 350.165 ;
      RECT 12074.56 189.04 12079.185 350.165 ;
      RECT 12074.56 189.04 12100.515 228.875 ;
      RECT 12074.56 189.04 12102.56 195.075 ;
      RECT 12059.04 307.445 12072.04 350.165 ;
      RECT 12069.035 194.37 12072.04 350.165 ;
      RECT 12059.04 189.04 12064.125 350.165 ;
      RECT 12059.04 228.445 12072.04 291.075 ;
      RECT 12059.04 194.37 12072.04 212.075 ;
      RECT 12059.04 189.04 12067.37 212.075 ;
      RECT 12059.04 189.04 12072.04 190.17 ;
      RECT 12042.06 307.445 12055.06 330.165 ;
      RECT 12046.705 189.04 12055.06 330.165 ;
      RECT 12046.54 228.445 12055.06 330.165 ;
      RECT 12042.06 228.445 12055.06 291.075 ;
      RECT 12042.06 189.04 12055.06 212.075 ;
      RECT 12025.08 324.445 12038.08 350.165 ;
      RECT 12025.08 189.04 12037.125 350.165 ;
      RECT 12025.08 211.445 12038.08 308.075 ;
      RECT 12025.08 189.04 12038.08 195.075 ;
      RECT 11994.56 324.445 12022.56 350.165 ;
      RECT 12020.705 189.04 12022.56 350.165 ;
      RECT 11994.56 228.445 12015.795 350.165 ;
      RECT 12018.115 189.04 12022.56 308.075 ;
      RECT 12001.11 211.445 12022.56 308.075 ;
      RECT 11994.56 189.04 12013.205 212.075 ;
      RECT 11994.56 189.04 12022.56 195.075 ;
      RECT 11979.04 290.445 11992.04 350.165 ;
      RECT 11991.425 194.42 11992.04 350.165 ;
      RECT 11979.04 189.04 11983.675 350.165 ;
      RECT 11979.04 194.42 11992.04 259.875 ;
      RECT 11979.04 189.04 11990.41 259.875 ;
      RECT 11979.04 189.04 11992.04 190.125 ;
      RECT 11962.06 211.445 11975.06 330.165 ;
      RECT 11965.425 189.04 11975.06 330.165 ;
      RECT 11962.06 189.04 11975.06 195.075 ;
      RECT 11945.08 259.445 11958.08 350.165 ;
      RECT 11946.935 189.04 11958.08 350.165 ;
      RECT 11945.08 189.04 11958.08 228.875 ;
      RECT 11914.56 307.445 11942.56 350.165 ;
      RECT 11929.035 259.445 11942.56 350.165 ;
      RECT 11914.56 189.04 11924.125 350.165 ;
      RECT 11914.56 228.445 11939.185 291.075 ;
      RECT 11933.09 189.04 11942.56 228.875 ;
      RECT 11929.035 194.37 11942.56 228.875 ;
      RECT 11914.56 194.37 11942.56 212.075 ;
      RECT 11914.56 189.04 11927.37 212.075 ;
      RECT 11914.56 189.04 11942.56 190.17 ;
      RECT 11899.04 324.445 11912.04 350.165 ;
      RECT 11906.705 189.04 11912.04 350.165 ;
      RECT 11902.035 307.445 11912.04 350.165 ;
      RECT 11899.04 307.445 11912.04 308.075 ;
      RECT 11899.04 211.445 11901.795 308.075 ;
      RECT 11899.04 228.445 11912.04 291.075 ;
      RECT 11899.04 211.445 11912.04 212.075 ;
      RECT 11902.035 189.04 11912.04 212.075 ;
      RECT 11899.04 189.04 11912.04 195.075 ;
      RECT 11865.08 324.445 11878.08 350.165 ;
      RECT 11865.08 228.445 11875.795 350.165 ;
      RECT 11870.31 211.445 11878.08 308.075 ;
      RECT 11865.08 189.04 11873.125 212.075 ;
      RECT 11865.08 189.04 11878.08 195.075 ;
      RECT 11834.56 290.445 11862.56 350.165 ;
      RECT 11853.19 189.04 11862.56 350.165 ;
      RECT 11851.425 194.425 11862.56 350.165 ;
      RECT 11834.56 189.04 11843.675 350.165 ;
      RECT 11834.56 194.425 11862.56 259.875 ;
      RECT 11834.56 189.04 11850.41 259.875 ;
      RECT 11834.56 189.04 11862.56 190.125 ;
      RECT 11819.04 211.445 11832.04 350.165 ;
      RECT 11825.425 189.04 11832.04 350.165 ;
      RECT 11819.04 189.04 11820.515 350.165 ;
      RECT 11819.04 189.04 11832.04 195.075 ;
      RECT 11802.06 259.445 11815.06 330.165 ;
      RECT 11806.935 189.04 11815.06 330.165 ;
      RECT 11802.06 189.04 11815.06 228.875 ;
      RECT 11785.08 307.445 11798.08 350.165 ;
      RECT 11793.09 189.04 11798.08 350.165 ;
      RECT 11789.035 194.37 11798.08 350.165 ;
      RECT 11785.08 228.445 11798.08 291.075 ;
      RECT 11785.08 194.37 11798.08 212.075 ;
      RECT 11785.08 189.04 11787.37 212.075 ;
      RECT 11785.08 189.04 11798.08 190.38 ;
      RECT 11754.56 324.445 11782.56 350.165 ;
      RECT 11766.705 189.04 11782.56 350.165 ;
      RECT 11762.035 307.445 11782.56 350.165 ;
      RECT 11754.56 189.04 11757.125 350.165 ;
      RECT 11754.56 307.445 11782.56 308.075 ;
      RECT 11754.56 211.445 11761.795 308.075 ;
      RECT 11754.56 228.445 11782.56 291.075 ;
      RECT 11754.56 211.445 11782.56 212.075 ;
      RECT 11762.035 189.04 11782.56 212.075 ;
      RECT 11754.56 189.04 11782.56 195.075 ;
      RECT 11739.04 324.445 11752.04 350.165 ;
      RECT 11740.705 189.04 11752.04 350.165 ;
      RECT 11739.04 189.04 11752.04 308.075 ;
      RECT 11722.06 228.445 11735.06 330.165 ;
      RECT 11728.69 211.445 11735.06 330.165 ;
      RECT 11722.06 189.04 11732.015 212.075 ;
      RECT 11722.06 189.04 11735.06 195.075 ;
      RECT 11705.08 290.445 11718.08 350.165 ;
      RECT 11713.19 189.04 11718.08 350.165 ;
      RECT 11711.425 194.425 11718.08 350.165 ;
      RECT 11705.08 194.425 11718.08 259.875 ;
      RECT 11705.08 189.04 11710.41 259.875 ;
      RECT 11705.08 189.04 11718.08 190.125 ;
      RECT 11674.56 211.445 11702.56 350.165 ;
      RECT 11685.425 189.04 11702.56 350.165 ;
      RECT 11674.56 189.04 11680.515 350.165 ;
      RECT 11674.56 189.04 11702.56 195.075 ;
      RECT 11659.04 259.445 11672.04 350.165 ;
      RECT 11666.935 189.04 11672.04 350.165 ;
      RECT 11659.04 189.04 11672.04 228.875 ;
      RECT 11642.06 307.445 11655.06 330.165 ;
      RECT 11652.99 189.04 11655.06 330.165 ;
      RECT 11649.035 194.37 11655.06 330.165 ;
      RECT 11642.06 189.04 11644.125 330.165 ;
      RECT 11642.06 228.445 11655.06 291.075 ;
      RECT 11642.06 194.37 11655.06 212.075 ;
      RECT 11642.06 189.04 11647.37 212.075 ;
      RECT 11642.06 189.04 11655.06 190.17 ;
      RECT 11625.08 307.445 11638.08 350.165 ;
      RECT 11626.705 189.04 11638.08 350.165 ;
      RECT 11625.08 228.445 11638.08 291.075 ;
      RECT 11625.08 189.04 11638.08 212.075 ;
      RECT 11594.56 324.445 11622.56 350.165 ;
      RECT 11600.705 189.04 11617.125 350.165 ;
      RECT 11594.56 211.445 11595.795 350.165 ;
      RECT 11594.56 211.445 11621.795 308.075 ;
      RECT 11594.56 228.445 11622.56 291.075 ;
      RECT 11596.925 189.04 11617.125 308.075 ;
      RECT 11594.56 189.04 11622.56 195.075 ;
      RECT 11579.04 228.445 11592.04 350.165 ;
      RECT 11579.04 189.04 11585.395 350.165 ;
      RECT 11579.04 189.04 11592.04 212.075 ;
      RECT 11562.06 290.445 11575.06 330.165 ;
      RECT 11573.19 189.04 11575.06 330.165 ;
      RECT 11571.425 194.425 11575.06 330.165 ;
      RECT 11562.06 189.04 11563.675 330.165 ;
      RECT 11562.06 194.425 11575.06 259.875 ;
      RECT 11562.06 189.04 11570.41 259.875 ;
      RECT 11562.06 189.04 11575.06 190.125 ;
      RECT 11545.08 211.445 11558.08 350.165 ;
      RECT 11545.425 189.04 11558.08 350.165 ;
      RECT 11545.08 189.04 11558.08 195.075 ;
      RECT 11514.56 259.445 11542.56 350.165 ;
      RECT 11526.935 211.445 11542.56 350.165 ;
      RECT 11514.56 189.04 11519.185 350.165 ;
      RECT 11514.56 189.04 11540.515 228.875 ;
      RECT 11514.56 189.04 11542.56 195.075 ;
      RECT 11499.04 307.445 11512.04 350.165 ;
      RECT 11509.035 194.37 11512.04 350.165 ;
      RECT 11499.04 189.04 11504.125 350.165 ;
      RECT 11499.04 228.445 11512.04 291.075 ;
      RECT 11499.04 194.37 11512.04 212.075 ;
      RECT 11499.04 189.04 11507.37 212.075 ;
      RECT 11499.04 189.04 11512.04 190.17 ;
      RECT 11482.06 307.445 11495.06 330.165 ;
      RECT 11486.705 189.04 11495.06 330.165 ;
      RECT 11486.54 228.445 11495.06 330.165 ;
      RECT 11482.06 228.445 11495.06 291.075 ;
      RECT 11482.06 189.04 11495.06 212.075 ;
      RECT 11465.08 324.445 11478.08 350.165 ;
      RECT 11465.08 189.04 11477.125 350.165 ;
      RECT 11465.08 211.445 11478.08 308.075 ;
      RECT 11465.08 189.04 11478.08 195.075 ;
      RECT 11434.56 324.445 11462.56 350.165 ;
      RECT 11460.705 189.04 11462.56 350.165 ;
      RECT 11434.56 228.445 11455.795 350.165 ;
      RECT 11458.115 189.04 11462.56 308.075 ;
      RECT 11441.11 211.445 11462.56 308.075 ;
      RECT 11434.56 189.04 11453.205 212.075 ;
      RECT 11434.56 189.04 11462.56 195.075 ;
      RECT 11419.04 290.445 11432.04 350.165 ;
      RECT 11431.425 194.42 11432.04 350.165 ;
      RECT 11419.04 189.04 11423.675 350.165 ;
      RECT 11419.04 194.42 11432.04 259.875 ;
      RECT 11419.04 189.04 11430.41 259.875 ;
      RECT 11419.04 189.04 11432.04 190.125 ;
      RECT 11402.06 211.445 11415.06 330.165 ;
      RECT 11405.425 189.04 11415.06 330.165 ;
      RECT 11402.06 189.04 11415.06 195.075 ;
      RECT 11385.08 259.445 11398.08 350.165 ;
      RECT 11386.935 189.04 11398.08 350.165 ;
      RECT 11385.08 189.04 11398.08 228.875 ;
      RECT 11354.56 307.445 11382.56 350.165 ;
      RECT 11369.035 259.445 11382.56 350.165 ;
      RECT 11354.56 189.04 11364.125 350.165 ;
      RECT 11354.56 228.445 11379.185 291.075 ;
      RECT 11373.09 189.04 11382.56 228.875 ;
      RECT 11369.035 194.37 11382.56 228.875 ;
      RECT 11354.56 194.37 11382.56 212.075 ;
      RECT 11354.56 189.04 11367.37 212.075 ;
      RECT 11354.56 189.04 11382.56 190.17 ;
      RECT 11339.04 324.445 11352.04 350.165 ;
      RECT 11346.705 189.04 11352.04 350.165 ;
      RECT 11342.035 307.445 11352.04 350.165 ;
      RECT 11339.04 307.445 11352.04 308.075 ;
      RECT 11339.04 211.445 11341.795 308.075 ;
      RECT 11339.04 228.445 11352.04 291.075 ;
      RECT 11339.04 211.445 11352.04 212.075 ;
      RECT 11342.035 189.04 11352.04 212.075 ;
      RECT 11339.04 189.04 11352.04 195.075 ;
      RECT 11305.08 324.445 11318.08 350.165 ;
      RECT 11305.08 228.445 11315.795 350.165 ;
      RECT 11310.31 211.445 11318.08 308.075 ;
      RECT 11305.08 189.04 11313.125 212.075 ;
      RECT 11305.08 189.04 11318.08 195.075 ;
      RECT 11274.56 290.445 11302.56 350.165 ;
      RECT 11293.19 189.04 11302.56 350.165 ;
      RECT 11291.425 194.425 11302.56 350.165 ;
      RECT 11274.56 189.04 11283.675 350.165 ;
      RECT 11274.56 194.425 11302.56 259.875 ;
      RECT 11274.56 189.04 11290.41 259.875 ;
      RECT 11274.56 189.04 11302.56 190.125 ;
      RECT 11259.04 211.445 11272.04 350.165 ;
      RECT 11265.425 189.04 11272.04 350.165 ;
      RECT 11259.04 189.04 11260.515 350.165 ;
      RECT 11259.04 189.04 11272.04 195.075 ;
      RECT 11242.06 259.445 11255.06 330.165 ;
      RECT 11246.935 189.04 11255.06 330.165 ;
      RECT 11242.06 189.04 11255.06 228.875 ;
      RECT 11225.08 307.445 11238.08 350.165 ;
      RECT 11233.09 189.04 11238.08 350.165 ;
      RECT 11229.035 194.37 11238.08 350.165 ;
      RECT 11225.08 228.445 11238.08 291.075 ;
      RECT 11225.08 194.37 11238.08 212.075 ;
      RECT 11225.08 189.04 11227.37 212.075 ;
      RECT 11225.08 189.04 11238.08 190.38 ;
      RECT 11194.56 324.445 11222.56 350.165 ;
      RECT 11206.705 189.04 11222.56 350.165 ;
      RECT 11202.035 307.445 11222.56 350.165 ;
      RECT 11194.56 189.04 11197.125 350.165 ;
      RECT 11194.56 307.445 11222.56 308.075 ;
      RECT 11194.56 211.445 11201.795 308.075 ;
      RECT 11194.56 228.445 11222.56 291.075 ;
      RECT 11194.56 211.445 11222.56 212.075 ;
      RECT 11202.035 189.04 11222.56 212.075 ;
      RECT 11194.56 189.04 11222.56 195.075 ;
      RECT 11179.04 324.445 11192.04 350.165 ;
      RECT 11180.705 189.04 11192.04 350.165 ;
      RECT 11179.04 189.04 11192.04 308.075 ;
      RECT 11162.06 228.445 11175.06 330.165 ;
      RECT 11168.69 211.445 11175.06 330.165 ;
      RECT 11162.06 189.04 11172.015 212.075 ;
      RECT 11162.06 189.04 11175.06 195.075 ;
      RECT 11145.08 290.445 11158.08 350.165 ;
      RECT 11153.19 189.04 11158.08 350.165 ;
      RECT 11151.425 194.425 11158.08 350.165 ;
      RECT 11145.08 194.425 11158.08 259.875 ;
      RECT 11145.08 189.04 11150.41 259.875 ;
      RECT 11145.08 189.04 11158.08 190.125 ;
      RECT 11114.56 211.445 11142.56 350.165 ;
      RECT 11125.425 189.04 11142.56 350.165 ;
      RECT 11114.56 189.04 11120.515 350.165 ;
      RECT 11114.56 189.04 11142.56 195.075 ;
      RECT 11099.04 259.445 11112.04 350.165 ;
      RECT 11106.935 189.04 11112.04 350.165 ;
      RECT 11099.04 189.04 11112.04 228.875 ;
      RECT 11082.06 307.445 11095.06 330.165 ;
      RECT 11092.99 189.04 11095.06 330.165 ;
      RECT 11089.035 194.37 11095.06 330.165 ;
      RECT 11082.06 189.04 11084.125 330.165 ;
      RECT 11082.06 228.445 11095.06 291.075 ;
      RECT 11082.06 194.37 11095.06 212.075 ;
      RECT 11082.06 189.04 11087.37 212.075 ;
      RECT 11082.06 189.04 11095.06 190.17 ;
      RECT 11065.08 307.445 11078.08 350.165 ;
      RECT 11066.705 189.04 11078.08 350.165 ;
      RECT 11065.08 228.445 11078.08 291.075 ;
      RECT 11065.08 189.04 11078.08 212.075 ;
      RECT 11034.56 324.445 11062.56 350.165 ;
      RECT 11040.705 189.04 11057.125 350.165 ;
      RECT 11034.56 211.445 11035.795 350.165 ;
      RECT 11034.56 211.445 11061.795 308.075 ;
      RECT 11034.56 228.445 11062.56 291.075 ;
      RECT 11036.925 189.04 11057.125 308.075 ;
      RECT 11034.56 189.04 11062.56 195.075 ;
      RECT 11019.04 228.445 11032.04 350.165 ;
      RECT 11019.04 189.04 11025.395 350.165 ;
      RECT 11019.04 189.04 11032.04 212.075 ;
      RECT 11002.06 290.445 11015.06 330.165 ;
      RECT 11013.19 189.04 11015.06 330.165 ;
      RECT 11011.425 194.425 11015.06 330.165 ;
      RECT 11002.06 189.04 11003.675 330.165 ;
      RECT 11002.06 194.425 11015.06 259.875 ;
      RECT 11002.06 189.04 11010.41 259.875 ;
      RECT 11002.06 189.04 11015.06 190.125 ;
      RECT 10985.08 211.445 10998.08 350.165 ;
      RECT 10985.425 189.04 10998.08 350.165 ;
      RECT 10985.08 189.04 10998.08 195.075 ;
      RECT 10954.56 259.445 10982.56 350.165 ;
      RECT 10966.935 211.445 10982.56 350.165 ;
      RECT 10954.56 189.04 10959.185 350.165 ;
      RECT 10954.56 189.04 10980.515 228.875 ;
      RECT 10954.56 189.04 10982.56 195.075 ;
      RECT 10939.04 307.445 10952.04 350.165 ;
      RECT 10949.035 194.37 10952.04 350.165 ;
      RECT 10939.04 189.04 10944.125 350.165 ;
      RECT 10939.04 228.445 10952.04 291.075 ;
      RECT 10939.04 194.37 10952.04 212.075 ;
      RECT 10939.04 189.04 10947.37 212.075 ;
      RECT 10939.04 189.04 10952.04 190.17 ;
      RECT 10922.06 307.445 10935.06 330.165 ;
      RECT 10926.705 189.04 10935.06 330.165 ;
      RECT 10926.54 228.445 10935.06 330.165 ;
      RECT 10922.06 228.445 10935.06 291.075 ;
      RECT 10922.06 189.04 10935.06 212.075 ;
      RECT 10905.08 324.445 10918.08 350.165 ;
      RECT 10905.08 189.04 10917.125 350.165 ;
      RECT 10905.08 211.445 10918.08 308.075 ;
      RECT 10905.08 189.04 10918.08 195.075 ;
      RECT 10874.56 324.445 10902.56 350.165 ;
      RECT 10900.705 189.04 10902.56 350.165 ;
      RECT 10874.56 228.445 10895.795 350.165 ;
      RECT 10898.115 189.04 10902.56 308.075 ;
      RECT 10881.11 211.445 10902.56 308.075 ;
      RECT 10874.56 189.04 10893.205 212.075 ;
      RECT 10874.56 189.04 10902.56 195.075 ;
      RECT 10859.04 290.445 10872.04 350.165 ;
      RECT 10871.425 194.42 10872.04 350.165 ;
      RECT 10859.04 189.04 10863.675 350.165 ;
      RECT 10859.04 194.42 10872.04 259.875 ;
      RECT 10859.04 189.04 10870.41 259.875 ;
      RECT 10859.04 189.04 10872.04 190.125 ;
      RECT 10842.06 211.445 10855.06 330.165 ;
      RECT 10845.425 189.04 10855.06 330.165 ;
      RECT 10842.06 189.04 10855.06 195.075 ;
      RECT 10825.08 259.445 10838.08 350.165 ;
      RECT 10826.935 189.04 10838.08 350.165 ;
      RECT 10825.08 189.04 10838.08 228.875 ;
      RECT 10794.56 307.445 10822.56 350.165 ;
      RECT 10809.035 259.445 10822.56 350.165 ;
      RECT 10794.56 189.04 10804.125 350.165 ;
      RECT 10794.56 228.445 10819.185 291.075 ;
      RECT 10813.09 189.04 10822.56 228.875 ;
      RECT 10809.035 194.37 10822.56 228.875 ;
      RECT 10794.56 194.37 10822.56 212.075 ;
      RECT 10794.56 189.04 10807.37 212.075 ;
      RECT 10794.56 189.04 10822.56 190.17 ;
      RECT 10779.04 324.445 10792.04 350.165 ;
      RECT 10786.705 189.04 10792.04 350.165 ;
      RECT 10782.035 307.445 10792.04 350.165 ;
      RECT 10779.04 307.445 10792.04 308.075 ;
      RECT 10779.04 211.445 10781.795 308.075 ;
      RECT 10779.04 228.445 10792.04 291.075 ;
      RECT 10779.04 211.445 10792.04 212.075 ;
      RECT 10782.035 189.04 10792.04 212.075 ;
      RECT 10779.04 189.04 10792.04 195.075 ;
      RECT 10745.08 324.445 10758.08 350.165 ;
      RECT 10745.08 228.445 10755.795 350.165 ;
      RECT 10750.31 211.445 10758.08 308.075 ;
      RECT 10745.08 189.04 10753.125 212.075 ;
      RECT 10745.08 189.04 10758.08 195.075 ;
      RECT 10714.56 290.445 10742.56 350.165 ;
      RECT 10733.19 189.04 10742.56 350.165 ;
      RECT 10731.425 194.425 10742.56 350.165 ;
      RECT 10714.56 189.04 10723.675 350.165 ;
      RECT 10714.56 194.425 10742.56 259.875 ;
      RECT 10714.56 189.04 10730.41 259.875 ;
      RECT 10714.56 189.04 10742.56 190.125 ;
      RECT 10699.04 211.445 10712.04 350.165 ;
      RECT 10705.425 189.04 10712.04 350.165 ;
      RECT 10699.04 189.04 10700.515 350.165 ;
      RECT 10699.04 189.04 10712.04 195.075 ;
      RECT 10682.06 259.445 10695.06 330.165 ;
      RECT 10686.935 189.04 10695.06 330.165 ;
      RECT 10682.06 189.04 10695.06 228.875 ;
      RECT 10665.08 307.445 10678.08 350.165 ;
      RECT 10673.09 189.04 10678.08 350.165 ;
      RECT 10669.035 194.37 10678.08 350.165 ;
      RECT 10665.08 228.445 10678.08 291.075 ;
      RECT 10665.08 194.37 10678.08 212.075 ;
      RECT 10665.08 189.04 10667.37 212.075 ;
      RECT 10665.08 189.04 10678.08 190.38 ;
      RECT 10634.56 324.445 10662.56 350.165 ;
      RECT 10646.705 189.04 10662.56 350.165 ;
      RECT 10642.035 307.445 10662.56 350.165 ;
      RECT 10634.56 189.04 10637.125 350.165 ;
      RECT 10634.56 307.445 10662.56 308.075 ;
      RECT 10634.56 211.445 10641.795 308.075 ;
      RECT 10634.56 228.445 10662.56 291.075 ;
      RECT 10634.56 211.445 10662.56 212.075 ;
      RECT 10642.035 189.04 10662.56 212.075 ;
      RECT 10634.56 189.04 10662.56 195.075 ;
      RECT 10619.04 324.445 10632.04 350.165 ;
      RECT 10620.705 189.04 10632.04 350.165 ;
      RECT 10619.04 189.04 10632.04 308.075 ;
      RECT 10602.06 228.445 10615.06 330.165 ;
      RECT 10608.69 211.445 10615.06 330.165 ;
      RECT 10602.06 189.04 10612.015 212.075 ;
      RECT 10602.06 189.04 10615.06 195.075 ;
      RECT 10585.08 290.445 10598.08 350.165 ;
      RECT 10593.19 189.04 10598.08 350.165 ;
      RECT 10591.425 194.425 10598.08 350.165 ;
      RECT 10585.08 194.425 10598.08 259.875 ;
      RECT 10585.08 189.04 10590.41 259.875 ;
      RECT 10585.08 189.04 10598.08 190.125 ;
      RECT 10554.56 211.445 10582.56 350.165 ;
      RECT 10565.425 189.04 10582.56 350.165 ;
      RECT 10554.56 189.04 10560.515 350.165 ;
      RECT 10554.56 189.04 10582.56 195.075 ;
      RECT 10539.04 259.445 10552.04 350.165 ;
      RECT 10546.935 189.04 10552.04 350.165 ;
      RECT 10539.04 189.04 10552.04 228.875 ;
      RECT 10522.06 307.445 10535.06 330.165 ;
      RECT 10532.99 189.04 10535.06 330.165 ;
      RECT 10529.035 194.37 10535.06 330.165 ;
      RECT 10522.06 189.04 10524.125 330.165 ;
      RECT 10522.06 228.445 10535.06 291.075 ;
      RECT 10522.06 194.37 10535.06 212.075 ;
      RECT 10522.06 189.04 10527.37 212.075 ;
      RECT 10522.06 189.04 10535.06 190.17 ;
      RECT 10505.08 307.445 10518.08 350.165 ;
      RECT 10506.705 189.04 10518.08 350.165 ;
      RECT 10505.08 228.445 10518.08 291.075 ;
      RECT 10505.08 189.04 10518.08 212.075 ;
      RECT 10474.56 324.445 10502.56 350.165 ;
      RECT 10480.705 189.04 10497.125 350.165 ;
      RECT 10474.56 211.445 10475.795 350.165 ;
      RECT 10474.56 211.445 10501.795 308.075 ;
      RECT 10474.56 228.445 10502.56 291.075 ;
      RECT 10476.925 189.04 10497.125 308.075 ;
      RECT 10474.56 189.04 10502.56 195.075 ;
      RECT 10459.04 228.445 10472.04 350.165 ;
      RECT 10459.04 189.04 10465.395 350.165 ;
      RECT 10459.04 189.04 10472.04 212.075 ;
      RECT 10442.06 290.445 10455.06 330.165 ;
      RECT 10453.19 189.04 10455.06 330.165 ;
      RECT 10451.425 194.425 10455.06 330.165 ;
      RECT 10442.06 189.04 10443.675 330.165 ;
      RECT 10442.06 194.425 10455.06 259.875 ;
      RECT 10442.06 189.04 10450.41 259.875 ;
      RECT 10442.06 189.04 10455.06 190.125 ;
      RECT 10425.08 211.445 10438.08 350.165 ;
      RECT 10425.425 189.04 10438.08 350.165 ;
      RECT 10425.08 189.04 10438.08 195.075 ;
      RECT 10394.56 259.445 10422.56 350.165 ;
      RECT 10406.935 211.445 10422.56 350.165 ;
      RECT 10394.56 189.04 10399.185 350.165 ;
      RECT 10394.56 189.04 10420.515 228.875 ;
      RECT 10394.56 189.04 10422.56 195.075 ;
      RECT 10379.04 307.445 10392.04 350.165 ;
      RECT 10389.035 194.37 10392.04 350.165 ;
      RECT 10379.04 189.04 10384.125 350.165 ;
      RECT 10379.04 228.445 10392.04 291.075 ;
      RECT 10379.04 194.37 10392.04 212.075 ;
      RECT 10379.04 189.04 10387.37 212.075 ;
      RECT 10379.04 189.04 10392.04 190.17 ;
      RECT 10362.06 307.445 10375.06 330.165 ;
      RECT 10366.705 189.04 10375.06 330.165 ;
      RECT 10366.54 228.445 10375.06 330.165 ;
      RECT 10362.06 228.445 10375.06 291.075 ;
      RECT 10362.06 189.04 10375.06 212.075 ;
      RECT 10345.08 324.445 10358.08 350.165 ;
      RECT 10345.08 189.04 10357.125 350.165 ;
      RECT 10345.08 211.445 10358.08 308.075 ;
      RECT 10345.08 189.04 10358.08 195.075 ;
      RECT 10314.56 324.445 10342.56 350.165 ;
      RECT 10340.705 189.04 10342.56 350.165 ;
      RECT 10314.56 228.445 10335.795 350.165 ;
      RECT 10338.115 189.04 10342.56 308.075 ;
      RECT 10321.11 211.445 10342.56 308.075 ;
      RECT 10314.56 189.04 10333.205 212.075 ;
      RECT 10314.56 189.04 10342.56 195.075 ;
      RECT 10299.04 290.445 10312.04 350.165 ;
      RECT 10311.425 194.42 10312.04 350.165 ;
      RECT 10299.04 189.04 10303.675 350.165 ;
      RECT 10299.04 194.42 10312.04 259.875 ;
      RECT 10299.04 189.04 10310.41 259.875 ;
      RECT 10299.04 189.04 10312.04 190.125 ;
      RECT 10282.06 211.445 10295.06 330.165 ;
      RECT 10285.425 189.04 10295.06 330.165 ;
      RECT 10282.06 189.04 10295.06 195.075 ;
      RECT 10265.08 259.445 10278.08 350.165 ;
      RECT 10266.935 189.04 10278.08 350.165 ;
      RECT 10265.08 189.04 10278.08 228.875 ;
      RECT 10234.56 307.445 10262.56 350.165 ;
      RECT 10249.035 259.445 10262.56 350.165 ;
      RECT 10234.56 189.04 10244.125 350.165 ;
      RECT 10234.56 228.445 10259.185 291.075 ;
      RECT 10253.09 189.04 10262.56 228.875 ;
      RECT 10249.035 194.37 10262.56 228.875 ;
      RECT 10234.56 194.37 10262.56 212.075 ;
      RECT 10234.56 189.04 10247.37 212.075 ;
      RECT 10234.56 189.04 10262.56 190.17 ;
      RECT 10219.04 324.445 10232.04 350.165 ;
      RECT 10226.705 189.04 10232.04 350.165 ;
      RECT 10222.035 307.445 10232.04 350.165 ;
      RECT 10219.04 307.445 10232.04 308.075 ;
      RECT 10219.04 211.445 10221.795 308.075 ;
      RECT 10219.04 228.445 10232.04 291.075 ;
      RECT 10219.04 211.445 10232.04 212.075 ;
      RECT 10222.035 189.04 10232.04 212.075 ;
      RECT 10219.04 189.04 10232.04 195.075 ;
      RECT 10185.08 324.445 10198.08 350.165 ;
      RECT 10185.08 228.445 10195.795 350.165 ;
      RECT 10190.31 211.445 10198.08 308.075 ;
      RECT 10185.08 189.04 10193.125 212.075 ;
      RECT 10185.08 189.04 10198.08 195.075 ;
      RECT 10154.56 290.445 10182.56 350.165 ;
      RECT 10173.19 189.04 10182.56 350.165 ;
      RECT 10171.425 194.425 10182.56 350.165 ;
      RECT 10154.56 189.04 10163.675 350.165 ;
      RECT 10154.56 194.425 10182.56 259.875 ;
      RECT 10154.56 189.04 10170.41 259.875 ;
      RECT 10154.56 189.04 10182.56 190.125 ;
      RECT 10139.04 211.445 10152.04 350.165 ;
      RECT 10145.425 189.04 10152.04 350.165 ;
      RECT 10139.04 189.04 10140.515 350.165 ;
      RECT 10139.04 189.04 10152.04 195.075 ;
      RECT 10122.06 259.445 10135.06 330.165 ;
      RECT 10126.935 189.04 10135.06 330.165 ;
      RECT 10122.06 189.04 10135.06 228.875 ;
      RECT 10105.08 307.445 10118.08 350.165 ;
      RECT 10113.09 189.04 10118.08 350.165 ;
      RECT 10109.035 194.37 10118.08 350.165 ;
      RECT 10105.08 228.445 10118.08 291.075 ;
      RECT 10105.08 194.37 10118.08 212.075 ;
      RECT 10105.08 189.04 10107.37 212.075 ;
      RECT 10105.08 189.04 10118.08 190.38 ;
      RECT 10074.56 324.445 10102.56 350.165 ;
      RECT 10086.705 189.04 10102.56 350.165 ;
      RECT 10082.035 307.445 10102.56 350.165 ;
      RECT 10074.56 189.04 10077.125 350.165 ;
      RECT 10074.56 307.445 10102.56 308.075 ;
      RECT 10074.56 211.445 10081.795 308.075 ;
      RECT 10074.56 228.445 10102.56 291.075 ;
      RECT 10074.56 211.445 10102.56 212.075 ;
      RECT 10082.035 189.04 10102.56 212.075 ;
      RECT 10074.56 189.04 10102.56 195.075 ;
      RECT 10059.04 324.445 10072.04 350.165 ;
      RECT 10060.705 189.04 10072.04 350.165 ;
      RECT 10059.04 189.04 10072.04 308.075 ;
      RECT 10042.06 228.445 10055.06 330.165 ;
      RECT 10048.69 211.445 10055.06 330.165 ;
      RECT 10042.06 189.04 10052.015 212.075 ;
      RECT 10042.06 189.04 10055.06 195.075 ;
      RECT 10025.08 290.445 10038.08 350.165 ;
      RECT 10033.19 189.04 10038.08 350.165 ;
      RECT 10031.425 194.425 10038.08 350.165 ;
      RECT 10025.08 194.425 10038.08 259.875 ;
      RECT 10025.08 189.04 10030.41 259.875 ;
      RECT 10025.08 189.04 10038.08 190.125 ;
      RECT 9994.56 211.445 10022.56 350.165 ;
      RECT 10005.425 189.04 10022.56 350.165 ;
      RECT 9994.56 189.04 10000.515 350.165 ;
      RECT 9994.56 189.04 10022.56 195.075 ;
      RECT 9979.04 259.445 9992.04 350.165 ;
      RECT 9986.935 189.04 9992.04 350.165 ;
      RECT 9979.04 189.04 9992.04 228.875 ;
      RECT 9962.06 307.445 9975.06 330.165 ;
      RECT 9972.99 189.04 9975.06 330.165 ;
      RECT 9969.035 194.37 9975.06 330.165 ;
      RECT 9962.06 189.04 9964.125 330.165 ;
      RECT 9962.06 228.445 9975.06 291.075 ;
      RECT 9962.06 194.37 9975.06 212.075 ;
      RECT 9962.06 189.04 9967.37 212.075 ;
      RECT 9962.06 189.04 9975.06 190.17 ;
      RECT 9945.08 307.445 9958.08 350.165 ;
      RECT 9946.705 189.04 9958.08 350.165 ;
      RECT 9945.08 228.445 9958.08 291.075 ;
      RECT 9945.08 189.04 9958.08 212.075 ;
      RECT 9914.56 324.445 9942.56 350.165 ;
      RECT 9920.705 189.04 9937.125 350.165 ;
      RECT 9914.56 211.445 9915.795 350.165 ;
      RECT 9914.56 211.445 9941.795 308.075 ;
      RECT 9914.56 228.445 9942.56 291.075 ;
      RECT 9916.925 189.04 9937.125 308.075 ;
      RECT 9914.56 189.04 9942.56 195.075 ;
      RECT 9899.04 228.445 9912.04 350.165 ;
      RECT 9899.04 189.04 9905.395 350.165 ;
      RECT 9899.04 189.04 9912.04 212.075 ;
      RECT 9882.06 290.445 9895.06 330.165 ;
      RECT 9893.19 189.04 9895.06 330.165 ;
      RECT 9891.425 194.425 9895.06 330.165 ;
      RECT 9882.06 189.04 9883.675 330.165 ;
      RECT 9882.06 194.425 9895.06 259.875 ;
      RECT 9882.06 189.04 9890.41 259.875 ;
      RECT 9882.06 189.04 9895.06 190.125 ;
      RECT 9865.08 211.445 9878.08 350.165 ;
      RECT 9865.425 189.04 9878.08 350.165 ;
      RECT 9865.08 189.04 9878.08 195.075 ;
      RECT 9834.56 259.445 9862.56 350.165 ;
      RECT 9846.935 211.445 9862.56 350.165 ;
      RECT 9834.56 189.04 9839.185 350.165 ;
      RECT 9834.56 189.04 9860.515 228.875 ;
      RECT 9834.56 189.04 9862.56 195.075 ;
      RECT 9819.04 307.445 9832.04 350.165 ;
      RECT 9829.035 194.37 9832.04 350.165 ;
      RECT 9819.04 189.04 9824.125 350.165 ;
      RECT 9819.04 228.445 9832.04 291.075 ;
      RECT 9819.04 194.37 9832.04 212.075 ;
      RECT 9819.04 189.04 9827.37 212.075 ;
      RECT 9819.04 189.04 9832.04 190.17 ;
      RECT 9802.06 307.445 9815.06 330.165 ;
      RECT 9806.705 189.04 9815.06 330.165 ;
      RECT 9806.54 228.445 9815.06 330.165 ;
      RECT 9802.06 228.445 9815.06 291.075 ;
      RECT 9802.06 189.04 9815.06 212.075 ;
      RECT 9785.08 324.445 9798.08 350.165 ;
      RECT 9785.08 189.04 9797.125 350.165 ;
      RECT 9785.08 211.445 9798.08 308.075 ;
      RECT 9785.08 189.04 9798.08 195.075 ;
      RECT 9754.56 324.445 9782.56 350.165 ;
      RECT 9780.705 189.04 9782.56 350.165 ;
      RECT 9754.56 228.445 9775.795 350.165 ;
      RECT 9778.115 189.04 9782.56 308.075 ;
      RECT 9761.11 211.445 9782.56 308.075 ;
      RECT 9754.56 189.04 9773.205 212.075 ;
      RECT 9754.56 189.04 9782.56 195.075 ;
      RECT 9739.04 290.445 9752.04 350.165 ;
      RECT 9751.425 194.42 9752.04 350.165 ;
      RECT 9739.04 189.04 9743.675 350.165 ;
      RECT 9739.04 194.42 9752.04 259.875 ;
      RECT 9739.04 189.04 9750.41 259.875 ;
      RECT 9739.04 189.04 9752.04 190.125 ;
      RECT 9722.06 211.445 9735.06 330.165 ;
      RECT 9725.425 189.04 9735.06 330.165 ;
      RECT 9722.06 189.04 9735.06 195.075 ;
      RECT 9705.08 259.445 9718.08 350.165 ;
      RECT 9706.935 189.04 9718.08 350.165 ;
      RECT 9705.08 189.04 9718.08 228.875 ;
      RECT 9674.56 307.445 9702.56 350.165 ;
      RECT 9689.035 259.445 9702.56 350.165 ;
      RECT 9674.56 189.04 9684.125 350.165 ;
      RECT 9674.56 228.445 9699.185 291.075 ;
      RECT 9693.09 189.04 9702.56 228.875 ;
      RECT 9689.035 194.37 9702.56 228.875 ;
      RECT 9674.56 194.37 9702.56 212.075 ;
      RECT 9674.56 189.04 9687.37 212.075 ;
      RECT 9674.56 189.04 9702.56 190.17 ;
      RECT 9659.04 324.445 9672.04 350.165 ;
      RECT 9666.705 189.04 9672.04 350.165 ;
      RECT 9662.035 307.445 9672.04 350.165 ;
      RECT 9659.04 307.445 9672.04 308.075 ;
      RECT 9659.04 211.445 9661.795 308.075 ;
      RECT 9659.04 228.445 9672.04 291.075 ;
      RECT 9659.04 211.445 9672.04 212.075 ;
      RECT 9662.035 189.04 9672.04 212.075 ;
      RECT 9659.04 189.04 9672.04 195.075 ;
      RECT 9625.08 324.445 9638.08 350.165 ;
      RECT 9625.08 228.445 9635.795 350.165 ;
      RECT 9630.31 211.445 9638.08 308.075 ;
      RECT 9625.08 189.04 9633.125 212.075 ;
      RECT 9625.08 189.04 9638.08 195.075 ;
      RECT 9594.56 290.445 9622.56 350.165 ;
      RECT 9613.19 189.04 9622.56 350.165 ;
      RECT 9611.425 194.425 9622.56 350.165 ;
      RECT 9594.56 189.04 9603.675 350.165 ;
      RECT 9594.56 194.425 9622.56 259.875 ;
      RECT 9594.56 189.04 9610.41 259.875 ;
      RECT 9594.56 189.04 9622.56 190.125 ;
      RECT 9579.04 211.445 9592.04 350.165 ;
      RECT 9585.425 189.04 9592.04 350.165 ;
      RECT 9579.04 189.04 9580.515 350.165 ;
      RECT 9579.04 189.04 9592.04 195.075 ;
      RECT 9562.06 259.445 9575.06 330.165 ;
      RECT 9566.935 189.04 9575.06 330.165 ;
      RECT 9562.06 189.04 9575.06 228.875 ;
      RECT 9545.08 307.445 9558.08 350.165 ;
      RECT 9553.09 189.04 9558.08 350.165 ;
      RECT 9549.035 194.37 9558.08 350.165 ;
      RECT 9545.08 228.445 9558.08 291.075 ;
      RECT 9545.08 194.37 9558.08 212.075 ;
      RECT 9545.08 189.04 9547.37 212.075 ;
      RECT 9545.08 189.04 9558.08 190.38 ;
      RECT 9514.56 324.445 9542.56 350.165 ;
      RECT 9526.705 189.04 9542.56 350.165 ;
      RECT 9522.035 307.445 9542.56 350.165 ;
      RECT 9514.56 189.04 9517.125 350.165 ;
      RECT 9514.56 307.445 9542.56 308.075 ;
      RECT 9514.56 211.445 9521.795 308.075 ;
      RECT 9514.56 228.445 9542.56 291.075 ;
      RECT 9514.56 211.445 9542.56 212.075 ;
      RECT 9522.035 189.04 9542.56 212.075 ;
      RECT 9514.56 189.04 9542.56 195.075 ;
      RECT 9499.04 324.445 9512.04 350.165 ;
      RECT 9500.705 189.04 9512.04 350.165 ;
      RECT 9499.04 189.04 9512.04 308.075 ;
      RECT 9482.06 228.445 9495.06 330.165 ;
      RECT 9488.69 211.445 9495.06 330.165 ;
      RECT 9482.06 189.04 9492.015 212.075 ;
      RECT 9482.06 189.04 9495.06 195.075 ;
      RECT 9465.08 290.445 9478.08 350.165 ;
      RECT 9473.19 189.04 9478.08 350.165 ;
      RECT 9471.425 194.425 9478.08 350.165 ;
      RECT 9465.08 194.425 9478.08 259.875 ;
      RECT 9465.08 189.04 9470.41 259.875 ;
      RECT 9465.08 189.04 9478.08 190.125 ;
      RECT 9434.56 211.445 9462.56 350.165 ;
      RECT 9445.425 189.04 9462.56 350.165 ;
      RECT 9434.56 189.04 9440.515 350.165 ;
      RECT 9434.56 189.04 9462.56 195.075 ;
      RECT 9419.04 259.445 9432.04 350.165 ;
      RECT 9426.935 189.04 9432.04 350.165 ;
      RECT 9419.04 189.04 9432.04 228.875 ;
      RECT 9402.06 307.445 9415.06 330.165 ;
      RECT 9412.99 189.04 9415.06 330.165 ;
      RECT 9409.035 194.37 9415.06 330.165 ;
      RECT 9402.06 189.04 9404.125 330.165 ;
      RECT 9402.06 228.445 9415.06 291.075 ;
      RECT 9402.06 194.37 9415.06 212.075 ;
      RECT 9402.06 189.04 9407.37 212.075 ;
      RECT 9402.06 189.04 9415.06 190.17 ;
      RECT 9385.08 307.445 9398.08 350.165 ;
      RECT 9386.705 189.04 9398.08 350.165 ;
      RECT 9385.08 228.445 9398.08 291.075 ;
      RECT 9385.08 189.04 9398.08 212.075 ;
      RECT 9354.56 324.445 9382.56 350.165 ;
      RECT 9360.705 189.04 9377.125 350.165 ;
      RECT 9354.56 211.445 9355.795 350.165 ;
      RECT 9354.56 211.445 9381.795 308.075 ;
      RECT 9354.56 228.445 9382.56 291.075 ;
      RECT 9356.925 189.04 9377.125 308.075 ;
      RECT 9354.56 189.04 9382.56 195.075 ;
      RECT 9339.04 228.445 9352.04 350.165 ;
      RECT 9339.04 189.04 9345.395 350.165 ;
      RECT 9339.04 189.04 9352.04 212.075 ;
      RECT 9322.06 290.445 9335.06 330.165 ;
      RECT 9333.19 189.04 9335.06 330.165 ;
      RECT 9331.425 194.425 9335.06 330.165 ;
      RECT 9322.06 189.04 9323.675 330.165 ;
      RECT 9322.06 194.425 9335.06 259.875 ;
      RECT 9322.06 189.04 9330.41 259.875 ;
      RECT 9322.06 189.04 9335.06 190.125 ;
      RECT 9305.08 211.445 9318.08 350.165 ;
      RECT 9305.425 189.04 9318.08 350.165 ;
      RECT 9305.08 189.04 9318.08 195.075 ;
      RECT 9274.56 259.445 9302.56 350.165 ;
      RECT 9286.935 211.445 9302.56 350.165 ;
      RECT 9274.56 189.04 9279.185 350.165 ;
      RECT 9274.56 189.04 9300.515 228.875 ;
      RECT 9274.56 189.04 9302.56 195.075 ;
      RECT 9259.04 307.445 9272.04 350.165 ;
      RECT 9269.035 194.37 9272.04 350.165 ;
      RECT 9259.04 189.04 9264.125 350.165 ;
      RECT 9259.04 228.445 9272.04 291.075 ;
      RECT 9259.04 194.37 9272.04 212.075 ;
      RECT 9259.04 189.04 9267.37 212.075 ;
      RECT 9259.04 189.04 9272.04 190.17 ;
      RECT 9242.06 307.445 9255.06 330.165 ;
      RECT 9246.705 189.04 9255.06 330.165 ;
      RECT 9246.54 228.445 9255.06 330.165 ;
      RECT 9242.06 228.445 9255.06 291.075 ;
      RECT 9242.06 189.04 9255.06 212.075 ;
      RECT 9225.08 324.445 9238.08 350.165 ;
      RECT 9225.08 189.04 9237.125 350.165 ;
      RECT 9225.08 211.445 9238.08 308.075 ;
      RECT 9225.08 189.04 9238.08 195.075 ;
      RECT 9194.56 324.445 9222.56 350.165 ;
      RECT 9220.705 189.04 9222.56 350.165 ;
      RECT 9194.56 228.445 9215.795 350.165 ;
      RECT 9218.115 189.04 9222.56 308.075 ;
      RECT 9201.11 211.445 9222.56 308.075 ;
      RECT 9194.56 189.04 9213.205 212.075 ;
      RECT 9194.56 189.04 9222.56 195.075 ;
      RECT 9179.04 290.445 9192.04 350.165 ;
      RECT 9191.425 194.42 9192.04 350.165 ;
      RECT 9179.04 189.04 9183.675 350.165 ;
      RECT 9179.04 194.42 9192.04 259.875 ;
      RECT 9179.04 189.04 9190.41 259.875 ;
      RECT 9179.04 189.04 9192.04 190.125 ;
      RECT 9162.06 211.445 9175.06 330.165 ;
      RECT 9165.425 189.04 9175.06 330.165 ;
      RECT 9162.06 189.04 9175.06 195.075 ;
      RECT 9145.08 259.445 9158.08 350.165 ;
      RECT 9146.935 189.04 9158.08 350.165 ;
      RECT 9145.08 189.04 9158.08 228.875 ;
      RECT 9114.56 307.445 9142.56 350.165 ;
      RECT 9129.035 259.445 9142.56 350.165 ;
      RECT 9114.56 189.04 9124.125 350.165 ;
      RECT 9114.56 228.445 9139.185 291.075 ;
      RECT 9133.09 189.04 9142.56 228.875 ;
      RECT 9129.035 194.37 9142.56 228.875 ;
      RECT 9114.56 194.37 9142.56 212.075 ;
      RECT 9114.56 189.04 9127.37 212.075 ;
      RECT 9114.56 189.04 9142.56 190.17 ;
      RECT 9099.04 324.445 9112.04 350.165 ;
      RECT 9106.705 189.04 9112.04 350.165 ;
      RECT 9102.035 307.445 9112.04 350.165 ;
      RECT 9099.04 307.445 9112.04 308.075 ;
      RECT 9099.04 211.445 9101.795 308.075 ;
      RECT 9099.04 228.445 9112.04 291.075 ;
      RECT 9099.04 211.445 9112.04 212.075 ;
      RECT 9102.035 189.04 9112.04 212.075 ;
      RECT 9099.04 189.04 9112.04 195.075 ;
      RECT 9065.08 324.445 9078.08 350.165 ;
      RECT 9065.08 228.445 9075.795 350.165 ;
      RECT 9070.31 211.445 9078.08 308.075 ;
      RECT 9065.08 189.04 9073.125 212.075 ;
      RECT 9065.08 189.04 9078.08 195.075 ;
      RECT 9034.56 290.445 9062.56 350.165 ;
      RECT 9053.19 189.04 9062.56 350.165 ;
      RECT 9051.425 194.425 9062.56 350.165 ;
      RECT 9034.56 189.04 9043.675 350.165 ;
      RECT 9034.56 194.425 9062.56 259.875 ;
      RECT 9034.56 189.04 9050.41 259.875 ;
      RECT 9034.56 189.04 9062.56 190.125 ;
      RECT 9019.04 211.445 9032.04 350.165 ;
      RECT 9025.425 189.04 9032.04 350.165 ;
      RECT 9019.04 189.04 9020.515 350.165 ;
      RECT 9019.04 189.04 9032.04 195.075 ;
      RECT 9002.06 259.445 9015.06 330.165 ;
      RECT 9006.935 189.04 9015.06 330.165 ;
      RECT 9002.06 189.04 9015.06 228.875 ;
      RECT 8985.08 307.445 8998.08 350.165 ;
      RECT 8993.09 189.04 8998.08 350.165 ;
      RECT 8989.035 194.37 8998.08 350.165 ;
      RECT 8985.08 228.445 8998.08 291.075 ;
      RECT 8985.08 194.37 8998.08 212.075 ;
      RECT 8985.08 189.04 8987.37 212.075 ;
      RECT 8985.08 189.04 8998.08 190.38 ;
      RECT 8954.56 324.445 8982.56 350.165 ;
      RECT 8966.705 189.04 8982.56 350.165 ;
      RECT 8962.035 307.445 8982.56 350.165 ;
      RECT 8954.56 189.04 8957.125 350.165 ;
      RECT 8954.56 307.445 8982.56 308.075 ;
      RECT 8954.56 211.445 8961.795 308.075 ;
      RECT 8954.56 228.445 8982.56 291.075 ;
      RECT 8954.56 211.445 8982.56 212.075 ;
      RECT 8962.035 189.04 8982.56 212.075 ;
      RECT 8954.56 189.04 8982.56 195.075 ;
      RECT 8939.04 324.445 8952.04 350.165 ;
      RECT 8940.705 189.04 8952.04 350.165 ;
      RECT 8939.04 189.04 8952.04 308.075 ;
      RECT 8922.06 228.445 8935.06 330.165 ;
      RECT 8928.69 211.445 8935.06 330.165 ;
      RECT 8922.06 189.04 8932.015 212.075 ;
      RECT 8922.06 189.04 8935.06 195.075 ;
      RECT 8905.08 290.445 8918.08 350.165 ;
      RECT 8913.19 189.04 8918.08 350.165 ;
      RECT 8911.425 194.425 8918.08 350.165 ;
      RECT 8905.08 194.425 8918.08 259.875 ;
      RECT 8905.08 189.04 8910.41 259.875 ;
      RECT 8905.08 189.04 8918.08 190.125 ;
      RECT 8874.56 211.445 8902.56 350.165 ;
      RECT 8885.425 189.04 8902.56 350.165 ;
      RECT 8874.56 189.04 8880.515 350.165 ;
      RECT 8874.56 189.04 8902.56 195.075 ;
      RECT 8859.04 259.445 8872.04 350.165 ;
      RECT 8866.935 189.04 8872.04 350.165 ;
      RECT 8859.04 189.04 8872.04 228.875 ;
      RECT 8842.06 307.445 8855.06 330.165 ;
      RECT 8852.99 189.04 8855.06 330.165 ;
      RECT 8849.035 194.37 8855.06 330.165 ;
      RECT 8842.06 189.04 8844.125 330.165 ;
      RECT 8842.06 228.445 8855.06 291.075 ;
      RECT 8842.06 194.37 8855.06 212.075 ;
      RECT 8842.06 189.04 8847.37 212.075 ;
      RECT 8842.06 189.04 8855.06 190.17 ;
      RECT 8825.08 307.445 8838.08 350.165 ;
      RECT 8826.705 189.04 8838.08 350.165 ;
      RECT 8825.08 228.445 8838.08 291.075 ;
      RECT 8825.08 189.04 8838.08 212.075 ;
      RECT 8794.56 324.445 8822.56 350.165 ;
      RECT 8800.705 189.04 8817.125 350.165 ;
      RECT 8794.56 211.445 8795.795 350.165 ;
      RECT 8794.56 211.445 8821.795 308.075 ;
      RECT 8794.56 228.445 8822.56 291.075 ;
      RECT 8796.925 189.04 8817.125 308.075 ;
      RECT 8794.56 189.04 8822.56 195.075 ;
      RECT 8779.04 228.445 8792.04 350.165 ;
      RECT 8779.04 189.04 8785.395 350.165 ;
      RECT 8779.04 189.04 8792.04 212.075 ;
      RECT 8762.06 290.445 8775.06 330.165 ;
      RECT 8773.19 189.04 8775.06 330.165 ;
      RECT 8771.425 194.425 8775.06 330.165 ;
      RECT 8762.06 189.04 8763.675 330.165 ;
      RECT 8762.06 194.425 8775.06 259.875 ;
      RECT 8762.06 189.04 8770.41 259.875 ;
      RECT 8762.06 189.04 8775.06 190.125 ;
      RECT 8745.08 211.445 8758.08 350.165 ;
      RECT 8745.425 189.04 8758.08 350.165 ;
      RECT 8745.08 189.04 8758.08 195.075 ;
      RECT 8714.56 259.445 8742.56 350.165 ;
      RECT 8726.935 211.445 8742.56 350.165 ;
      RECT 8714.56 189.04 8719.185 350.165 ;
      RECT 8714.56 189.04 8740.515 228.875 ;
      RECT 8714.56 189.04 8742.56 195.075 ;
      RECT 8699.04 307.445 8712.04 350.165 ;
      RECT 8709.035 194.37 8712.04 350.165 ;
      RECT 8699.04 189.04 8704.125 350.165 ;
      RECT 8699.04 228.445 8712.04 291.075 ;
      RECT 8699.04 194.37 8712.04 212.075 ;
      RECT 8699.04 189.04 8707.37 212.075 ;
      RECT 8699.04 189.04 8712.04 190.17 ;
      RECT 8682.06 307.445 8695.06 330.165 ;
      RECT 8686.705 189.04 8695.06 330.165 ;
      RECT 8686.54 228.445 8695.06 330.165 ;
      RECT 8682.06 228.445 8695.06 291.075 ;
      RECT 8682.06 189.04 8695.06 212.075 ;
      RECT 8665.08 324.445 8678.08 350.165 ;
      RECT 8665.08 189.04 8677.125 350.165 ;
      RECT 8665.08 211.445 8678.08 308.075 ;
      RECT 8665.08 189.04 8678.08 195.075 ;
      RECT 8634.56 324.445 8662.56 350.165 ;
      RECT 8660.705 189.04 8662.56 350.165 ;
      RECT 8634.56 228.445 8655.795 350.165 ;
      RECT 8658.115 189.04 8662.56 308.075 ;
      RECT 8641.11 211.445 8662.56 308.075 ;
      RECT 8634.56 189.04 8653.205 212.075 ;
      RECT 8634.56 189.04 8662.56 195.075 ;
      RECT 8619.04 290.445 8632.04 350.165 ;
      RECT 8631.425 194.42 8632.04 350.165 ;
      RECT 8619.04 189.04 8623.675 350.165 ;
      RECT 8619.04 194.42 8632.04 259.875 ;
      RECT 8619.04 189.04 8630.41 259.875 ;
      RECT 8619.04 189.04 8632.04 190.125 ;
      RECT 8602.06 211.445 8615.06 330.165 ;
      RECT 8605.425 189.04 8615.06 330.165 ;
      RECT 8602.06 189.04 8615.06 195.075 ;
      RECT 8585.08 259.445 8598.08 350.165 ;
      RECT 8586.935 189.04 8598.08 350.165 ;
      RECT 8585.08 189.04 8598.08 228.875 ;
      RECT 8554.56 307.445 8582.56 350.165 ;
      RECT 8569.035 259.445 8582.56 350.165 ;
      RECT 8554.56 189.04 8564.125 350.165 ;
      RECT 8554.56 228.445 8579.185 291.075 ;
      RECT 8573.09 189.04 8582.56 228.875 ;
      RECT 8569.035 194.37 8582.56 228.875 ;
      RECT 8554.56 194.37 8582.56 212.075 ;
      RECT 8554.56 189.04 8567.37 212.075 ;
      RECT 8554.56 189.04 8582.56 190.17 ;
      RECT 8539.04 324.445 8552.04 350.165 ;
      RECT 8546.705 189.04 8552.04 350.165 ;
      RECT 8542.035 307.445 8552.04 350.165 ;
      RECT 8539.04 307.445 8552.04 308.075 ;
      RECT 8539.04 211.445 8541.795 308.075 ;
      RECT 8539.04 228.445 8552.04 291.075 ;
      RECT 8539.04 211.445 8552.04 212.075 ;
      RECT 8542.035 189.04 8552.04 212.075 ;
      RECT 8539.04 189.04 8552.04 195.075 ;
      RECT 8505.08 324.445 8518.08 350.165 ;
      RECT 8505.08 228.445 8515.795 350.165 ;
      RECT 8510.31 211.445 8518.08 308.075 ;
      RECT 8505.08 189.04 8513.125 212.075 ;
      RECT 8505.08 189.04 8518.08 195.075 ;
      RECT 8474.56 290.445 8502.56 350.165 ;
      RECT 8493.19 189.04 8502.56 350.165 ;
      RECT 8491.425 194.425 8502.56 350.165 ;
      RECT 8474.56 189.04 8483.675 350.165 ;
      RECT 8474.56 194.425 8502.56 259.875 ;
      RECT 8474.56 189.04 8490.41 259.875 ;
      RECT 8474.56 189.04 8502.56 190.125 ;
      RECT 8459.04 211.445 8472.04 350.165 ;
      RECT 8465.425 189.04 8472.04 350.165 ;
      RECT 8459.04 189.04 8460.515 350.165 ;
      RECT 8459.04 189.04 8472.04 195.075 ;
      RECT 8442.06 259.445 8455.06 330.165 ;
      RECT 8446.935 189.04 8455.06 330.165 ;
      RECT 8442.06 189.04 8455.06 228.875 ;
      RECT 8425.08 307.445 8438.08 350.165 ;
      RECT 8433.09 189.04 8438.08 350.165 ;
      RECT 8429.035 194.37 8438.08 350.165 ;
      RECT 8425.08 228.445 8438.08 291.075 ;
      RECT 8425.08 194.37 8438.08 212.075 ;
      RECT 8425.08 189.04 8427.37 212.075 ;
      RECT 8425.08 189.04 8438.08 190.38 ;
      RECT 8394.56 324.445 8422.56 350.165 ;
      RECT 8406.705 189.04 8422.56 350.165 ;
      RECT 8402.035 307.445 8422.56 350.165 ;
      RECT 8394.56 189.04 8397.125 350.165 ;
      RECT 8394.56 307.445 8422.56 308.075 ;
      RECT 8394.56 211.445 8401.795 308.075 ;
      RECT 8394.56 228.445 8422.56 291.075 ;
      RECT 8394.56 211.445 8422.56 212.075 ;
      RECT 8402.035 189.04 8422.56 212.075 ;
      RECT 8394.56 189.04 8422.56 195.075 ;
      RECT 8379.04 324.445 8392.04 350.165 ;
      RECT 8380.705 189.04 8392.04 350.165 ;
      RECT 8379.04 189.04 8392.04 308.075 ;
      RECT 8362.06 228.445 8375.06 330.165 ;
      RECT 8368.69 211.445 8375.06 330.165 ;
      RECT 8362.06 189.04 8372.015 212.075 ;
      RECT 8362.06 189.04 8375.06 195.075 ;
      RECT 8345.08 290.445 8358.08 350.165 ;
      RECT 8353.19 189.04 8358.08 350.165 ;
      RECT 8351.425 194.425 8358.08 350.165 ;
      RECT 8345.08 194.425 8358.08 259.875 ;
      RECT 8345.08 189.04 8350.41 259.875 ;
      RECT 8345.08 189.04 8358.08 190.125 ;
      RECT 8314.56 211.445 8342.56 350.165 ;
      RECT 8325.425 189.04 8342.56 350.165 ;
      RECT 8314.56 189.04 8320.515 350.165 ;
      RECT 8314.56 189.04 8342.56 195.075 ;
      RECT 8299.04 259.445 8312.04 350.165 ;
      RECT 8306.935 189.04 8312.04 350.165 ;
      RECT 8299.04 189.04 8312.04 228.875 ;
      RECT 8282.06 307.445 8295.06 330.165 ;
      RECT 8292.99 189.04 8295.06 330.165 ;
      RECT 8289.035 194.37 8295.06 330.165 ;
      RECT 8282.06 189.04 8284.125 330.165 ;
      RECT 8282.06 228.445 8295.06 291.075 ;
      RECT 8282.06 194.37 8295.06 212.075 ;
      RECT 8282.06 189.04 8287.37 212.075 ;
      RECT 8282.06 189.04 8295.06 190.17 ;
      RECT 8265.08 307.445 8278.08 350.165 ;
      RECT 8266.705 189.04 8278.08 350.165 ;
      RECT 8265.08 228.445 8278.08 291.075 ;
      RECT 8265.08 189.04 8278.08 212.075 ;
      RECT 8234.56 324.445 8262.56 350.165 ;
      RECT 8240.705 189.04 8257.125 350.165 ;
      RECT 8234.56 211.445 8235.795 350.165 ;
      RECT 8234.56 211.445 8261.795 308.075 ;
      RECT 8234.56 228.445 8262.56 291.075 ;
      RECT 8236.925 189.04 8257.125 308.075 ;
      RECT 8234.56 189.04 8262.56 195.075 ;
      RECT 8219.04 228.445 8232.04 350.165 ;
      RECT 8219.04 189.04 8225.395 350.165 ;
      RECT 8219.04 189.04 8232.04 212.075 ;
      RECT 8202.06 290.445 8215.06 330.165 ;
      RECT 8213.19 189.04 8215.06 330.165 ;
      RECT 8211.425 194.425 8215.06 330.165 ;
      RECT 8202.06 189.04 8203.675 330.165 ;
      RECT 8202.06 194.425 8215.06 259.875 ;
      RECT 8202.06 189.04 8210.41 259.875 ;
      RECT 8202.06 189.04 8215.06 190.125 ;
      RECT 8185.08 211.445 8198.08 350.165 ;
      RECT 8185.425 189.04 8198.08 350.165 ;
      RECT 8185.08 189.04 8198.08 195.075 ;
      RECT 8154.56 259.445 8182.56 350.165 ;
      RECT 8166.935 211.445 8182.56 350.165 ;
      RECT 8154.56 189.04 8159.185 350.165 ;
      RECT 8154.56 189.04 8180.515 228.875 ;
      RECT 8154.56 189.04 8182.56 195.075 ;
      RECT 8139.04 307.445 8152.04 350.165 ;
      RECT 8149.035 194.37 8152.04 350.165 ;
      RECT 8139.04 189.04 8144.125 350.165 ;
      RECT 8139.04 228.445 8152.04 291.075 ;
      RECT 8139.04 194.37 8152.04 212.075 ;
      RECT 8139.04 189.04 8147.37 212.075 ;
      RECT 8139.04 189.04 8152.04 190.17 ;
      RECT 8122.06 307.445 8135.06 330.165 ;
      RECT 8126.705 189.04 8135.06 330.165 ;
      RECT 8126.54 228.445 8135.06 330.165 ;
      RECT 8122.06 228.445 8135.06 291.075 ;
      RECT 8122.06 189.04 8135.06 212.075 ;
      RECT 8105.08 324.445 8118.08 350.165 ;
      RECT 8105.08 189.04 8117.125 350.165 ;
      RECT 8105.08 211.445 8118.08 308.075 ;
      RECT 8105.08 189.04 8118.08 195.075 ;
      RECT 8074.56 324.445 8102.56 350.165 ;
      RECT 8100.705 189.04 8102.56 350.165 ;
      RECT 8074.56 228.445 8095.795 350.165 ;
      RECT 8098.115 189.04 8102.56 308.075 ;
      RECT 8081.11 211.445 8102.56 308.075 ;
      RECT 8074.56 189.04 8093.205 212.075 ;
      RECT 8074.56 189.04 8102.56 195.075 ;
      RECT 8059.04 290.445 8072.04 350.165 ;
      RECT 8071.425 194.42 8072.04 350.165 ;
      RECT 8059.04 189.04 8063.675 350.165 ;
      RECT 8059.04 194.42 8072.04 259.875 ;
      RECT 8059.04 189.04 8070.41 259.875 ;
      RECT 8059.04 189.04 8072.04 190.125 ;
      RECT 8042.06 211.445 8055.06 330.165 ;
      RECT 8045.425 189.04 8055.06 330.165 ;
      RECT 8042.06 189.04 8055.06 195.075 ;
      RECT 8025.08 259.445 8038.08 350.165 ;
      RECT 8026.935 189.04 8038.08 350.165 ;
      RECT 8025.08 189.04 8038.08 228.875 ;
      RECT 7994.56 307.445 8022.56 350.165 ;
      RECT 8009.035 259.445 8022.56 350.165 ;
      RECT 7994.56 189.04 8004.125 350.165 ;
      RECT 7994.56 228.445 8019.185 291.075 ;
      RECT 8013.09 189.04 8022.56 228.875 ;
      RECT 8009.035 194.37 8022.56 228.875 ;
      RECT 7994.56 194.37 8022.56 212.075 ;
      RECT 7994.56 189.04 8007.37 212.075 ;
      RECT 7994.56 189.04 8022.56 190.17 ;
      RECT 7979.04 324.445 7992.04 350.165 ;
      RECT 7986.705 189.04 7992.04 350.165 ;
      RECT 7982.035 307.445 7992.04 350.165 ;
      RECT 7979.04 307.445 7992.04 308.075 ;
      RECT 7979.04 211.445 7981.795 308.075 ;
      RECT 7979.04 228.445 7992.04 291.075 ;
      RECT 7979.04 211.445 7992.04 212.075 ;
      RECT 7982.035 189.04 7992.04 212.075 ;
      RECT 7979.04 189.04 7992.04 195.075 ;
      RECT 7945.08 324.445 7958.08 350.165 ;
      RECT 7945.08 228.445 7955.795 350.165 ;
      RECT 7950.31 211.445 7958.08 308.075 ;
      RECT 7945.08 189.04 7953.125 212.075 ;
      RECT 7945.08 189.04 7958.08 195.075 ;
      RECT 7914.56 290.445 7942.56 350.165 ;
      RECT 7933.19 189.04 7942.56 350.165 ;
      RECT 7931.425 194.425 7942.56 350.165 ;
      RECT 7914.56 189.04 7923.675 350.165 ;
      RECT 7914.56 194.425 7942.56 259.875 ;
      RECT 7914.56 189.04 7930.41 259.875 ;
      RECT 7914.56 189.04 7942.56 190.125 ;
      RECT 7899.04 211.445 7912.04 350.165 ;
      RECT 7905.425 189.04 7912.04 350.165 ;
      RECT 7899.04 189.04 7900.515 350.165 ;
      RECT 7899.04 189.04 7912.04 195.075 ;
      RECT 7882.06 259.445 7895.06 330.165 ;
      RECT 7886.935 189.04 7895.06 330.165 ;
      RECT 7882.06 189.04 7895.06 228.875 ;
      RECT 7865.08 307.445 7878.08 350.165 ;
      RECT 7873.09 189.04 7878.08 350.165 ;
      RECT 7869.035 194.37 7878.08 350.165 ;
      RECT 7865.08 228.445 7878.08 291.075 ;
      RECT 7865.08 194.37 7878.08 212.075 ;
      RECT 7865.08 189.04 7867.37 212.075 ;
      RECT 7865.08 189.04 7878.08 190.38 ;
      RECT 7834.56 324.445 7862.56 350.165 ;
      RECT 7846.705 189.04 7862.56 350.165 ;
      RECT 7842.035 307.445 7862.56 350.165 ;
      RECT 7834.56 189.04 7837.125 350.165 ;
      RECT 7834.56 307.445 7862.56 308.075 ;
      RECT 7834.56 211.445 7841.795 308.075 ;
      RECT 7834.56 228.445 7862.56 291.075 ;
      RECT 7834.56 211.445 7862.56 212.075 ;
      RECT 7842.035 189.04 7862.56 212.075 ;
      RECT 7834.56 189.04 7862.56 195.075 ;
      RECT 7819.04 324.445 7832.04 350.165 ;
      RECT 7820.705 189.04 7832.04 350.165 ;
      RECT 7819.04 189.04 7832.04 308.075 ;
      RECT 7802.06 228.445 7815.06 330.165 ;
      RECT 7808.69 211.445 7815.06 330.165 ;
      RECT 7802.06 189.04 7812.015 212.075 ;
      RECT 7802.06 189.04 7815.06 195.075 ;
      RECT 7785.08 290.445 7798.08 350.165 ;
      RECT 7793.19 189.04 7798.08 350.165 ;
      RECT 7791.425 194.425 7798.08 350.165 ;
      RECT 7785.08 194.425 7798.08 259.875 ;
      RECT 7785.08 189.04 7790.41 259.875 ;
      RECT 7785.08 189.04 7798.08 190.125 ;
      RECT 7754.56 211.445 7782.56 350.165 ;
      RECT 7765.425 189.04 7782.56 350.165 ;
      RECT 7754.56 189.04 7760.515 350.165 ;
      RECT 7754.56 189.04 7782.56 195.075 ;
      RECT 7739.04 259.445 7752.04 350.165 ;
      RECT 7746.935 189.04 7752.04 350.165 ;
      RECT 7739.04 189.04 7752.04 228.875 ;
      RECT 7722.06 307.445 7735.06 330.165 ;
      RECT 7732.99 189.04 7735.06 330.165 ;
      RECT 7729.035 194.37 7735.06 330.165 ;
      RECT 7722.06 189.04 7724.125 330.165 ;
      RECT 7722.06 228.445 7735.06 291.075 ;
      RECT 7722.06 194.37 7735.06 212.075 ;
      RECT 7722.06 189.04 7727.37 212.075 ;
      RECT 7722.06 189.04 7735.06 190.17 ;
      RECT 7705.08 307.445 7718.08 350.165 ;
      RECT 7706.705 189.04 7718.08 350.165 ;
      RECT 7705.08 228.445 7718.08 291.075 ;
      RECT 7705.08 189.04 7718.08 212.075 ;
      RECT 7674.56 324.445 7702.56 350.165 ;
      RECT 7680.705 189.04 7697.125 350.165 ;
      RECT 7674.56 211.445 7675.795 350.165 ;
      RECT 7674.56 211.445 7701.795 308.075 ;
      RECT 7674.56 228.445 7702.56 291.075 ;
      RECT 7676.925 189.04 7697.125 308.075 ;
      RECT 7674.56 189.04 7702.56 195.075 ;
      RECT 7659.04 228.445 7672.04 350.165 ;
      RECT 7659.04 189.04 7665.395 350.165 ;
      RECT 7659.04 189.04 7672.04 212.075 ;
      RECT 7642.06 290.445 7655.06 330.165 ;
      RECT 7653.19 189.04 7655.06 330.165 ;
      RECT 7651.425 194.425 7655.06 330.165 ;
      RECT 7642.06 189.04 7643.675 330.165 ;
      RECT 7642.06 194.425 7655.06 259.875 ;
      RECT 7642.06 189.04 7650.41 259.875 ;
      RECT 7642.06 189.04 7655.06 190.125 ;
      RECT 7625.08 211.445 7638.08 350.165 ;
      RECT 7625.425 189.04 7638.08 350.165 ;
      RECT 7625.08 189.04 7638.08 195.075 ;
      RECT 7594.56 259.445 7622.56 350.165 ;
      RECT 7606.935 211.445 7622.56 350.165 ;
      RECT 7594.56 189.04 7599.185 350.165 ;
      RECT 7594.56 189.04 7620.515 228.875 ;
      RECT 7594.56 189.04 7622.56 195.075 ;
      RECT 7579.04 307.445 7592.04 350.165 ;
      RECT 7589.035 194.37 7592.04 350.165 ;
      RECT 7579.04 189.04 7584.125 350.165 ;
      RECT 7579.04 228.445 7592.04 291.075 ;
      RECT 7579.04 194.37 7592.04 212.075 ;
      RECT 7579.04 189.04 7587.37 212.075 ;
      RECT 7579.04 189.04 7592.04 190.17 ;
      RECT 7562.06 307.445 7575.06 330.165 ;
      RECT 7566.705 189.04 7575.06 330.165 ;
      RECT 7566.54 228.445 7575.06 330.165 ;
      RECT 7562.06 228.445 7575.06 291.075 ;
      RECT 7562.06 189.04 7575.06 212.075 ;
      RECT 7545.08 324.445 7558.08 350.165 ;
      RECT 7545.08 189.04 7557.125 350.165 ;
      RECT 7545.08 211.445 7558.08 308.075 ;
      RECT 7545.08 189.04 7558.08 195.075 ;
      RECT 7514.56 324.445 7542.56 350.165 ;
      RECT 7540.705 189.04 7542.56 350.165 ;
      RECT 7514.56 228.445 7535.795 350.165 ;
      RECT 7538.115 189.04 7542.56 308.075 ;
      RECT 7521.11 211.445 7542.56 308.075 ;
      RECT 7514.56 189.04 7533.205 212.075 ;
      RECT 7514.56 189.04 7542.56 195.075 ;
      RECT 7499.04 290.445 7512.04 350.165 ;
      RECT 7511.425 194.42 7512.04 350.165 ;
      RECT 7499.04 189.04 7503.675 350.165 ;
      RECT 7499.04 194.42 7512.04 259.875 ;
      RECT 7499.04 189.04 7510.41 259.875 ;
      RECT 7499.04 189.04 7512.04 190.125 ;
      RECT 7482.06 211.445 7495.06 330.165 ;
      RECT 7485.425 189.04 7495.06 330.165 ;
      RECT 7482.06 189.04 7495.06 195.075 ;
      RECT 7465.08 259.445 7478.08 350.165 ;
      RECT 7466.935 189.04 7478.08 350.165 ;
      RECT 7465.08 189.04 7478.08 228.875 ;
      RECT 7434.56 307.445 7462.56 350.165 ;
      RECT 7449.035 259.445 7462.56 350.165 ;
      RECT 7434.56 189.04 7444.125 350.165 ;
      RECT 7434.56 228.445 7459.185 291.075 ;
      RECT 7453.09 189.04 7462.56 228.875 ;
      RECT 7449.035 194.37 7462.56 228.875 ;
      RECT 7434.56 194.37 7462.56 212.075 ;
      RECT 7434.56 189.04 7447.37 212.075 ;
      RECT 7434.56 189.04 7462.56 190.17 ;
      RECT 7419.04 324.445 7432.04 350.165 ;
      RECT 7426.705 189.04 7432.04 350.165 ;
      RECT 7422.035 307.445 7432.04 350.165 ;
      RECT 7419.04 307.445 7432.04 308.075 ;
      RECT 7419.04 211.445 7421.795 308.075 ;
      RECT 7419.04 228.445 7432.04 291.075 ;
      RECT 7419.04 211.445 7432.04 212.075 ;
      RECT 7422.035 189.04 7432.04 212.075 ;
      RECT 7419.04 189.04 7432.04 195.075 ;
      RECT 7385.08 324.445 7398.08 350.165 ;
      RECT 7385.08 228.445 7395.795 350.165 ;
      RECT 7390.31 211.445 7398.08 308.075 ;
      RECT 7385.08 189.04 7393.125 212.075 ;
      RECT 7385.08 189.04 7398.08 195.075 ;
      RECT 7354.56 290.445 7382.56 350.165 ;
      RECT 7373.19 189.04 7382.56 350.165 ;
      RECT 7371.425 194.425 7382.56 350.165 ;
      RECT 7354.56 189.04 7363.675 350.165 ;
      RECT 7354.56 194.425 7382.56 259.875 ;
      RECT 7354.56 189.04 7370.41 259.875 ;
      RECT 7354.56 189.04 7382.56 190.125 ;
      RECT 7339.04 211.445 7352.04 350.165 ;
      RECT 7345.425 189.04 7352.04 350.165 ;
      RECT 7339.04 189.04 7340.515 350.165 ;
      RECT 7339.04 189.04 7352.04 195.075 ;
      RECT 7322.06 259.445 7335.06 330.165 ;
      RECT 7326.935 189.04 7335.06 330.165 ;
      RECT 7322.06 189.04 7335.06 228.875 ;
      RECT 7305.08 307.445 7318.08 350.165 ;
      RECT 7313.09 189.04 7318.08 350.165 ;
      RECT 7309.035 194.37 7318.08 350.165 ;
      RECT 7305.08 228.445 7318.08 291.075 ;
      RECT 7305.08 194.37 7318.08 212.075 ;
      RECT 7305.08 189.04 7307.37 212.075 ;
      RECT 7305.08 189.04 7318.08 190.38 ;
      RECT 7274.56 324.445 7302.56 350.165 ;
      RECT 7286.705 189.04 7302.56 350.165 ;
      RECT 7282.035 307.445 7302.56 350.165 ;
      RECT 7274.56 189.04 7277.125 350.165 ;
      RECT 7274.56 307.445 7302.56 308.075 ;
      RECT 7274.56 211.445 7281.795 308.075 ;
      RECT 7274.56 228.445 7302.56 291.075 ;
      RECT 7274.56 211.445 7302.56 212.075 ;
      RECT 7282.035 189.04 7302.56 212.075 ;
      RECT 7274.56 189.04 7302.56 195.075 ;
      RECT 7259.04 324.445 7272.04 350.165 ;
      RECT 7260.705 189.04 7272.04 350.165 ;
      RECT 7259.04 189.04 7272.04 308.075 ;
      RECT 7242.06 228.445 7255.06 330.165 ;
      RECT 7248.69 211.445 7255.06 330.165 ;
      RECT 7242.06 189.04 7252.015 212.075 ;
      RECT 7242.06 189.04 7255.06 195.075 ;
      RECT 7225.08 290.445 7238.08 350.165 ;
      RECT 7233.19 189.04 7238.08 350.165 ;
      RECT 7231.425 194.425 7238.08 350.165 ;
      RECT 7225.08 194.425 7238.08 259.875 ;
      RECT 7225.08 189.04 7230.41 259.875 ;
      RECT 7225.08 189.04 7238.08 190.125 ;
      RECT 7194.56 211.445 7222.56 350.165 ;
      RECT 7205.425 189.04 7222.56 350.165 ;
      RECT 7194.56 189.04 7200.515 350.165 ;
      RECT 7194.56 189.04 7222.56 195.075 ;
      RECT 7179.04 259.445 7192.04 350.165 ;
      RECT 7186.935 189.04 7192.04 350.165 ;
      RECT 7179.04 189.04 7192.04 228.875 ;
      RECT 7162.06 307.445 7175.06 330.165 ;
      RECT 7172.99 189.04 7175.06 330.165 ;
      RECT 7169.035 194.37 7175.06 330.165 ;
      RECT 7162.06 189.04 7164.125 330.165 ;
      RECT 7162.06 228.445 7175.06 291.075 ;
      RECT 7162.06 194.37 7175.06 212.075 ;
      RECT 7162.06 189.04 7167.37 212.075 ;
      RECT 7162.06 189.04 7175.06 190.17 ;
      RECT 7145.08 307.445 7158.08 350.165 ;
      RECT 7146.705 189.04 7158.08 350.165 ;
      RECT 7145.08 228.445 7158.08 291.075 ;
      RECT 7145.08 189.04 7158.08 212.075 ;
      RECT 7114.56 324.445 7142.56 350.165 ;
      RECT 7120.705 189.04 7137.125 350.165 ;
      RECT 7114.56 211.445 7115.795 350.165 ;
      RECT 7114.56 211.445 7141.795 308.075 ;
      RECT 7114.56 228.445 7142.56 291.075 ;
      RECT 7116.925 189.04 7137.125 308.075 ;
      RECT 7114.56 189.04 7142.56 195.075 ;
      RECT 7099.04 228.445 7112.04 350.165 ;
      RECT 7099.04 189.04 7105.395 350.165 ;
      RECT 7099.04 189.04 7112.04 212.075 ;
      RECT 7082.06 290.445 7095.06 330.165 ;
      RECT 7093.19 189.04 7095.06 330.165 ;
      RECT 7091.425 194.425 7095.06 330.165 ;
      RECT 7082.06 189.04 7083.675 330.165 ;
      RECT 7082.06 194.425 7095.06 259.875 ;
      RECT 7082.06 189.04 7090.41 259.875 ;
      RECT 7082.06 189.04 7095.06 190.125 ;
      RECT 7065.08 211.445 7078.08 350.165 ;
      RECT 7065.425 189.04 7078.08 350.165 ;
      RECT 7065.08 189.04 7078.08 195.075 ;
      RECT 7034.56 259.445 7062.56 350.165 ;
      RECT 7046.935 211.445 7062.56 350.165 ;
      RECT 7034.56 189.04 7039.185 350.165 ;
      RECT 7034.56 189.04 7060.515 228.875 ;
      RECT 7034.56 189.04 7062.56 195.075 ;
      RECT 7019.04 307.445 7032.04 350.165 ;
      RECT 7029.035 194.37 7032.04 350.165 ;
      RECT 7019.04 189.04 7024.125 350.165 ;
      RECT 7019.04 228.445 7032.04 291.075 ;
      RECT 7019.04 194.37 7032.04 212.075 ;
      RECT 7019.04 189.04 7027.37 212.075 ;
      RECT 7019.04 189.04 7032.04 190.17 ;
      RECT 7002.06 307.445 7015.06 330.165 ;
      RECT 7006.705 189.04 7015.06 330.165 ;
      RECT 7006.54 228.445 7015.06 330.165 ;
      RECT 7002.06 228.445 7015.06 291.075 ;
      RECT 7002.06 189.04 7015.06 212.075 ;
      RECT 6985.08 324.445 6998.08 350.165 ;
      RECT 6985.08 189.04 6997.125 350.165 ;
      RECT 6985.08 211.445 6998.08 308.075 ;
      RECT 6985.08 189.04 6998.08 195.075 ;
      RECT 6954.56 324.445 6982.56 350.165 ;
      RECT 6980.705 189.04 6982.56 350.165 ;
      RECT 6954.56 228.445 6975.795 350.165 ;
      RECT 6978.115 189.04 6982.56 308.075 ;
      RECT 6961.11 211.445 6982.56 308.075 ;
      RECT 6954.56 189.04 6973.205 212.075 ;
      RECT 6954.56 189.04 6982.56 195.075 ;
      RECT 6939.04 290.445 6952.04 350.165 ;
      RECT 6951.425 194.42 6952.04 350.165 ;
      RECT 6939.04 189.04 6943.675 350.165 ;
      RECT 6939.04 194.42 6952.04 259.875 ;
      RECT 6939.04 189.04 6950.41 259.875 ;
      RECT 6939.04 189.04 6952.04 190.125 ;
      RECT 6922.06 211.445 6935.06 330.165 ;
      RECT 6925.425 189.04 6935.06 330.165 ;
      RECT 6922.06 189.04 6935.06 195.075 ;
      RECT 6905.08 259.445 6918.08 350.165 ;
      RECT 6906.935 189.04 6918.08 350.165 ;
      RECT 6905.08 189.04 6918.08 228.875 ;
      RECT 6874.56 307.445 6902.56 350.165 ;
      RECT 6889.035 259.445 6902.56 350.165 ;
      RECT 6874.56 189.04 6884.125 350.165 ;
      RECT 6874.56 228.445 6899.185 291.075 ;
      RECT 6893.09 189.04 6902.56 228.875 ;
      RECT 6889.035 194.37 6902.56 228.875 ;
      RECT 6874.56 194.37 6902.56 212.075 ;
      RECT 6874.56 189.04 6887.37 212.075 ;
      RECT 6874.56 189.04 6902.56 190.17 ;
      RECT 6859.04 324.445 6872.04 350.165 ;
      RECT 6866.705 189.04 6872.04 350.165 ;
      RECT 6862.035 307.445 6872.04 350.165 ;
      RECT 6859.04 307.445 6872.04 308.075 ;
      RECT 6859.04 211.445 6861.795 308.075 ;
      RECT 6859.04 228.445 6872.04 291.075 ;
      RECT 6859.04 211.445 6872.04 212.075 ;
      RECT 6862.035 189.04 6872.04 212.075 ;
      RECT 6859.04 189.04 6872.04 195.075 ;
      RECT 6825.08 324.445 6838.08 350.165 ;
      RECT 6825.08 228.445 6835.795 350.165 ;
      RECT 6830.31 211.445 6838.08 308.075 ;
      RECT 6825.08 189.04 6833.125 212.075 ;
      RECT 6825.08 189.04 6838.08 195.075 ;
      RECT 6794.56 290.445 6822.56 350.165 ;
      RECT 6813.19 189.04 6822.56 350.165 ;
      RECT 6811.425 194.425 6822.56 350.165 ;
      RECT 6794.56 189.04 6803.675 350.165 ;
      RECT 6794.56 194.425 6822.56 259.875 ;
      RECT 6794.56 189.04 6810.41 259.875 ;
      RECT 6794.56 189.04 6822.56 190.125 ;
      RECT 6779.04 211.445 6792.04 350.165 ;
      RECT 6785.425 189.04 6792.04 350.165 ;
      RECT 6779.04 189.04 6780.515 350.165 ;
      RECT 6779.04 189.04 6792.04 195.075 ;
      RECT 6762.06 259.445 6775.06 330.165 ;
      RECT 6766.935 189.04 6775.06 330.165 ;
      RECT 6762.06 189.04 6775.06 228.875 ;
      RECT 6745.08 307.445 6758.08 350.165 ;
      RECT 6753.09 189.04 6758.08 350.165 ;
      RECT 6749.035 194.37 6758.08 350.165 ;
      RECT 6745.08 228.445 6758.08 291.075 ;
      RECT 6745.08 194.37 6758.08 212.075 ;
      RECT 6745.08 189.04 6747.37 212.075 ;
      RECT 6745.08 189.04 6758.08 190.38 ;
      RECT 6714.56 324.445 6742.56 350.165 ;
      RECT 6726.705 189.04 6742.56 350.165 ;
      RECT 6722.035 307.445 6742.56 350.165 ;
      RECT 6714.56 189.04 6717.125 350.165 ;
      RECT 6714.56 307.445 6742.56 308.075 ;
      RECT 6714.56 211.445 6721.795 308.075 ;
      RECT 6714.56 228.445 6742.56 291.075 ;
      RECT 6714.56 211.445 6742.56 212.075 ;
      RECT 6722.035 189.04 6742.56 212.075 ;
      RECT 6714.56 189.04 6742.56 195.075 ;
      RECT 6699.04 324.445 6712.04 350.165 ;
      RECT 6700.705 189.04 6712.04 350.165 ;
      RECT 6699.04 189.04 6712.04 308.075 ;
      RECT 6682.06 228.445 6695.06 330.165 ;
      RECT 6688.69 211.445 6695.06 330.165 ;
      RECT 6682.06 189.04 6692.015 212.075 ;
      RECT 6682.06 189.04 6695.06 195.075 ;
      RECT 6665.08 290.445 6678.08 350.165 ;
      RECT 6673.19 189.04 6678.08 350.165 ;
      RECT 6671.425 194.425 6678.08 350.165 ;
      RECT 6665.08 194.425 6678.08 259.875 ;
      RECT 6665.08 189.04 6670.41 259.875 ;
      RECT 6665.08 189.04 6678.08 190.125 ;
      RECT 6634.56 211.445 6662.56 350.165 ;
      RECT 6645.425 189.04 6662.56 350.165 ;
      RECT 6634.56 189.04 6640.515 350.165 ;
      RECT 6634.56 189.04 6662.56 195.075 ;
      RECT 6619.04 259.445 6632.04 350.165 ;
      RECT 6626.935 189.04 6632.04 350.165 ;
      RECT 6619.04 189.04 6632.04 228.875 ;
      RECT 6602.06 307.445 6615.06 330.165 ;
      RECT 6612.99 189.04 6615.06 330.165 ;
      RECT 6609.035 194.37 6615.06 330.165 ;
      RECT 6602.06 189.04 6604.125 330.165 ;
      RECT 6602.06 228.445 6615.06 291.075 ;
      RECT 6602.06 194.37 6615.06 212.075 ;
      RECT 6602.06 189.04 6607.37 212.075 ;
      RECT 6602.06 189.04 6615.06 190.17 ;
      RECT 6585.08 307.445 6598.08 350.165 ;
      RECT 6586.705 189.04 6598.08 350.165 ;
      RECT 6585.08 228.445 6598.08 291.075 ;
      RECT 6585.08 189.04 6598.08 212.075 ;
      RECT 6554.56 324.445 6582.56 350.165 ;
      RECT 6560.705 189.04 6577.125 350.165 ;
      RECT 6554.56 211.445 6555.795 350.165 ;
      RECT 6554.56 211.445 6581.795 308.075 ;
      RECT 6554.56 228.445 6582.56 291.075 ;
      RECT 6556.925 189.04 6577.125 308.075 ;
      RECT 6554.56 189.04 6582.56 195.075 ;
      RECT 6539.04 228.445 6552.04 350.165 ;
      RECT 6539.04 189.04 6545.395 350.165 ;
      RECT 6539.04 189.04 6552.04 212.075 ;
      RECT 6522.06 290.445 6535.06 330.165 ;
      RECT 6533.19 189.04 6535.06 330.165 ;
      RECT 6531.425 194.425 6535.06 330.165 ;
      RECT 6522.06 189.04 6523.675 330.165 ;
      RECT 6522.06 194.425 6535.06 259.875 ;
      RECT 6522.06 189.04 6530.41 259.875 ;
      RECT 6522.06 189.04 6535.06 190.125 ;
      RECT 6505.08 211.445 6518.08 350.165 ;
      RECT 6505.425 189.04 6518.08 350.165 ;
      RECT 6505.08 189.04 6518.08 195.075 ;
      RECT 6474.56 259.445 6502.56 350.165 ;
      RECT 6486.935 211.445 6502.56 350.165 ;
      RECT 6474.56 189.04 6479.185 350.165 ;
      RECT 6474.56 189.04 6500.515 228.875 ;
      RECT 6474.56 189.04 6502.56 195.075 ;
      RECT 6459.04 307.445 6472.04 350.165 ;
      RECT 6469.035 194.37 6472.04 350.165 ;
      RECT 6459.04 189.04 6464.125 350.165 ;
      RECT 6459.04 228.445 6472.04 291.075 ;
      RECT 6459.04 194.37 6472.04 212.075 ;
      RECT 6459.04 189.04 6467.37 212.075 ;
      RECT 6459.04 189.04 6472.04 190.17 ;
      RECT 6442.06 307.445 6455.06 330.165 ;
      RECT 6446.705 189.04 6455.06 330.165 ;
      RECT 6446.54 228.445 6455.06 330.165 ;
      RECT 6442.06 228.445 6455.06 291.075 ;
      RECT 6442.06 189.04 6455.06 212.075 ;
      RECT 6425.08 324.445 6438.08 350.165 ;
      RECT 6425.08 189.04 6437.125 350.165 ;
      RECT 6425.08 211.445 6438.08 308.075 ;
      RECT 6425.08 189.04 6438.08 195.075 ;
      RECT 6394.56 324.445 6422.56 350.165 ;
      RECT 6420.705 189.04 6422.56 350.165 ;
      RECT 6394.56 228.445 6415.795 350.165 ;
      RECT 6418.115 189.04 6422.56 308.075 ;
      RECT 6401.11 211.445 6422.56 308.075 ;
      RECT 6394.56 189.04 6413.205 212.075 ;
      RECT 6394.56 189.04 6422.56 195.075 ;
      RECT 6379.04 290.445 6392.04 350.165 ;
      RECT 6391.425 194.42 6392.04 350.165 ;
      RECT 6379.04 189.04 6383.675 350.165 ;
      RECT 6379.04 194.42 6392.04 259.875 ;
      RECT 6379.04 189.04 6390.41 259.875 ;
      RECT 6379.04 189.04 6392.04 190.125 ;
      RECT 6362.06 211.445 6375.06 330.165 ;
      RECT 6365.425 189.04 6375.06 330.165 ;
      RECT 6362.06 189.04 6375.06 195.075 ;
      RECT 6345.08 259.445 6358.08 350.165 ;
      RECT 6346.935 189.04 6358.08 350.165 ;
      RECT 6345.08 189.04 6358.08 228.875 ;
      RECT 6314.56 307.445 6342.56 350.165 ;
      RECT 6329.035 259.445 6342.56 350.165 ;
      RECT 6314.56 189.04 6324.125 350.165 ;
      RECT 6314.56 228.445 6339.185 291.075 ;
      RECT 6333.09 189.04 6342.56 228.875 ;
      RECT 6329.035 194.37 6342.56 228.875 ;
      RECT 6314.56 194.37 6342.56 212.075 ;
      RECT 6314.56 189.04 6327.37 212.075 ;
      RECT 6314.56 189.04 6342.56 190.17 ;
      RECT 6299.04 324.445 6312.04 350.165 ;
      RECT 6306.705 189.04 6312.04 350.165 ;
      RECT 6302.035 307.445 6312.04 350.165 ;
      RECT 6299.04 307.445 6312.04 308.075 ;
      RECT 6299.04 211.445 6301.795 308.075 ;
      RECT 6299.04 228.445 6312.04 291.075 ;
      RECT 6299.04 211.445 6312.04 212.075 ;
      RECT 6302.035 189.04 6312.04 212.075 ;
      RECT 6299.04 189.04 6312.04 195.075 ;
      RECT 6265.08 324.445 6278.08 350.165 ;
      RECT 6265.08 228.445 6275.795 350.165 ;
      RECT 6270.31 211.445 6278.08 308.075 ;
      RECT 6265.08 189.04 6273.125 212.075 ;
      RECT 6265.08 189.04 6278.08 195.075 ;
      RECT 6234.56 290.445 6262.56 350.165 ;
      RECT 6253.19 189.04 6262.56 350.165 ;
      RECT 6251.425 194.425 6262.56 350.165 ;
      RECT 6234.56 189.04 6243.675 350.165 ;
      RECT 6234.56 194.425 6262.56 259.875 ;
      RECT 6234.56 189.04 6250.41 259.875 ;
      RECT 6234.56 189.04 6262.56 190.125 ;
      RECT 6219.04 211.445 6232.04 350.165 ;
      RECT 6225.425 189.04 6232.04 350.165 ;
      RECT 6219.04 189.04 6220.515 350.165 ;
      RECT 6219.04 189.04 6232.04 195.075 ;
      RECT 6202.06 259.445 6215.06 330.165 ;
      RECT 6206.935 189.04 6215.06 330.165 ;
      RECT 6202.06 189.04 6215.06 228.875 ;
      RECT 6185.08 307.445 6198.08 350.165 ;
      RECT 6193.09 189.04 6198.08 350.165 ;
      RECT 6189.035 194.37 6198.08 350.165 ;
      RECT 6185.08 228.445 6198.08 291.075 ;
      RECT 6185.08 194.37 6198.08 212.075 ;
      RECT 6185.08 189.04 6187.37 212.075 ;
      RECT 6185.08 189.04 6198.08 190.38 ;
      RECT 6154.56 324.445 6182.56 350.165 ;
      RECT 6166.705 189.04 6182.56 350.165 ;
      RECT 6162.035 307.445 6182.56 350.165 ;
      RECT 6154.56 189.04 6157.125 350.165 ;
      RECT 6154.56 307.445 6182.56 308.075 ;
      RECT 6154.56 211.445 6161.795 308.075 ;
      RECT 6154.56 228.445 6182.56 291.075 ;
      RECT 6154.56 211.445 6182.56 212.075 ;
      RECT 6162.035 189.04 6182.56 212.075 ;
      RECT 6154.56 189.04 6182.56 195.075 ;
      RECT 6139.04 324.445 6152.04 350.165 ;
      RECT 6140.705 189.04 6152.04 350.165 ;
      RECT 6139.04 189.04 6152.04 308.075 ;
      RECT 6122.06 228.445 6135.06 330.165 ;
      RECT 6128.69 211.445 6135.06 330.165 ;
      RECT 6122.06 189.04 6132.015 212.075 ;
      RECT 6122.06 189.04 6135.06 195.075 ;
      RECT 6105.08 290.445 6118.08 350.165 ;
      RECT 6113.19 189.04 6118.08 350.165 ;
      RECT 6111.425 194.425 6118.08 350.165 ;
      RECT 6105.08 194.425 6118.08 259.875 ;
      RECT 6105.08 189.04 6110.41 259.875 ;
      RECT 6105.08 189.04 6118.08 190.125 ;
      RECT 6074.56 211.445 6102.56 350.165 ;
      RECT 6085.425 189.04 6102.56 350.165 ;
      RECT 6074.56 189.04 6080.515 350.165 ;
      RECT 6074.56 189.04 6102.56 195.075 ;
      RECT 6059.04 259.445 6072.04 350.165 ;
      RECT 6066.935 189.04 6072.04 350.165 ;
      RECT 6059.04 189.04 6072.04 228.875 ;
      RECT 6042.06 307.445 6055.06 330.165 ;
      RECT 6052.99 189.04 6055.06 330.165 ;
      RECT 6049.035 194.37 6055.06 330.165 ;
      RECT 6042.06 189.04 6044.125 330.165 ;
      RECT 6042.06 228.445 6055.06 291.075 ;
      RECT 6042.06 194.37 6055.06 212.075 ;
      RECT 6042.06 189.04 6047.37 212.075 ;
      RECT 6042.06 189.04 6055.06 190.17 ;
      RECT 6025.08 307.445 6038.08 350.165 ;
      RECT 6026.705 189.04 6038.08 350.165 ;
      RECT 6025.08 228.445 6038.08 291.075 ;
      RECT 6025.08 189.04 6038.08 212.075 ;
      RECT 5994.56 324.445 6022.56 350.165 ;
      RECT 6000.705 189.04 6017.125 350.165 ;
      RECT 5994.56 211.445 5995.795 350.165 ;
      RECT 5994.56 211.445 6021.795 308.075 ;
      RECT 5994.56 228.445 6022.56 291.075 ;
      RECT 5996.925 189.04 6017.125 308.075 ;
      RECT 5994.56 189.04 6022.56 195.075 ;
      RECT 5979.04 228.445 5992.04 350.165 ;
      RECT 5979.04 189.04 5985.395 350.165 ;
      RECT 5979.04 189.04 5992.04 212.075 ;
      RECT 5962.06 290.445 5975.06 330.165 ;
      RECT 5973.19 189.04 5975.06 330.165 ;
      RECT 5971.425 194.425 5975.06 330.165 ;
      RECT 5962.06 189.04 5963.675 330.165 ;
      RECT 5962.06 194.425 5975.06 259.875 ;
      RECT 5962.06 189.04 5970.41 259.875 ;
      RECT 5962.06 189.04 5975.06 190.125 ;
      RECT 5945.08 211.445 5958.08 350.165 ;
      RECT 5945.425 189.04 5958.08 350.165 ;
      RECT 5945.08 189.04 5958.08 195.075 ;
      RECT 5914.56 259.445 5942.56 350.165 ;
      RECT 5926.935 211.445 5942.56 350.165 ;
      RECT 5914.56 189.04 5919.185 350.165 ;
      RECT 5914.56 189.04 5940.515 228.875 ;
      RECT 5914.56 189.04 5942.56 195.075 ;
      RECT 5899.04 307.445 5912.04 350.165 ;
      RECT 5909.035 194.37 5912.04 350.165 ;
      RECT 5899.04 189.04 5904.125 350.165 ;
      RECT 5899.04 228.445 5912.04 291.075 ;
      RECT 5899.04 194.37 5912.04 212.075 ;
      RECT 5899.04 189.04 5907.37 212.075 ;
      RECT 5899.04 189.04 5912.04 190.17 ;
      RECT 5882.06 307.445 5895.06 330.165 ;
      RECT 5886.705 189.04 5895.06 330.165 ;
      RECT 5886.54 228.445 5895.06 330.165 ;
      RECT 5882.06 228.445 5895.06 291.075 ;
      RECT 5882.06 189.04 5895.06 212.075 ;
      RECT 5865.08 324.445 5878.08 350.165 ;
      RECT 5865.08 189.04 5877.125 350.165 ;
      RECT 5865.08 211.445 5878.08 308.075 ;
      RECT 5865.08 189.04 5878.08 195.075 ;
      RECT 5834.56 324.445 5862.56 350.165 ;
      RECT 5860.705 189.04 5862.56 350.165 ;
      RECT 5834.56 228.445 5855.795 350.165 ;
      RECT 5858.115 189.04 5862.56 308.075 ;
      RECT 5841.11 211.445 5862.56 308.075 ;
      RECT 5834.56 189.04 5853.205 212.075 ;
      RECT 5834.56 189.04 5862.56 195.075 ;
      RECT 5819.04 290.445 5832.04 350.165 ;
      RECT 5831.425 194.42 5832.04 350.165 ;
      RECT 5819.04 189.04 5823.675 350.165 ;
      RECT 5819.04 194.42 5832.04 259.875 ;
      RECT 5819.04 189.04 5830.41 259.875 ;
      RECT 5819.04 189.04 5832.04 190.125 ;
      RECT 5802.06 211.445 5815.06 330.165 ;
      RECT 5805.425 189.04 5815.06 330.165 ;
      RECT 5802.06 189.04 5815.06 195.075 ;
      RECT 5785.08 259.445 5798.08 350.165 ;
      RECT 5786.935 189.04 5798.08 350.165 ;
      RECT 5785.08 189.04 5798.08 228.875 ;
      RECT 5754.56 307.445 5782.56 350.165 ;
      RECT 5769.035 259.445 5782.56 350.165 ;
      RECT 5754.56 189.04 5764.125 350.165 ;
      RECT 5754.56 228.445 5779.185 291.075 ;
      RECT 5773.09 189.04 5782.56 228.875 ;
      RECT 5769.035 194.37 5782.56 228.875 ;
      RECT 5754.56 194.37 5782.56 212.075 ;
      RECT 5754.56 189.04 5767.37 212.075 ;
      RECT 5754.56 189.04 5782.56 190.17 ;
      RECT 5739.04 324.445 5752.04 350.165 ;
      RECT 5746.705 189.04 5752.04 350.165 ;
      RECT 5742.035 307.445 5752.04 350.165 ;
      RECT 5739.04 307.445 5752.04 308.075 ;
      RECT 5739.04 211.445 5741.795 308.075 ;
      RECT 5739.04 228.445 5752.04 291.075 ;
      RECT 5739.04 211.445 5752.04 212.075 ;
      RECT 5742.035 189.04 5752.04 212.075 ;
      RECT 5739.04 189.04 5752.04 195.075 ;
      RECT 5705.08 324.445 5718.08 350.165 ;
      RECT 5705.08 228.445 5715.795 350.165 ;
      RECT 5710.31 211.445 5718.08 308.075 ;
      RECT 5705.08 189.04 5713.125 212.075 ;
      RECT 5705.08 189.04 5718.08 195.075 ;
      RECT 5674.56 290.445 5702.56 350.165 ;
      RECT 5693.19 189.04 5702.56 350.165 ;
      RECT 5691.425 194.425 5702.56 350.165 ;
      RECT 5674.56 189.04 5683.675 350.165 ;
      RECT 5674.56 194.425 5702.56 259.875 ;
      RECT 5674.56 189.04 5690.41 259.875 ;
      RECT 5674.56 189.04 5702.56 190.125 ;
      RECT 5659.04 211.445 5672.04 350.165 ;
      RECT 5665.425 189.04 5672.04 350.165 ;
      RECT 5659.04 189.04 5660.515 350.165 ;
      RECT 5659.04 189.04 5672.04 195.075 ;
      RECT 5642.06 259.445 5655.06 330.165 ;
      RECT 5646.935 189.04 5655.06 330.165 ;
      RECT 5642.06 189.04 5655.06 228.875 ;
      RECT 5625.08 307.445 5638.08 350.165 ;
      RECT 5633.09 189.04 5638.08 350.165 ;
      RECT 5629.035 194.37 5638.08 350.165 ;
      RECT 5625.08 228.445 5638.08 291.075 ;
      RECT 5625.08 194.37 5638.08 212.075 ;
      RECT 5625.08 189.04 5627.37 212.075 ;
      RECT 5625.08 189.04 5638.08 190.38 ;
      RECT 5594.56 324.445 5622.56 350.165 ;
      RECT 5606.705 189.04 5622.56 350.165 ;
      RECT 5602.035 307.445 5622.56 350.165 ;
      RECT 5594.56 189.04 5597.125 350.165 ;
      RECT 5594.56 307.445 5622.56 308.075 ;
      RECT 5594.56 211.445 5601.795 308.075 ;
      RECT 5594.56 228.445 5622.56 291.075 ;
      RECT 5594.56 211.445 5622.56 212.075 ;
      RECT 5602.035 189.04 5622.56 212.075 ;
      RECT 5594.56 189.04 5622.56 195.075 ;
      RECT 5579.04 324.445 5592.04 350.165 ;
      RECT 5580.705 189.04 5592.04 350.165 ;
      RECT 5579.04 189.04 5592.04 308.075 ;
      RECT 5562.06 228.445 5575.06 330.165 ;
      RECT 5568.69 211.445 5575.06 330.165 ;
      RECT 5562.06 189.04 5572.015 212.075 ;
      RECT 5562.06 189.04 5575.06 195.075 ;
      RECT 5545.08 290.445 5558.08 350.165 ;
      RECT 5553.19 189.04 5558.08 350.165 ;
      RECT 5551.425 194.425 5558.08 350.165 ;
      RECT 5545.08 194.425 5558.08 259.875 ;
      RECT 5545.08 189.04 5550.41 259.875 ;
      RECT 5545.08 189.04 5558.08 190.125 ;
      RECT 5514.56 211.445 5542.56 350.165 ;
      RECT 5525.425 189.04 5542.56 350.165 ;
      RECT 5514.56 189.04 5520.515 350.165 ;
      RECT 5514.56 189.04 5542.56 195.075 ;
      RECT 5499.04 259.445 5512.04 350.165 ;
      RECT 5506.935 189.04 5512.04 350.165 ;
      RECT 5499.04 189.04 5512.04 228.875 ;
      RECT 5482.06 307.445 5495.06 330.165 ;
      RECT 5492.99 189.04 5495.06 330.165 ;
      RECT 5489.035 194.37 5495.06 330.165 ;
      RECT 5482.06 189.04 5484.125 330.165 ;
      RECT 5482.06 228.445 5495.06 291.075 ;
      RECT 5482.06 194.37 5495.06 212.075 ;
      RECT 5482.06 189.04 5487.37 212.075 ;
      RECT 5482.06 189.04 5495.06 190.17 ;
      RECT 5465.08 307.445 5478.08 350.165 ;
      RECT 5466.705 189.04 5478.08 350.165 ;
      RECT 5465.08 228.445 5478.08 291.075 ;
      RECT 5465.08 189.04 5478.08 212.075 ;
      RECT 5434.56 324.445 5462.56 350.165 ;
      RECT 5440.705 189.04 5457.125 350.165 ;
      RECT 5434.56 211.445 5435.795 350.165 ;
      RECT 5434.56 211.445 5461.795 308.075 ;
      RECT 5434.56 228.445 5462.56 291.075 ;
      RECT 5436.925 189.04 5457.125 308.075 ;
      RECT 5434.56 189.04 5462.56 195.075 ;
      RECT 5419.04 228.445 5432.04 350.165 ;
      RECT 5419.04 189.04 5425.395 350.165 ;
      RECT 5419.04 189.04 5432.04 212.075 ;
      RECT 5402.06 290.445 5415.06 330.165 ;
      RECT 5413.19 189.04 5415.06 330.165 ;
      RECT 5411.425 194.425 5415.06 330.165 ;
      RECT 5402.06 189.04 5403.675 330.165 ;
      RECT 5402.06 194.425 5415.06 259.875 ;
      RECT 5402.06 189.04 5410.41 259.875 ;
      RECT 5402.06 189.04 5415.06 190.125 ;
      RECT 5385.08 211.445 5398.08 350.165 ;
      RECT 5385.425 189.04 5398.08 350.165 ;
      RECT 5385.08 189.04 5398.08 195.075 ;
      RECT 5354.56 259.445 5382.56 350.165 ;
      RECT 5366.935 211.445 5382.56 350.165 ;
      RECT 5354.56 189.04 5359.185 350.165 ;
      RECT 5354.56 189.04 5380.515 228.875 ;
      RECT 5354.56 189.04 5382.56 195.075 ;
      RECT 5339.04 307.445 5352.04 350.165 ;
      RECT 5349.035 194.37 5352.04 350.165 ;
      RECT 5339.04 189.04 5344.125 350.165 ;
      RECT 5339.04 228.445 5352.04 291.075 ;
      RECT 5339.04 194.37 5352.04 212.075 ;
      RECT 5339.04 189.04 5347.37 212.075 ;
      RECT 5339.04 189.04 5352.04 190.17 ;
      RECT 5322.06 307.445 5335.06 330.165 ;
      RECT 5326.705 189.04 5335.06 330.165 ;
      RECT 5326.54 228.445 5335.06 330.165 ;
      RECT 5322.06 228.445 5335.06 291.075 ;
      RECT 5322.06 189.04 5335.06 212.075 ;
      RECT 5305.08 324.445 5318.08 350.165 ;
      RECT 5305.08 189.04 5317.125 350.165 ;
      RECT 5305.08 211.445 5318.08 308.075 ;
      RECT 5305.08 189.04 5318.08 195.075 ;
      RECT 5274.56 324.445 5302.56 350.165 ;
      RECT 5300.705 189.04 5302.56 350.165 ;
      RECT 5274.56 228.445 5295.795 350.165 ;
      RECT 5298.115 189.04 5302.56 308.075 ;
      RECT 5281.11 211.445 5302.56 308.075 ;
      RECT 5274.56 189.04 5293.205 212.075 ;
      RECT 5274.56 189.04 5302.56 195.075 ;
      RECT 5259.04 290.445 5272.04 350.165 ;
      RECT 5271.425 194.42 5272.04 350.165 ;
      RECT 5259.04 189.04 5263.675 350.165 ;
      RECT 5259.04 194.42 5272.04 259.875 ;
      RECT 5259.04 189.04 5270.41 259.875 ;
      RECT 5259.04 189.04 5272.04 190.125 ;
      RECT 5242.06 211.445 5255.06 330.165 ;
      RECT 5245.425 189.04 5255.06 330.165 ;
      RECT 5242.06 189.04 5255.06 195.075 ;
      RECT 5225.08 259.445 5238.08 350.165 ;
      RECT 5226.935 189.04 5238.08 350.165 ;
      RECT 5225.08 189.04 5238.08 228.875 ;
      RECT 5194.56 307.445 5222.56 350.165 ;
      RECT 5209.035 259.445 5222.56 350.165 ;
      RECT 5194.56 189.04 5204.125 350.165 ;
      RECT 5194.56 228.445 5219.185 291.075 ;
      RECT 5213.09 189.04 5222.56 228.875 ;
      RECT 5209.035 194.37 5222.56 228.875 ;
      RECT 5194.56 194.37 5222.56 212.075 ;
      RECT 5194.56 189.04 5207.37 212.075 ;
      RECT 5194.56 189.04 5222.56 190.17 ;
      RECT 5179.04 324.445 5192.04 350.165 ;
      RECT 5186.705 189.04 5192.04 350.165 ;
      RECT 5182.035 307.445 5192.04 350.165 ;
      RECT 5179.04 307.445 5192.04 308.075 ;
      RECT 5179.04 211.445 5181.795 308.075 ;
      RECT 5179.04 228.445 5192.04 291.075 ;
      RECT 5179.04 211.445 5192.04 212.075 ;
      RECT 5182.035 189.04 5192.04 212.075 ;
      RECT 5179.04 189.04 5192.04 195.075 ;
      RECT 5145.08 324.445 5158.08 350.165 ;
      RECT 5145.08 228.445 5155.795 350.165 ;
      RECT 5150.31 211.445 5158.08 308.075 ;
      RECT 5145.08 189.04 5153.125 212.075 ;
      RECT 5145.08 189.04 5158.08 195.075 ;
      RECT 5114.56 290.445 5142.56 350.165 ;
      RECT 5133.19 189.04 5142.56 350.165 ;
      RECT 5131.425 194.425 5142.56 350.165 ;
      RECT 5114.56 189.04 5123.675 350.165 ;
      RECT 5114.56 194.425 5142.56 259.875 ;
      RECT 5114.56 189.04 5130.41 259.875 ;
      RECT 5114.56 189.04 5142.56 190.125 ;
      RECT 5099.04 211.445 5112.04 350.165 ;
      RECT 5105.425 189.04 5112.04 350.165 ;
      RECT 5099.04 189.04 5100.515 350.165 ;
      RECT 5099.04 189.04 5112.04 195.075 ;
      RECT 5082.06 259.445 5095.06 330.165 ;
      RECT 5086.935 189.04 5095.06 330.165 ;
      RECT 5082.06 189.04 5095.06 228.875 ;
      RECT 5065.08 307.445 5078.08 350.165 ;
      RECT 5073.09 189.04 5078.08 350.165 ;
      RECT 5069.035 194.37 5078.08 350.165 ;
      RECT 5065.08 228.445 5078.08 291.075 ;
      RECT 5065.08 194.37 5078.08 212.075 ;
      RECT 5065.08 189.04 5067.37 212.075 ;
      RECT 5065.08 189.04 5078.08 190.38 ;
      RECT 5034.56 324.445 5062.56 350.165 ;
      RECT 5046.705 189.04 5062.56 350.165 ;
      RECT 5042.035 307.445 5062.56 350.165 ;
      RECT 5034.56 189.04 5037.125 350.165 ;
      RECT 5034.56 307.445 5062.56 308.075 ;
      RECT 5034.56 211.445 5041.795 308.075 ;
      RECT 5034.56 228.445 5062.56 291.075 ;
      RECT 5034.56 211.445 5062.56 212.075 ;
      RECT 5042.035 189.04 5062.56 212.075 ;
      RECT 5034.56 189.04 5062.56 195.075 ;
      RECT 5019.04 324.445 5032.04 350.165 ;
      RECT 5020.705 189.04 5032.04 350.165 ;
      RECT 5019.04 189.04 5032.04 308.075 ;
      RECT 5002.06 228.445 5015.06 330.165 ;
      RECT 5008.69 211.445 5015.06 330.165 ;
      RECT 5002.06 189.04 5012.015 212.075 ;
      RECT 5002.06 189.04 5015.06 195.075 ;
      RECT 4985.08 290.445 4998.08 350.165 ;
      RECT 4993.19 189.04 4998.08 350.165 ;
      RECT 4991.425 194.425 4998.08 350.165 ;
      RECT 4985.08 194.425 4998.08 259.875 ;
      RECT 4985.08 189.04 4990.41 259.875 ;
      RECT 4985.08 189.04 4998.08 190.125 ;
      RECT 4954.56 211.445 4982.56 350.165 ;
      RECT 4965.425 189.04 4982.56 350.165 ;
      RECT 4954.56 189.04 4960.515 350.165 ;
      RECT 4954.56 189.04 4982.56 195.075 ;
      RECT 4939.04 259.445 4952.04 350.165 ;
      RECT 4946.935 189.04 4952.04 350.165 ;
      RECT 4939.04 189.04 4952.04 228.875 ;
      RECT 4922.06 307.445 4935.06 330.165 ;
      RECT 4932.99 189.04 4935.06 330.165 ;
      RECT 4929.035 194.37 4935.06 330.165 ;
      RECT 4922.06 189.04 4924.125 330.165 ;
      RECT 4922.06 228.445 4935.06 291.075 ;
      RECT 4922.06 194.37 4935.06 212.075 ;
      RECT 4922.06 189.04 4927.37 212.075 ;
      RECT 4922.06 189.04 4935.06 190.17 ;
      RECT 4905.08 307.445 4918.08 350.165 ;
      RECT 4906.705 189.04 4918.08 350.165 ;
      RECT 4905.08 228.445 4918.08 291.075 ;
      RECT 4905.08 189.04 4918.08 212.075 ;
      RECT 4874.56 324.445 4902.56 350.165 ;
      RECT 4880.705 189.04 4897.125 350.165 ;
      RECT 4874.56 211.445 4875.795 350.165 ;
      RECT 4874.56 211.445 4901.795 308.075 ;
      RECT 4874.56 228.445 4902.56 291.075 ;
      RECT 4876.925 189.04 4897.125 308.075 ;
      RECT 4874.56 189.04 4902.56 195.075 ;
      RECT 4859.04 228.445 4872.04 350.165 ;
      RECT 4859.04 189.04 4865.395 350.165 ;
      RECT 4859.04 189.04 4872.04 212.075 ;
      RECT 4842.06 290.445 4855.06 330.165 ;
      RECT 4853.19 189.04 4855.06 330.165 ;
      RECT 4851.425 194.425 4855.06 330.165 ;
      RECT 4842.06 189.04 4843.675 330.165 ;
      RECT 4842.06 194.425 4855.06 259.875 ;
      RECT 4842.06 189.04 4850.41 259.875 ;
      RECT 4842.06 189.04 4855.06 190.125 ;
      RECT 4825.08 211.445 4838.08 350.165 ;
      RECT 4825.425 189.04 4838.08 350.165 ;
      RECT 4825.08 189.04 4838.08 195.075 ;
      RECT 4794.56 259.445 4822.56 350.165 ;
      RECT 4806.935 211.445 4822.56 350.165 ;
      RECT 4794.56 189.04 4799.185 350.165 ;
      RECT 4794.56 189.04 4820.515 228.875 ;
      RECT 4794.56 189.04 4822.56 195.075 ;
      RECT 4779.04 307.445 4792.04 350.165 ;
      RECT 4789.035 194.37 4792.04 350.165 ;
      RECT 4779.04 189.04 4784.125 350.165 ;
      RECT 4779.04 228.445 4792.04 291.075 ;
      RECT 4779.04 194.37 4792.04 212.075 ;
      RECT 4779.04 189.04 4787.37 212.075 ;
      RECT 4779.04 189.04 4792.04 190.17 ;
      RECT 4762.06 307.445 4775.06 330.165 ;
      RECT 4766.705 189.04 4775.06 330.165 ;
      RECT 4766.54 228.445 4775.06 330.165 ;
      RECT 4762.06 228.445 4775.06 291.075 ;
      RECT 4762.06 189.04 4775.06 212.075 ;
      RECT 4745.08 324.445 4758.08 350.165 ;
      RECT 4745.08 189.04 4757.125 350.165 ;
      RECT 4745.08 211.445 4758.08 308.075 ;
      RECT 4745.08 189.04 4758.08 195.075 ;
      RECT 4714.56 324.445 4742.56 350.165 ;
      RECT 4740.705 189.04 4742.56 350.165 ;
      RECT 4714.56 228.445 4735.795 350.165 ;
      RECT 4738.115 189.04 4742.56 308.075 ;
      RECT 4721.11 211.445 4742.56 308.075 ;
      RECT 4714.56 189.04 4733.205 212.075 ;
      RECT 4714.56 189.04 4742.56 195.075 ;
      RECT 4699.04 290.445 4712.04 350.165 ;
      RECT 4711.425 194.42 4712.04 350.165 ;
      RECT 4699.04 189.04 4703.675 350.165 ;
      RECT 4699.04 194.42 4712.04 259.875 ;
      RECT 4699.04 189.04 4710.41 259.875 ;
      RECT 4699.04 189.04 4712.04 190.125 ;
      RECT 4682.06 211.445 4695.06 330.165 ;
      RECT 4685.425 189.04 4695.06 330.165 ;
      RECT 4682.06 189.04 4695.06 195.075 ;
      RECT 4665.08 259.445 4678.08 350.165 ;
      RECT 4666.935 189.04 4678.08 350.165 ;
      RECT 4665.08 189.04 4678.08 228.875 ;
      RECT 4634.56 307.445 4662.56 350.165 ;
      RECT 4649.035 259.445 4662.56 350.165 ;
      RECT 4634.56 189.04 4644.125 350.165 ;
      RECT 4634.56 228.445 4659.185 291.075 ;
      RECT 4653.09 189.04 4662.56 228.875 ;
      RECT 4649.035 194.37 4662.56 228.875 ;
      RECT 4634.56 194.37 4662.56 212.075 ;
      RECT 4634.56 189.04 4647.37 212.075 ;
      RECT 4634.56 189.04 4662.56 190.17 ;
      RECT 4619.04 324.445 4632.04 350.165 ;
      RECT 4626.705 189.04 4632.04 350.165 ;
      RECT 4622.035 307.445 4632.04 350.165 ;
      RECT 4619.04 307.445 4632.04 308.075 ;
      RECT 4619.04 211.445 4621.795 308.075 ;
      RECT 4619.04 228.445 4632.04 291.075 ;
      RECT 4619.04 211.445 4632.04 212.075 ;
      RECT 4622.035 189.04 4632.04 212.075 ;
      RECT 4619.04 189.04 4632.04 195.075 ;
      RECT 4585.08 324.445 4598.08 350.165 ;
      RECT 4585.08 228.445 4595.795 350.165 ;
      RECT 4590.31 211.445 4598.08 308.075 ;
      RECT 4585.08 189.04 4593.125 212.075 ;
      RECT 4585.08 189.04 4598.08 195.075 ;
      RECT 4554.56 290.445 4582.56 350.165 ;
      RECT 4573.19 189.04 4582.56 350.165 ;
      RECT 4571.425 194.425 4582.56 350.165 ;
      RECT 4554.56 189.04 4563.675 350.165 ;
      RECT 4554.56 194.425 4582.56 259.875 ;
      RECT 4554.56 189.04 4570.41 259.875 ;
      RECT 4554.56 189.04 4582.56 190.125 ;
      RECT 4539.04 211.445 4552.04 350.165 ;
      RECT 4545.425 189.04 4552.04 350.165 ;
      RECT 4539.04 189.04 4540.515 350.165 ;
      RECT 4539.04 189.04 4552.04 195.075 ;
      RECT 4522.06 259.445 4535.06 330.165 ;
      RECT 4526.935 189.04 4535.06 330.165 ;
      RECT 4522.06 189.04 4535.06 228.875 ;
      RECT 4505.08 307.445 4518.08 350.165 ;
      RECT 4513.09 189.04 4518.08 350.165 ;
      RECT 4509.035 194.37 4518.08 350.165 ;
      RECT 4505.08 228.445 4518.08 291.075 ;
      RECT 4505.08 194.37 4518.08 212.075 ;
      RECT 4505.08 189.04 4507.37 212.075 ;
      RECT 4505.08 189.04 4518.08 190.38 ;
      RECT 4474.56 324.445 4502.56 350.165 ;
      RECT 4486.705 189.04 4502.56 350.165 ;
      RECT 4482.035 307.445 4502.56 350.165 ;
      RECT 4474.56 189.04 4477.125 350.165 ;
      RECT 4474.56 307.445 4502.56 308.075 ;
      RECT 4474.56 211.445 4481.795 308.075 ;
      RECT 4474.56 228.445 4502.56 291.075 ;
      RECT 4474.56 211.445 4502.56 212.075 ;
      RECT 4482.035 189.04 4502.56 212.075 ;
      RECT 4474.56 189.04 4502.56 195.075 ;
      RECT 4459.04 324.445 4472.04 350.165 ;
      RECT 4460.705 189.04 4472.04 350.165 ;
      RECT 4459.04 189.04 4472.04 308.075 ;
      RECT 4442.06 228.445 4455.06 330.165 ;
      RECT 4448.69 211.445 4455.06 330.165 ;
      RECT 4442.06 189.04 4452.015 212.075 ;
      RECT 4442.06 189.04 4455.06 195.075 ;
      RECT 4425.08 290.445 4438.08 350.165 ;
      RECT 4433.19 189.04 4438.08 350.165 ;
      RECT 4431.425 194.425 4438.08 350.165 ;
      RECT 4425.08 194.425 4438.08 259.875 ;
      RECT 4425.08 189.04 4430.41 259.875 ;
      RECT 4425.08 189.04 4438.08 190.125 ;
      RECT 4394.56 211.445 4422.56 350.165 ;
      RECT 4405.425 189.04 4422.56 350.165 ;
      RECT 4394.56 189.04 4400.515 350.165 ;
      RECT 4394.56 189.04 4422.56 195.075 ;
      RECT 4379.04 259.445 4392.04 350.165 ;
      RECT 4386.935 189.04 4392.04 350.165 ;
      RECT 4379.04 189.04 4392.04 228.875 ;
      RECT 4362.06 307.445 4375.06 330.165 ;
      RECT 4372.99 189.04 4375.06 330.165 ;
      RECT 4369.035 194.37 4375.06 330.165 ;
      RECT 4362.06 189.04 4364.125 330.165 ;
      RECT 4362.06 228.445 4375.06 291.075 ;
      RECT 4362.06 194.37 4375.06 212.075 ;
      RECT 4362.06 189.04 4367.37 212.075 ;
      RECT 4362.06 189.04 4375.06 190.17 ;
      RECT 4345.08 307.445 4358.08 350.165 ;
      RECT 4346.705 189.04 4358.08 350.165 ;
      RECT 4345.08 228.445 4358.08 291.075 ;
      RECT 4345.08 189.04 4358.08 212.075 ;
      RECT 4314.56 324.445 4342.56 350.165 ;
      RECT 4320.705 189.04 4337.125 350.165 ;
      RECT 4314.56 211.445 4315.795 350.165 ;
      RECT 4314.56 211.445 4341.795 308.075 ;
      RECT 4314.56 228.445 4342.56 291.075 ;
      RECT 4316.925 189.04 4337.125 308.075 ;
      RECT 4314.56 189.04 4342.56 195.075 ;
      RECT 4299.04 228.445 4312.04 350.165 ;
      RECT 4299.04 189.04 4305.395 350.165 ;
      RECT 4299.04 189.04 4312.04 212.075 ;
      RECT 4282.06 290.445 4295.06 330.165 ;
      RECT 4293.19 189.04 4295.06 330.165 ;
      RECT 4291.425 194.425 4295.06 330.165 ;
      RECT 4282.06 189.04 4283.675 330.165 ;
      RECT 4282.06 194.425 4295.06 259.875 ;
      RECT 4282.06 189.04 4290.41 259.875 ;
      RECT 4282.06 189.04 4295.06 190.125 ;
      RECT 4265.08 211.445 4278.08 350.165 ;
      RECT 4265.425 189.04 4278.08 350.165 ;
      RECT 4265.08 189.04 4278.08 195.075 ;
      RECT 4234.56 259.445 4262.56 350.165 ;
      RECT 4246.935 211.445 4262.56 350.165 ;
      RECT 4234.56 189.04 4239.185 350.165 ;
      RECT 4234.56 189.04 4260.515 228.875 ;
      RECT 4234.56 189.04 4262.56 195.075 ;
      RECT 4219.04 307.445 4232.04 350.165 ;
      RECT 4229.035 194.37 4232.04 350.165 ;
      RECT 4219.04 189.04 4224.125 350.165 ;
      RECT 4219.04 228.445 4232.04 291.075 ;
      RECT 4219.04 194.37 4232.04 212.075 ;
      RECT 4219.04 189.04 4227.37 212.075 ;
      RECT 4219.04 189.04 4232.04 190.17 ;
      RECT 4202.06 307.445 4215.06 330.165 ;
      RECT 4206.705 189.04 4215.06 330.165 ;
      RECT 4206.54 228.445 4215.06 330.165 ;
      RECT 4202.06 228.445 4215.06 291.075 ;
      RECT 4202.06 189.04 4215.06 212.075 ;
      RECT 4185.08 324.445 4198.08 350.165 ;
      RECT 4185.08 189.04 4197.125 350.165 ;
      RECT 4185.08 211.445 4198.08 308.075 ;
      RECT 4185.08 189.04 4198.08 195.075 ;
      RECT 4154.56 324.445 4182.56 350.165 ;
      RECT 4180.705 189.04 4182.56 350.165 ;
      RECT 4154.56 228.445 4175.795 350.165 ;
      RECT 4178.115 189.04 4182.56 308.075 ;
      RECT 4161.11 211.445 4182.56 308.075 ;
      RECT 4154.56 189.04 4173.205 212.075 ;
      RECT 4154.56 189.04 4182.56 195.075 ;
      RECT 4139.04 290.445 4152.04 350.165 ;
      RECT 4151.425 194.42 4152.04 350.165 ;
      RECT 4139.04 189.04 4143.675 350.165 ;
      RECT 4139.04 194.42 4152.04 259.875 ;
      RECT 4139.04 189.04 4150.41 259.875 ;
      RECT 4139.04 189.04 4152.04 190.125 ;
      RECT 4122.06 211.445 4135.06 330.165 ;
      RECT 4125.425 189.04 4135.06 330.165 ;
      RECT 4122.06 189.04 4135.06 195.075 ;
      RECT 4105.08 259.445 4118.08 350.165 ;
      RECT 4106.935 189.04 4118.08 350.165 ;
      RECT 4105.08 189.04 4118.08 228.875 ;
      RECT 4074.56 307.445 4102.56 350.165 ;
      RECT 4089.035 259.445 4102.56 350.165 ;
      RECT 4074.56 189.04 4084.125 350.165 ;
      RECT 4074.56 228.445 4099.185 291.075 ;
      RECT 4093.09 189.04 4102.56 228.875 ;
      RECT 4089.035 194.37 4102.56 228.875 ;
      RECT 4074.56 194.37 4102.56 212.075 ;
      RECT 4074.56 189.04 4087.37 212.075 ;
      RECT 4074.56 189.04 4102.56 190.17 ;
      RECT 4059.04 324.445 4072.04 350.165 ;
      RECT 4066.705 189.04 4072.04 350.165 ;
      RECT 4062.035 307.445 4072.04 350.165 ;
      RECT 4059.04 307.445 4072.04 308.075 ;
      RECT 4059.04 211.445 4061.795 308.075 ;
      RECT 4059.04 228.445 4072.04 291.075 ;
      RECT 4059.04 211.445 4072.04 212.075 ;
      RECT 4062.035 189.04 4072.04 212.075 ;
      RECT 4059.04 189.04 4072.04 195.075 ;
      RECT 4025.08 324.445 4038.08 350.165 ;
      RECT 4025.08 228.445 4035.795 350.165 ;
      RECT 4030.31 211.445 4038.08 308.075 ;
      RECT 4025.08 189.04 4033.125 212.075 ;
      RECT 4025.08 189.04 4038.08 195.075 ;
      RECT 3994.56 290.445 4022.56 350.165 ;
      RECT 4013.19 189.04 4022.56 350.165 ;
      RECT 4011.425 194.425 4022.56 350.165 ;
      RECT 3994.56 189.04 4003.675 350.165 ;
      RECT 3994.56 194.425 4022.56 259.875 ;
      RECT 3994.56 189.04 4010.41 259.875 ;
      RECT 3994.56 189.04 4022.56 190.125 ;
      RECT 3979.04 211.445 3992.04 350.165 ;
      RECT 3985.425 189.04 3992.04 350.165 ;
      RECT 3979.04 189.04 3980.515 350.165 ;
      RECT 3979.04 189.04 3992.04 195.075 ;
      RECT 3962.06 259.445 3975.06 330.165 ;
      RECT 3966.935 189.04 3975.06 330.165 ;
      RECT 3962.06 189.04 3975.06 228.875 ;
      RECT 3945.08 307.445 3958.08 350.165 ;
      RECT 3953.09 189.04 3958.08 350.165 ;
      RECT 3949.035 194.37 3958.08 350.165 ;
      RECT 3945.08 228.445 3958.08 291.075 ;
      RECT 3945.08 194.37 3958.08 212.075 ;
      RECT 3945.08 189.04 3947.37 212.075 ;
      RECT 3945.08 189.04 3958.08 190.38 ;
      RECT 3914.56 324.445 3942.56 350.165 ;
      RECT 3926.705 189.04 3942.56 350.165 ;
      RECT 3922.035 307.445 3942.56 350.165 ;
      RECT 3914.56 189.04 3917.125 350.165 ;
      RECT 3914.56 307.445 3942.56 308.075 ;
      RECT 3914.56 211.445 3921.795 308.075 ;
      RECT 3914.56 228.445 3942.56 291.075 ;
      RECT 3914.56 211.445 3942.56 212.075 ;
      RECT 3922.035 189.04 3942.56 212.075 ;
      RECT 3914.56 189.04 3942.56 195.075 ;
      RECT 3899.04 324.445 3912.04 350.165 ;
      RECT 3900.705 189.04 3912.04 350.165 ;
      RECT 3899.04 189.04 3912.04 308.075 ;
      RECT 3882.06 228.445 3895.06 330.165 ;
      RECT 3888.69 211.445 3895.06 330.165 ;
      RECT 3882.06 189.04 3892.015 212.075 ;
      RECT 3882.06 189.04 3895.06 195.075 ;
      RECT 3865.08 290.445 3878.08 350.165 ;
      RECT 3873.19 189.04 3878.08 350.165 ;
      RECT 3871.425 194.425 3878.08 350.165 ;
      RECT 3865.08 194.425 3878.08 259.875 ;
      RECT 3865.08 189.04 3870.41 259.875 ;
      RECT 3865.08 189.04 3878.08 190.125 ;
      RECT 3834.56 211.445 3862.56 350.165 ;
      RECT 3845.425 189.04 3862.56 350.165 ;
      RECT 3834.56 189.04 3840.515 350.165 ;
      RECT 3834.56 189.04 3862.56 195.075 ;
      RECT 3819.04 259.445 3832.04 350.165 ;
      RECT 3826.935 189.04 3832.04 350.165 ;
      RECT 3819.04 189.04 3832.04 228.875 ;
      RECT 3802.06 307.445 3815.06 330.165 ;
      RECT 3812.99 189.04 3815.06 330.165 ;
      RECT 3809.035 194.37 3815.06 330.165 ;
      RECT 3802.06 189.04 3804.125 330.165 ;
      RECT 3802.06 228.445 3815.06 291.075 ;
      RECT 3802.06 194.37 3815.06 212.075 ;
      RECT 3802.06 189.04 3807.37 212.075 ;
      RECT 3802.06 189.04 3815.06 190.17 ;
      RECT 3785.08 307.445 3798.08 350.165 ;
      RECT 3786.705 189.04 3798.08 350.165 ;
      RECT 3785.08 228.445 3798.08 291.075 ;
      RECT 3785.08 189.04 3798.08 212.075 ;
      RECT 3754.56 324.445 3782.56 350.165 ;
      RECT 3760.705 189.04 3777.125 350.165 ;
      RECT 3754.56 211.445 3755.795 350.165 ;
      RECT 3754.56 211.445 3781.795 308.075 ;
      RECT 3754.56 228.445 3782.56 291.075 ;
      RECT 3756.925 189.04 3777.125 308.075 ;
      RECT 3754.56 189.04 3782.56 195.075 ;
      RECT 3739.04 228.445 3752.04 350.165 ;
      RECT 3739.04 189.04 3745.395 350.165 ;
      RECT 3739.04 189.04 3752.04 212.075 ;
      RECT 3722.06 290.445 3735.06 330.165 ;
      RECT 3733.19 189.04 3735.06 330.165 ;
      RECT 3731.425 194.425 3735.06 330.165 ;
      RECT 3722.06 189.04 3723.675 330.165 ;
      RECT 3722.06 194.425 3735.06 259.875 ;
      RECT 3722.06 189.04 3730.41 259.875 ;
      RECT 3722.06 189.04 3735.06 190.125 ;
      RECT 3705.08 211.445 3718.08 350.165 ;
      RECT 3705.425 189.04 3718.08 350.165 ;
      RECT 3705.08 189.04 3718.08 195.075 ;
      RECT 3674.56 259.445 3702.56 350.165 ;
      RECT 3686.935 211.445 3702.56 350.165 ;
      RECT 3674.56 189.04 3679.185 350.165 ;
      RECT 3674.56 189.04 3700.515 228.875 ;
      RECT 3674.56 189.04 3702.56 195.075 ;
      RECT 3659.04 307.445 3672.04 350.165 ;
      RECT 3669.035 194.37 3672.04 350.165 ;
      RECT 3659.04 189.04 3664.125 350.165 ;
      RECT 3659.04 228.445 3672.04 291.075 ;
      RECT 3659.04 194.37 3672.04 212.075 ;
      RECT 3659.04 189.04 3667.37 212.075 ;
      RECT 3659.04 189.04 3672.04 190.17 ;
      RECT 3642.06 307.445 3655.06 330.165 ;
      RECT 3646.705 189.04 3655.06 330.165 ;
      RECT 3646.54 228.445 3655.06 330.165 ;
      RECT 3642.06 228.445 3655.06 291.075 ;
      RECT 3642.06 189.04 3655.06 212.075 ;
      RECT 3625.08 324.445 3638.08 350.165 ;
      RECT 3625.08 189.04 3637.125 350.165 ;
      RECT 3625.08 211.445 3638.08 308.075 ;
      RECT 3625.08 189.04 3638.08 195.075 ;
      RECT 3594.56 324.445 3622.56 350.165 ;
      RECT 3620.705 189.04 3622.56 350.165 ;
      RECT 3594.56 228.445 3615.795 350.165 ;
      RECT 3618.115 189.04 3622.56 308.075 ;
      RECT 3601.11 211.445 3622.56 308.075 ;
      RECT 3594.56 189.04 3613.205 212.075 ;
      RECT 3594.56 189.04 3622.56 195.075 ;
      RECT 3579.04 290.445 3592.04 350.165 ;
      RECT 3591.425 194.42 3592.04 350.165 ;
      RECT 3579.04 189.04 3583.675 350.165 ;
      RECT 3579.04 194.42 3592.04 259.875 ;
      RECT 3579.04 189.04 3590.41 259.875 ;
      RECT 3579.04 189.04 3592.04 190.125 ;
      RECT 3562.06 211.445 3575.06 330.165 ;
      RECT 3565.425 189.04 3575.06 330.165 ;
      RECT 3562.06 189.04 3575.06 195.075 ;
      RECT 3545.08 259.445 3558.08 350.165 ;
      RECT 3546.935 189.04 3558.08 350.165 ;
      RECT 3545.08 189.04 3558.08 228.875 ;
      RECT 3514.56 307.445 3542.56 350.165 ;
      RECT 3529.035 259.445 3542.56 350.165 ;
      RECT 3514.56 189.04 3524.125 350.165 ;
      RECT 3514.56 228.445 3539.185 291.075 ;
      RECT 3533.09 189.04 3542.56 228.875 ;
      RECT 3529.035 194.37 3542.56 228.875 ;
      RECT 3514.56 194.37 3542.56 212.075 ;
      RECT 3514.56 189.04 3527.37 212.075 ;
      RECT 3514.56 189.04 3542.56 190.17 ;
      RECT 3499.04 324.445 3512.04 350.165 ;
      RECT 3506.705 189.04 3512.04 350.165 ;
      RECT 3502.035 307.445 3512.04 350.165 ;
      RECT 3499.04 307.445 3512.04 308.075 ;
      RECT 3499.04 211.445 3501.795 308.075 ;
      RECT 3499.04 228.445 3512.04 291.075 ;
      RECT 3499.04 211.445 3512.04 212.075 ;
      RECT 3502.035 189.04 3512.04 212.075 ;
      RECT 3499.04 189.04 3512.04 195.075 ;
      RECT 3465.08 324.445 3478.08 350.165 ;
      RECT 3465.08 228.445 3475.795 350.165 ;
      RECT 3470.31 211.445 3478.08 308.075 ;
      RECT 3465.08 189.04 3473.125 212.075 ;
      RECT 3465.08 189.04 3478.08 195.075 ;
      RECT 3434.56 290.445 3462.56 350.165 ;
      RECT 3453.19 189.04 3462.56 350.165 ;
      RECT 3451.425 194.425 3462.56 350.165 ;
      RECT 3434.56 189.04 3443.675 350.165 ;
      RECT 3434.56 194.425 3462.56 259.875 ;
      RECT 3434.56 189.04 3450.41 259.875 ;
      RECT 3434.56 189.04 3462.56 190.125 ;
      RECT 3419.04 211.445 3432.04 350.165 ;
      RECT 3425.425 189.04 3432.04 350.165 ;
      RECT 3419.04 189.04 3420.515 350.165 ;
      RECT 3419.04 189.04 3432.04 195.075 ;
      RECT 3402.06 259.445 3415.06 330.165 ;
      RECT 3406.935 189.04 3415.06 330.165 ;
      RECT 3402.06 189.04 3415.06 228.875 ;
      RECT 3385.08 307.445 3398.08 350.165 ;
      RECT 3393.09 189.04 3398.08 350.165 ;
      RECT 3389.035 194.37 3398.08 350.165 ;
      RECT 3385.08 228.445 3398.08 291.075 ;
      RECT 3385.08 194.37 3398.08 212.075 ;
      RECT 3385.08 189.04 3387.37 212.075 ;
      RECT 3385.08 189.04 3398.08 190.38 ;
      RECT 3354.56 324.445 3382.56 350.165 ;
      RECT 3366.705 189.04 3382.56 350.165 ;
      RECT 3362.035 307.445 3382.56 350.165 ;
      RECT 3354.56 189.04 3357.125 350.165 ;
      RECT 3354.56 307.445 3382.56 308.075 ;
      RECT 3354.56 211.445 3361.795 308.075 ;
      RECT 3354.56 228.445 3382.56 291.075 ;
      RECT 3354.56 211.445 3382.56 212.075 ;
      RECT 3362.035 189.04 3382.56 212.075 ;
      RECT 3354.56 189.04 3382.56 195.075 ;
      RECT 3339.04 324.445 3352.04 350.165 ;
      RECT 3340.705 189.04 3352.04 350.165 ;
      RECT 3339.04 189.04 3352.04 308.075 ;
      RECT 3322.06 228.445 3335.06 330.165 ;
      RECT 3328.69 211.445 3335.06 330.165 ;
      RECT 3322.06 189.04 3332.015 212.075 ;
      RECT 3322.06 189.04 3335.06 195.075 ;
      RECT 3305.08 290.445 3318.08 350.165 ;
      RECT 3313.19 189.04 3318.08 350.165 ;
      RECT 3311.425 194.425 3318.08 350.165 ;
      RECT 3305.08 194.425 3318.08 259.875 ;
      RECT 3305.08 189.04 3310.41 259.875 ;
      RECT 3305.08 189.04 3318.08 190.125 ;
      RECT 3274.56 211.445 3302.56 350.165 ;
      RECT 3285.425 189.04 3302.56 350.165 ;
      RECT 3274.56 189.04 3280.515 350.165 ;
      RECT 3274.56 189.04 3302.56 195.075 ;
      RECT 3259.04 259.445 3272.04 350.165 ;
      RECT 3266.935 189.04 3272.04 350.165 ;
      RECT 3259.04 189.04 3272.04 228.875 ;
      RECT 3242.06 307.445 3255.06 330.165 ;
      RECT 3252.99 189.04 3255.06 330.165 ;
      RECT 3249.035 194.37 3255.06 330.165 ;
      RECT 3242.06 189.04 3244.125 330.165 ;
      RECT 3242.06 228.445 3255.06 291.075 ;
      RECT 3242.06 194.37 3255.06 212.075 ;
      RECT 3242.06 189.04 3247.37 212.075 ;
      RECT 3242.06 189.04 3255.06 190.17 ;
      RECT 3225.08 307.445 3238.08 350.165 ;
      RECT 3226.705 189.04 3238.08 350.165 ;
      RECT 3225.08 228.445 3238.08 291.075 ;
      RECT 3225.08 189.04 3238.08 212.075 ;
      RECT 3194.56 324.445 3222.56 350.165 ;
      RECT 3200.705 189.04 3217.125 350.165 ;
      RECT 3194.56 211.445 3195.795 350.165 ;
      RECT 3194.56 211.445 3221.795 308.075 ;
      RECT 3194.56 228.445 3222.56 291.075 ;
      RECT 3196.925 189.04 3217.125 308.075 ;
      RECT 3194.56 189.04 3222.56 195.075 ;
      RECT 3179.04 228.445 3192.04 350.165 ;
      RECT 3179.04 189.04 3185.395 350.165 ;
      RECT 3179.04 189.04 3192.04 212.075 ;
      RECT 3162.06 290.445 3175.06 330.165 ;
      RECT 3173.19 189.04 3175.06 330.165 ;
      RECT 3171.425 194.425 3175.06 330.165 ;
      RECT 3162.06 189.04 3163.675 330.165 ;
      RECT 3162.06 194.425 3175.06 259.875 ;
      RECT 3162.06 189.04 3170.41 259.875 ;
      RECT 3162.06 189.04 3175.06 190.125 ;
      RECT 3145.08 211.445 3158.08 350.165 ;
      RECT 3145.425 189.04 3158.08 350.165 ;
      RECT 3145.08 189.04 3158.08 195.075 ;
      RECT 3114.56 259.445 3142.56 350.165 ;
      RECT 3126.935 211.445 3142.56 350.165 ;
      RECT 3114.56 189.04 3119.185 350.165 ;
      RECT 3114.56 189.04 3140.515 228.875 ;
      RECT 3114.56 189.04 3142.56 195.075 ;
      RECT 3099.04 307.445 3112.04 350.165 ;
      RECT 3109.035 194.37 3112.04 350.165 ;
      RECT 3099.04 189.04 3104.125 350.165 ;
      RECT 3099.04 228.445 3112.04 291.075 ;
      RECT 3099.04 194.37 3112.04 212.075 ;
      RECT 3099.04 189.04 3107.37 212.075 ;
      RECT 3099.04 189.04 3112.04 190.17 ;
      RECT 3082.06 307.445 3095.06 330.165 ;
      RECT 3086.705 189.04 3095.06 330.165 ;
      RECT 3086.54 228.445 3095.06 330.165 ;
      RECT 3082.06 228.445 3095.06 291.075 ;
      RECT 3082.06 189.04 3095.06 212.075 ;
      RECT 3065.08 324.445 3078.08 350.165 ;
      RECT 3065.08 189.04 3077.125 350.165 ;
      RECT 3065.08 211.445 3078.08 308.075 ;
      RECT 3065.08 189.04 3078.08 195.075 ;
      RECT 3034.56 324.445 3062.56 350.165 ;
      RECT 3060.705 189.04 3062.56 350.165 ;
      RECT 3034.56 228.445 3055.795 350.165 ;
      RECT 3058.115 189.04 3062.56 308.075 ;
      RECT 3041.11 211.445 3062.56 308.075 ;
      RECT 3034.56 189.04 3053.205 212.075 ;
      RECT 3034.56 189.04 3062.56 195.075 ;
      RECT 3019.04 290.445 3032.04 350.165 ;
      RECT 3031.425 194.42 3032.04 350.165 ;
      RECT 3019.04 189.04 3023.675 350.165 ;
      RECT 3019.04 194.42 3032.04 259.875 ;
      RECT 3019.04 189.04 3030.41 259.875 ;
      RECT 3019.04 189.04 3032.04 190.125 ;
      RECT 3002.06 211.445 3015.06 330.165 ;
      RECT 3005.425 189.04 3015.06 330.165 ;
      RECT 3002.06 189.04 3015.06 195.075 ;
      RECT 2985.08 259.445 2998.08 350.165 ;
      RECT 2986.935 189.04 2998.08 350.165 ;
      RECT 2985.08 189.04 2998.08 228.875 ;
      RECT 2954.56 307.445 2982.56 350.165 ;
      RECT 2969.035 259.445 2982.56 350.165 ;
      RECT 2954.56 189.04 2964.125 350.165 ;
      RECT 2954.56 228.445 2979.185 291.075 ;
      RECT 2973.09 189.04 2982.56 228.875 ;
      RECT 2969.035 194.37 2982.56 228.875 ;
      RECT 2954.56 194.37 2982.56 212.075 ;
      RECT 2954.56 189.04 2967.37 212.075 ;
      RECT 2954.56 189.04 2982.56 190.17 ;
      RECT 2939.04 324.445 2952.04 350.165 ;
      RECT 2946.705 189.04 2952.04 350.165 ;
      RECT 2942.035 307.445 2952.04 350.165 ;
      RECT 2939.04 307.445 2952.04 308.075 ;
      RECT 2939.04 211.445 2941.795 308.075 ;
      RECT 2939.04 228.445 2952.04 291.075 ;
      RECT 2939.04 211.445 2952.04 212.075 ;
      RECT 2942.035 189.04 2952.04 212.075 ;
      RECT 2939.04 189.04 2952.04 195.075 ;
      RECT 2905.08 324.445 2918.08 350.165 ;
      RECT 2905.08 228.445 2915.795 350.165 ;
      RECT 2910.31 211.445 2918.08 308.075 ;
      RECT 2905.08 189.04 2913.125 212.075 ;
      RECT 2905.08 189.04 2918.08 195.075 ;
      RECT 2874.56 290.445 2902.56 350.165 ;
      RECT 2893.19 189.04 2902.56 350.165 ;
      RECT 2891.425 194.425 2902.56 350.165 ;
      RECT 2874.56 189.04 2883.675 350.165 ;
      RECT 2874.56 194.425 2902.56 259.875 ;
      RECT 2874.56 189.04 2890.41 259.875 ;
      RECT 2874.56 189.04 2902.56 190.125 ;
      RECT 2859.04 211.445 2872.04 350.165 ;
      RECT 2865.425 189.04 2872.04 350.165 ;
      RECT 2859.04 189.04 2860.515 350.165 ;
      RECT 2859.04 189.04 2872.04 195.075 ;
      RECT 2842.06 259.445 2855.06 330.165 ;
      RECT 2846.935 189.04 2855.06 330.165 ;
      RECT 2842.06 189.04 2855.06 228.875 ;
      RECT 2825.08 307.445 2838.08 350.165 ;
      RECT 2833.09 189.04 2838.08 350.165 ;
      RECT 2829.035 194.37 2838.08 350.165 ;
      RECT 2825.08 228.445 2838.08 291.075 ;
      RECT 2825.08 194.37 2838.08 212.075 ;
      RECT 2825.08 189.04 2827.37 212.075 ;
      RECT 2825.08 189.04 2838.08 190.38 ;
      RECT 2794.56 324.445 2822.56 350.165 ;
      RECT 2806.705 189.04 2822.56 350.165 ;
      RECT 2802.035 307.445 2822.56 350.165 ;
      RECT 2794.56 189.04 2797.125 350.165 ;
      RECT 2794.56 307.445 2822.56 308.075 ;
      RECT 2794.56 211.445 2801.795 308.075 ;
      RECT 2794.56 228.445 2822.56 291.075 ;
      RECT 2794.56 211.445 2822.56 212.075 ;
      RECT 2802.035 189.04 2822.56 212.075 ;
      RECT 2794.56 189.04 2822.56 195.075 ;
      RECT 2779.04 324.445 2792.04 350.165 ;
      RECT 2780.705 189.04 2792.04 350.165 ;
      RECT 2779.04 189.04 2792.04 308.075 ;
      RECT 2762.06 228.445 2775.06 330.165 ;
      RECT 2768.69 211.445 2775.06 330.165 ;
      RECT 2762.06 189.04 2772.015 212.075 ;
      RECT 2762.06 189.04 2775.06 195.075 ;
      RECT 2745.08 290.445 2758.08 350.165 ;
      RECT 2753.19 189.04 2758.08 350.165 ;
      RECT 2751.425 194.425 2758.08 350.165 ;
      RECT 2745.08 194.425 2758.08 259.875 ;
      RECT 2745.08 189.04 2750.41 259.875 ;
      RECT 2745.08 189.04 2758.08 190.125 ;
      RECT 2714.56 211.445 2742.56 350.165 ;
      RECT 2725.425 189.04 2742.56 350.165 ;
      RECT 2714.56 189.04 2720.515 350.165 ;
      RECT 2714.56 189.04 2742.56 195.075 ;
      RECT 2699.04 259.445 2712.04 350.165 ;
      RECT 2706.935 189.04 2712.04 350.165 ;
      RECT 2699.04 189.04 2712.04 228.875 ;
      RECT 2682.06 307.445 2695.06 330.165 ;
      RECT 2692.99 189.04 2695.06 330.165 ;
      RECT 2689.035 194.37 2695.06 330.165 ;
      RECT 2682.06 189.04 2684.125 330.165 ;
      RECT 2682.06 228.445 2695.06 291.075 ;
      RECT 2682.06 194.37 2695.06 212.075 ;
      RECT 2682.06 189.04 2687.37 212.075 ;
      RECT 2682.06 189.04 2695.06 190.17 ;
      RECT 2665.08 307.445 2678.08 350.165 ;
      RECT 2666.705 189.04 2678.08 350.165 ;
      RECT 2665.08 228.445 2678.08 291.075 ;
      RECT 2665.08 189.04 2678.08 212.075 ;
      RECT 2634.56 324.445 2662.56 350.165 ;
      RECT 2640.705 189.04 2657.125 350.165 ;
      RECT 2634.56 211.445 2635.795 350.165 ;
      RECT 2634.56 211.445 2661.795 308.075 ;
      RECT 2634.56 228.445 2662.56 291.075 ;
      RECT 2636.925 189.04 2657.125 308.075 ;
      RECT 2634.56 189.04 2662.56 195.075 ;
      RECT 2619.04 228.445 2632.04 350.165 ;
      RECT 2619.04 189.04 2625.395 350.165 ;
      RECT 2619.04 189.04 2632.04 212.075 ;
      RECT 2602.06 290.445 2615.06 330.165 ;
      RECT 2613.19 189.04 2615.06 330.165 ;
      RECT 2611.425 194.425 2615.06 330.165 ;
      RECT 2602.06 189.04 2603.675 330.165 ;
      RECT 2602.06 194.425 2615.06 259.875 ;
      RECT 2602.06 189.04 2610.41 259.875 ;
      RECT 2602.06 189.04 2615.06 190.125 ;
      RECT 2585.08 211.445 2598.08 350.165 ;
      RECT 2585.425 189.04 2598.08 350.165 ;
      RECT 2585.08 189.04 2598.08 195.075 ;
      RECT 2554.56 259.445 2582.56 350.165 ;
      RECT 2566.935 211.445 2582.56 350.165 ;
      RECT 2554.56 189.04 2559.185 350.165 ;
      RECT 2554.56 189.04 2580.515 228.875 ;
      RECT 2554.56 189.04 2582.56 195.075 ;
      RECT 2539.04 307.445 2552.04 350.165 ;
      RECT 2549.035 194.37 2552.04 350.165 ;
      RECT 2539.04 189.04 2544.125 350.165 ;
      RECT 2539.04 228.445 2552.04 291.075 ;
      RECT 2539.04 194.37 2552.04 212.075 ;
      RECT 2539.04 189.04 2547.37 212.075 ;
      RECT 2539.04 189.04 2552.04 190.17 ;
      RECT 2522.06 307.445 2535.06 330.165 ;
      RECT 2526.705 189.04 2535.06 330.165 ;
      RECT 2526.54 228.445 2535.06 330.165 ;
      RECT 2522.06 228.445 2535.06 291.075 ;
      RECT 2522.06 189.04 2535.06 212.075 ;
      RECT 2505.08 324.445 2518.08 350.165 ;
      RECT 2505.08 189.04 2517.125 350.165 ;
      RECT 2505.08 211.445 2518.08 308.075 ;
      RECT 2505.08 189.04 2518.08 195.075 ;
      RECT 2474.56 324.445 2502.56 350.165 ;
      RECT 2500.705 189.04 2502.56 350.165 ;
      RECT 2474.56 228.445 2495.795 350.165 ;
      RECT 2498.115 189.04 2502.56 308.075 ;
      RECT 2481.11 211.445 2502.56 308.075 ;
      RECT 2474.56 189.04 2493.205 212.075 ;
      RECT 2474.56 189.04 2502.56 195.075 ;
      RECT 2459.04 290.445 2472.04 350.165 ;
      RECT 2471.425 194.42 2472.04 350.165 ;
      RECT 2459.04 189.04 2463.675 350.165 ;
      RECT 2459.04 194.42 2472.04 259.875 ;
      RECT 2459.04 189.04 2470.41 259.875 ;
      RECT 2459.04 189.04 2472.04 190.125 ;
      RECT 2442.06 211.445 2455.06 330.165 ;
      RECT 2445.425 189.04 2455.06 330.165 ;
      RECT 2442.06 189.04 2455.06 195.075 ;
      RECT 2425.08 259.445 2438.08 350.165 ;
      RECT 2426.935 189.04 2438.08 350.165 ;
      RECT 2425.08 189.04 2438.08 228.875 ;
      RECT 2394.56 307.445 2422.56 350.165 ;
      RECT 2409.035 259.445 2422.56 350.165 ;
      RECT 2394.56 189.04 2404.125 350.165 ;
      RECT 2394.56 228.445 2419.185 291.075 ;
      RECT 2413.09 189.04 2422.56 228.875 ;
      RECT 2409.035 194.37 2422.56 228.875 ;
      RECT 2394.56 194.37 2422.56 212.075 ;
      RECT 2394.56 189.04 2407.37 212.075 ;
      RECT 2394.56 189.04 2422.56 190.17 ;
      RECT 2379.04 324.445 2392.04 350.165 ;
      RECT 2386.705 189.04 2392.04 350.165 ;
      RECT 2382.035 307.445 2392.04 350.165 ;
      RECT 2379.04 307.445 2392.04 308.075 ;
      RECT 2379.04 211.445 2381.795 308.075 ;
      RECT 2379.04 228.445 2392.04 291.075 ;
      RECT 2379.04 211.445 2392.04 212.075 ;
      RECT 2382.035 189.04 2392.04 212.075 ;
      RECT 2379.04 189.04 2392.04 195.075 ;
      RECT 2345.08 324.445 2358.08 350.165 ;
      RECT 2345.08 228.445 2355.795 350.165 ;
      RECT 2350.31 211.445 2358.08 308.075 ;
      RECT 2345.08 189.04 2353.125 212.075 ;
      RECT 2345.08 189.04 2358.08 195.075 ;
      RECT 2314.56 290.445 2342.56 350.165 ;
      RECT 2333.19 189.04 2342.56 350.165 ;
      RECT 2331.425 194.425 2342.56 350.165 ;
      RECT 2314.56 189.04 2323.675 350.165 ;
      RECT 2314.56 194.425 2342.56 259.875 ;
      RECT 2314.56 189.04 2330.41 259.875 ;
      RECT 2314.56 189.04 2342.56 190.125 ;
      RECT 2299.04 211.445 2312.04 350.165 ;
      RECT 2305.425 189.04 2312.04 350.165 ;
      RECT 2299.04 189.04 2300.515 350.165 ;
      RECT 2299.04 189.04 2312.04 195.075 ;
      RECT 2282.06 259.445 2295.06 330.165 ;
      RECT 2286.935 189.04 2295.06 330.165 ;
      RECT 2282.06 189.04 2295.06 228.875 ;
      RECT 2265.08 307.445 2278.08 350.165 ;
      RECT 2273.09 189.04 2278.08 350.165 ;
      RECT 2269.035 194.37 2278.08 350.165 ;
      RECT 2265.08 228.445 2278.08 291.075 ;
      RECT 2265.08 194.37 2278.08 212.075 ;
      RECT 2265.08 189.04 2267.37 212.075 ;
      RECT 2265.08 189.04 2278.08 190.38 ;
      RECT 2234.56 324.445 2262.56 350.165 ;
      RECT 2246.705 189.04 2262.56 350.165 ;
      RECT 2242.035 307.445 2262.56 350.165 ;
      RECT 2234.56 189.04 2237.125 350.165 ;
      RECT 2234.56 307.445 2262.56 308.075 ;
      RECT 2234.56 211.445 2241.795 308.075 ;
      RECT 2234.56 228.445 2262.56 291.075 ;
      RECT 2234.56 211.445 2262.56 212.075 ;
      RECT 2242.035 189.04 2262.56 212.075 ;
      RECT 2234.56 189.04 2262.56 195.075 ;
      RECT 2219.04 324.445 2232.04 350.165 ;
      RECT 2220.705 189.04 2232.04 350.165 ;
      RECT 2219.04 189.04 2232.04 308.075 ;
      RECT 2202.06 228.445 2215.06 330.165 ;
      RECT 2208.69 211.445 2215.06 330.165 ;
      RECT 2202.06 189.04 2212.015 212.075 ;
      RECT 2202.06 189.04 2215.06 195.075 ;
      RECT 2185.08 290.445 2198.08 350.165 ;
      RECT 2193.19 189.04 2198.08 350.165 ;
      RECT 2191.425 194.425 2198.08 350.165 ;
      RECT 2185.08 194.425 2198.08 259.875 ;
      RECT 2185.08 189.04 2190.41 259.875 ;
      RECT 2185.08 189.04 2198.08 190.125 ;
      RECT 2154.56 211.445 2182.56 350.165 ;
      RECT 2165.425 189.04 2182.56 350.165 ;
      RECT 2154.56 189.04 2160.515 350.165 ;
      RECT 2154.56 189.04 2182.56 195.075 ;
      RECT 2139.04 259.445 2152.04 350.165 ;
      RECT 2146.935 189.04 2152.04 350.165 ;
      RECT 2139.04 189.04 2152.04 228.875 ;
      RECT 2122.06 307.445 2135.06 330.165 ;
      RECT 2132.99 189.04 2135.06 330.165 ;
      RECT 2129.035 194.37 2135.06 330.165 ;
      RECT 2122.06 189.04 2124.125 330.165 ;
      RECT 2122.06 228.445 2135.06 291.075 ;
      RECT 2122.06 194.37 2135.06 212.075 ;
      RECT 2122.06 189.04 2127.37 212.075 ;
      RECT 2122.06 189.04 2135.06 190.17 ;
      RECT 2105.08 307.445 2118.08 350.165 ;
      RECT 2106.705 189.04 2118.08 350.165 ;
      RECT 2105.08 228.445 2118.08 291.075 ;
      RECT 2105.08 189.04 2118.08 212.075 ;
      RECT 2074.56 324.445 2102.56 350.165 ;
      RECT 2080.705 189.04 2097.125 350.165 ;
      RECT 2074.56 211.445 2075.795 350.165 ;
      RECT 2074.56 211.445 2101.795 308.075 ;
      RECT 2074.56 228.445 2102.56 291.075 ;
      RECT 2076.925 189.04 2097.125 308.075 ;
      RECT 2074.56 189.04 2102.56 195.075 ;
      RECT 2059.04 228.445 2072.04 350.165 ;
      RECT 2059.04 189.04 2065.395 350.165 ;
      RECT 2059.04 189.04 2072.04 212.075 ;
      RECT 2042.06 290.445 2055.06 330.165 ;
      RECT 2053.19 189.04 2055.06 330.165 ;
      RECT 2051.425 194.425 2055.06 330.165 ;
      RECT 2042.06 189.04 2043.675 330.165 ;
      RECT 2042.06 194.425 2055.06 259.875 ;
      RECT 2042.06 189.04 2050.41 259.875 ;
      RECT 2042.06 189.04 2055.06 190.125 ;
      RECT 2025.08 211.445 2038.08 350.165 ;
      RECT 2025.425 189.04 2038.08 350.165 ;
      RECT 2025.08 189.04 2038.08 195.075 ;
      RECT 1994.56 259.445 2022.56 350.165 ;
      RECT 2006.935 211.445 2022.56 350.165 ;
      RECT 1994.56 189.04 1999.185 350.165 ;
      RECT 1994.56 189.04 2020.515 228.875 ;
      RECT 1994.56 189.04 2022.56 195.075 ;
      RECT 1979.04 307.445 1992.04 350.165 ;
      RECT 1989.035 194.37 1992.04 350.165 ;
      RECT 1979.04 189.04 1984.125 350.165 ;
      RECT 1979.04 228.445 1992.04 291.075 ;
      RECT 1979.04 194.37 1992.04 212.075 ;
      RECT 1979.04 189.04 1987.37 212.075 ;
      RECT 1979.04 189.04 1992.04 190.17 ;
      RECT 1962.06 307.445 1975.06 330.165 ;
      RECT 1966.705 189.04 1975.06 330.165 ;
      RECT 1966.54 228.445 1975.06 330.165 ;
      RECT 1962.06 228.445 1975.06 291.075 ;
      RECT 1962.06 189.04 1975.06 212.075 ;
      RECT 1945.08 324.445 1958.08 350.165 ;
      RECT 1945.08 189.04 1957.125 350.165 ;
      RECT 1945.08 211.445 1958.08 308.075 ;
      RECT 1945.08 189.04 1958.08 195.075 ;
      RECT 1914.56 324.445 1942.56 350.165 ;
      RECT 1940.705 189.04 1942.56 350.165 ;
      RECT 1914.56 228.445 1935.795 350.165 ;
      RECT 1938.115 189.04 1942.56 308.075 ;
      RECT 1921.11 211.445 1942.56 308.075 ;
      RECT 1914.56 189.04 1933.205 212.075 ;
      RECT 1914.56 189.04 1942.56 195.075 ;
      RECT 1899.04 290.445 1912.04 350.165 ;
      RECT 1911.425 194.42 1912.04 350.165 ;
      RECT 1899.04 189.04 1903.675 350.165 ;
      RECT 1899.04 194.42 1912.04 259.875 ;
      RECT 1899.04 189.04 1910.41 259.875 ;
      RECT 1899.04 189.04 1912.04 190.125 ;
      RECT 1882.06 211.445 1895.06 330.165 ;
      RECT 1885.425 189.04 1895.06 330.165 ;
      RECT 1882.06 189.04 1895.06 195.075 ;
      RECT 1865.08 259.445 1878.08 350.165 ;
      RECT 1866.935 189.04 1878.08 350.165 ;
      RECT 1865.08 189.04 1878.08 228.875 ;
      RECT 1834.56 307.445 1862.56 350.165 ;
      RECT 1849.035 259.445 1862.56 350.165 ;
      RECT 1834.56 189.04 1844.125 350.165 ;
      RECT 1834.56 228.445 1859.185 291.075 ;
      RECT 1853.09 189.04 1862.56 228.875 ;
      RECT 1849.035 194.37 1862.56 228.875 ;
      RECT 1834.56 194.37 1862.56 212.075 ;
      RECT 1834.56 189.04 1847.37 212.075 ;
      RECT 1834.56 189.04 1862.56 190.17 ;
      RECT 1819.04 324.445 1832.04 350.165 ;
      RECT 1826.705 189.04 1832.04 350.165 ;
      RECT 1822.035 307.445 1832.04 350.165 ;
      RECT 1819.04 307.445 1832.04 308.075 ;
      RECT 1819.04 211.445 1821.795 308.075 ;
      RECT 1819.04 228.445 1832.04 291.075 ;
      RECT 1819.04 211.445 1832.04 212.075 ;
      RECT 1822.035 189.04 1832.04 212.075 ;
      RECT 1819.04 189.04 1832.04 195.075 ;
      RECT 1785.08 324.445 1798.08 350.165 ;
      RECT 1785.08 228.445 1795.795 350.165 ;
      RECT 1790.31 211.445 1798.08 308.075 ;
      RECT 1785.08 189.04 1793.125 212.075 ;
      RECT 1785.08 189.04 1798.08 195.075 ;
      RECT 1754.56 290.445 1782.56 350.165 ;
      RECT 1773.19 189.04 1782.56 350.165 ;
      RECT 1771.425 194.425 1782.56 350.165 ;
      RECT 1754.56 189.04 1763.675 350.165 ;
      RECT 1754.56 194.425 1782.56 259.875 ;
      RECT 1754.56 189.04 1770.41 259.875 ;
      RECT 1754.56 189.04 1782.56 190.125 ;
      RECT 1739.04 211.445 1752.04 350.165 ;
      RECT 1745.425 189.04 1752.04 350.165 ;
      RECT 1739.04 189.04 1740.515 350.165 ;
      RECT 1739.04 189.04 1752.04 195.075 ;
      RECT 1722.06 259.445 1735.06 330.165 ;
      RECT 1726.935 189.04 1735.06 330.165 ;
      RECT 1722.06 189.04 1735.06 228.875 ;
      RECT 1705.08 307.445 1718.08 350.165 ;
      RECT 1713.09 189.04 1718.08 350.165 ;
      RECT 1709.035 194.37 1718.08 350.165 ;
      RECT 1705.08 228.445 1718.08 291.075 ;
      RECT 1705.08 194.37 1718.08 212.075 ;
      RECT 1705.08 189.04 1707.37 212.075 ;
      RECT 1705.08 189.04 1718.08 190.38 ;
      RECT 1674.56 324.445 1702.56 350.165 ;
      RECT 1686.705 189.04 1702.56 350.165 ;
      RECT 1682.035 307.445 1702.56 350.165 ;
      RECT 1674.56 189.04 1677.125 350.165 ;
      RECT 1674.56 307.445 1702.56 308.075 ;
      RECT 1674.56 211.445 1681.795 308.075 ;
      RECT 1674.56 228.445 1702.56 291.075 ;
      RECT 1674.56 211.445 1702.56 212.075 ;
      RECT 1682.035 189.04 1702.56 212.075 ;
      RECT 1674.56 189.04 1702.56 195.075 ;
      RECT 1659.04 324.445 1672.04 350.165 ;
      RECT 1660.705 189.04 1672.04 350.165 ;
      RECT 1659.04 189.04 1672.04 308.075 ;
      RECT 1642.06 228.445 1655.06 330.165 ;
      RECT 1648.69 211.445 1655.06 330.165 ;
      RECT 1642.06 189.04 1652.015 212.075 ;
      RECT 1642.06 189.04 1655.06 195.075 ;
      RECT 1625.08 290.445 1638.08 350.165 ;
      RECT 1633.19 189.04 1638.08 350.165 ;
      RECT 1631.425 194.425 1638.08 350.165 ;
      RECT 1625.08 194.425 1638.08 259.875 ;
      RECT 1625.08 189.04 1630.41 259.875 ;
      RECT 1625.08 189.04 1638.08 190.125 ;
      RECT 1594.56 211.445 1622.56 350.165 ;
      RECT 1605.425 189.04 1622.56 350.165 ;
      RECT 1594.56 189.04 1600.515 350.165 ;
      RECT 1594.56 189.04 1622.56 195.075 ;
      RECT 1579.04 259.445 1592.04 350.165 ;
      RECT 1586.935 189.04 1592.04 350.165 ;
      RECT 1579.04 189.04 1592.04 228.875 ;
      RECT 1562.06 307.445 1575.06 330.165 ;
      RECT 1572.99 189.04 1575.06 330.165 ;
      RECT 1569.035 194.37 1575.06 330.165 ;
      RECT 1562.06 189.04 1564.125 330.165 ;
      RECT 1562.06 228.445 1575.06 291.075 ;
      RECT 1562.06 194.37 1575.06 212.075 ;
      RECT 1562.06 189.04 1567.37 212.075 ;
      RECT 1562.06 189.04 1575.06 190.17 ;
      RECT 1545.08 307.445 1558.08 350.165 ;
      RECT 1546.705 189.04 1558.08 350.165 ;
      RECT 1545.08 228.445 1558.08 291.075 ;
      RECT 1545.08 189.04 1558.08 212.075 ;
      RECT 1514.56 324.445 1542.56 350.165 ;
      RECT 1520.705 189.04 1537.125 350.165 ;
      RECT 1514.56 211.445 1515.795 350.165 ;
      RECT 1514.56 211.445 1541.795 308.075 ;
      RECT 1514.56 228.445 1542.56 291.075 ;
      RECT 1516.925 189.04 1537.125 308.075 ;
      RECT 1514.56 189.04 1542.56 195.075 ;
      RECT 1499.04 228.445 1512.04 350.165 ;
      RECT 1499.04 189.04 1505.395 350.165 ;
      RECT 1499.04 189.04 1512.04 212.075 ;
      RECT 1482.06 290.445 1495.06 330.165 ;
      RECT 1493.19 189.04 1495.06 330.165 ;
      RECT 1491.425 194.425 1495.06 330.165 ;
      RECT 1482.06 189.04 1483.675 330.165 ;
      RECT 1482.06 194.425 1495.06 259.875 ;
      RECT 1482.06 189.04 1490.41 259.875 ;
      RECT 1482.06 189.04 1495.06 190.125 ;
      RECT 1465.08 211.445 1478.08 350.165 ;
      RECT 1465.425 189.04 1478.08 350.165 ;
      RECT 1465.08 189.04 1478.08 195.075 ;
      RECT 1434.56 259.445 1462.56 350.165 ;
      RECT 1446.935 211.445 1462.56 350.165 ;
      RECT 1434.56 189.04 1439.185 350.165 ;
      RECT 1434.56 189.04 1460.515 228.875 ;
      RECT 1434.56 189.04 1462.56 195.075 ;
      RECT 1419.04 307.445 1432.04 350.165 ;
      RECT 1429.035 194.37 1432.04 350.165 ;
      RECT 1419.04 189.04 1424.125 350.165 ;
      RECT 1419.04 228.445 1432.04 291.075 ;
      RECT 1419.04 194.37 1432.04 212.075 ;
      RECT 1419.04 189.04 1427.37 212.075 ;
      RECT 1419.04 189.04 1432.04 190.17 ;
      RECT 1402.06 307.445 1415.06 330.165 ;
      RECT 1406.705 189.04 1415.06 330.165 ;
      RECT 1406.54 228.445 1415.06 330.165 ;
      RECT 1402.06 228.445 1415.06 291.075 ;
      RECT 1402.06 189.04 1415.06 212.075 ;
      RECT 1385.08 324.445 1398.08 350.165 ;
      RECT 1385.08 189.04 1397.125 350.165 ;
      RECT 1385.08 211.445 1398.08 308.075 ;
      RECT 1385.08 189.04 1398.08 195.075 ;
      RECT 1354.56 324.445 1382.56 350.165 ;
      RECT 1380.705 189.04 1382.56 350.165 ;
      RECT 1354.56 228.445 1375.795 350.165 ;
      RECT 1378.115 189.04 1382.56 308.075 ;
      RECT 1361.11 211.445 1382.56 308.075 ;
      RECT 1354.56 189.04 1373.205 212.075 ;
      RECT 1354.56 189.04 1382.56 195.075 ;
      RECT 1339.04 290.445 1352.04 350.165 ;
      RECT 1351.425 194.42 1352.04 350.165 ;
      RECT 1339.04 189.04 1343.675 350.165 ;
      RECT 1339.04 194.42 1352.04 259.875 ;
      RECT 1339.04 189.04 1350.41 259.875 ;
      RECT 1339.04 189.04 1352.04 190.125 ;
      RECT 1322.06 211.445 1335.06 330.165 ;
      RECT 1325.425 189.04 1335.06 330.165 ;
      RECT 1322.06 189.04 1335.06 195.075 ;
      RECT 1305.08 259.445 1318.08 350.165 ;
      RECT 1306.935 189.04 1318.08 350.165 ;
      RECT 1305.08 189.04 1318.08 228.875 ;
      RECT 1274.56 307.445 1302.56 350.165 ;
      RECT 1289.035 259.445 1302.56 350.165 ;
      RECT 1274.56 189.04 1284.125 350.165 ;
      RECT 1274.56 228.445 1299.185 291.075 ;
      RECT 1293.09 189.04 1302.56 228.875 ;
      RECT 1289.035 194.37 1302.56 228.875 ;
      RECT 1274.56 194.37 1302.56 212.075 ;
      RECT 1274.56 189.04 1287.37 212.075 ;
      RECT 1274.56 189.04 1302.56 190.17 ;
      RECT 1259.04 324.445 1272.04 350.165 ;
      RECT 1266.705 189.04 1272.04 350.165 ;
      RECT 1262.035 307.445 1272.04 350.165 ;
      RECT 1259.04 307.445 1272.04 308.075 ;
      RECT 1259.04 211.445 1261.795 308.075 ;
      RECT 1259.04 228.445 1272.04 291.075 ;
      RECT 1259.04 211.445 1272.04 212.075 ;
      RECT 1262.035 189.04 1272.04 212.075 ;
      RECT 1259.04 189.04 1272.04 195.075 ;
      RECT 1225.08 324.445 1238.08 350.165 ;
      RECT 1225.08 228.445 1235.795 350.165 ;
      RECT 1230.31 211.445 1238.08 308.075 ;
      RECT 1225.08 189.04 1233.125 212.075 ;
      RECT 1225.08 189.04 1238.08 195.075 ;
      RECT 1194.56 290.445 1222.56 350.165 ;
      RECT 1213.19 189.04 1222.56 350.165 ;
      RECT 1211.425 194.425 1222.56 350.165 ;
      RECT 1194.56 189.04 1203.675 350.165 ;
      RECT 1194.56 194.425 1222.56 259.875 ;
      RECT 1194.56 189.04 1210.41 259.875 ;
      RECT 1194.56 189.04 1222.56 190.125 ;
      RECT 1179.04 211.445 1192.04 350.165 ;
      RECT 1185.425 189.04 1192.04 350.165 ;
      RECT 1179.04 189.04 1180.515 350.165 ;
      RECT 1179.04 189.04 1192.04 195.075 ;
      RECT 1162.06 259.445 1175.06 330.165 ;
      RECT 1166.935 189.04 1175.06 330.165 ;
      RECT 1162.06 189.04 1175.06 228.875 ;
      RECT 1145.08 307.445 1158.08 350.165 ;
      RECT 1153.09 189.04 1158.08 350.165 ;
      RECT 1149.035 194.37 1158.08 350.165 ;
      RECT 1145.08 228.445 1158.08 291.075 ;
      RECT 1145.08 194.37 1158.08 212.075 ;
      RECT 1145.08 189.04 1147.37 212.075 ;
      RECT 1145.08 189.04 1158.08 190.38 ;
      RECT 1114.56 324.445 1142.56 350.165 ;
      RECT 1126.705 189.04 1142.56 350.165 ;
      RECT 1122.035 307.445 1142.56 350.165 ;
      RECT 1114.56 189.04 1117.125 350.165 ;
      RECT 1114.56 307.445 1142.56 308.075 ;
      RECT 1114.56 211.445 1121.795 308.075 ;
      RECT 1114.56 228.445 1142.56 291.075 ;
      RECT 1114.56 211.445 1142.56 212.075 ;
      RECT 1122.035 189.04 1142.56 212.075 ;
      RECT 1114.56 189.04 1142.56 195.075 ;
      RECT 1099.04 324.445 1112.04 350.165 ;
      RECT 1100.705 189.04 1112.04 350.165 ;
      RECT 1099.04 189.04 1112.04 308.075 ;
      RECT 1082.06 228.445 1095.06 330.165 ;
      RECT 1088.69 211.445 1095.06 330.165 ;
      RECT 1082.06 189.04 1092.015 212.075 ;
      RECT 1082.06 189.04 1095.06 195.075 ;
      RECT 1065.08 290.445 1078.08 350.165 ;
      RECT 1073.19 189.04 1078.08 350.165 ;
      RECT 1071.425 194.425 1078.08 350.165 ;
      RECT 1065.08 194.425 1078.08 259.875 ;
      RECT 1065.08 189.04 1070.41 259.875 ;
      RECT 1065.08 189.04 1078.08 190.125 ;
      RECT 1034.56 211.445 1062.56 350.165 ;
      RECT 1045.425 189.04 1062.56 350.165 ;
      RECT 1034.56 189.04 1040.515 350.165 ;
      RECT 1034.56 189.04 1062.56 195.075 ;
      RECT 1019.04 259.445 1032.04 350.165 ;
      RECT 1026.935 189.04 1032.04 350.165 ;
      RECT 1019.04 189.04 1032.04 228.875 ;
      RECT 1002.06 307.445 1015.06 330.165 ;
      RECT 1012.99 189.04 1015.06 330.165 ;
      RECT 1009.035 194.37 1015.06 330.165 ;
      RECT 1002.06 189.04 1004.125 330.165 ;
      RECT 1002.06 228.445 1015.06 291.075 ;
      RECT 1002.06 194.37 1015.06 212.075 ;
      RECT 1002.06 189.04 1007.37 212.075 ;
      RECT 1002.06 189.04 1015.06 190.17 ;
      RECT 985.08 307.445 998.08 350.165 ;
      RECT 986.705 189.04 998.08 350.165 ;
      RECT 985.08 228.445 998.08 291.075 ;
      RECT 985.08 189.04 998.08 212.075 ;
      RECT 954.56 324.445 982.56 350.165 ;
      RECT 960.705 189.04 977.125 350.165 ;
      RECT 954.56 211.445 955.795 350.165 ;
      RECT 954.56 211.445 981.795 308.075 ;
      RECT 954.56 228.445 982.56 291.075 ;
      RECT 956.925 189.04 977.125 308.075 ;
      RECT 954.56 189.04 982.56 195.075 ;
      RECT 939.04 228.445 952.04 350.165 ;
      RECT 939.04 189.04 945.395 350.165 ;
      RECT 939.04 189.04 952.04 212.075 ;
      RECT 922.06 290.445 935.06 330.165 ;
      RECT 933.19 189.04 935.06 330.165 ;
      RECT 931.425 194.425 935.06 330.165 ;
      RECT 922.06 189.04 923.675 330.165 ;
      RECT 922.06 194.425 935.06 259.875 ;
      RECT 922.06 189.04 930.41 259.875 ;
      RECT 922.06 189.04 935.06 190.125 ;
      RECT 905.08 211.445 918.08 350.165 ;
      RECT 905.425 189.04 918.08 350.165 ;
      RECT 905.08 189.04 918.08 195.075 ;
      RECT 874.56 259.445 902.56 350.165 ;
      RECT 886.935 211.445 902.56 350.165 ;
      RECT 874.56 189.04 879.185 350.165 ;
      RECT 874.56 189.04 900.515 228.875 ;
      RECT 874.56 189.04 902.56 195.075 ;
      RECT 859.04 307.445 872.04 350.165 ;
      RECT 869.035 194.37 872.04 350.165 ;
      RECT 859.04 189.04 864.125 350.165 ;
      RECT 859.04 228.445 872.04 291.075 ;
      RECT 859.04 194.37 872.04 212.075 ;
      RECT 859.04 189.04 867.37 212.075 ;
      RECT 859.04 189.04 872.04 190.17 ;
      RECT 842.06 307.445 855.06 330.165 ;
      RECT 846.705 189.04 855.06 330.165 ;
      RECT 846.54 228.445 855.06 330.165 ;
      RECT 842.06 228.445 855.06 291.075 ;
      RECT 842.06 189.04 855.06 212.075 ;
      RECT 825.08 324.445 838.08 350.165 ;
      RECT 825.08 189.04 837.125 350.165 ;
      RECT 825.08 211.445 838.08 308.075 ;
      RECT 825.08 189.04 838.08 195.075 ;
      RECT 794.56 324.445 822.56 350.165 ;
      RECT 820.705 189.04 822.56 350.165 ;
      RECT 794.56 228.445 815.795 350.165 ;
      RECT 818.115 189.04 822.56 308.075 ;
      RECT 801.11 211.445 822.56 308.075 ;
      RECT 794.56 189.04 813.205 212.075 ;
      RECT 794.56 189.04 822.56 195.075 ;
      RECT 779.04 290.445 792.04 350.165 ;
      RECT 791.425 194.42 792.04 350.165 ;
      RECT 779.04 189.04 783.675 350.165 ;
      RECT 779.04 194.42 792.04 259.875 ;
      RECT 779.04 189.04 790.41 259.875 ;
      RECT 779.04 189.04 792.04 190.125 ;
      RECT 762.06 211.445 775.06 330.165 ;
      RECT 765.425 189.04 775.06 330.165 ;
      RECT 762.06 189.04 775.06 195.075 ;
      RECT 745.08 259.445 758.08 350.165 ;
      RECT 746.935 189.04 758.08 350.165 ;
      RECT 745.08 189.04 758.08 228.875 ;
      RECT 714.56 307.445 742.56 350.165 ;
      RECT 729.035 259.445 742.56 350.165 ;
      RECT 714.56 189.04 724.125 350.165 ;
      RECT 714.56 228.445 739.185 291.075 ;
      RECT 733.09 189.04 742.56 228.875 ;
      RECT 729.035 194.37 742.56 228.875 ;
      RECT 714.56 194.37 742.56 212.075 ;
      RECT 714.56 189.04 727.37 212.075 ;
      RECT 714.56 189.04 742.56 190.17 ;
      RECT 699.04 324.445 712.04 350.165 ;
      RECT 706.705 189.04 712.04 350.165 ;
      RECT 702.035 307.445 712.04 350.165 ;
      RECT 699.04 307.445 712.04 308.075 ;
      RECT 699.04 211.445 701.795 308.075 ;
      RECT 699.04 228.445 712.04 291.075 ;
      RECT 699.04 211.445 712.04 212.075 ;
      RECT 702.035 189.04 712.04 212.075 ;
      RECT 699.04 189.04 712.04 195.075 ;
      RECT 665.08 324.445 678.08 350.165 ;
      RECT 665.08 228.445 675.795 350.165 ;
      RECT 670.31 211.445 678.08 308.075 ;
      RECT 665.08 189.04 673.125 212.075 ;
      RECT 665.08 189.04 678.08 195.075 ;
      RECT 634.56 290.445 662.56 350.165 ;
      RECT 653.19 189.04 662.56 350.165 ;
      RECT 651.425 194.425 662.56 350.165 ;
      RECT 634.56 189.04 643.675 350.165 ;
      RECT 634.56 194.425 662.56 259.875 ;
      RECT 634.56 189.04 650.41 259.875 ;
      RECT 634.56 189.04 662.56 190.125 ;
      RECT 619.04 211.445 632.04 350.165 ;
      RECT 625.425 189.04 632.04 350.165 ;
      RECT 619.04 189.04 620.515 350.165 ;
      RECT 619.04 189.04 632.04 195.075 ;
      RECT 602.06 259.445 615.06 330.165 ;
      RECT 606.935 189.04 615.06 330.165 ;
      RECT 602.06 189.04 615.06 228.875 ;
      RECT 585.08 307.445 598.08 350.165 ;
      RECT 593.09 189.04 598.08 350.165 ;
      RECT 589.035 194.37 598.08 350.165 ;
      RECT 585.08 228.445 598.08 291.075 ;
      RECT 585.08 194.37 598.08 212.075 ;
      RECT 585.08 189.04 587.37 212.075 ;
      RECT 585.08 189.04 598.08 190.38 ;
      RECT 554.56 324.445 582.56 350.165 ;
      RECT 566.705 189.04 582.56 350.165 ;
      RECT 562.035 307.445 582.56 350.165 ;
      RECT 554.56 189.04 557.125 350.165 ;
      RECT 554.56 307.445 582.56 308.075 ;
      RECT 554.56 211.445 561.795 308.075 ;
      RECT 554.56 228.445 582.56 291.075 ;
      RECT 554.56 211.445 582.56 212.075 ;
      RECT 562.035 189.04 582.56 212.075 ;
      RECT 554.56 189.04 582.56 195.075 ;
      RECT 539.04 324.445 552.04 350.165 ;
      RECT 540.705 189.04 552.04 350.165 ;
      RECT 539.04 189.04 552.04 308.075 ;
      RECT 522.06 228.445 535.06 330.165 ;
      RECT 528.69 211.445 535.06 330.165 ;
      RECT 522.06 189.04 532.015 212.075 ;
      RECT 522.06 189.04 535.06 195.075 ;
      RECT 505.08 290.445 518.08 350.165 ;
      RECT 513.19 189.04 518.08 350.165 ;
      RECT 511.425 194.425 518.08 350.165 ;
      RECT 505.08 194.425 518.08 259.875 ;
      RECT 505.08 189.04 510.41 259.875 ;
      RECT 505.08 189.04 518.08 190.125 ;
      RECT 474.56 211.445 502.56 350.165 ;
      RECT 485.425 189.04 502.56 350.165 ;
      RECT 474.56 189.04 480.515 350.165 ;
      RECT 474.56 189.04 502.56 195.075 ;
      RECT 459.04 259.445 472.04 350.165 ;
      RECT 466.935 189.04 472.04 350.165 ;
      RECT 459.04 189.04 472.04 228.875 ;
      RECT 18440.77 258.23 18490.46 258.79 ;
      RECT 18438.37 259.99 18488.86 261.19 ;
      RECT 18435.97 262.39 18488.86 263.59 ;
      RECT 18433.57 264.79 18488.86 265.99 ;
      RECT 18431.17 267.19 18488.86 268.39 ;
      RECT 18455.125 511.37 18460.125 8613.565 ;
      RECT 18042.06 189.04 18055.06 330.165 ;
      RECT 17482.06 189.04 17495.06 330.165 ;
      RECT 16922.06 189.04 16935.06 330.165 ;
      RECT 16362.06 189.04 16375.06 330.165 ;
      RECT 15802.06 189.04 15815.06 330.165 ;
      RECT 15242.06 189.04 15255.06 330.165 ;
      RECT 14682.06 189.04 14695.06 330.165 ;
      RECT 14122.06 189.04 14135.06 330.165 ;
      RECT 13562.06 189.04 13575.06 330.165 ;
      RECT 13002.06 189.04 13015.06 330.165 ;
      RECT 12442.06 189.04 12455.06 330.165 ;
      RECT 11882.06 189.04 11895.06 330.165 ;
      RECT 11322.06 189.04 11335.06 330.165 ;
      RECT 10762.06 189.04 10775.06 330.165 ;
      RECT 10202.06 189.04 10215.06 330.165 ;
      RECT 9642.06 189.04 9655.06 330.165 ;
      RECT 9082.06 189.04 9095.06 330.165 ;
      RECT 8522.06 189.04 8535.06 330.165 ;
      RECT 7962.06 189.04 7975.06 330.165 ;
      RECT 7402.06 189.04 7415.06 330.165 ;
      RECT 6842.06 189.04 6855.06 330.165 ;
      RECT 6282.06 189.04 6295.06 330.165 ;
      RECT 5722.06 189.04 5735.06 330.165 ;
      RECT 5162.06 189.04 5175.06 330.165 ;
      RECT 4602.06 189.04 4615.06 330.165 ;
      RECT 4042.06 189.04 4055.06 330.165 ;
      RECT 3482.06 189.04 3495.06 330.165 ;
      RECT 2922.06 189.04 2935.06 330.165 ;
      RECT 2362.06 189.04 2375.06 330.165 ;
      RECT 1802.06 189.04 1815.06 330.165 ;
      RECT 1242.06 189.04 1255.06 330.165 ;
      RECT 682.06 189.04 695.06 330.165 ;
      RECT 326.66 255.83 453.68 256.39 ;
      RECT 328.26 257.59 449.785 258.79 ;
      RECT 328.26 259.99 449.785 261.19 ;
      RECT 328.26 267.19 449.785 268.39 ;
      RECT 328.26 262.39 438.95 263.59 ;
      RECT 328.26 264.79 438.95 265.99 ;
      RECT 356.995 511.82 361.995 8613.565 ;
    LAYER M5 SPACING 0.28 ;
      RECT 326.66 8583.935 18490.46 8613.565 ;
      RECT 328.08 268.86 18489.04 8613.565 ;
      RECT 326.66 8545.42 18490.46 8581.675 ;
      RECT 326.66 8511.935 18490.46 8543.16 ;
      RECT 326.66 8473.42 18490.46 8509.675 ;
      RECT 326.66 8439.935 18490.46 8471.16 ;
      RECT 326.66 8401.42 18490.46 8437.675 ;
      RECT 326.66 268.86 18490.46 8399.16 ;
      RECT 328.13 188.91 18488.99 8613.565 ;
      RECT 18375.53 187.44 18490.46 259.52 ;
      RECT 326.66 187.44 458.57 257.12 ;
      RECT 18358.55 188.86 18361.59 8613.565 ;
      RECT 18343.03 187.44 18344.61 8613.565 ;
      RECT 18312.51 187.44 18314.09 8613.565 ;
      RECT 18295.53 187.44 18298.57 8613.565 ;
      RECT 18278.55 188.86 18281.59 8613.565 ;
      RECT 18263.03 187.44 18264.61 8613.565 ;
      RECT 18232.51 187.44 18234.09 8613.565 ;
      RECT 18215.53 188.86 18218.57 8613.565 ;
      RECT 18198.55 187.44 18201.59 8613.565 ;
      RECT 18183.03 188.86 18184.61 8613.565 ;
      RECT 18152.51 187.44 18154.09 8613.565 ;
      RECT 18135.53 188.86 18138.57 8613.565 ;
      RECT 18118.55 188.86 18121.59 8613.565 ;
      RECT 18120.965 187.44 18121.59 8613.565 ;
      RECT 18103.03 187.44 18104.61 8613.565 ;
      RECT 18072.51 188.86 18074.09 8613.565 ;
      RECT 18055.53 187.44 18058.57 8613.565 ;
      RECT 18038.55 187.44 18041.59 8613.565 ;
      RECT 18023.03 187.44 18024.61 8613.565 ;
      RECT 17992.51 188.86 17994.09 8613.565 ;
      RECT 17975.53 188.86 17978.57 8613.565 ;
      RECT 17958.55 187.44 17961.59 8613.565 ;
      RECT 17943.03 187.44 17944.61 8613.565 ;
      RECT 17912.51 188.86 17914.09 8613.565 ;
      RECT 17895.53 187.44 17898.57 8613.565 ;
      RECT 17878.55 187.44 17881.59 8613.565 ;
      RECT 17863.03 187.44 17864.61 8613.565 ;
      RECT 17832.51 188.86 17834.09 8613.565 ;
      RECT 17815.53 187.44 17818.57 8613.565 ;
      RECT 17798.55 188.86 17801.59 8613.565 ;
      RECT 17801.205 187.44 17801.59 8613.565 ;
      RECT 17783.03 187.44 17784.61 8613.565 ;
      RECT 17752.51 187.44 17754.09 8613.565 ;
      RECT 17735.53 187.44 17738.57 8613.565 ;
      RECT 17718.55 188.86 17721.59 8613.565 ;
      RECT 17703.03 187.44 17704.61 8613.565 ;
      RECT 17672.51 187.44 17674.09 8613.565 ;
      RECT 17655.53 188.86 17658.57 8613.565 ;
      RECT 17638.55 187.44 17641.59 8613.565 ;
      RECT 17623.03 188.86 17624.61 8613.565 ;
      RECT 17592.51 187.44 17594.09 8613.565 ;
      RECT 17575.53 188.86 17578.57 8613.565 ;
      RECT 17558.55 188.86 17561.59 8613.565 ;
      RECT 17560.965 187.44 17561.59 8613.565 ;
      RECT 17543.03 187.44 17544.61 8613.565 ;
      RECT 17512.51 188.86 17514.09 8613.565 ;
      RECT 17495.53 187.44 17498.57 8613.565 ;
      RECT 17478.55 187.44 17481.59 8613.565 ;
      RECT 17463.03 187.44 17464.61 8613.565 ;
      RECT 17432.51 188.86 17434.09 8613.565 ;
      RECT 17415.53 188.86 17418.57 8613.565 ;
      RECT 17398.55 187.44 17401.59 8613.565 ;
      RECT 17383.03 187.44 17384.61 8613.565 ;
      RECT 17352.51 188.86 17354.09 8613.565 ;
      RECT 17335.53 187.44 17338.57 8613.565 ;
      RECT 17318.55 187.44 17321.59 8613.565 ;
      RECT 17303.03 187.44 17304.61 8613.565 ;
      RECT 17272.51 188.86 17274.09 8613.565 ;
      RECT 17255.53 187.44 17258.57 8613.565 ;
      RECT 17238.55 188.86 17241.59 8613.565 ;
      RECT 17241.205 187.44 17241.59 8613.565 ;
      RECT 17223.03 187.44 17224.61 8613.565 ;
      RECT 17192.51 187.44 17194.09 8613.565 ;
      RECT 17175.53 187.44 17178.57 8613.565 ;
      RECT 17158.55 188.86 17161.59 8613.565 ;
      RECT 17143.03 187.44 17144.61 8613.565 ;
      RECT 17112.51 187.44 17114.09 8613.565 ;
      RECT 17095.53 188.86 17098.57 8613.565 ;
      RECT 17078.55 187.44 17081.59 8613.565 ;
      RECT 17063.03 188.86 17064.61 8613.565 ;
      RECT 17032.51 187.44 17034.09 8613.565 ;
      RECT 17015.53 188.86 17018.57 8613.565 ;
      RECT 16998.55 188.86 17001.59 8613.565 ;
      RECT 17000.965 187.44 17001.59 8613.565 ;
      RECT 16983.03 187.44 16984.61 8613.565 ;
      RECT 16952.51 188.86 16954.09 8613.565 ;
      RECT 16935.53 187.44 16938.57 8613.565 ;
      RECT 16918.55 187.44 16921.59 8613.565 ;
      RECT 16903.03 187.44 16904.61 8613.565 ;
      RECT 16872.51 188.86 16874.09 8613.565 ;
      RECT 16855.53 188.86 16858.57 8613.565 ;
      RECT 16838.55 187.44 16841.59 8613.565 ;
      RECT 16823.03 187.44 16824.61 8613.565 ;
      RECT 16792.51 188.86 16794.09 8613.565 ;
      RECT 16775.53 187.44 16778.57 8613.565 ;
      RECT 16758.55 187.44 16761.59 8613.565 ;
      RECT 16743.03 187.44 16744.61 8613.565 ;
      RECT 16712.51 188.86 16714.09 8613.565 ;
      RECT 16695.53 187.44 16698.57 8613.565 ;
      RECT 16678.55 188.86 16681.59 8613.565 ;
      RECT 16681.205 187.44 16681.59 8613.565 ;
      RECT 16663.03 187.44 16664.61 8613.565 ;
      RECT 16632.51 187.44 16634.09 8613.565 ;
      RECT 16615.53 187.44 16618.57 8613.565 ;
      RECT 16598.55 188.86 16601.59 8613.565 ;
      RECT 16583.03 187.44 16584.61 8613.565 ;
      RECT 16552.51 187.44 16554.09 8613.565 ;
      RECT 16535.53 188.86 16538.57 8613.565 ;
      RECT 16518.55 187.44 16521.59 8613.565 ;
      RECT 16503.03 188.86 16504.61 8613.565 ;
      RECT 16472.51 187.44 16474.09 8613.565 ;
      RECT 16455.53 188.86 16458.57 8613.565 ;
      RECT 16438.55 188.86 16441.59 8613.565 ;
      RECT 16440.965 187.44 16441.59 8613.565 ;
      RECT 16423.03 187.44 16424.61 8613.565 ;
      RECT 16392.51 188.86 16394.09 8613.565 ;
      RECT 16375.53 187.44 16378.57 8613.565 ;
      RECT 16358.55 187.44 16361.59 8613.565 ;
      RECT 16343.03 187.44 16344.61 8613.565 ;
      RECT 16312.51 188.86 16314.09 8613.565 ;
      RECT 16295.53 188.86 16298.57 8613.565 ;
      RECT 16278.55 187.44 16281.59 8613.565 ;
      RECT 16263.03 187.44 16264.61 8613.565 ;
      RECT 16232.51 188.86 16234.09 8613.565 ;
      RECT 16215.53 187.44 16218.57 8613.565 ;
      RECT 16198.55 187.44 16201.59 8613.565 ;
      RECT 16183.03 187.44 16184.61 8613.565 ;
      RECT 16152.51 188.86 16154.09 8613.565 ;
      RECT 16135.53 187.44 16138.57 8613.565 ;
      RECT 16118.55 188.86 16121.59 8613.565 ;
      RECT 16121.205 187.44 16121.59 8613.565 ;
      RECT 16103.03 187.44 16104.61 8613.565 ;
      RECT 16072.51 187.44 16074.09 8613.565 ;
      RECT 16055.53 187.44 16058.57 8613.565 ;
      RECT 16038.55 188.86 16041.59 8613.565 ;
      RECT 16023.03 187.44 16024.61 8613.565 ;
      RECT 15992.51 187.44 15994.09 8613.565 ;
      RECT 15975.53 188.86 15978.57 8613.565 ;
      RECT 15958.55 187.44 15961.59 8613.565 ;
      RECT 15943.03 188.86 15944.61 8613.565 ;
      RECT 15912.51 187.44 15914.09 8613.565 ;
      RECT 15895.53 188.86 15898.57 8613.565 ;
      RECT 15878.55 188.86 15881.59 8613.565 ;
      RECT 15880.965 187.44 15881.59 8613.565 ;
      RECT 15863.03 187.44 15864.61 8613.565 ;
      RECT 15832.51 188.86 15834.09 8613.565 ;
      RECT 15815.53 187.44 15818.57 8613.565 ;
      RECT 15798.55 187.44 15801.59 8613.565 ;
      RECT 15783.03 187.44 15784.61 8613.565 ;
      RECT 15752.51 188.86 15754.09 8613.565 ;
      RECT 15735.53 188.86 15738.57 8613.565 ;
      RECT 15718.55 187.44 15721.59 8613.565 ;
      RECT 15703.03 187.44 15704.61 8613.565 ;
      RECT 15672.51 188.86 15674.09 8613.565 ;
      RECT 15655.53 187.44 15658.57 8613.565 ;
      RECT 15638.55 187.44 15641.59 8613.565 ;
      RECT 15623.03 187.44 15624.61 8613.565 ;
      RECT 15592.51 188.86 15594.09 8613.565 ;
      RECT 15575.53 187.44 15578.57 8613.565 ;
      RECT 15558.55 188.86 15561.59 8613.565 ;
      RECT 15561.205 187.44 15561.59 8613.565 ;
      RECT 15543.03 187.44 15544.61 8613.565 ;
      RECT 15512.51 187.44 15514.09 8613.565 ;
      RECT 15495.53 187.44 15498.57 8613.565 ;
      RECT 15478.55 188.86 15481.59 8613.565 ;
      RECT 15463.03 187.44 15464.61 8613.565 ;
      RECT 15432.51 187.44 15434.09 8613.565 ;
      RECT 15415.53 188.86 15418.57 8613.565 ;
      RECT 15398.55 187.44 15401.59 8613.565 ;
      RECT 15383.03 188.86 15384.61 8613.565 ;
      RECT 15352.51 187.44 15354.09 8613.565 ;
      RECT 15335.53 188.86 15338.57 8613.565 ;
      RECT 15318.55 188.86 15321.59 8613.565 ;
      RECT 15320.965 187.44 15321.59 8613.565 ;
      RECT 15303.03 187.44 15304.61 8613.565 ;
      RECT 15272.51 188.86 15274.09 8613.565 ;
      RECT 15255.53 187.44 15258.57 8613.565 ;
      RECT 15238.55 187.44 15241.59 8613.565 ;
      RECT 15223.03 187.44 15224.61 8613.565 ;
      RECT 15192.51 188.86 15194.09 8613.565 ;
      RECT 15175.53 188.86 15178.57 8613.565 ;
      RECT 15158.55 187.44 15161.59 8613.565 ;
      RECT 15143.03 187.44 15144.61 8613.565 ;
      RECT 15112.51 188.86 15114.09 8613.565 ;
      RECT 15095.53 187.44 15098.57 8613.565 ;
      RECT 15078.55 187.44 15081.59 8613.565 ;
      RECT 15063.03 187.44 15064.61 8613.565 ;
      RECT 15032.51 188.86 15034.09 8613.565 ;
      RECT 15015.53 187.44 15018.57 8613.565 ;
      RECT 14998.55 188.86 15001.59 8613.565 ;
      RECT 15001.205 187.44 15001.59 8613.565 ;
      RECT 14983.03 187.44 14984.61 8613.565 ;
      RECT 14952.51 187.44 14954.09 8613.565 ;
      RECT 14935.53 187.44 14938.57 8613.565 ;
      RECT 14918.55 188.86 14921.59 8613.565 ;
      RECT 14903.03 187.44 14904.61 8613.565 ;
      RECT 14872.51 187.44 14874.09 8613.565 ;
      RECT 14855.53 188.86 14858.57 8613.565 ;
      RECT 14838.55 187.44 14841.59 8613.565 ;
      RECT 14823.03 188.86 14824.61 8613.565 ;
      RECT 14792.51 187.44 14794.09 8613.565 ;
      RECT 14775.53 188.86 14778.57 8613.565 ;
      RECT 14758.55 188.86 14761.59 8613.565 ;
      RECT 14760.965 187.44 14761.59 8613.565 ;
      RECT 14743.03 187.44 14744.61 8613.565 ;
      RECT 14712.51 188.86 14714.09 8613.565 ;
      RECT 14695.53 187.44 14698.57 8613.565 ;
      RECT 14678.55 187.44 14681.59 8613.565 ;
      RECT 14663.03 187.44 14664.61 8613.565 ;
      RECT 14632.51 188.86 14634.09 8613.565 ;
      RECT 14615.53 188.86 14618.57 8613.565 ;
      RECT 14598.55 187.44 14601.59 8613.565 ;
      RECT 14583.03 187.44 14584.61 8613.565 ;
      RECT 14552.51 188.86 14554.09 8613.565 ;
      RECT 14535.53 187.44 14538.57 8613.565 ;
      RECT 14518.55 187.44 14521.59 8613.565 ;
      RECT 14503.03 187.44 14504.61 8613.565 ;
      RECT 14472.51 188.86 14474.09 8613.565 ;
      RECT 14455.53 187.44 14458.57 8613.565 ;
      RECT 14438.55 188.86 14441.59 8613.565 ;
      RECT 14441.205 187.44 14441.59 8613.565 ;
      RECT 14423.03 187.44 14424.61 8613.565 ;
      RECT 14392.51 187.44 14394.09 8613.565 ;
      RECT 14375.53 187.44 14378.57 8613.565 ;
      RECT 14358.55 188.86 14361.59 8613.565 ;
      RECT 14343.03 187.44 14344.61 8613.565 ;
      RECT 14312.51 187.44 14314.09 8613.565 ;
      RECT 14295.53 188.86 14298.57 8613.565 ;
      RECT 14278.55 187.44 14281.59 8613.565 ;
      RECT 14263.03 188.86 14264.61 8613.565 ;
      RECT 14232.51 187.44 14234.09 8613.565 ;
      RECT 14215.53 188.86 14218.57 8613.565 ;
      RECT 14198.55 188.86 14201.59 8613.565 ;
      RECT 14200.965 187.44 14201.59 8613.565 ;
      RECT 14183.03 187.44 14184.61 8613.565 ;
      RECT 14152.51 188.86 14154.09 8613.565 ;
      RECT 14135.53 187.44 14138.57 8613.565 ;
      RECT 14118.55 187.44 14121.59 8613.565 ;
      RECT 14103.03 187.44 14104.61 8613.565 ;
      RECT 14072.51 188.86 14074.09 8613.565 ;
      RECT 14055.53 188.86 14058.57 8613.565 ;
      RECT 14038.55 187.44 14041.59 8613.565 ;
      RECT 14023.03 187.44 14024.61 8613.565 ;
      RECT 13992.51 188.86 13994.09 8613.565 ;
      RECT 13975.53 187.44 13978.57 8613.565 ;
      RECT 13958.55 187.44 13961.59 8613.565 ;
      RECT 13943.03 187.44 13944.61 8613.565 ;
      RECT 13912.51 188.86 13914.09 8613.565 ;
      RECT 13895.53 187.44 13898.57 8613.565 ;
      RECT 13878.55 188.86 13881.59 8613.565 ;
      RECT 13881.205 187.44 13881.59 8613.565 ;
      RECT 13863.03 187.44 13864.61 8613.565 ;
      RECT 13832.51 187.44 13834.09 8613.565 ;
      RECT 13815.53 187.44 13818.57 8613.565 ;
      RECT 13798.55 188.86 13801.59 8613.565 ;
      RECT 13783.03 187.44 13784.61 8613.565 ;
      RECT 13752.51 187.44 13754.09 8613.565 ;
      RECT 13735.53 188.86 13738.57 8613.565 ;
      RECT 13718.55 187.44 13721.59 8613.565 ;
      RECT 13703.03 188.86 13704.61 8613.565 ;
      RECT 13672.51 187.44 13674.09 8613.565 ;
      RECT 13655.53 188.86 13658.57 8613.565 ;
      RECT 13638.55 188.86 13641.59 8613.565 ;
      RECT 13640.965 187.44 13641.59 8613.565 ;
      RECT 13623.03 187.44 13624.61 8613.565 ;
      RECT 13592.51 188.86 13594.09 8613.565 ;
      RECT 13575.53 187.44 13578.57 8613.565 ;
      RECT 13558.55 187.44 13561.59 8613.565 ;
      RECT 13543.03 187.44 13544.61 8613.565 ;
      RECT 13512.51 188.86 13514.09 8613.565 ;
      RECT 13495.53 188.86 13498.57 8613.565 ;
      RECT 13478.55 187.44 13481.59 8613.565 ;
      RECT 13463.03 187.44 13464.61 8613.565 ;
      RECT 13432.51 188.86 13434.09 8613.565 ;
      RECT 13415.53 187.44 13418.57 8613.565 ;
      RECT 13398.55 187.44 13401.59 8613.565 ;
      RECT 13383.03 187.44 13384.61 8613.565 ;
      RECT 13352.51 188.86 13354.09 8613.565 ;
      RECT 13335.53 187.44 13338.57 8613.565 ;
      RECT 13318.55 188.86 13321.59 8613.565 ;
      RECT 13321.205 187.44 13321.59 8613.565 ;
      RECT 13303.03 187.44 13304.61 8613.565 ;
      RECT 13272.51 187.44 13274.09 8613.565 ;
      RECT 13255.53 187.44 13258.57 8613.565 ;
      RECT 13238.55 188.86 13241.59 8613.565 ;
      RECT 13223.03 187.44 13224.61 8613.565 ;
      RECT 13192.51 187.44 13194.09 8613.565 ;
      RECT 13175.53 188.86 13178.57 8613.565 ;
      RECT 13158.55 187.44 13161.59 8613.565 ;
      RECT 13143.03 188.86 13144.61 8613.565 ;
      RECT 13112.51 187.44 13114.09 8613.565 ;
      RECT 13095.53 188.86 13098.57 8613.565 ;
      RECT 13078.55 188.86 13081.59 8613.565 ;
      RECT 13080.965 187.44 13081.59 8613.565 ;
      RECT 13063.03 187.44 13064.61 8613.565 ;
      RECT 13032.51 188.86 13034.09 8613.565 ;
      RECT 13015.53 187.44 13018.57 8613.565 ;
      RECT 12998.55 187.44 13001.59 8613.565 ;
      RECT 12983.03 187.44 12984.61 8613.565 ;
      RECT 12952.51 188.86 12954.09 8613.565 ;
      RECT 12935.53 188.86 12938.57 8613.565 ;
      RECT 12918.55 187.44 12921.59 8613.565 ;
      RECT 12903.03 187.44 12904.61 8613.565 ;
      RECT 12872.51 188.86 12874.09 8613.565 ;
      RECT 12855.53 187.44 12858.57 8613.565 ;
      RECT 12838.55 187.44 12841.59 8613.565 ;
      RECT 12823.03 187.44 12824.61 8613.565 ;
      RECT 12792.51 188.86 12794.09 8613.565 ;
      RECT 12775.53 187.44 12778.57 8613.565 ;
      RECT 12758.55 188.86 12761.59 8613.565 ;
      RECT 12761.205 187.44 12761.59 8613.565 ;
      RECT 12743.03 187.44 12744.61 8613.565 ;
      RECT 12712.51 187.44 12714.09 8613.565 ;
      RECT 12695.53 187.44 12698.57 8613.565 ;
      RECT 12678.55 188.86 12681.59 8613.565 ;
      RECT 12663.03 187.44 12664.61 8613.565 ;
      RECT 12632.51 187.44 12634.09 8613.565 ;
      RECT 12615.53 188.86 12618.57 8613.565 ;
      RECT 12598.55 187.44 12601.59 8613.565 ;
      RECT 12583.03 188.86 12584.61 8613.565 ;
      RECT 12552.51 187.44 12554.09 8613.565 ;
      RECT 12535.53 188.86 12538.57 8613.565 ;
      RECT 12518.55 188.86 12521.59 8613.565 ;
      RECT 12520.965 187.44 12521.59 8613.565 ;
      RECT 12503.03 187.44 12504.61 8613.565 ;
      RECT 12472.51 188.86 12474.09 8613.565 ;
      RECT 12455.53 187.44 12458.57 8613.565 ;
      RECT 12438.55 187.44 12441.59 8613.565 ;
      RECT 12423.03 187.44 12424.61 8613.565 ;
      RECT 12392.51 188.86 12394.09 8613.565 ;
      RECT 12375.53 188.86 12378.57 8613.565 ;
      RECT 12358.55 187.44 12361.59 8613.565 ;
      RECT 12343.03 187.44 12344.61 8613.565 ;
      RECT 12312.51 188.86 12314.09 8613.565 ;
      RECT 12295.53 187.44 12298.57 8613.565 ;
      RECT 12278.55 187.44 12281.59 8613.565 ;
      RECT 12263.03 187.44 12264.61 8613.565 ;
      RECT 12232.51 188.86 12234.09 8613.565 ;
      RECT 12215.53 187.44 12218.57 8613.565 ;
      RECT 12198.55 188.86 12201.59 8613.565 ;
      RECT 12201.205 187.44 12201.59 8613.565 ;
      RECT 12183.03 187.44 12184.61 8613.565 ;
      RECT 12152.51 187.44 12154.09 8613.565 ;
      RECT 12135.53 187.44 12138.57 8613.565 ;
      RECT 12118.55 188.86 12121.59 8613.565 ;
      RECT 12103.03 187.44 12104.61 8613.565 ;
      RECT 12072.51 187.44 12074.09 8613.565 ;
      RECT 12055.53 188.86 12058.57 8613.565 ;
      RECT 12038.55 187.44 12041.59 8613.565 ;
      RECT 12023.03 188.86 12024.61 8613.565 ;
      RECT 11992.51 187.44 11994.09 8613.565 ;
      RECT 11975.53 188.86 11978.57 8613.565 ;
      RECT 11958.55 188.86 11961.59 8613.565 ;
      RECT 11960.965 187.44 11961.59 8613.565 ;
      RECT 11943.03 187.44 11944.61 8613.565 ;
      RECT 11912.51 188.86 11914.09 8613.565 ;
      RECT 11895.53 187.44 11898.57 8613.565 ;
      RECT 11878.55 187.44 11881.59 8613.565 ;
      RECT 11863.03 187.44 11864.61 8613.565 ;
      RECT 11832.51 188.86 11834.09 8613.565 ;
      RECT 11815.53 188.86 11818.57 8613.565 ;
      RECT 11798.55 187.44 11801.59 8613.565 ;
      RECT 11783.03 187.44 11784.61 8613.565 ;
      RECT 11752.51 188.86 11754.09 8613.565 ;
      RECT 11735.53 187.44 11738.57 8613.565 ;
      RECT 11718.55 187.44 11721.59 8613.565 ;
      RECT 11703.03 187.44 11704.61 8613.565 ;
      RECT 11672.51 188.86 11674.09 8613.565 ;
      RECT 11655.53 187.44 11658.57 8613.565 ;
      RECT 11638.55 188.86 11641.59 8613.565 ;
      RECT 11641.205 187.44 11641.59 8613.565 ;
      RECT 11623.03 187.44 11624.61 8613.565 ;
      RECT 11592.51 187.44 11594.09 8613.565 ;
      RECT 11575.53 187.44 11578.57 8613.565 ;
      RECT 11558.55 188.86 11561.59 8613.565 ;
      RECT 11543.03 187.44 11544.61 8613.565 ;
      RECT 11512.51 187.44 11514.09 8613.565 ;
      RECT 11495.53 188.86 11498.57 8613.565 ;
      RECT 11478.55 187.44 11481.59 8613.565 ;
      RECT 11463.03 188.86 11464.61 8613.565 ;
      RECT 11432.51 187.44 11434.09 8613.565 ;
      RECT 11415.53 188.86 11418.57 8613.565 ;
      RECT 11398.55 188.86 11401.59 8613.565 ;
      RECT 11400.965 187.44 11401.59 8613.565 ;
      RECT 11383.03 187.44 11384.61 8613.565 ;
      RECT 11352.51 188.86 11354.09 8613.565 ;
      RECT 11335.53 187.44 11338.57 8613.565 ;
      RECT 11318.55 187.44 11321.59 8613.565 ;
      RECT 11303.03 187.44 11304.61 8613.565 ;
      RECT 11272.51 188.86 11274.09 8613.565 ;
      RECT 11255.53 188.86 11258.57 8613.565 ;
      RECT 11238.55 187.44 11241.59 8613.565 ;
      RECT 11223.03 187.44 11224.61 8613.565 ;
      RECT 11192.51 188.86 11194.09 8613.565 ;
      RECT 11175.53 187.44 11178.57 8613.565 ;
      RECT 11158.55 187.44 11161.59 8613.565 ;
      RECT 11143.03 187.44 11144.61 8613.565 ;
      RECT 11112.51 188.86 11114.09 8613.565 ;
      RECT 11095.53 187.44 11098.57 8613.565 ;
      RECT 11078.55 188.86 11081.59 8613.565 ;
      RECT 11081.205 187.44 11081.59 8613.565 ;
      RECT 11063.03 187.44 11064.61 8613.565 ;
      RECT 11032.51 187.44 11034.09 8613.565 ;
      RECT 11015.53 187.44 11018.57 8613.565 ;
      RECT 10998.55 188.86 11001.59 8613.565 ;
      RECT 10983.03 187.44 10984.61 8613.565 ;
      RECT 10952.51 187.44 10954.09 8613.565 ;
      RECT 10935.53 188.86 10938.57 8613.565 ;
      RECT 10918.55 187.44 10921.59 8613.565 ;
      RECT 10903.03 188.86 10904.61 8613.565 ;
      RECT 10872.51 187.44 10874.09 8613.565 ;
      RECT 10855.53 188.86 10858.57 8613.565 ;
      RECT 10838.55 188.86 10841.59 8613.565 ;
      RECT 10840.965 187.44 10841.59 8613.565 ;
      RECT 10823.03 187.44 10824.61 8613.565 ;
      RECT 10792.51 188.86 10794.09 8613.565 ;
      RECT 10775.53 187.44 10778.57 8613.565 ;
      RECT 10758.55 187.44 10761.59 8613.565 ;
      RECT 10743.03 187.44 10744.61 8613.565 ;
      RECT 10712.51 188.86 10714.09 8613.565 ;
      RECT 10695.53 188.86 10698.57 8613.565 ;
      RECT 10678.55 187.44 10681.59 8613.565 ;
      RECT 10663.03 187.44 10664.61 8613.565 ;
      RECT 10632.51 188.86 10634.09 8613.565 ;
      RECT 10615.53 187.44 10618.57 8613.565 ;
      RECT 10598.55 187.44 10601.59 8613.565 ;
      RECT 10583.03 187.44 10584.61 8613.565 ;
      RECT 10552.51 188.86 10554.09 8613.565 ;
      RECT 10535.53 187.44 10538.57 8613.565 ;
      RECT 10518.55 188.86 10521.59 8613.565 ;
      RECT 10521.205 187.44 10521.59 8613.565 ;
      RECT 10503.03 187.44 10504.61 8613.565 ;
      RECT 10472.51 187.44 10474.09 8613.565 ;
      RECT 10455.53 187.44 10458.57 8613.565 ;
      RECT 10438.55 188.86 10441.59 8613.565 ;
      RECT 10423.03 187.44 10424.61 8613.565 ;
      RECT 10392.51 187.44 10394.09 8613.565 ;
      RECT 10375.53 188.86 10378.57 8613.565 ;
      RECT 10358.55 187.44 10361.59 8613.565 ;
      RECT 10343.03 188.86 10344.61 8613.565 ;
      RECT 10312.51 187.44 10314.09 8613.565 ;
      RECT 10295.53 188.86 10298.57 8613.565 ;
      RECT 10278.55 188.86 10281.59 8613.565 ;
      RECT 10280.965 187.44 10281.59 8613.565 ;
      RECT 10263.03 187.44 10264.61 8613.565 ;
      RECT 10232.51 188.86 10234.09 8613.565 ;
      RECT 10215.53 187.44 10218.57 8613.565 ;
      RECT 10198.55 187.44 10201.59 8613.565 ;
      RECT 10183.03 187.44 10184.61 8613.565 ;
      RECT 10152.51 188.86 10154.09 8613.565 ;
      RECT 10135.53 188.86 10138.57 8613.565 ;
      RECT 10118.55 187.44 10121.59 8613.565 ;
      RECT 10103.03 187.44 10104.61 8613.565 ;
      RECT 10072.51 188.86 10074.09 8613.565 ;
      RECT 10055.53 187.44 10058.57 8613.565 ;
      RECT 10038.55 187.44 10041.59 8613.565 ;
      RECT 10023.03 187.44 10024.61 8613.565 ;
      RECT 9992.51 188.86 9994.09 8613.565 ;
      RECT 9975.53 187.44 9978.57 8613.565 ;
      RECT 9958.55 188.86 9961.59 8613.565 ;
      RECT 9961.205 187.44 9961.59 8613.565 ;
      RECT 9943.03 187.44 9944.61 8613.565 ;
      RECT 9912.51 187.44 9914.09 8613.565 ;
      RECT 9895.53 187.44 9898.57 8613.565 ;
      RECT 9878.55 188.86 9881.59 8613.565 ;
      RECT 9863.03 187.44 9864.61 8613.565 ;
      RECT 9832.51 187.44 9834.09 8613.565 ;
      RECT 9815.53 188.86 9818.57 8613.565 ;
      RECT 9798.55 187.44 9801.59 8613.565 ;
      RECT 9783.03 188.86 9784.61 8613.565 ;
      RECT 9752.51 187.44 9754.09 8613.565 ;
      RECT 9735.53 188.86 9738.57 8613.565 ;
      RECT 9718.55 188.86 9721.59 8613.565 ;
      RECT 9720.965 187.44 9721.59 8613.565 ;
      RECT 9703.03 187.44 9704.61 8613.565 ;
      RECT 9672.51 188.86 9674.09 8613.565 ;
      RECT 9655.53 187.44 9658.57 8613.565 ;
      RECT 9638.55 187.44 9641.59 8613.565 ;
      RECT 9623.03 187.44 9624.61 8613.565 ;
      RECT 9592.51 188.86 9594.09 8613.565 ;
      RECT 9575.53 188.86 9578.57 8613.565 ;
      RECT 9558.55 187.44 9561.59 8613.565 ;
      RECT 9543.03 187.44 9544.61 8613.565 ;
      RECT 9512.51 188.86 9514.09 8613.565 ;
      RECT 9495.53 187.44 9498.57 8613.565 ;
      RECT 9478.55 187.44 9481.59 8613.565 ;
      RECT 9463.03 187.44 9464.61 8613.565 ;
      RECT 9432.51 188.86 9434.09 8613.565 ;
      RECT 9415.53 187.44 9418.57 8613.565 ;
      RECT 9398.55 188.86 9401.59 8613.565 ;
      RECT 9401.205 187.44 9401.59 8613.565 ;
      RECT 9383.03 187.44 9384.61 8613.565 ;
      RECT 9352.51 187.44 9354.09 8613.565 ;
      RECT 9335.53 187.44 9338.57 8613.565 ;
      RECT 9318.55 188.86 9321.59 8613.565 ;
      RECT 9303.03 187.44 9304.61 8613.565 ;
      RECT 9272.51 187.44 9274.09 8613.565 ;
      RECT 9255.53 188.86 9258.57 8613.565 ;
      RECT 9238.55 187.44 9241.59 8613.565 ;
      RECT 9223.03 188.86 9224.61 8613.565 ;
      RECT 9192.51 187.44 9194.09 8613.565 ;
      RECT 9175.53 188.86 9178.57 8613.565 ;
      RECT 9158.55 188.86 9161.59 8613.565 ;
      RECT 9160.965 187.44 9161.59 8613.565 ;
      RECT 9143.03 187.44 9144.61 8613.565 ;
      RECT 9112.51 188.86 9114.09 8613.565 ;
      RECT 9095.53 187.44 9098.57 8613.565 ;
      RECT 9078.55 187.44 9081.59 8613.565 ;
      RECT 9063.03 187.44 9064.61 8613.565 ;
      RECT 9032.51 188.86 9034.09 8613.565 ;
      RECT 9015.53 188.86 9018.57 8613.565 ;
      RECT 8998.55 187.44 9001.59 8613.565 ;
      RECT 8983.03 187.44 8984.61 8613.565 ;
      RECT 8952.51 188.86 8954.09 8613.565 ;
      RECT 8935.53 187.44 8938.57 8613.565 ;
      RECT 8918.55 187.44 8921.59 8613.565 ;
      RECT 8903.03 187.44 8904.61 8613.565 ;
      RECT 8872.51 188.86 8874.09 8613.565 ;
      RECT 8855.53 187.44 8858.57 8613.565 ;
      RECT 8838.55 188.86 8841.59 8613.565 ;
      RECT 8841.205 187.44 8841.59 8613.565 ;
      RECT 8823.03 187.44 8824.61 8613.565 ;
      RECT 8792.51 187.44 8794.09 8613.565 ;
      RECT 8775.53 187.44 8778.57 8613.565 ;
      RECT 8758.55 188.86 8761.59 8613.565 ;
      RECT 8743.03 187.44 8744.61 8613.565 ;
      RECT 8712.51 187.44 8714.09 8613.565 ;
      RECT 8695.53 188.86 8698.57 8613.565 ;
      RECT 8678.55 187.44 8681.59 8613.565 ;
      RECT 8663.03 188.86 8664.61 8613.565 ;
      RECT 8632.51 187.44 8634.09 8613.565 ;
      RECT 8615.53 188.86 8618.57 8613.565 ;
      RECT 8598.55 188.86 8601.59 8613.565 ;
      RECT 8600.965 187.44 8601.59 8613.565 ;
      RECT 8583.03 187.44 8584.61 8613.565 ;
      RECT 8552.51 188.86 8554.09 8613.565 ;
      RECT 8535.53 187.44 8538.57 8613.565 ;
      RECT 8518.55 187.44 8521.59 8613.565 ;
      RECT 8503.03 187.44 8504.61 8613.565 ;
      RECT 8472.51 188.86 8474.09 8613.565 ;
      RECT 8455.53 188.86 8458.57 8613.565 ;
      RECT 8438.55 187.44 8441.59 8613.565 ;
      RECT 8423.03 187.44 8424.61 8613.565 ;
      RECT 8392.51 188.86 8394.09 8613.565 ;
      RECT 8375.53 187.44 8378.57 8613.565 ;
      RECT 8358.55 187.44 8361.59 8613.565 ;
      RECT 8343.03 187.44 8344.61 8613.565 ;
      RECT 8312.51 188.86 8314.09 8613.565 ;
      RECT 8295.53 187.44 8298.57 8613.565 ;
      RECT 8278.55 188.86 8281.59 8613.565 ;
      RECT 8281.205 187.44 8281.59 8613.565 ;
      RECT 8263.03 187.44 8264.61 8613.565 ;
      RECT 8232.51 187.44 8234.09 8613.565 ;
      RECT 8215.53 187.44 8218.57 8613.565 ;
      RECT 8198.55 188.86 8201.59 8613.565 ;
      RECT 8183.03 187.44 8184.61 8613.565 ;
      RECT 8152.51 187.44 8154.09 8613.565 ;
      RECT 8135.53 188.86 8138.57 8613.565 ;
      RECT 8118.55 187.44 8121.59 8613.565 ;
      RECT 8103.03 188.86 8104.61 8613.565 ;
      RECT 8072.51 187.44 8074.09 8613.565 ;
      RECT 8055.53 188.86 8058.57 8613.565 ;
      RECT 8038.55 188.86 8041.59 8613.565 ;
      RECT 8040.965 187.44 8041.59 8613.565 ;
      RECT 8023.03 187.44 8024.61 8613.565 ;
      RECT 7992.51 188.86 7994.09 8613.565 ;
      RECT 7975.53 187.44 7978.57 8613.565 ;
      RECT 7958.55 187.44 7961.59 8613.565 ;
      RECT 7943.03 187.44 7944.61 8613.565 ;
      RECT 7912.51 188.86 7914.09 8613.565 ;
      RECT 7895.53 188.86 7898.57 8613.565 ;
      RECT 7878.55 187.44 7881.59 8613.565 ;
      RECT 7863.03 187.44 7864.61 8613.565 ;
      RECT 7832.51 188.86 7834.09 8613.565 ;
      RECT 7815.53 187.44 7818.57 8613.565 ;
      RECT 7798.55 187.44 7801.59 8613.565 ;
      RECT 7783.03 187.44 7784.61 8613.565 ;
      RECT 7752.51 188.86 7754.09 8613.565 ;
      RECT 7735.53 187.44 7738.57 8613.565 ;
      RECT 7718.55 188.86 7721.59 8613.565 ;
      RECT 7721.205 187.44 7721.59 8613.565 ;
      RECT 7703.03 187.44 7704.61 8613.565 ;
      RECT 7672.51 187.44 7674.09 8613.565 ;
      RECT 7655.53 187.44 7658.57 8613.565 ;
      RECT 7638.55 188.86 7641.59 8613.565 ;
      RECT 7623.03 187.44 7624.61 8613.565 ;
      RECT 7592.51 187.44 7594.09 8613.565 ;
      RECT 7575.53 188.86 7578.57 8613.565 ;
      RECT 7558.55 187.44 7561.59 8613.565 ;
      RECT 7543.03 188.86 7544.61 8613.565 ;
      RECT 7512.51 187.44 7514.09 8613.565 ;
      RECT 7495.53 188.86 7498.57 8613.565 ;
      RECT 7478.55 188.86 7481.59 8613.565 ;
      RECT 7480.965 187.44 7481.59 8613.565 ;
      RECT 7463.03 187.44 7464.61 8613.565 ;
      RECT 7432.51 188.86 7434.09 8613.565 ;
      RECT 7415.53 187.44 7418.57 8613.565 ;
      RECT 7398.55 187.44 7401.59 8613.565 ;
      RECT 7383.03 187.44 7384.61 8613.565 ;
      RECT 7352.51 188.86 7354.09 8613.565 ;
      RECT 7335.53 188.86 7338.57 8613.565 ;
      RECT 7318.55 187.44 7321.59 8613.565 ;
      RECT 7303.03 187.44 7304.61 8613.565 ;
      RECT 7272.51 188.86 7274.09 8613.565 ;
      RECT 7255.53 187.44 7258.57 8613.565 ;
      RECT 7238.55 187.44 7241.59 8613.565 ;
      RECT 7223.03 187.44 7224.61 8613.565 ;
      RECT 7192.51 188.86 7194.09 8613.565 ;
      RECT 7175.53 187.44 7178.57 8613.565 ;
      RECT 7158.55 188.86 7161.59 8613.565 ;
      RECT 7161.205 187.44 7161.59 8613.565 ;
      RECT 7143.03 187.44 7144.61 8613.565 ;
      RECT 7112.51 187.44 7114.09 8613.565 ;
      RECT 7095.53 187.44 7098.57 8613.565 ;
      RECT 7078.55 188.86 7081.59 8613.565 ;
      RECT 7063.03 187.44 7064.61 8613.565 ;
      RECT 7032.51 187.44 7034.09 8613.565 ;
      RECT 7015.53 188.86 7018.57 8613.565 ;
      RECT 6998.55 187.44 7001.59 8613.565 ;
      RECT 6983.03 188.86 6984.61 8613.565 ;
      RECT 6952.51 187.44 6954.09 8613.565 ;
      RECT 6935.53 188.86 6938.57 8613.565 ;
      RECT 6918.55 188.86 6921.59 8613.565 ;
      RECT 6920.965 187.44 6921.59 8613.565 ;
      RECT 6903.03 187.44 6904.61 8613.565 ;
      RECT 6872.51 188.86 6874.09 8613.565 ;
      RECT 6855.53 187.44 6858.57 8613.565 ;
      RECT 6838.55 187.44 6841.59 8613.565 ;
      RECT 6823.03 187.44 6824.61 8613.565 ;
      RECT 6792.51 188.86 6794.09 8613.565 ;
      RECT 6775.53 188.86 6778.57 8613.565 ;
      RECT 6758.55 187.44 6761.59 8613.565 ;
      RECT 6743.03 187.44 6744.61 8613.565 ;
      RECT 6712.51 188.86 6714.09 8613.565 ;
      RECT 6695.53 187.44 6698.57 8613.565 ;
      RECT 6678.55 187.44 6681.59 8613.565 ;
      RECT 6663.03 187.44 6664.61 8613.565 ;
      RECT 6632.51 188.86 6634.09 8613.565 ;
      RECT 6615.53 187.44 6618.57 8613.565 ;
      RECT 6598.55 188.86 6601.59 8613.565 ;
      RECT 6601.205 187.44 6601.59 8613.565 ;
      RECT 6583.03 187.44 6584.61 8613.565 ;
      RECT 6552.51 187.44 6554.09 8613.565 ;
      RECT 6535.53 187.44 6538.57 8613.565 ;
      RECT 6518.55 188.86 6521.59 8613.565 ;
      RECT 6503.03 187.44 6504.61 8613.565 ;
      RECT 6472.51 187.44 6474.09 8613.565 ;
      RECT 6455.53 188.86 6458.57 8613.565 ;
      RECT 6438.55 187.44 6441.59 8613.565 ;
      RECT 6423.03 188.86 6424.61 8613.565 ;
      RECT 6392.51 187.44 6394.09 8613.565 ;
      RECT 6375.53 188.86 6378.57 8613.565 ;
      RECT 6358.55 188.86 6361.59 8613.565 ;
      RECT 6360.965 187.44 6361.59 8613.565 ;
      RECT 6343.03 187.44 6344.61 8613.565 ;
      RECT 6312.51 188.86 6314.09 8613.565 ;
      RECT 6295.53 187.44 6298.57 8613.565 ;
      RECT 6278.55 187.44 6281.59 8613.565 ;
      RECT 6263.03 187.44 6264.61 8613.565 ;
      RECT 6232.51 188.86 6234.09 8613.565 ;
      RECT 6215.53 188.86 6218.57 8613.565 ;
      RECT 6198.55 187.44 6201.59 8613.565 ;
      RECT 6183.03 187.44 6184.61 8613.565 ;
      RECT 6152.51 188.86 6154.09 8613.565 ;
      RECT 6135.53 187.44 6138.57 8613.565 ;
      RECT 6118.55 187.44 6121.59 8613.565 ;
      RECT 6103.03 187.44 6104.61 8613.565 ;
      RECT 6072.51 188.86 6074.09 8613.565 ;
      RECT 6055.53 187.44 6058.57 8613.565 ;
      RECT 6038.55 188.86 6041.59 8613.565 ;
      RECT 6041.205 187.44 6041.59 8613.565 ;
      RECT 6023.03 187.44 6024.61 8613.565 ;
      RECT 5992.51 187.44 5994.09 8613.565 ;
      RECT 5975.53 187.44 5978.57 8613.565 ;
      RECT 5958.55 188.86 5961.59 8613.565 ;
      RECT 5943.03 187.44 5944.61 8613.565 ;
      RECT 5912.51 187.44 5914.09 8613.565 ;
      RECT 5895.53 188.86 5898.57 8613.565 ;
      RECT 5878.55 187.44 5881.59 8613.565 ;
      RECT 5863.03 188.86 5864.61 8613.565 ;
      RECT 5832.51 187.44 5834.09 8613.565 ;
      RECT 5815.53 188.86 5818.57 8613.565 ;
      RECT 5798.55 188.86 5801.59 8613.565 ;
      RECT 5800.965 187.44 5801.59 8613.565 ;
      RECT 5783.03 187.44 5784.61 8613.565 ;
      RECT 5752.51 188.86 5754.09 8613.565 ;
      RECT 5735.53 187.44 5738.57 8613.565 ;
      RECT 5718.55 187.44 5721.59 8613.565 ;
      RECT 5703.03 187.44 5704.61 8613.565 ;
      RECT 5672.51 188.86 5674.09 8613.565 ;
      RECT 5655.53 188.86 5658.57 8613.565 ;
      RECT 5638.55 187.44 5641.59 8613.565 ;
      RECT 5623.03 187.44 5624.61 8613.565 ;
      RECT 5592.51 188.86 5594.09 8613.565 ;
      RECT 5575.53 187.44 5578.57 8613.565 ;
      RECT 5558.55 187.44 5561.59 8613.565 ;
      RECT 5543.03 187.44 5544.61 8613.565 ;
      RECT 5512.51 188.86 5514.09 8613.565 ;
      RECT 5495.53 187.44 5498.57 8613.565 ;
      RECT 5478.55 188.86 5481.59 8613.565 ;
      RECT 5481.205 187.44 5481.59 8613.565 ;
      RECT 5463.03 187.44 5464.61 8613.565 ;
      RECT 5432.51 187.44 5434.09 8613.565 ;
      RECT 5415.53 187.44 5418.57 8613.565 ;
      RECT 5398.55 188.86 5401.59 8613.565 ;
      RECT 5383.03 187.44 5384.61 8613.565 ;
      RECT 5352.51 187.44 5354.09 8613.565 ;
      RECT 5335.53 188.86 5338.57 8613.565 ;
      RECT 5318.55 187.44 5321.59 8613.565 ;
      RECT 5303.03 188.86 5304.61 8613.565 ;
      RECT 5272.51 187.44 5274.09 8613.565 ;
      RECT 5255.53 188.86 5258.57 8613.565 ;
      RECT 5238.55 188.86 5241.59 8613.565 ;
      RECT 5240.965 187.44 5241.59 8613.565 ;
      RECT 5223.03 187.44 5224.61 8613.565 ;
      RECT 5192.51 188.86 5194.09 8613.565 ;
      RECT 5175.53 187.44 5178.57 8613.565 ;
      RECT 5158.55 187.44 5161.59 8613.565 ;
      RECT 5143.03 187.44 5144.61 8613.565 ;
      RECT 5112.51 188.86 5114.09 8613.565 ;
      RECT 5095.53 188.86 5098.57 8613.565 ;
      RECT 5078.55 187.44 5081.59 8613.565 ;
      RECT 5063.03 187.44 5064.61 8613.565 ;
      RECT 5032.51 188.86 5034.09 8613.565 ;
      RECT 5015.53 187.44 5018.57 8613.565 ;
      RECT 4998.55 187.44 5001.59 8613.565 ;
      RECT 4983.03 187.44 4984.61 8613.565 ;
      RECT 4952.51 188.86 4954.09 8613.565 ;
      RECT 4935.53 187.44 4938.57 8613.565 ;
      RECT 4918.55 188.86 4921.59 8613.565 ;
      RECT 4921.205 187.44 4921.59 8613.565 ;
      RECT 4903.03 187.44 4904.61 8613.565 ;
      RECT 4872.51 187.44 4874.09 8613.565 ;
      RECT 4855.53 187.44 4858.57 8613.565 ;
      RECT 4838.55 188.86 4841.59 8613.565 ;
      RECT 4823.03 187.44 4824.61 8613.565 ;
      RECT 4792.51 187.44 4794.09 8613.565 ;
      RECT 4775.53 188.86 4778.57 8613.565 ;
      RECT 4758.55 187.44 4761.59 8613.565 ;
      RECT 4743.03 188.86 4744.61 8613.565 ;
      RECT 4712.51 187.44 4714.09 8613.565 ;
      RECT 4695.53 188.86 4698.57 8613.565 ;
      RECT 4678.55 188.86 4681.59 8613.565 ;
      RECT 4680.965 187.44 4681.59 8613.565 ;
      RECT 4663.03 187.44 4664.61 8613.565 ;
      RECT 4632.51 188.86 4634.09 8613.565 ;
      RECT 4615.53 187.44 4618.57 8613.565 ;
      RECT 4598.55 187.44 4601.59 8613.565 ;
      RECT 4583.03 187.44 4584.61 8613.565 ;
      RECT 4552.51 188.86 4554.09 8613.565 ;
      RECT 4535.53 188.86 4538.57 8613.565 ;
      RECT 4518.55 187.44 4521.59 8613.565 ;
      RECT 4503.03 187.44 4504.61 8613.565 ;
      RECT 4472.51 188.86 4474.09 8613.565 ;
      RECT 4455.53 187.44 4458.57 8613.565 ;
      RECT 4438.55 187.44 4441.59 8613.565 ;
      RECT 4423.03 187.44 4424.61 8613.565 ;
      RECT 4392.51 188.86 4394.09 8613.565 ;
      RECT 4375.53 187.44 4378.57 8613.565 ;
      RECT 4358.55 188.86 4361.59 8613.565 ;
      RECT 4361.205 187.44 4361.59 8613.565 ;
      RECT 4343.03 187.44 4344.61 8613.565 ;
      RECT 4312.51 187.44 4314.09 8613.565 ;
      RECT 4295.53 187.44 4298.57 8613.565 ;
      RECT 4278.55 188.86 4281.59 8613.565 ;
      RECT 4263.03 187.44 4264.61 8613.565 ;
      RECT 4232.51 187.44 4234.09 8613.565 ;
      RECT 4215.53 188.86 4218.57 8613.565 ;
      RECT 4198.55 187.44 4201.59 8613.565 ;
      RECT 4183.03 188.86 4184.61 8613.565 ;
      RECT 4152.51 187.44 4154.09 8613.565 ;
      RECT 4135.53 188.86 4138.57 8613.565 ;
      RECT 4118.55 188.86 4121.59 8613.565 ;
      RECT 4120.965 187.44 4121.59 8613.565 ;
      RECT 4103.03 187.44 4104.61 8613.565 ;
      RECT 4072.51 188.86 4074.09 8613.565 ;
      RECT 4055.53 187.44 4058.57 8613.565 ;
      RECT 4038.55 187.44 4041.59 8613.565 ;
      RECT 4023.03 187.44 4024.61 8613.565 ;
      RECT 3992.51 188.86 3994.09 8613.565 ;
      RECT 3975.53 188.86 3978.57 8613.565 ;
      RECT 3958.55 187.44 3961.59 8613.565 ;
      RECT 3943.03 187.44 3944.61 8613.565 ;
      RECT 3912.51 188.86 3914.09 8613.565 ;
      RECT 3895.53 187.44 3898.57 8613.565 ;
      RECT 3878.55 187.44 3881.59 8613.565 ;
      RECT 3863.03 187.44 3864.61 8613.565 ;
      RECT 3832.51 188.86 3834.09 8613.565 ;
      RECT 3815.53 187.44 3818.57 8613.565 ;
      RECT 3798.55 188.86 3801.59 8613.565 ;
      RECT 3801.205 187.44 3801.59 8613.565 ;
      RECT 3783.03 187.44 3784.61 8613.565 ;
      RECT 3752.51 187.44 3754.09 8613.565 ;
      RECT 3735.53 187.44 3738.57 8613.565 ;
      RECT 3718.55 188.86 3721.59 8613.565 ;
      RECT 3703.03 187.44 3704.61 8613.565 ;
      RECT 3672.51 187.44 3674.09 8613.565 ;
      RECT 3655.53 188.86 3658.57 8613.565 ;
      RECT 3638.55 187.44 3641.59 8613.565 ;
      RECT 3623.03 188.86 3624.61 8613.565 ;
      RECT 3592.51 187.44 3594.09 8613.565 ;
      RECT 3575.53 188.86 3578.57 8613.565 ;
      RECT 3558.55 188.86 3561.59 8613.565 ;
      RECT 3560.965 187.44 3561.59 8613.565 ;
      RECT 3543.03 187.44 3544.61 8613.565 ;
      RECT 3512.51 188.86 3514.09 8613.565 ;
      RECT 3495.53 187.44 3498.57 8613.565 ;
      RECT 3478.55 187.44 3481.59 8613.565 ;
      RECT 3463.03 187.44 3464.61 8613.565 ;
      RECT 3432.51 188.86 3434.09 8613.565 ;
      RECT 3415.53 188.86 3418.57 8613.565 ;
      RECT 3398.55 187.44 3401.59 8613.565 ;
      RECT 3383.03 187.44 3384.61 8613.565 ;
      RECT 3352.51 188.86 3354.09 8613.565 ;
      RECT 3335.53 187.44 3338.57 8613.565 ;
      RECT 3318.55 187.44 3321.59 8613.565 ;
      RECT 3303.03 187.44 3304.61 8613.565 ;
      RECT 3272.51 188.86 3274.09 8613.565 ;
      RECT 3255.53 187.44 3258.57 8613.565 ;
      RECT 3238.55 188.86 3241.59 8613.565 ;
      RECT 3241.205 187.44 3241.59 8613.565 ;
      RECT 3223.03 187.44 3224.61 8613.565 ;
      RECT 3192.51 187.44 3194.09 8613.565 ;
      RECT 3175.53 187.44 3178.57 8613.565 ;
      RECT 3158.55 188.86 3161.59 8613.565 ;
      RECT 3143.03 187.44 3144.61 8613.565 ;
      RECT 3112.51 187.44 3114.09 8613.565 ;
      RECT 3095.53 188.86 3098.57 8613.565 ;
      RECT 3078.55 187.44 3081.59 8613.565 ;
      RECT 3063.03 188.86 3064.61 8613.565 ;
      RECT 3032.51 187.44 3034.09 8613.565 ;
      RECT 3015.53 188.86 3018.57 8613.565 ;
      RECT 2998.55 188.86 3001.59 8613.565 ;
      RECT 3000.965 187.44 3001.59 8613.565 ;
      RECT 2983.03 187.44 2984.61 8613.565 ;
      RECT 2952.51 188.86 2954.09 8613.565 ;
      RECT 2935.53 187.44 2938.57 8613.565 ;
      RECT 2918.55 187.44 2921.59 8613.565 ;
      RECT 2903.03 187.44 2904.61 8613.565 ;
      RECT 2872.51 188.86 2874.09 8613.565 ;
      RECT 2855.53 188.86 2858.57 8613.565 ;
      RECT 2838.55 187.44 2841.59 8613.565 ;
      RECT 2823.03 187.44 2824.61 8613.565 ;
      RECT 2792.51 188.86 2794.09 8613.565 ;
      RECT 2775.53 187.44 2778.57 8613.565 ;
      RECT 2758.55 187.44 2761.59 8613.565 ;
      RECT 2743.03 187.44 2744.61 8613.565 ;
      RECT 2712.51 188.86 2714.09 8613.565 ;
      RECT 2695.53 187.44 2698.57 8613.565 ;
      RECT 2678.55 188.86 2681.59 8613.565 ;
      RECT 2681.205 187.44 2681.59 8613.565 ;
      RECT 2663.03 187.44 2664.61 8613.565 ;
      RECT 2632.51 187.44 2634.09 8613.565 ;
      RECT 2615.53 187.44 2618.57 8613.565 ;
      RECT 2598.55 188.86 2601.59 8613.565 ;
      RECT 2583.03 187.44 2584.61 8613.565 ;
      RECT 2552.51 187.44 2554.09 8613.565 ;
      RECT 2535.53 188.86 2538.57 8613.565 ;
      RECT 2518.55 187.44 2521.59 8613.565 ;
      RECT 2503.03 188.86 2504.61 8613.565 ;
      RECT 2472.51 187.44 2474.09 8613.565 ;
      RECT 2455.53 188.86 2458.57 8613.565 ;
      RECT 2438.55 188.86 2441.59 8613.565 ;
      RECT 2440.965 187.44 2441.59 8613.565 ;
      RECT 2423.03 187.44 2424.61 8613.565 ;
      RECT 2392.51 188.86 2394.09 8613.565 ;
      RECT 2375.53 187.44 2378.57 8613.565 ;
      RECT 2358.55 187.44 2361.59 8613.565 ;
      RECT 2343.03 187.44 2344.61 8613.565 ;
      RECT 2312.51 188.86 2314.09 8613.565 ;
      RECT 2295.53 188.86 2298.57 8613.565 ;
      RECT 2278.55 187.44 2281.59 8613.565 ;
      RECT 2263.03 187.44 2264.61 8613.565 ;
      RECT 2232.51 188.86 2234.09 8613.565 ;
      RECT 2215.53 187.44 2218.57 8613.565 ;
      RECT 2198.55 187.44 2201.59 8613.565 ;
      RECT 2183.03 187.44 2184.61 8613.565 ;
      RECT 2152.51 188.86 2154.09 8613.565 ;
      RECT 2135.53 187.44 2138.57 8613.565 ;
      RECT 2118.55 188.86 2121.59 8613.565 ;
      RECT 2121.205 187.44 2121.59 8613.565 ;
      RECT 2103.03 187.44 2104.61 8613.565 ;
      RECT 2072.51 187.44 2074.09 8613.565 ;
      RECT 2055.53 187.44 2058.57 8613.565 ;
      RECT 2038.55 188.86 2041.59 8613.565 ;
      RECT 2023.03 187.44 2024.61 8613.565 ;
      RECT 1992.51 187.44 1994.09 8613.565 ;
      RECT 1975.53 188.86 1978.57 8613.565 ;
      RECT 1958.55 187.44 1961.59 8613.565 ;
      RECT 1943.03 188.86 1944.61 8613.565 ;
      RECT 1912.51 187.44 1914.09 8613.565 ;
      RECT 1895.53 188.86 1898.57 8613.565 ;
      RECT 1878.55 188.86 1881.59 8613.565 ;
      RECT 1880.965 187.44 1881.59 8613.565 ;
      RECT 1863.03 187.44 1864.61 8613.565 ;
      RECT 1832.51 188.86 1834.09 8613.565 ;
      RECT 1815.53 187.44 1818.57 8613.565 ;
      RECT 1798.55 187.44 1801.59 8613.565 ;
      RECT 1783.03 187.44 1784.61 8613.565 ;
      RECT 1752.51 188.86 1754.09 8613.565 ;
      RECT 1735.53 188.86 1738.57 8613.565 ;
      RECT 1718.55 187.44 1721.59 8613.565 ;
      RECT 1703.03 187.44 1704.61 8613.565 ;
      RECT 1672.51 188.86 1674.09 8613.565 ;
      RECT 1655.53 187.44 1658.57 8613.565 ;
      RECT 1638.55 187.44 1641.59 8613.565 ;
      RECT 1623.03 187.44 1624.61 8613.565 ;
      RECT 1592.51 188.86 1594.09 8613.565 ;
      RECT 1575.53 187.44 1578.57 8613.565 ;
      RECT 1558.55 188.86 1561.59 8613.565 ;
      RECT 1561.205 187.44 1561.59 8613.565 ;
      RECT 1543.03 187.44 1544.61 8613.565 ;
      RECT 1512.51 187.44 1514.09 8613.565 ;
      RECT 1495.53 187.44 1498.57 8613.565 ;
      RECT 1478.55 188.86 1481.59 8613.565 ;
      RECT 1463.03 187.44 1464.61 8613.565 ;
      RECT 1432.51 187.44 1434.09 8613.565 ;
      RECT 1415.53 188.86 1418.57 8613.565 ;
      RECT 1398.55 187.44 1401.59 8613.565 ;
      RECT 1383.03 188.86 1384.61 8613.565 ;
      RECT 1352.51 187.44 1354.09 8613.565 ;
      RECT 1335.53 188.86 1338.57 8613.565 ;
      RECT 1318.55 188.86 1321.59 8613.565 ;
      RECT 1320.965 187.44 1321.59 8613.565 ;
      RECT 1303.03 187.44 1304.61 8613.565 ;
      RECT 1272.51 188.86 1274.09 8613.565 ;
      RECT 1255.53 187.44 1258.57 8613.565 ;
      RECT 1238.55 187.44 1241.59 8613.565 ;
      RECT 1223.03 187.44 1224.61 8613.565 ;
      RECT 1192.51 188.86 1194.09 8613.565 ;
      RECT 1175.53 188.86 1178.57 8613.565 ;
      RECT 1158.55 187.44 1161.59 8613.565 ;
      RECT 1143.03 187.44 1144.61 8613.565 ;
      RECT 1112.51 188.86 1114.09 8613.565 ;
      RECT 1095.53 187.44 1098.57 8613.565 ;
      RECT 1078.55 187.44 1081.59 8613.565 ;
      RECT 1063.03 187.44 1064.61 8613.565 ;
      RECT 1032.51 188.86 1034.09 8613.565 ;
      RECT 1015.53 187.44 1018.57 8613.565 ;
      RECT 998.55 188.86 1001.59 8613.565 ;
      RECT 1001.205 187.44 1001.59 8613.565 ;
      RECT 983.03 187.44 984.61 8613.565 ;
      RECT 952.51 187.44 954.09 8613.565 ;
      RECT 935.53 187.44 938.57 8613.565 ;
      RECT 918.55 188.86 921.59 8613.565 ;
      RECT 903.03 187.44 904.61 8613.565 ;
      RECT 872.51 187.44 874.09 8613.565 ;
      RECT 855.53 188.86 858.57 8613.565 ;
      RECT 838.55 187.44 841.59 8613.565 ;
      RECT 823.03 188.86 824.61 8613.565 ;
      RECT 792.51 187.44 794.09 8613.565 ;
      RECT 775.53 188.86 778.57 8613.565 ;
      RECT 758.55 188.86 761.59 8613.565 ;
      RECT 760.965 187.44 761.59 8613.565 ;
      RECT 743.03 187.44 744.61 8613.565 ;
      RECT 712.51 188.86 714.09 8613.565 ;
      RECT 695.53 187.44 698.57 8613.565 ;
      RECT 678.55 187.44 681.59 8613.565 ;
      RECT 663.03 187.44 664.61 8613.565 ;
      RECT 632.51 188.86 634.09 8613.565 ;
      RECT 615.53 188.86 618.57 8613.565 ;
      RECT 598.55 187.44 601.59 8613.565 ;
      RECT 583.03 187.44 584.61 8613.565 ;
      RECT 552.51 188.86 554.09 8613.565 ;
      RECT 535.53 187.44 538.57 8613.565 ;
      RECT 518.55 187.44 521.59 8613.565 ;
      RECT 503.03 187.44 504.61 8613.565 ;
      RECT 472.51 188.86 474.09 8613.565 ;
      RECT 17832.51 187.44 17833.125 8613.565 ;
      RECT 17272.51 187.44 17273.125 8613.565 ;
      RECT 16712.51 187.44 16713.125 8613.565 ;
      RECT 16152.51 187.44 16153.125 8613.565 ;
      RECT 15592.51 187.44 15593.125 8613.565 ;
      RECT 15032.51 187.44 15033.125 8613.565 ;
      RECT 14472.51 187.44 14473.125 8613.565 ;
      RECT 13912.51 187.44 13913.125 8613.565 ;
      RECT 13352.51 187.44 13353.125 8613.565 ;
      RECT 12792.51 187.44 12793.125 8613.565 ;
      RECT 12232.51 187.44 12233.125 8613.565 ;
      RECT 11672.51 187.44 11673.125 8613.565 ;
      RECT 11112.51 187.44 11113.125 8613.565 ;
      RECT 10552.51 187.44 10553.125 8613.565 ;
      RECT 9992.51 187.44 9993.125 8613.565 ;
      RECT 9432.51 187.44 9433.125 8613.565 ;
      RECT 8872.51 187.44 8873.125 8613.565 ;
      RECT 8312.51 187.44 8313.125 8613.565 ;
      RECT 7752.51 187.44 7753.125 8613.565 ;
      RECT 7192.51 187.44 7193.125 8613.565 ;
      RECT 6632.51 187.44 6633.125 8613.565 ;
      RECT 6072.51 187.44 6073.125 8613.565 ;
      RECT 5512.51 187.44 5513.125 8613.565 ;
      RECT 4952.51 187.44 4953.125 8613.565 ;
      RECT 4392.51 187.44 4393.125 8613.565 ;
      RECT 3832.51 187.44 3833.125 8613.565 ;
      RECT 3272.51 187.44 3273.125 8613.565 ;
      RECT 2712.51 187.44 2713.125 8613.565 ;
      RECT 2152.51 187.44 2153.125 8613.565 ;
      RECT 1592.51 187.44 1593.125 8613.565 ;
      RECT 1032.51 187.44 1033.125 8613.565 ;
      RECT 472.51 187.44 473.125 8613.565 ;
    LAYER TOP_M ;
      RECT 18368.56 339.555 18490.46 372.555 ;
      RECT 18368.56 382.555 18490.46 415.555 ;
      RECT 18368.56 425.555 18490.46 458.555 ;
      RECT 18368.56 468.555 18490.46 501.555 ;
      RECT 18370 191.275 18488.86 193.275 ;
      RECT 18368.56 196.245 18488.86 210.275 ;
      RECT 18368.56 213.245 18488.86 227.275 ;
      RECT 18368.56 230.245 18488.86 258.275 ;
      RECT 18368.56 261.245 18488.86 289.275 ;
      RECT 18368.56 292.245 18488.86 306.275 ;
      RECT 18368.56 309.245 18488.86 323.275 ;
      RECT 18368.99 505.445 18488.86 506.445 ;
      RECT 18368.99 508.445 18488.86 509.445 ;
      RECT 18368.17 512.265 18488.86 514.265 ;
      RECT 18465.79 521.56 18488.86 522.68 ;
      RECT 18465.79 535.975 18488.86 540.585 ;
      RECT 18465.79 542.585 18488.86 547.195 ;
      RECT 18465.79 549.195 18488.86 550.315 ;
      RECT 18465.79 558.435 18488.86 564.205 ;
      RECT 18465.79 566.205 18488.86 577.745 ;
      RECT 18465.79 579.745 18488.86 585.515 ;
      RECT 18465.79 593.635 18488.86 594.755 ;
      RECT 18465.79 596.755 18488.86 601.365 ;
      RECT 18465.79 603.365 18488.86 612.585 ;
      RECT 18465.79 614.585 18488.86 619.195 ;
      RECT 18465.79 621.195 18488.86 622.315 ;
      RECT 18465.79 630.435 18488.86 636.205 ;
      RECT 18465.79 638.205 18488.86 649.745 ;
      RECT 18465.79 651.745 18488.86 657.515 ;
      RECT 18465.79 665.635 18488.86 666.755 ;
      RECT 18465.79 668.755 18488.86 673.365 ;
      RECT 18465.79 675.365 18488.86 684.585 ;
      RECT 18465.79 686.585 18488.86 691.195 ;
      RECT 18465.79 693.195 18488.86 694.315 ;
      RECT 18465.79 702.435 18488.86 708.205 ;
      RECT 18465.79 710.205 18488.86 721.745 ;
      RECT 18465.79 723.745 18488.86 729.515 ;
      RECT 18465.79 737.635 18488.86 738.755 ;
      RECT 18465.79 740.755 18488.86 745.365 ;
      RECT 18465.79 747.365 18488.86 756.585 ;
      RECT 18465.79 758.585 18488.86 763.195 ;
      RECT 18465.79 765.195 18488.86 766.315 ;
      RECT 18465.79 774.435 18488.86 780.205 ;
      RECT 18465.79 782.205 18488.86 793.745 ;
      RECT 18465.79 795.745 18488.86 801.515 ;
      RECT 18465.79 809.635 18488.86 810.755 ;
      RECT 18465.79 812.755 18488.86 817.365 ;
      RECT 18465.79 819.365 18488.86 828.585 ;
      RECT 18465.79 830.585 18488.86 835.195 ;
      RECT 18465.79 837.195 18488.86 838.315 ;
      RECT 18465.79 846.435 18488.86 852.205 ;
      RECT 18465.79 854.205 18488.86 865.745 ;
      RECT 18465.79 867.745 18488.86 873.515 ;
      RECT 18465.79 881.635 18488.86 882.755 ;
      RECT 18465.79 884.755 18488.86 889.365 ;
      RECT 18465.79 891.365 18488.86 900.585 ;
      RECT 18465.79 902.585 18488.86 907.195 ;
      RECT 18465.79 909.195 18488.86 910.315 ;
      RECT 18465.79 918.435 18488.86 924.205 ;
      RECT 18465.79 926.205 18488.86 937.745 ;
      RECT 18465.79 939.745 18488.86 945.515 ;
      RECT 18465.79 953.635 18488.86 954.755 ;
      RECT 18465.79 956.755 18488.86 961.365 ;
      RECT 18465.79 963.365 18488.86 972.585 ;
      RECT 18465.79 974.585 18488.86 979.195 ;
      RECT 18465.79 981.195 18488.86 982.315 ;
      RECT 18465.79 990.435 18488.86 996.205 ;
      RECT 18465.79 998.205 18488.86 1009.745 ;
      RECT 18465.79 1011.745 18488.86 1017.515 ;
      RECT 18465.79 1025.635 18488.86 1026.755 ;
      RECT 18465.79 1028.755 18488.86 1033.365 ;
      RECT 18465.79 1035.365 18488.86 1044.585 ;
      RECT 18465.79 1046.585 18488.86 1051.195 ;
      RECT 18465.79 1053.195 18488.86 1054.315 ;
      RECT 18465.79 1062.435 18488.86 1068.205 ;
      RECT 18465.79 1070.205 18488.86 1081.745 ;
      RECT 18465.79 1083.745 18488.86 1089.515 ;
      RECT 18465.79 1097.635 18488.86 1098.755 ;
      RECT 18465.79 1100.755 18488.86 1105.365 ;
      RECT 18465.79 1107.365 18488.86 1116.585 ;
      RECT 18465.79 1118.585 18488.86 1123.195 ;
      RECT 18465.79 1125.195 18488.86 1126.315 ;
      RECT 18465.79 1134.435 18488.86 1140.205 ;
      RECT 18465.79 1142.205 18488.86 1153.745 ;
      RECT 18465.79 1155.745 18488.86 1161.515 ;
      RECT 18465.79 1169.635 18488.86 1170.755 ;
      RECT 18465.79 1172.755 18488.86 1177.365 ;
      RECT 18465.79 1179.365 18488.86 1188.585 ;
      RECT 18465.79 1190.585 18488.86 1195.195 ;
      RECT 18465.79 1197.195 18488.86 1198.315 ;
      RECT 18465.79 1206.435 18488.86 1212.205 ;
      RECT 18465.79 1214.205 18488.86 1225.745 ;
      RECT 18465.79 1227.745 18488.86 1233.515 ;
      RECT 18465.79 1241.635 18488.86 1242.755 ;
      RECT 18465.79 1244.755 18488.86 1249.365 ;
      RECT 18465.79 1251.365 18488.86 1260.585 ;
      RECT 18465.79 1262.585 18488.86 1267.195 ;
      RECT 18465.79 1269.195 18488.86 1270.315 ;
      RECT 18465.79 1278.435 18488.86 1284.205 ;
      RECT 18465.79 1286.205 18488.86 1297.745 ;
      RECT 18465.79 1299.745 18488.86 1305.515 ;
      RECT 18465.79 1313.635 18488.86 1314.755 ;
      RECT 18465.79 1316.755 18488.86 1321.365 ;
      RECT 18465.79 1323.365 18488.86 1332.585 ;
      RECT 18465.79 1334.585 18488.86 1339.195 ;
      RECT 18465.79 1341.195 18488.86 1342.315 ;
      RECT 18465.79 1350.435 18488.86 1356.205 ;
      RECT 18465.79 1358.205 18488.86 1369.745 ;
      RECT 18465.79 1371.745 18488.86 1377.515 ;
      RECT 18465.79 1385.635 18488.86 1386.755 ;
      RECT 18465.79 1388.755 18488.86 1393.365 ;
      RECT 18465.79 1395.365 18488.86 1404.585 ;
      RECT 18465.79 1406.585 18488.86 1411.195 ;
      RECT 18465.79 1413.195 18488.86 1414.315 ;
      RECT 18465.79 1422.435 18488.86 1428.205 ;
      RECT 18465.79 1430.205 18488.86 1441.745 ;
      RECT 18465.79 1443.745 18488.86 1449.515 ;
      RECT 18465.79 1457.635 18488.86 1458.755 ;
      RECT 18465.79 1460.755 18488.86 1465.365 ;
      RECT 18465.79 1467.365 18488.86 1476.585 ;
      RECT 18465.79 1478.585 18488.86 1483.195 ;
      RECT 18465.79 1485.195 18488.86 1486.315 ;
      RECT 18465.79 1494.435 18488.86 1500.205 ;
      RECT 18465.79 1502.205 18488.86 1513.745 ;
      RECT 18465.79 1515.745 18488.86 1521.515 ;
      RECT 18465.79 1529.635 18488.86 1530.755 ;
      RECT 18465.79 1532.755 18488.86 1537.365 ;
      RECT 18465.79 1539.365 18488.86 1548.585 ;
      RECT 18465.79 1550.585 18488.86 1555.195 ;
      RECT 18465.79 1557.195 18488.86 1558.315 ;
      RECT 18465.79 1566.435 18488.86 1572.205 ;
      RECT 18465.79 1574.205 18488.86 1585.745 ;
      RECT 18465.79 1587.745 18488.86 1593.515 ;
      RECT 18465.79 1601.635 18488.86 1602.755 ;
      RECT 18465.79 1604.755 18488.86 1609.365 ;
      RECT 18465.79 1611.365 18488.86 1620.585 ;
      RECT 18465.79 1622.585 18488.86 1627.195 ;
      RECT 18465.79 1629.195 18488.86 1630.315 ;
      RECT 18465.79 1638.435 18488.86 1644.205 ;
      RECT 18465.79 1646.205 18488.86 1657.745 ;
      RECT 18465.79 1659.745 18488.86 1665.515 ;
      RECT 18465.79 1673.635 18488.86 1674.755 ;
      RECT 18465.79 1676.755 18488.86 1681.365 ;
      RECT 18465.79 1683.365 18488.86 1692.585 ;
      RECT 18465.79 1694.585 18488.86 1699.195 ;
      RECT 18465.79 1701.195 18488.86 1702.315 ;
      RECT 18465.79 1710.435 18488.86 1716.205 ;
      RECT 18465.79 1718.205 18488.86 1729.745 ;
      RECT 18465.79 1731.745 18488.86 1737.515 ;
      RECT 18465.79 1745.635 18488.86 1746.755 ;
      RECT 18465.79 1748.755 18488.86 1753.365 ;
      RECT 18465.79 1755.365 18488.86 1764.585 ;
      RECT 18465.79 1766.585 18488.86 1771.195 ;
      RECT 18465.79 1773.195 18488.86 1774.315 ;
      RECT 18465.79 1782.435 18488.86 1788.205 ;
      RECT 18465.79 1790.205 18488.86 1801.745 ;
      RECT 18465.79 1803.745 18488.86 1809.515 ;
      RECT 18465.79 1817.635 18488.86 1818.755 ;
      RECT 18465.79 1820.755 18488.86 1825.365 ;
      RECT 18465.79 1827.365 18488.86 1836.585 ;
      RECT 18465.79 1838.585 18488.86 1843.195 ;
      RECT 18465.79 1845.195 18488.86 1846.315 ;
      RECT 18465.79 1854.435 18488.86 1860.205 ;
      RECT 18465.79 1862.205 18488.86 1873.745 ;
      RECT 18465.79 1875.745 18488.86 1881.515 ;
      RECT 18465.79 1889.635 18488.86 1890.755 ;
      RECT 18465.79 1892.755 18488.86 1897.365 ;
      RECT 18465.79 1899.365 18488.86 1908.585 ;
      RECT 18465.79 1910.585 18488.86 1915.195 ;
      RECT 18465.79 1917.195 18488.86 1918.315 ;
      RECT 18465.79 1926.435 18488.86 1932.205 ;
      RECT 18465.79 1934.205 18488.86 1945.745 ;
      RECT 18465.79 1947.745 18488.86 1953.515 ;
      RECT 18465.79 1961.635 18488.86 1962.755 ;
      RECT 18465.79 1964.755 18488.86 1969.365 ;
      RECT 18465.79 1971.365 18488.86 1980.585 ;
      RECT 18465.79 1982.585 18488.86 1987.195 ;
      RECT 18465.79 1989.195 18488.86 1990.315 ;
      RECT 18465.79 1998.435 18488.86 2004.205 ;
      RECT 18465.79 2006.205 18488.86 2017.745 ;
      RECT 18465.79 2019.745 18488.86 2025.515 ;
      RECT 18465.79 2033.635 18488.86 2034.755 ;
      RECT 18465.79 2036.755 18488.86 2041.365 ;
      RECT 18465.79 2043.365 18488.86 2052.585 ;
      RECT 18465.79 2054.585 18488.86 2059.195 ;
      RECT 18465.79 2061.195 18488.86 2062.315 ;
      RECT 18465.79 2070.435 18488.86 2076.205 ;
      RECT 18465.79 2078.205 18488.86 2089.745 ;
      RECT 18465.79 2091.745 18488.86 2097.515 ;
      RECT 18465.79 2105.635 18488.86 2106.755 ;
      RECT 18465.79 2108.755 18488.86 2113.365 ;
      RECT 18465.79 2115.365 18488.86 2124.585 ;
      RECT 18465.79 2126.585 18488.86 2131.195 ;
      RECT 18465.79 2133.195 18488.86 2134.315 ;
      RECT 18465.79 2142.435 18488.86 2148.205 ;
      RECT 18465.79 2150.205 18488.86 2161.745 ;
      RECT 18465.79 2163.745 18488.86 2169.515 ;
      RECT 18465.79 2177.635 18488.86 2178.755 ;
      RECT 18465.79 2180.755 18488.86 2185.365 ;
      RECT 18465.79 2187.365 18488.86 2196.585 ;
      RECT 18465.79 2198.585 18488.86 2203.195 ;
      RECT 18465.79 2205.195 18488.86 2206.315 ;
      RECT 18465.79 2214.435 18488.86 2220.205 ;
      RECT 18465.79 2222.205 18488.86 2233.745 ;
      RECT 18465.79 2235.745 18488.86 2241.515 ;
      RECT 18465.79 2249.635 18488.86 2250.755 ;
      RECT 18465.79 2252.755 18488.86 2257.365 ;
      RECT 18465.79 2259.365 18488.86 2268.585 ;
      RECT 18465.79 2270.585 18488.86 2275.195 ;
      RECT 18465.79 2277.195 18488.86 2278.315 ;
      RECT 18465.79 2286.435 18488.86 2292.205 ;
      RECT 18465.79 2294.205 18488.86 2305.745 ;
      RECT 18465.79 2307.745 18488.86 2313.515 ;
      RECT 18465.79 2321.635 18488.86 2322.755 ;
      RECT 18465.79 2324.755 18488.86 2329.365 ;
      RECT 18465.79 2331.365 18488.86 2340.585 ;
      RECT 18465.79 2342.585 18488.86 2347.195 ;
      RECT 18465.79 2349.195 18488.86 2350.315 ;
      RECT 18465.79 2358.435 18488.86 2364.205 ;
      RECT 18465.79 2366.205 18488.86 2377.745 ;
      RECT 18465.79 2379.745 18488.86 2385.515 ;
      RECT 18465.79 2393.635 18488.86 2394.755 ;
      RECT 18465.79 2396.755 18488.86 2401.365 ;
      RECT 18465.79 2403.365 18488.86 2412.585 ;
      RECT 18465.79 2414.585 18488.86 2419.195 ;
      RECT 18465.79 2421.195 18488.86 2422.315 ;
      RECT 18465.79 2430.435 18488.86 2436.205 ;
      RECT 18465.79 2438.205 18488.86 2449.745 ;
      RECT 18465.79 2451.745 18488.86 2457.515 ;
      RECT 18465.79 2465.635 18488.86 2466.755 ;
      RECT 18465.79 2468.755 18488.86 2473.365 ;
      RECT 18465.79 2475.365 18488.86 2484.585 ;
      RECT 18465.79 2486.585 18488.86 2491.195 ;
      RECT 18465.79 2493.195 18488.86 2494.315 ;
      RECT 18465.79 2502.435 18488.86 2508.205 ;
      RECT 18465.79 2510.205 18488.86 2521.745 ;
      RECT 18465.79 2523.745 18488.86 2529.515 ;
      RECT 18465.79 2537.635 18488.86 2538.755 ;
      RECT 18465.79 2540.755 18488.86 2545.365 ;
      RECT 18465.79 2547.365 18488.86 2556.585 ;
      RECT 18465.79 2558.585 18488.86 2563.195 ;
      RECT 18465.79 2565.195 18488.86 2566.315 ;
      RECT 18465.79 2574.435 18488.86 2580.205 ;
      RECT 18465.79 2582.205 18488.86 2593.745 ;
      RECT 18465.79 2595.745 18488.86 2601.515 ;
      RECT 18465.79 2609.635 18488.86 2610.755 ;
      RECT 18465.79 2612.755 18488.86 2617.365 ;
      RECT 18465.79 2619.365 18488.86 2628.585 ;
      RECT 18465.79 2630.585 18488.86 2635.195 ;
      RECT 18465.79 2637.195 18488.86 2638.315 ;
      RECT 18465.79 2646.435 18488.86 2652.205 ;
      RECT 18465.79 2654.205 18488.86 2665.745 ;
      RECT 18465.79 2667.745 18488.86 2673.515 ;
      RECT 18465.79 2681.635 18488.86 2682.755 ;
      RECT 18465.79 2684.755 18488.86 2689.365 ;
      RECT 18465.79 2691.365 18488.86 2700.585 ;
      RECT 18465.79 2702.585 18488.86 2707.195 ;
      RECT 18465.79 2709.195 18488.86 2710.315 ;
      RECT 18465.79 2718.435 18488.86 2724.205 ;
      RECT 18465.79 2726.205 18488.86 2737.745 ;
      RECT 18465.79 2739.745 18488.86 2745.515 ;
      RECT 18465.79 2753.635 18488.86 2754.755 ;
      RECT 18465.79 2756.755 18488.86 2761.365 ;
      RECT 18465.79 2763.365 18488.86 2772.585 ;
      RECT 18465.79 2774.585 18488.86 2779.195 ;
      RECT 18465.79 2781.195 18488.86 2782.315 ;
      RECT 18465.79 2790.435 18488.86 2796.205 ;
      RECT 18465.79 2798.205 18488.86 2809.745 ;
      RECT 18465.79 2811.745 18488.86 2817.515 ;
      RECT 18465.79 2825.635 18488.86 2826.755 ;
      RECT 18465.79 2828.755 18488.86 2833.365 ;
      RECT 18465.79 2835.365 18488.86 2844.585 ;
      RECT 18465.79 2846.585 18488.86 2851.195 ;
      RECT 18465.79 2853.195 18488.86 2854.315 ;
      RECT 18465.79 2862.435 18488.86 2868.205 ;
      RECT 18465.79 2870.205 18488.86 2881.745 ;
      RECT 18465.79 2883.745 18488.86 2889.515 ;
      RECT 18465.79 2897.635 18488.86 2898.755 ;
      RECT 18465.79 2900.755 18488.86 2905.365 ;
      RECT 18465.79 2907.365 18488.86 2916.585 ;
      RECT 18465.79 2918.585 18488.86 2923.195 ;
      RECT 18465.79 2925.195 18488.86 2926.315 ;
      RECT 18465.79 2934.435 18488.86 2940.205 ;
      RECT 18465.79 2942.205 18488.86 2953.745 ;
      RECT 18465.79 2955.745 18488.86 2961.515 ;
      RECT 18465.79 2969.635 18488.86 2970.755 ;
      RECT 18465.79 2972.755 18488.86 2977.365 ;
      RECT 18465.79 2979.365 18488.86 2988.585 ;
      RECT 18465.79 2990.585 18488.86 2995.195 ;
      RECT 18465.79 2997.195 18488.86 2998.315 ;
      RECT 18465.79 3006.435 18488.86 3012.205 ;
      RECT 18465.79 3014.205 18488.86 3025.745 ;
      RECT 18465.79 3027.745 18488.86 3033.515 ;
      RECT 18465.79 3041.635 18488.86 3042.755 ;
      RECT 18465.79 3044.755 18488.86 3049.365 ;
      RECT 18465.79 3051.365 18488.86 3060.585 ;
      RECT 18465.79 3062.585 18488.86 3067.195 ;
      RECT 18465.79 3069.195 18488.86 3070.315 ;
      RECT 18465.79 3078.435 18488.86 3084.205 ;
      RECT 18465.79 3086.205 18488.86 3097.745 ;
      RECT 18465.79 3099.745 18488.86 3105.515 ;
      RECT 18465.79 3113.635 18488.86 3114.755 ;
      RECT 18465.79 3116.755 18488.86 3121.365 ;
      RECT 18465.79 3123.365 18488.86 3132.585 ;
      RECT 18465.79 3134.585 18488.86 3139.195 ;
      RECT 18465.79 3141.195 18488.86 3142.315 ;
      RECT 18465.79 3150.435 18488.86 3156.205 ;
      RECT 18465.79 3158.205 18488.86 3169.745 ;
      RECT 18465.79 3171.745 18488.86 3177.515 ;
      RECT 18465.79 3185.635 18488.86 3186.755 ;
      RECT 18465.79 3188.755 18488.86 3193.365 ;
      RECT 18465.79 3195.365 18488.86 3204.585 ;
      RECT 18465.79 3206.585 18488.86 3211.195 ;
      RECT 18465.79 3213.195 18488.86 3214.315 ;
      RECT 18465.79 3222.435 18488.86 3228.205 ;
      RECT 18465.79 3230.205 18488.86 3241.745 ;
      RECT 18465.79 3243.745 18488.86 3249.515 ;
      RECT 18465.79 3257.635 18488.86 3258.755 ;
      RECT 18465.79 3260.755 18488.86 3265.365 ;
      RECT 18465.79 3267.365 18488.86 3276.585 ;
      RECT 18465.79 3278.585 18488.86 3283.195 ;
      RECT 18465.79 3285.195 18488.86 3286.315 ;
      RECT 18465.79 3294.435 18488.86 3300.205 ;
      RECT 18465.79 3302.205 18488.86 3313.745 ;
      RECT 18465.79 3315.745 18488.86 3321.515 ;
      RECT 18465.79 3329.635 18488.86 3330.755 ;
      RECT 18465.79 3332.755 18488.86 3337.365 ;
      RECT 18465.79 3339.365 18488.86 3348.585 ;
      RECT 18465.79 3350.585 18488.86 3355.195 ;
      RECT 18465.79 3357.195 18488.86 3358.315 ;
      RECT 18465.79 3366.435 18488.86 3372.205 ;
      RECT 18465.79 3374.205 18488.86 3385.745 ;
      RECT 18465.79 3387.745 18488.86 3393.515 ;
      RECT 18465.79 3401.635 18488.86 3402.755 ;
      RECT 18465.79 3404.755 18488.86 3409.365 ;
      RECT 18465.79 3411.365 18488.86 3420.585 ;
      RECT 18465.79 3422.585 18488.86 3427.195 ;
      RECT 18465.79 3429.195 18488.86 3430.315 ;
      RECT 18465.79 3438.435 18488.86 3444.205 ;
      RECT 18465.79 3446.205 18488.86 3457.745 ;
      RECT 18465.79 3459.745 18488.86 3465.515 ;
      RECT 18465.79 3473.635 18488.86 3474.755 ;
      RECT 18465.79 3476.755 18488.86 3481.365 ;
      RECT 18465.79 3483.365 18488.86 3492.585 ;
      RECT 18465.79 3494.585 18488.86 3499.195 ;
      RECT 18465.79 3501.195 18488.86 3502.315 ;
      RECT 18465.79 3510.435 18488.86 3516.205 ;
      RECT 18465.79 3518.205 18488.86 3529.745 ;
      RECT 18465.79 3531.745 18488.86 3537.515 ;
      RECT 18465.79 3545.635 18488.86 3546.755 ;
      RECT 18465.79 3548.755 18488.86 3553.365 ;
      RECT 18465.79 3555.365 18488.86 3564.585 ;
      RECT 18465.79 3566.585 18488.86 3571.195 ;
      RECT 18465.79 3573.195 18488.86 3574.315 ;
      RECT 18465.79 3582.435 18488.86 3588.205 ;
      RECT 18465.79 3590.205 18488.86 3601.745 ;
      RECT 18465.79 3603.745 18488.86 3609.515 ;
      RECT 18465.79 3617.635 18488.86 3618.755 ;
      RECT 18465.79 3620.755 18488.86 3625.365 ;
      RECT 18465.79 3627.365 18488.86 3636.585 ;
      RECT 18465.79 3638.585 18488.86 3643.195 ;
      RECT 18465.79 3645.195 18488.86 3646.315 ;
      RECT 18465.79 3654.435 18488.86 3660.205 ;
      RECT 18465.79 3662.205 18488.86 3673.745 ;
      RECT 18465.79 3675.745 18488.86 3681.515 ;
      RECT 18465.79 3689.635 18488.86 3690.755 ;
      RECT 18465.79 3692.755 18488.86 3697.365 ;
      RECT 18465.79 3699.365 18488.86 3708.585 ;
      RECT 18465.79 3710.585 18488.86 3715.195 ;
      RECT 18465.79 3717.195 18488.86 3718.315 ;
      RECT 18465.79 3726.435 18488.86 3732.205 ;
      RECT 18465.79 3734.205 18488.86 3745.745 ;
      RECT 18465.79 3747.745 18488.86 3753.515 ;
      RECT 18465.79 3761.635 18488.86 3762.755 ;
      RECT 18465.79 3764.755 18488.86 3769.365 ;
      RECT 18465.79 3771.365 18488.86 3780.585 ;
      RECT 18465.79 3782.585 18488.86 3787.195 ;
      RECT 18465.79 3789.195 18488.86 3790.315 ;
      RECT 18465.79 3798.435 18488.86 3804.205 ;
      RECT 18465.79 3806.205 18488.86 3817.745 ;
      RECT 18465.79 3819.745 18488.86 3825.515 ;
      RECT 18465.79 3833.635 18488.86 3834.755 ;
      RECT 18465.79 3836.755 18488.86 3841.365 ;
      RECT 18465.79 3843.365 18488.86 3852.585 ;
      RECT 18465.79 3854.585 18488.86 3859.195 ;
      RECT 18465.79 3861.195 18488.86 3862.315 ;
      RECT 18465.79 3870.435 18488.86 3876.205 ;
      RECT 18465.79 3878.205 18488.86 3889.745 ;
      RECT 18465.79 3891.745 18488.86 3897.515 ;
      RECT 18465.79 3905.635 18488.86 3906.755 ;
      RECT 18465.79 3908.755 18488.86 3913.365 ;
      RECT 18465.79 3915.365 18488.86 3924.585 ;
      RECT 18465.79 3926.585 18488.86 3931.195 ;
      RECT 18465.79 3933.195 18488.86 3934.315 ;
      RECT 18465.79 3942.435 18488.86 3948.205 ;
      RECT 18465.79 3950.205 18488.86 3961.745 ;
      RECT 18465.79 3963.745 18488.86 3969.515 ;
      RECT 18465.79 3977.635 18488.86 3978.755 ;
      RECT 18465.79 3980.755 18488.86 3985.365 ;
      RECT 18465.79 3987.365 18488.86 3996.585 ;
      RECT 18465.79 3998.585 18488.86 4003.195 ;
      RECT 18465.79 4005.195 18488.86 4006.315 ;
      RECT 18465.79 4014.435 18488.86 4020.205 ;
      RECT 18465.79 4022.205 18488.86 4033.745 ;
      RECT 18465.79 4035.745 18488.86 4041.515 ;
      RECT 18465.79 4049.635 18488.86 4050.755 ;
      RECT 18465.79 4052.755 18488.86 4057.365 ;
      RECT 18465.79 4059.365 18488.86 4068.585 ;
      RECT 18465.79 4070.585 18488.86 4075.195 ;
      RECT 18465.79 4077.195 18488.86 4078.315 ;
      RECT 18465.79 4086.435 18488.86 4092.205 ;
      RECT 18465.79 4094.205 18488.86 4105.745 ;
      RECT 18465.79 4107.745 18488.86 4113.515 ;
      RECT 18465.79 4121.635 18488.86 4122.755 ;
      RECT 18465.79 4124.755 18488.86 4129.365 ;
      RECT 18465.79 4131.365 18488.86 4140.585 ;
      RECT 18465.79 4142.585 18488.86 4147.195 ;
      RECT 18465.79 4149.195 18488.86 4150.315 ;
      RECT 18465.79 4158.435 18488.86 4164.205 ;
      RECT 18465.79 4166.205 18488.86 4177.745 ;
      RECT 18465.79 4179.745 18488.86 4185.515 ;
      RECT 18465.79 4193.635 18488.86 4194.755 ;
      RECT 18465.79 4196.755 18488.86 4201.365 ;
      RECT 18465.79 4203.365 18488.86 4212.585 ;
      RECT 18465.79 4214.585 18488.86 4219.195 ;
      RECT 18465.79 4221.195 18488.86 4222.315 ;
      RECT 18465.79 4230.435 18488.86 4236.205 ;
      RECT 18465.79 4238.205 18488.86 4249.745 ;
      RECT 18465.79 4251.745 18488.86 4257.515 ;
      RECT 18465.79 4265.635 18488.86 4266.755 ;
      RECT 18465.79 4268.755 18488.86 4273.365 ;
      RECT 18465.79 4275.365 18488.86 4284.585 ;
      RECT 18465.79 4286.585 18488.86 4291.195 ;
      RECT 18465.79 4293.195 18488.86 4294.315 ;
      RECT 18465.79 4302.435 18488.86 4308.205 ;
      RECT 18465.79 4310.205 18488.86 4321.745 ;
      RECT 18465.79 4323.745 18488.86 4329.515 ;
      RECT 18465.79 4337.635 18488.86 4338.755 ;
      RECT 18465.79 4340.755 18488.86 4345.365 ;
      RECT 18465.79 4347.365 18488.86 4356.585 ;
      RECT 18465.79 4358.585 18488.86 4363.195 ;
      RECT 18465.79 4365.195 18488.86 4366.315 ;
      RECT 18465.79 4374.435 18488.86 4380.205 ;
      RECT 18465.79 4382.205 18488.86 4393.745 ;
      RECT 18465.79 4395.745 18488.86 4401.515 ;
      RECT 18465.79 4409.635 18488.86 4410.755 ;
      RECT 18465.79 4412.755 18488.86 4417.365 ;
      RECT 18465.79 4419.365 18488.86 4428.585 ;
      RECT 18465.79 4430.585 18488.86 4435.195 ;
      RECT 18465.79 4437.195 18488.86 4438.315 ;
      RECT 18465.79 4446.435 18488.86 4452.205 ;
      RECT 18465.79 4454.205 18488.86 4465.745 ;
      RECT 18465.79 4467.745 18488.86 4473.515 ;
      RECT 18465.79 4481.635 18488.86 4482.755 ;
      RECT 18465.79 4484.755 18488.86 4489.365 ;
      RECT 18465.79 4491.365 18488.86 4500.585 ;
      RECT 18465.79 4502.585 18488.86 4507.195 ;
      RECT 18465.79 4509.195 18488.86 4510.315 ;
      RECT 18465.79 4518.435 18488.86 4524.205 ;
      RECT 18465.79 4526.205 18488.86 4537.745 ;
      RECT 18465.79 4539.745 18488.86 4545.515 ;
      RECT 18465.79 4553.635 18488.86 4554.755 ;
      RECT 18465.79 4556.755 18488.86 4561.365 ;
      RECT 18465.79 4563.365 18488.86 4572.585 ;
      RECT 18465.79 4574.585 18488.86 4579.195 ;
      RECT 18465.79 4581.195 18488.86 4582.315 ;
      RECT 18465.79 4590.435 18488.86 4596.205 ;
      RECT 18465.79 4598.205 18488.86 4609.745 ;
      RECT 18465.79 4611.745 18488.86 4617.515 ;
      RECT 18465.79 4625.635 18488.86 4626.755 ;
      RECT 18465.79 4628.755 18488.86 4633.365 ;
      RECT 18465.79 4635.365 18488.86 4644.585 ;
      RECT 18465.79 4646.585 18488.86 4651.195 ;
      RECT 18465.79 4653.195 18488.86 4654.315 ;
      RECT 18465.79 4662.435 18488.86 4668.205 ;
      RECT 18465.79 4670.205 18488.86 4681.745 ;
      RECT 18465.79 4683.745 18488.86 4689.515 ;
      RECT 18465.79 4697.635 18488.86 4698.755 ;
      RECT 18465.79 4700.755 18488.86 4705.365 ;
      RECT 18465.79 4707.365 18488.86 4716.585 ;
      RECT 18465.79 4718.585 18488.86 4723.195 ;
      RECT 18465.79 4725.195 18488.86 4726.315 ;
      RECT 18465.79 4734.435 18488.86 4740.205 ;
      RECT 18465.79 4742.205 18488.86 4753.745 ;
      RECT 18465.79 4755.745 18488.86 4761.515 ;
      RECT 18465.79 4769.635 18488.86 4770.755 ;
      RECT 18465.79 4772.755 18488.86 4777.365 ;
      RECT 18465.79 4779.365 18488.86 4788.585 ;
      RECT 18465.79 4790.585 18488.86 4795.195 ;
      RECT 18465.79 4797.195 18488.86 4798.315 ;
      RECT 18465.79 4806.435 18488.86 4812.205 ;
      RECT 18465.79 4814.205 18488.86 4825.745 ;
      RECT 18465.79 4827.745 18488.86 4833.515 ;
      RECT 18465.79 4841.635 18488.86 4842.755 ;
      RECT 18465.79 4844.755 18488.86 4849.365 ;
      RECT 18465.79 4851.365 18488.86 4860.585 ;
      RECT 18465.79 4862.585 18488.86 4867.195 ;
      RECT 18465.79 4869.195 18488.86 4870.315 ;
      RECT 18465.79 4878.435 18488.86 4884.205 ;
      RECT 18465.79 4886.205 18488.86 4897.745 ;
      RECT 18465.79 4899.745 18488.86 4905.515 ;
      RECT 18465.79 4913.635 18488.86 4914.755 ;
      RECT 18465.79 4916.755 18488.86 4921.365 ;
      RECT 18465.79 4923.365 18488.86 4932.585 ;
      RECT 18465.79 4934.585 18488.86 4939.195 ;
      RECT 18465.79 4941.195 18488.86 4942.315 ;
      RECT 18465.79 4950.435 18488.86 4956.205 ;
      RECT 18465.79 4958.205 18488.86 4969.745 ;
      RECT 18465.79 4971.745 18488.86 4977.515 ;
      RECT 18465.79 4985.635 18488.86 4986.755 ;
      RECT 18465.79 4988.755 18488.86 4993.365 ;
      RECT 18465.79 4995.365 18488.86 5004.585 ;
      RECT 18465.79 5006.585 18488.86 5011.195 ;
      RECT 18465.79 5013.195 18488.86 5014.315 ;
      RECT 18465.79 5022.435 18488.86 5028.205 ;
      RECT 18465.79 5030.205 18488.86 5041.745 ;
      RECT 18465.79 5043.745 18488.86 5049.515 ;
      RECT 18465.79 5057.635 18488.86 5058.755 ;
      RECT 18465.79 5060.755 18488.86 5065.365 ;
      RECT 18465.79 5067.365 18488.86 5076.585 ;
      RECT 18465.79 5078.585 18488.86 5083.195 ;
      RECT 18465.79 5085.195 18488.86 5086.315 ;
      RECT 18465.79 5094.435 18488.86 5100.205 ;
      RECT 18465.79 5102.205 18488.86 5113.745 ;
      RECT 18465.79 5115.745 18488.86 5121.515 ;
      RECT 18465.79 5129.635 18488.86 5130.755 ;
      RECT 18465.79 5132.755 18488.86 5137.365 ;
      RECT 18465.79 5139.365 18488.86 5148.585 ;
      RECT 18465.79 5150.585 18488.86 5155.195 ;
      RECT 18465.79 5157.195 18488.86 5158.315 ;
      RECT 18465.79 5166.435 18488.86 5172.205 ;
      RECT 18465.79 5174.205 18488.86 5185.745 ;
      RECT 18465.79 5187.745 18488.86 5193.515 ;
      RECT 18465.79 5201.635 18488.86 5202.755 ;
      RECT 18465.79 5204.755 18488.86 5209.365 ;
      RECT 18465.79 5211.365 18488.86 5220.585 ;
      RECT 18465.79 5222.585 18488.86 5227.195 ;
      RECT 18465.79 5229.195 18488.86 5230.315 ;
      RECT 18465.79 5238.435 18488.86 5244.205 ;
      RECT 18465.79 5246.205 18488.86 5257.745 ;
      RECT 18465.79 5259.745 18488.86 5265.515 ;
      RECT 18465.79 5273.635 18488.86 5274.755 ;
      RECT 18465.79 5276.755 18488.86 5281.365 ;
      RECT 18465.79 5283.365 18488.86 5292.585 ;
      RECT 18465.79 5294.585 18488.86 5299.195 ;
      RECT 18465.79 5301.195 18488.86 5302.315 ;
      RECT 18465.79 5310.435 18488.86 5316.205 ;
      RECT 18465.79 5318.205 18488.86 5329.745 ;
      RECT 18465.79 5331.745 18488.86 5337.515 ;
      RECT 18465.79 5345.635 18488.86 5346.755 ;
      RECT 18465.79 5348.755 18488.86 5353.365 ;
      RECT 18465.79 5355.365 18488.86 5364.585 ;
      RECT 18465.79 5366.585 18488.86 5371.195 ;
      RECT 18465.79 5373.195 18488.86 5374.315 ;
      RECT 18465.79 5382.435 18488.86 5388.205 ;
      RECT 18465.79 5390.205 18488.86 5401.745 ;
      RECT 18465.79 5403.745 18488.86 5409.515 ;
      RECT 18465.79 5417.635 18488.86 5418.755 ;
      RECT 18465.79 5420.755 18488.86 5425.365 ;
      RECT 18465.79 5427.365 18488.86 5436.585 ;
      RECT 18465.79 5438.585 18488.86 5443.195 ;
      RECT 18465.79 5445.195 18488.86 5446.315 ;
      RECT 18465.79 5454.435 18488.86 5460.205 ;
      RECT 18465.79 5462.205 18488.86 5473.745 ;
      RECT 18465.79 5475.745 18488.86 5481.515 ;
      RECT 18465.79 5489.635 18488.86 5490.755 ;
      RECT 18465.79 5492.755 18488.86 5497.365 ;
      RECT 18465.79 5499.365 18488.86 5508.585 ;
      RECT 18465.79 5510.585 18488.86 5515.195 ;
      RECT 18465.79 5517.195 18488.86 5518.315 ;
      RECT 18465.79 5526.435 18488.86 5532.205 ;
      RECT 18465.79 5534.205 18488.86 5545.745 ;
      RECT 18465.79 5547.745 18488.86 5553.515 ;
      RECT 18465.79 5561.635 18488.86 5562.755 ;
      RECT 18465.79 5564.755 18488.86 5569.365 ;
      RECT 18465.79 5571.365 18488.86 5580.585 ;
      RECT 18465.79 5582.585 18488.86 5587.195 ;
      RECT 18465.79 5589.195 18488.86 5590.315 ;
      RECT 18465.79 5598.435 18488.86 5604.205 ;
      RECT 18465.79 5606.205 18488.86 5617.745 ;
      RECT 18465.79 5619.745 18488.86 5625.515 ;
      RECT 18465.79 5633.635 18488.86 5634.755 ;
      RECT 18465.79 5636.755 18488.86 5641.365 ;
      RECT 18465.79 5643.365 18488.86 5652.585 ;
      RECT 18465.79 5654.585 18488.86 5659.195 ;
      RECT 18465.79 5661.195 18488.86 5662.315 ;
      RECT 18465.79 5670.435 18488.86 5676.205 ;
      RECT 18465.79 5678.205 18488.86 5689.745 ;
      RECT 18465.79 5691.745 18488.86 5697.515 ;
      RECT 18465.79 5705.635 18488.86 5706.755 ;
      RECT 18465.79 5708.755 18488.86 5713.365 ;
      RECT 18465.79 5715.365 18488.86 5724.585 ;
      RECT 18465.79 5726.585 18488.86 5731.195 ;
      RECT 18465.79 5733.195 18488.86 5734.315 ;
      RECT 18465.79 5742.435 18488.86 5748.205 ;
      RECT 18465.79 5750.205 18488.86 5761.745 ;
      RECT 18465.79 5763.745 18488.86 5769.515 ;
      RECT 18465.79 5777.635 18488.86 5778.755 ;
      RECT 18465.79 5780.755 18488.86 5785.365 ;
      RECT 18465.79 5787.365 18488.86 5796.585 ;
      RECT 18465.79 5798.585 18488.86 5803.195 ;
      RECT 18465.79 5805.195 18488.86 5806.315 ;
      RECT 18465.79 5814.435 18488.86 5820.205 ;
      RECT 18465.79 5822.205 18488.86 5833.745 ;
      RECT 18465.79 5835.745 18488.86 5841.515 ;
      RECT 18465.79 5849.635 18488.86 5850.755 ;
      RECT 18465.79 5852.755 18488.86 5857.365 ;
      RECT 18465.79 5859.365 18488.86 5868.585 ;
      RECT 18465.79 5870.585 18488.86 5875.195 ;
      RECT 18465.79 5877.195 18488.86 5878.315 ;
      RECT 18465.79 5886.435 18488.86 5892.205 ;
      RECT 18465.79 5894.205 18488.86 5905.745 ;
      RECT 18465.79 5907.745 18488.86 5913.515 ;
      RECT 18465.79 5921.635 18488.86 5922.755 ;
      RECT 18465.79 5924.755 18488.86 5929.365 ;
      RECT 18465.79 5931.365 18488.86 5940.585 ;
      RECT 18465.79 5942.585 18488.86 5947.195 ;
      RECT 18465.79 5949.195 18488.86 5950.315 ;
      RECT 18465.79 5958.435 18488.86 5964.205 ;
      RECT 18465.79 5966.205 18488.86 5977.745 ;
      RECT 18465.79 5979.745 18488.86 5985.515 ;
      RECT 18465.79 5993.635 18488.86 5994.755 ;
      RECT 18465.79 5996.755 18488.86 6001.365 ;
      RECT 18465.79 6003.365 18488.86 6012.585 ;
      RECT 18465.79 6014.585 18488.86 6019.195 ;
      RECT 18465.79 6021.195 18488.86 6022.315 ;
      RECT 18465.79 6030.435 18488.86 6036.205 ;
      RECT 18465.79 6038.205 18488.86 6049.745 ;
      RECT 18465.79 6051.745 18488.86 6057.515 ;
      RECT 18465.79 6065.635 18488.86 6066.755 ;
      RECT 18465.79 6068.755 18488.86 6073.365 ;
      RECT 18465.79 6075.365 18488.86 6084.585 ;
      RECT 18465.79 6086.585 18488.86 6091.195 ;
      RECT 18465.79 6093.195 18488.86 6094.315 ;
      RECT 18465.79 6102.435 18488.86 6108.205 ;
      RECT 18465.79 6110.205 18488.86 6121.745 ;
      RECT 18465.79 6123.745 18488.86 6129.515 ;
      RECT 18465.79 6137.635 18488.86 6138.755 ;
      RECT 18465.79 6140.755 18488.86 6145.365 ;
      RECT 18465.79 6147.365 18488.86 6156.585 ;
      RECT 18465.79 6158.585 18488.86 6163.195 ;
      RECT 18465.79 6165.195 18488.86 6166.315 ;
      RECT 18465.79 6174.435 18488.86 6180.205 ;
      RECT 18465.79 6182.205 18488.86 6193.745 ;
      RECT 18465.79 6195.745 18488.86 6201.515 ;
      RECT 18465.79 6209.635 18488.86 6210.755 ;
      RECT 18465.79 6212.755 18488.86 6217.365 ;
      RECT 18465.79 6219.365 18488.86 6228.585 ;
      RECT 18465.79 6230.585 18488.86 6235.195 ;
      RECT 18465.79 6237.195 18488.86 6238.315 ;
      RECT 18465.79 6246.435 18488.86 6252.205 ;
      RECT 18465.79 6254.205 18488.86 6265.745 ;
      RECT 18465.79 6267.745 18488.86 6273.515 ;
      RECT 18465.79 6281.635 18488.86 6282.755 ;
      RECT 18465.79 6284.755 18488.86 6289.365 ;
      RECT 18465.79 6291.365 18488.86 6300.585 ;
      RECT 18465.79 6302.585 18488.86 6307.195 ;
      RECT 18465.79 6309.195 18488.86 6310.315 ;
      RECT 18465.79 6318.435 18488.86 6324.205 ;
      RECT 18465.79 6326.205 18488.86 6337.745 ;
      RECT 18465.79 6339.745 18488.86 6345.515 ;
      RECT 18465.79 6353.635 18488.86 6354.755 ;
      RECT 18465.79 6356.755 18488.86 6361.365 ;
      RECT 18465.79 6363.365 18488.86 6372.585 ;
      RECT 18465.79 6374.585 18488.86 6379.195 ;
      RECT 18465.79 6381.195 18488.86 6382.315 ;
      RECT 18465.79 6390.435 18488.86 6396.205 ;
      RECT 18465.79 6398.205 18488.86 6409.745 ;
      RECT 18465.79 6411.745 18488.86 6417.515 ;
      RECT 18465.79 6425.635 18488.86 6426.755 ;
      RECT 18465.79 6428.755 18488.86 6433.365 ;
      RECT 18465.79 6435.365 18488.86 6444.585 ;
      RECT 18465.79 6446.585 18488.86 6451.195 ;
      RECT 18465.79 6453.195 18488.86 6454.315 ;
      RECT 18465.79 6462.435 18488.86 6468.205 ;
      RECT 18465.79 6470.205 18488.86 6481.745 ;
      RECT 18465.79 6483.745 18488.86 6489.515 ;
      RECT 18465.79 6497.635 18488.86 6498.755 ;
      RECT 18465.79 6500.755 18488.86 6505.365 ;
      RECT 18465.79 6507.365 18488.86 6516.585 ;
      RECT 18465.79 6518.585 18488.86 6523.195 ;
      RECT 18465.79 6525.195 18488.86 6526.315 ;
      RECT 18465.79 6534.435 18488.86 6540.205 ;
      RECT 18465.79 6542.205 18488.86 6553.745 ;
      RECT 18465.79 6555.745 18488.86 6561.515 ;
      RECT 18465.79 6569.635 18488.86 6570.755 ;
      RECT 18465.79 6572.755 18488.86 6577.365 ;
      RECT 18465.79 6579.365 18488.86 6588.585 ;
      RECT 18465.79 6590.585 18488.86 6595.195 ;
      RECT 18465.79 6597.195 18488.86 6598.315 ;
      RECT 18465.79 6606.435 18488.86 6612.205 ;
      RECT 18465.79 6614.205 18488.86 6625.745 ;
      RECT 18465.79 6627.745 18488.86 6633.515 ;
      RECT 18465.79 6641.635 18488.86 6642.755 ;
      RECT 18465.79 6644.755 18488.86 6649.365 ;
      RECT 18465.79 6651.365 18488.86 6660.585 ;
      RECT 18465.79 6662.585 18488.86 6667.195 ;
      RECT 18465.79 6669.195 18488.86 6670.315 ;
      RECT 18465.79 6678.435 18488.86 6684.205 ;
      RECT 18465.79 6686.205 18488.86 6697.745 ;
      RECT 18465.79 6699.745 18488.86 6705.515 ;
      RECT 18465.79 6713.635 18488.86 6714.755 ;
      RECT 18465.79 6716.755 18488.86 6721.365 ;
      RECT 18465.79 6723.365 18488.86 6732.585 ;
      RECT 18465.79 6734.585 18488.86 6739.195 ;
      RECT 18465.79 6741.195 18488.86 6742.315 ;
      RECT 18465.79 6750.435 18488.86 6756.205 ;
      RECT 18465.79 6758.205 18488.86 6769.745 ;
      RECT 18465.79 6771.745 18488.86 6777.515 ;
      RECT 18465.79 6785.635 18488.86 6786.755 ;
      RECT 18465.79 6788.755 18488.86 6793.365 ;
      RECT 18465.79 6795.365 18488.86 6804.585 ;
      RECT 18465.79 6806.585 18488.86 6811.195 ;
      RECT 18465.79 6813.195 18488.86 6814.315 ;
      RECT 18465.79 6822.435 18488.86 6828.205 ;
      RECT 18465.79 6830.205 18488.86 6841.745 ;
      RECT 18465.79 6843.745 18488.86 6849.515 ;
      RECT 18465.79 6857.635 18488.86 6858.755 ;
      RECT 18465.79 6860.755 18488.86 6865.365 ;
      RECT 18465.79 6867.365 18488.86 6876.585 ;
      RECT 18465.79 6878.585 18488.86 6883.195 ;
      RECT 18465.79 6885.195 18488.86 6886.315 ;
      RECT 18465.79 6894.435 18488.86 6900.205 ;
      RECT 18465.79 6902.205 18488.86 6913.745 ;
      RECT 18465.79 6915.745 18488.86 6921.515 ;
      RECT 18465.79 6929.635 18488.86 6930.755 ;
      RECT 18465.79 6932.755 18488.86 6937.365 ;
      RECT 18465.79 6939.365 18488.86 6948.585 ;
      RECT 18465.79 6950.585 18488.86 6955.195 ;
      RECT 18465.79 6957.195 18488.86 6958.315 ;
      RECT 18465.79 6966.435 18488.86 6972.205 ;
      RECT 18465.79 6974.205 18488.86 6985.745 ;
      RECT 18465.79 6987.745 18488.86 6993.515 ;
      RECT 18465.79 7001.635 18488.86 7002.755 ;
      RECT 18465.79 7004.755 18488.86 7009.365 ;
      RECT 18465.79 7011.365 18488.86 7020.585 ;
      RECT 18465.79 7022.585 18488.86 7027.195 ;
      RECT 18465.79 7029.195 18488.86 7030.315 ;
      RECT 18465.79 7038.435 18488.86 7044.205 ;
      RECT 18465.79 7046.205 18488.86 7057.745 ;
      RECT 18465.79 7059.745 18488.86 7065.515 ;
      RECT 18465.79 7073.635 18488.86 7074.755 ;
      RECT 18465.79 7076.755 18488.86 7081.365 ;
      RECT 18465.79 7083.365 18488.86 7092.585 ;
      RECT 18465.79 7094.585 18488.86 7099.195 ;
      RECT 18465.79 7101.195 18488.86 7102.315 ;
      RECT 18465.79 7110.435 18488.86 7116.205 ;
      RECT 18465.79 7118.205 18488.86 7129.745 ;
      RECT 18465.79 7131.745 18488.86 7137.515 ;
      RECT 18465.79 7145.635 18488.86 7146.755 ;
      RECT 18465.79 7148.755 18488.86 7153.365 ;
      RECT 18465.79 7155.365 18488.86 7164.585 ;
      RECT 18465.79 7166.585 18488.86 7171.195 ;
      RECT 18465.79 7173.195 18488.86 7174.315 ;
      RECT 18465.79 7182.435 18488.86 7188.205 ;
      RECT 18465.79 7190.205 18488.86 7201.745 ;
      RECT 18465.79 7203.745 18488.86 7209.515 ;
      RECT 18465.79 7217.635 18488.86 7218.755 ;
      RECT 18465.79 7220.755 18488.86 7225.365 ;
      RECT 18465.79 7227.365 18488.86 7236.585 ;
      RECT 18465.79 7238.585 18488.86 7243.195 ;
      RECT 18465.79 7245.195 18488.86 7246.315 ;
      RECT 18465.79 7254.435 18488.86 7260.205 ;
      RECT 18465.79 7262.205 18488.86 7273.745 ;
      RECT 18465.79 7275.745 18488.86 7281.515 ;
      RECT 18465.79 7289.635 18488.86 7290.755 ;
      RECT 18465.79 7292.755 18488.86 7297.365 ;
      RECT 18465.79 7299.365 18488.86 7308.585 ;
      RECT 18465.79 7310.585 18488.86 7315.195 ;
      RECT 18465.79 7317.195 18488.86 7318.315 ;
      RECT 18465.79 7326.435 18488.86 7332.205 ;
      RECT 18465.79 7334.205 18488.86 7345.745 ;
      RECT 18465.79 7347.745 18488.86 7353.515 ;
      RECT 18465.79 7361.635 18488.86 7362.755 ;
      RECT 18465.79 7364.755 18488.86 7369.365 ;
      RECT 18465.79 7371.365 18488.86 7380.585 ;
      RECT 18465.79 7382.585 18488.86 7387.195 ;
      RECT 18465.79 7389.195 18488.86 7390.315 ;
      RECT 18465.79 7398.435 18488.86 7404.205 ;
      RECT 18465.79 7406.205 18488.86 7417.745 ;
      RECT 18465.79 7419.745 18488.86 7425.515 ;
      RECT 18465.79 7433.635 18488.86 7434.755 ;
      RECT 18465.79 7436.755 18488.86 7441.365 ;
      RECT 18465.79 7443.365 18488.86 7452.585 ;
      RECT 18465.79 7454.585 18488.86 7459.195 ;
      RECT 18465.79 7461.195 18488.86 7462.315 ;
      RECT 18465.79 7470.435 18488.86 7476.205 ;
      RECT 18465.79 7478.205 18488.86 7489.745 ;
      RECT 18465.79 7491.745 18488.86 7497.515 ;
      RECT 18465.79 7505.635 18488.86 7506.755 ;
      RECT 18465.79 7508.755 18488.86 7513.365 ;
      RECT 18465.79 7515.365 18488.86 7524.585 ;
      RECT 18465.79 7526.585 18488.86 7531.195 ;
      RECT 18465.79 7533.195 18488.86 7534.315 ;
      RECT 18465.79 7542.435 18488.86 7548.205 ;
      RECT 18465.79 7550.205 18488.86 7561.745 ;
      RECT 18465.79 7563.745 18488.86 7569.515 ;
      RECT 18465.79 7577.635 18488.86 7578.755 ;
      RECT 18465.79 7580.755 18488.86 7585.365 ;
      RECT 18465.79 7587.365 18488.86 7596.585 ;
      RECT 18465.79 7598.585 18488.86 7603.195 ;
      RECT 18465.79 7605.195 18488.86 7606.315 ;
      RECT 18465.79 7614.435 18488.86 7620.205 ;
      RECT 18465.79 7622.205 18488.86 7633.745 ;
      RECT 18465.79 7635.745 18488.86 7641.515 ;
      RECT 18465.79 7649.635 18488.86 7650.755 ;
      RECT 18465.79 7652.755 18488.86 7657.365 ;
      RECT 18465.79 7659.365 18488.86 7668.585 ;
      RECT 18465.79 7670.585 18488.86 7675.195 ;
      RECT 18465.79 7677.195 18488.86 7678.315 ;
      RECT 18465.79 7686.435 18488.86 7692.205 ;
      RECT 18465.79 7694.205 18488.86 7705.745 ;
      RECT 18465.79 7707.745 18488.86 7713.515 ;
      RECT 18465.79 7721.635 18488.86 7722.755 ;
      RECT 18465.79 7724.755 18488.86 7729.365 ;
      RECT 18465.79 7731.365 18488.86 7740.585 ;
      RECT 18465.79 7742.585 18488.86 7747.195 ;
      RECT 18465.79 7749.195 18488.86 7750.315 ;
      RECT 18465.79 7758.435 18488.86 7764.205 ;
      RECT 18465.79 7766.205 18488.86 7777.745 ;
      RECT 18465.79 7779.745 18488.86 7785.515 ;
      RECT 18465.79 7793.635 18488.86 7794.755 ;
      RECT 18465.79 7796.755 18488.86 7801.365 ;
      RECT 18465.79 7803.365 18488.86 7812.585 ;
      RECT 18465.79 7814.585 18488.86 7819.195 ;
      RECT 18465.79 7821.195 18488.86 7822.315 ;
      RECT 18465.79 7830.435 18488.86 7836.205 ;
      RECT 18465.79 7838.205 18488.86 7849.745 ;
      RECT 18465.79 7851.745 18488.86 7857.515 ;
      RECT 18465.79 7865.635 18488.86 7866.755 ;
      RECT 18465.79 7868.755 18488.86 7873.365 ;
      RECT 18465.79 7875.365 18488.86 7884.585 ;
      RECT 18465.79 7886.585 18488.86 7891.195 ;
      RECT 18465.79 7893.195 18488.86 7894.315 ;
      RECT 18465.79 7902.435 18488.86 7908.205 ;
      RECT 18465.79 7910.205 18488.86 7921.745 ;
      RECT 18465.79 7923.745 18488.86 7929.515 ;
      RECT 18465.79 7937.635 18488.86 7938.755 ;
      RECT 18465.79 7940.755 18488.86 7945.365 ;
      RECT 18465.79 7947.365 18488.86 7956.585 ;
      RECT 18465.79 7958.585 18488.86 7963.195 ;
      RECT 18465.79 7965.195 18488.86 7966.315 ;
      RECT 18465.79 7974.435 18488.86 7980.205 ;
      RECT 18465.79 7982.205 18488.86 7993.745 ;
      RECT 18465.79 7995.745 18488.86 8001.515 ;
      RECT 18465.79 8009.635 18488.86 8010.755 ;
      RECT 18465.79 8012.755 18488.86 8017.365 ;
      RECT 18465.79 8019.365 18488.86 8028.585 ;
      RECT 18465.79 8030.585 18488.86 8035.195 ;
      RECT 18465.79 8037.195 18488.86 8038.315 ;
      RECT 18465.79 8046.435 18488.86 8052.205 ;
      RECT 18465.79 8054.205 18488.86 8065.745 ;
      RECT 18465.79 8067.745 18488.86 8073.515 ;
      RECT 18465.79 8081.635 18488.86 8082.755 ;
      RECT 18465.79 8084.755 18488.86 8089.365 ;
      RECT 18465.79 8091.365 18488.86 8100.585 ;
      RECT 18465.79 8102.585 18488.86 8107.195 ;
      RECT 18465.79 8109.195 18488.86 8110.315 ;
      RECT 18465.79 8118.435 18488.86 8124.205 ;
      RECT 18465.79 8126.205 18488.86 8137.745 ;
      RECT 18465.79 8139.745 18488.86 8145.515 ;
      RECT 18465.79 8153.635 18488.86 8154.755 ;
      RECT 18465.79 8156.755 18488.86 8161.365 ;
      RECT 18465.79 8163.365 18488.86 8172.585 ;
      RECT 18465.79 8174.585 18488.86 8179.195 ;
      RECT 18465.79 8181.195 18488.86 8182.315 ;
      RECT 18465.79 8190.435 18488.86 8196.205 ;
      RECT 18465.79 8198.205 18488.86 8209.745 ;
      RECT 18465.79 8211.745 18488.86 8217.515 ;
      RECT 18465.79 8225.635 18488.86 8226.755 ;
      RECT 18465.79 8228.755 18488.86 8233.365 ;
      RECT 18465.79 8235.365 18488.86 8244.585 ;
      RECT 18465.79 8246.585 18488.86 8251.195 ;
      RECT 18465.79 8253.195 18488.86 8254.315 ;
      RECT 18465.79 8262.435 18488.86 8268.205 ;
      RECT 18465.79 8270.205 18488.86 8281.745 ;
      RECT 18465.79 8283.745 18488.86 8289.515 ;
      RECT 18465.79 8297.635 18488.86 8298.755 ;
      RECT 18465.79 8300.755 18488.86 8305.365 ;
      RECT 18465.79 8307.365 18488.86 8316.585 ;
      RECT 18465.79 8318.585 18488.86 8323.195 ;
      RECT 18465.79 8325.195 18488.86 8326.315 ;
      RECT 18465.79 8334.435 18488.86 8340.205 ;
      RECT 18465.79 8342.205 18488.86 8353.745 ;
      RECT 18465.79 8355.745 18488.86 8361.515 ;
      RECT 18465.79 8369.635 18488.86 8370.755 ;
      RECT 18465.79 8372.755 18488.86 8377.365 ;
      RECT 18465.79 8379.365 18488.86 8388.585 ;
      RECT 18465.79 8390.585 18488.86 8395.195 ;
      RECT 18465.79 8397.195 18488.86 8398.315 ;
      RECT 18465.79 8406.435 18488.86 8412.205 ;
      RECT 18465.79 8414.205 18488.86 8425.745 ;
      RECT 18465.79 8427.745 18488.86 8433.515 ;
      RECT 18465.79 8441.635 18488.86 8442.755 ;
      RECT 18465.79 8444.755 18488.86 8449.365 ;
      RECT 18465.79 8451.365 18488.86 8460.585 ;
      RECT 18465.79 8462.585 18488.86 8467.195 ;
      RECT 18465.79 8469.195 18488.86 8470.315 ;
      RECT 18465.79 8478.435 18488.86 8484.205 ;
      RECT 18465.79 8486.205 18488.86 8497.745 ;
      RECT 18465.79 8499.745 18488.86 8505.515 ;
      RECT 18465.79 8513.635 18488.86 8514.755 ;
      RECT 18465.79 8516.755 18488.86 8521.365 ;
      RECT 18465.79 8523.365 18488.86 8532.585 ;
      RECT 18465.79 8534.585 18488.86 8539.195 ;
      RECT 18465.79 8541.195 18488.86 8542.315 ;
      RECT 18465.79 8550.435 18488.86 8556.205 ;
      RECT 18465.79 8558.205 18488.86 8569.745 ;
      RECT 18465.79 8571.745 18488.86 8577.515 ;
      RECT 18465.79 8585.635 18488.86 8586.755 ;
      RECT 18465.79 8588.755 18488.86 8593.365 ;
      RECT 18465.79 8595.365 18488.86 8599.975 ;
      RECT 18465.79 552.315 18488.36 552.875 ;
      RECT 18465.79 591.075 18488.36 591.635 ;
      RECT 18465.79 624.315 18488.36 624.875 ;
      RECT 18465.79 663.075 18488.36 663.635 ;
      RECT 18465.79 696.315 18488.36 696.875 ;
      RECT 18465.79 735.075 18488.36 735.635 ;
      RECT 18465.79 768.315 18488.36 768.875 ;
      RECT 18465.79 807.075 18488.36 807.635 ;
      RECT 18465.79 840.315 18488.36 840.875 ;
      RECT 18465.79 879.075 18488.36 879.635 ;
      RECT 18465.79 912.315 18488.36 912.875 ;
      RECT 18465.79 951.075 18488.36 951.635 ;
      RECT 18465.79 984.315 18488.36 984.875 ;
      RECT 18465.79 1023.075 18488.36 1023.635 ;
      RECT 18465.79 1056.315 18488.36 1056.875 ;
      RECT 18465.79 1095.075 18488.36 1095.635 ;
      RECT 18465.79 1128.315 18488.36 1128.875 ;
      RECT 18465.79 1167.075 18488.36 1167.635 ;
      RECT 18465.79 1200.315 18488.36 1200.875 ;
      RECT 18465.79 1239.075 18488.36 1239.635 ;
      RECT 18465.79 1272.315 18488.36 1272.875 ;
      RECT 18465.79 1311.075 18488.36 1311.635 ;
      RECT 18465.79 1344.315 18488.36 1344.875 ;
      RECT 18465.79 1383.075 18488.36 1383.635 ;
      RECT 18465.79 1416.315 18488.36 1416.875 ;
      RECT 18465.79 1455.075 18488.36 1455.635 ;
      RECT 18465.79 1488.315 18488.36 1488.875 ;
      RECT 18465.79 1527.075 18488.36 1527.635 ;
      RECT 18465.79 1560.315 18488.36 1560.875 ;
      RECT 18465.79 1599.075 18488.36 1599.635 ;
      RECT 18465.79 1632.315 18488.36 1632.875 ;
      RECT 18465.79 1671.075 18488.36 1671.635 ;
      RECT 18465.79 1704.315 18488.36 1704.875 ;
      RECT 18465.79 1743.075 18488.36 1743.635 ;
      RECT 18465.79 1776.315 18488.36 1776.875 ;
      RECT 18465.79 1815.075 18488.36 1815.635 ;
      RECT 18465.79 1848.315 18488.36 1848.875 ;
      RECT 18465.79 1887.075 18488.36 1887.635 ;
      RECT 18465.79 1920.315 18488.36 1920.875 ;
      RECT 18465.79 1959.075 18488.36 1959.635 ;
      RECT 18465.79 1992.315 18488.36 1992.875 ;
      RECT 18465.79 2031.075 18488.36 2031.635 ;
      RECT 18465.79 2064.315 18488.36 2064.875 ;
      RECT 18465.79 2103.075 18488.36 2103.635 ;
      RECT 18465.79 2136.315 18488.36 2136.875 ;
      RECT 18465.79 2175.075 18488.36 2175.635 ;
      RECT 18465.79 2208.315 18488.36 2208.875 ;
      RECT 18465.79 2247.075 18488.36 2247.635 ;
      RECT 18465.79 2280.315 18488.36 2280.875 ;
      RECT 18465.79 2319.075 18488.36 2319.635 ;
      RECT 18465.79 2352.315 18488.36 2352.875 ;
      RECT 18465.79 2391.075 18488.36 2391.635 ;
      RECT 18465.79 2424.315 18488.36 2424.875 ;
      RECT 18465.79 2463.075 18488.36 2463.635 ;
      RECT 18465.79 2496.315 18488.36 2496.875 ;
      RECT 18465.79 2535.075 18488.36 2535.635 ;
      RECT 18465.79 2568.315 18488.36 2568.875 ;
      RECT 18465.79 2607.075 18488.36 2607.635 ;
      RECT 18465.79 2640.315 18488.36 2640.875 ;
      RECT 18465.79 2679.075 18488.36 2679.635 ;
      RECT 18465.79 2712.315 18488.36 2712.875 ;
      RECT 18465.79 2751.075 18488.36 2751.635 ;
      RECT 18465.79 2784.315 18488.36 2784.875 ;
      RECT 18465.79 2823.075 18488.36 2823.635 ;
      RECT 18465.79 2856.315 18488.36 2856.875 ;
      RECT 18465.79 2895.075 18488.36 2895.635 ;
      RECT 18465.79 2928.315 18488.36 2928.875 ;
      RECT 18465.79 2967.075 18488.36 2967.635 ;
      RECT 18465.79 3000.315 18488.36 3000.875 ;
      RECT 18465.79 3039.075 18488.36 3039.635 ;
      RECT 18465.79 3072.315 18488.36 3072.875 ;
      RECT 18465.79 3111.075 18488.36 3111.635 ;
      RECT 18465.79 3144.315 18488.36 3144.875 ;
      RECT 18465.79 3183.075 18488.36 3183.635 ;
      RECT 18465.79 3216.315 18488.36 3216.875 ;
      RECT 18465.79 3255.075 18488.36 3255.635 ;
      RECT 18465.79 3288.315 18488.36 3288.875 ;
      RECT 18465.79 3327.075 18488.36 3327.635 ;
      RECT 18465.79 3360.315 18488.36 3360.875 ;
      RECT 18465.79 3399.075 18488.36 3399.635 ;
      RECT 18465.79 3432.315 18488.36 3432.875 ;
      RECT 18465.79 3471.075 18488.36 3471.635 ;
      RECT 18465.79 3504.315 18488.36 3504.875 ;
      RECT 18465.79 3543.075 18488.36 3543.635 ;
      RECT 18465.79 3576.315 18488.36 3576.875 ;
      RECT 18465.79 3615.075 18488.36 3615.635 ;
      RECT 18465.79 3648.315 18488.36 3648.875 ;
      RECT 18465.79 3687.075 18488.36 3687.635 ;
      RECT 18465.79 3720.315 18488.36 3720.875 ;
      RECT 18465.79 3759.075 18488.36 3759.635 ;
      RECT 18465.79 3792.315 18488.36 3792.875 ;
      RECT 18465.79 3831.075 18488.36 3831.635 ;
      RECT 18465.79 3864.315 18488.36 3864.875 ;
      RECT 18465.79 3903.075 18488.36 3903.635 ;
      RECT 18465.79 3936.315 18488.36 3936.875 ;
      RECT 18465.79 3975.075 18488.36 3975.635 ;
      RECT 18465.79 4008.315 18488.36 4008.875 ;
      RECT 18465.79 4047.075 18488.36 4047.635 ;
      RECT 18465.79 4080.315 18488.36 4080.875 ;
      RECT 18465.79 4119.075 18488.36 4119.635 ;
      RECT 18465.79 4152.315 18488.36 4152.875 ;
      RECT 18465.79 4191.075 18488.36 4191.635 ;
      RECT 18465.79 4224.315 18488.36 4224.875 ;
      RECT 18465.79 4263.075 18488.36 4263.635 ;
      RECT 18465.79 4296.315 18488.36 4296.875 ;
      RECT 18465.79 4335.075 18488.36 4335.635 ;
      RECT 18465.79 4368.315 18488.36 4368.875 ;
      RECT 18465.79 4407.075 18488.36 4407.635 ;
      RECT 18465.79 4440.315 18488.36 4440.875 ;
      RECT 18465.79 4479.075 18488.36 4479.635 ;
      RECT 18465.79 4512.315 18488.36 4512.875 ;
      RECT 18465.79 4551.075 18488.36 4551.635 ;
      RECT 18465.79 4584.315 18488.36 4584.875 ;
      RECT 18465.79 4623.075 18488.36 4623.635 ;
      RECT 18465.79 4656.315 18488.36 4656.875 ;
      RECT 18465.79 4695.075 18488.36 4695.635 ;
      RECT 18465.79 4728.315 18488.36 4728.875 ;
      RECT 18465.79 4767.075 18488.36 4767.635 ;
      RECT 18465.79 4800.315 18488.36 4800.875 ;
      RECT 18465.79 4839.075 18488.36 4839.635 ;
      RECT 18465.79 4872.315 18488.36 4872.875 ;
      RECT 18465.79 4911.075 18488.36 4911.635 ;
      RECT 18465.79 4944.315 18488.36 4944.875 ;
      RECT 18465.79 4983.075 18488.36 4983.635 ;
      RECT 18465.79 5016.315 18488.36 5016.875 ;
      RECT 18465.79 5055.075 18488.36 5055.635 ;
      RECT 18465.79 5088.315 18488.36 5088.875 ;
      RECT 18465.79 5127.075 18488.36 5127.635 ;
      RECT 18465.79 5160.315 18488.36 5160.875 ;
      RECT 18465.79 5199.075 18488.36 5199.635 ;
      RECT 18465.79 5232.315 18488.36 5232.875 ;
      RECT 18465.79 5271.075 18488.36 5271.635 ;
      RECT 18465.79 5304.315 18488.36 5304.875 ;
      RECT 18465.79 5343.075 18488.36 5343.635 ;
      RECT 18465.79 5376.315 18488.36 5376.875 ;
      RECT 18465.79 5415.075 18488.36 5415.635 ;
      RECT 18465.79 5448.315 18488.36 5448.875 ;
      RECT 18465.79 5487.075 18488.36 5487.635 ;
      RECT 18465.79 5520.315 18488.36 5520.875 ;
      RECT 18465.79 5559.075 18488.36 5559.635 ;
      RECT 18465.79 5592.315 18488.36 5592.875 ;
      RECT 18465.79 5631.075 18488.36 5631.635 ;
      RECT 18465.79 5664.315 18488.36 5664.875 ;
      RECT 18465.79 5703.075 18488.36 5703.635 ;
      RECT 18465.79 5736.315 18488.36 5736.875 ;
      RECT 18465.79 5775.075 18488.36 5775.635 ;
      RECT 18465.79 5808.315 18488.36 5808.875 ;
      RECT 18465.79 5847.075 18488.36 5847.635 ;
      RECT 18465.79 5880.315 18488.36 5880.875 ;
      RECT 18465.79 5919.075 18488.36 5919.635 ;
      RECT 18465.79 5952.315 18488.36 5952.875 ;
      RECT 18465.79 5991.075 18488.36 5991.635 ;
      RECT 18465.79 6024.315 18488.36 6024.875 ;
      RECT 18465.79 6063.075 18488.36 6063.635 ;
      RECT 18465.79 6096.315 18488.36 6096.875 ;
      RECT 18465.79 6135.075 18488.36 6135.635 ;
      RECT 18465.79 6168.315 18488.36 6168.875 ;
      RECT 18465.79 6207.075 18488.36 6207.635 ;
      RECT 18465.79 6240.315 18488.36 6240.875 ;
      RECT 18465.79 6279.075 18488.36 6279.635 ;
      RECT 18465.79 6312.315 18488.36 6312.875 ;
      RECT 18465.79 6351.075 18488.36 6351.635 ;
      RECT 18465.79 6384.315 18488.36 6384.875 ;
      RECT 18465.79 6423.075 18488.36 6423.635 ;
      RECT 18465.79 6456.315 18488.36 6456.875 ;
      RECT 18465.79 6495.075 18488.36 6495.635 ;
      RECT 18465.79 6528.315 18488.36 6528.875 ;
      RECT 18465.79 6567.075 18488.36 6567.635 ;
      RECT 18465.79 6600.315 18488.36 6600.875 ;
      RECT 18465.79 6639.075 18488.36 6639.635 ;
      RECT 18465.79 6672.315 18488.36 6672.875 ;
      RECT 18465.79 6711.075 18488.36 6711.635 ;
      RECT 18465.79 6744.315 18488.36 6744.875 ;
      RECT 18465.79 6783.075 18488.36 6783.635 ;
      RECT 18465.79 6816.315 18488.36 6816.875 ;
      RECT 18465.79 6855.075 18488.36 6855.635 ;
      RECT 18465.79 6888.315 18488.36 6888.875 ;
      RECT 18465.79 6927.075 18488.36 6927.635 ;
      RECT 18465.79 6960.315 18488.36 6960.875 ;
      RECT 18465.79 6999.075 18488.36 6999.635 ;
      RECT 18465.79 7032.315 18488.36 7032.875 ;
      RECT 18465.79 7071.075 18488.36 7071.635 ;
      RECT 18465.79 7104.315 18488.36 7104.875 ;
      RECT 18465.79 7143.075 18488.36 7143.635 ;
      RECT 18465.79 7176.315 18488.36 7176.875 ;
      RECT 18465.79 7215.075 18488.36 7215.635 ;
      RECT 18465.79 7248.315 18488.36 7248.875 ;
      RECT 18465.79 7287.075 18488.36 7287.635 ;
      RECT 18465.79 7320.315 18488.36 7320.875 ;
      RECT 18465.79 7359.075 18488.36 7359.635 ;
      RECT 18465.79 7392.315 18488.36 7392.875 ;
      RECT 18465.79 7431.075 18488.36 7431.635 ;
      RECT 18465.79 7464.315 18488.36 7464.875 ;
      RECT 18465.79 7503.075 18488.36 7503.635 ;
      RECT 18465.79 7536.315 18488.36 7536.875 ;
      RECT 18465.79 7575.075 18488.36 7575.635 ;
      RECT 18465.79 7608.315 18488.36 7608.875 ;
      RECT 18465.79 7647.075 18488.36 7647.635 ;
      RECT 18465.79 7680.315 18488.36 7680.875 ;
      RECT 18465.79 7719.075 18488.36 7719.635 ;
      RECT 18465.79 7752.315 18488.36 7752.875 ;
      RECT 18465.79 7791.075 18488.36 7791.635 ;
      RECT 18465.79 7824.315 18488.36 7824.875 ;
      RECT 18465.79 7863.075 18488.36 7863.635 ;
      RECT 18465.79 7896.315 18488.36 7896.875 ;
      RECT 18465.79 7935.075 18488.36 7935.635 ;
      RECT 18465.79 7968.315 18488.36 7968.875 ;
      RECT 18465.79 8007.075 18488.36 8007.635 ;
      RECT 18465.79 8040.315 18488.36 8040.875 ;
      RECT 18465.79 8079.075 18488.36 8079.635 ;
      RECT 18465.79 8112.315 18488.36 8112.875 ;
      RECT 18465.79 8151.075 18488.36 8151.635 ;
      RECT 18465.79 8184.315 18488.36 8184.875 ;
      RECT 18465.79 8223.075 18488.36 8223.635 ;
      RECT 18465.79 8256.315 18488.36 8256.875 ;
      RECT 18465.79 8295.075 18488.36 8295.635 ;
      RECT 18465.79 8328.315 18488.36 8328.875 ;
      RECT 18465.79 8367.075 18488.36 8367.635 ;
      RECT 18465.79 8400.315 18488.36 8400.875 ;
      RECT 18465.79 8439.075 18488.36 8439.635 ;
      RECT 18465.79 8472.315 18488.36 8472.875 ;
      RECT 18465.79 8511.075 18488.36 8511.635 ;
      RECT 18465.79 8544.315 18488.36 8544.875 ;
      RECT 18465.79 8583.075 18488.36 8583.635 ;
      RECT 328.26 500.265 448.95 510.265 ;
      RECT 328.26 512.265 448.95 514.265 ;
      RECT 328.26 191.275 448.56 193.275 ;
      RECT 328.26 196.245 448.56 210.275 ;
      RECT 328.26 213.245 448.56 227.275 ;
      RECT 328.26 230.245 448.56 258.275 ;
      RECT 328.26 261.245 448.56 289.275 ;
      RECT 328.26 292.245 448.56 306.275 ;
      RECT 328.26 309.245 448.56 323.275 ;
      RECT 326.66 339.555 448.56 372.555 ;
      RECT 326.66 382.555 448.56 415.555 ;
      RECT 326.66 425.555 448.56 458.555 ;
      RECT 326.66 468.555 448.56 496.265 ;
      RECT 328.26 521.56 351.33 522.68 ;
      RECT 328.26 535.975 351.33 540.585 ;
      RECT 328.26 542.585 351.33 547.195 ;
      RECT 328.26 549.195 351.33 550.315 ;
      RECT 328.26 558.435 351.33 564.205 ;
      RECT 328.26 566.205 351.33 577.745 ;
      RECT 328.26 579.745 351.33 585.515 ;
      RECT 328.26 593.635 351.33 594.755 ;
      RECT 328.26 596.755 351.33 601.365 ;
      RECT 328.26 603.365 351.33 612.585 ;
      RECT 328.26 614.585 351.33 619.195 ;
      RECT 328.26 621.195 351.33 622.315 ;
      RECT 328.26 630.435 351.33 636.205 ;
      RECT 328.26 638.205 351.33 649.745 ;
      RECT 328.26 651.745 351.33 657.515 ;
      RECT 328.26 665.635 351.33 666.755 ;
      RECT 328.26 668.755 351.33 673.365 ;
      RECT 328.26 675.365 351.33 684.585 ;
      RECT 328.26 686.585 351.33 691.195 ;
      RECT 328.26 693.195 351.33 694.315 ;
      RECT 328.26 702.435 351.33 708.205 ;
      RECT 328.26 710.205 351.33 721.745 ;
      RECT 328.26 723.745 351.33 729.515 ;
      RECT 328.26 737.635 351.33 738.755 ;
      RECT 328.26 740.755 351.33 745.365 ;
      RECT 328.26 747.365 351.33 756.585 ;
      RECT 328.26 758.585 351.33 763.195 ;
      RECT 328.26 765.195 351.33 766.315 ;
      RECT 328.26 774.435 351.33 780.205 ;
      RECT 328.26 782.205 351.33 793.745 ;
      RECT 328.26 795.745 351.33 801.515 ;
      RECT 328.26 809.635 351.33 810.755 ;
      RECT 328.26 812.755 351.33 817.365 ;
      RECT 328.26 819.365 351.33 828.585 ;
      RECT 328.26 830.585 351.33 835.195 ;
      RECT 328.26 837.195 351.33 838.315 ;
      RECT 328.26 846.435 351.33 852.205 ;
      RECT 328.26 854.205 351.33 865.745 ;
      RECT 328.26 867.745 351.33 873.515 ;
      RECT 328.26 881.635 351.33 882.755 ;
      RECT 328.26 884.755 351.33 889.365 ;
      RECT 328.26 891.365 351.33 900.585 ;
      RECT 328.26 902.585 351.33 907.195 ;
      RECT 328.26 909.195 351.33 910.315 ;
      RECT 328.26 918.435 351.33 924.205 ;
      RECT 328.26 926.205 351.33 937.745 ;
      RECT 328.26 939.745 351.33 945.515 ;
      RECT 328.26 953.635 351.33 954.755 ;
      RECT 328.26 956.755 351.33 961.365 ;
      RECT 328.26 963.365 351.33 972.585 ;
      RECT 328.26 974.585 351.33 979.195 ;
      RECT 328.26 981.195 351.33 982.315 ;
      RECT 328.26 990.435 351.33 996.205 ;
      RECT 328.26 998.205 351.33 1009.745 ;
      RECT 328.26 1011.745 351.33 1017.515 ;
      RECT 328.26 1025.635 351.33 1026.755 ;
      RECT 328.26 1028.755 351.33 1033.365 ;
      RECT 328.26 1035.365 351.33 1044.585 ;
      RECT 328.26 1046.585 351.33 1051.195 ;
      RECT 328.26 1053.195 351.33 1054.315 ;
      RECT 328.26 1062.435 351.33 1068.205 ;
      RECT 328.26 1070.205 351.33 1081.745 ;
      RECT 328.26 1083.745 351.33 1089.515 ;
      RECT 328.26 1097.635 351.33 1098.755 ;
      RECT 328.26 1100.755 351.33 1105.365 ;
      RECT 328.26 1107.365 351.33 1116.585 ;
      RECT 328.26 1118.585 351.33 1123.195 ;
      RECT 328.26 1125.195 351.33 1126.315 ;
      RECT 328.26 1134.435 351.33 1140.205 ;
      RECT 328.26 1142.205 351.33 1153.745 ;
      RECT 328.26 1155.745 351.33 1161.515 ;
      RECT 328.26 1169.635 351.33 1170.755 ;
      RECT 328.26 1172.755 351.33 1177.365 ;
      RECT 328.26 1179.365 351.33 1188.585 ;
      RECT 328.26 1190.585 351.33 1195.195 ;
      RECT 328.26 1197.195 351.33 1198.315 ;
      RECT 328.26 1206.435 351.33 1212.205 ;
      RECT 328.26 1214.205 351.33 1225.745 ;
      RECT 328.26 1227.745 351.33 1233.515 ;
      RECT 328.26 1241.635 351.33 1242.755 ;
      RECT 328.26 1244.755 351.33 1249.365 ;
      RECT 328.26 1251.365 351.33 1260.585 ;
      RECT 328.26 1262.585 351.33 1267.195 ;
      RECT 328.26 1269.195 351.33 1270.315 ;
      RECT 328.26 1278.435 351.33 1284.205 ;
      RECT 328.26 1286.205 351.33 1297.745 ;
      RECT 328.26 1299.745 351.33 1305.515 ;
      RECT 328.26 1313.635 351.33 1314.755 ;
      RECT 328.26 1316.755 351.33 1321.365 ;
      RECT 328.26 1323.365 351.33 1332.585 ;
      RECT 328.26 1334.585 351.33 1339.195 ;
      RECT 328.26 1341.195 351.33 1342.315 ;
      RECT 328.26 1350.435 351.33 1356.205 ;
      RECT 328.26 1358.205 351.33 1369.745 ;
      RECT 328.26 1371.745 351.33 1377.515 ;
      RECT 328.26 1385.635 351.33 1386.755 ;
      RECT 328.26 1388.755 351.33 1393.365 ;
      RECT 328.26 1395.365 351.33 1404.585 ;
      RECT 328.26 1406.585 351.33 1411.195 ;
      RECT 328.26 1413.195 351.33 1414.315 ;
      RECT 328.26 1422.435 351.33 1428.205 ;
      RECT 328.26 1430.205 351.33 1441.745 ;
      RECT 328.26 1443.745 351.33 1449.515 ;
      RECT 328.26 1457.635 351.33 1458.755 ;
      RECT 328.26 1460.755 351.33 1465.365 ;
      RECT 328.26 1467.365 351.33 1476.585 ;
      RECT 328.26 1478.585 351.33 1483.195 ;
      RECT 328.26 1485.195 351.33 1486.315 ;
      RECT 328.26 1494.435 351.33 1500.205 ;
      RECT 328.26 1502.205 351.33 1513.745 ;
      RECT 328.26 1515.745 351.33 1521.515 ;
      RECT 328.26 1529.635 351.33 1530.755 ;
      RECT 328.26 1532.755 351.33 1537.365 ;
      RECT 328.26 1539.365 351.33 1548.585 ;
      RECT 328.26 1550.585 351.33 1555.195 ;
      RECT 328.26 1557.195 351.33 1558.315 ;
      RECT 328.26 1566.435 351.33 1572.205 ;
      RECT 328.26 1574.205 351.33 1585.745 ;
      RECT 328.26 1587.745 351.33 1593.515 ;
      RECT 328.26 1601.635 351.33 1602.755 ;
      RECT 328.26 1604.755 351.33 1609.365 ;
      RECT 328.26 1611.365 351.33 1620.585 ;
      RECT 328.26 1622.585 351.33 1627.195 ;
      RECT 328.26 1629.195 351.33 1630.315 ;
      RECT 328.26 1638.435 351.33 1644.205 ;
      RECT 328.26 1646.205 351.33 1657.745 ;
      RECT 328.26 1659.745 351.33 1665.515 ;
      RECT 328.26 1673.635 351.33 1674.755 ;
      RECT 328.26 1676.755 351.33 1681.365 ;
      RECT 328.26 1683.365 351.33 1692.585 ;
      RECT 328.26 1694.585 351.33 1699.195 ;
      RECT 328.26 1701.195 351.33 1702.315 ;
      RECT 328.26 1710.435 351.33 1716.205 ;
      RECT 328.26 1718.205 351.33 1729.745 ;
      RECT 328.26 1731.745 351.33 1737.515 ;
      RECT 328.26 1745.635 351.33 1746.755 ;
      RECT 328.26 1748.755 351.33 1753.365 ;
      RECT 328.26 1755.365 351.33 1764.585 ;
      RECT 328.26 1766.585 351.33 1771.195 ;
      RECT 328.26 1773.195 351.33 1774.315 ;
      RECT 328.26 1782.435 351.33 1788.205 ;
      RECT 328.26 1790.205 351.33 1801.745 ;
      RECT 328.26 1803.745 351.33 1809.515 ;
      RECT 328.26 1817.635 351.33 1818.755 ;
      RECT 328.26 1820.755 351.33 1825.365 ;
      RECT 328.26 1827.365 351.33 1836.585 ;
      RECT 328.26 1838.585 351.33 1843.195 ;
      RECT 328.26 1845.195 351.33 1846.315 ;
      RECT 328.26 1854.435 351.33 1860.205 ;
      RECT 328.26 1862.205 351.33 1873.745 ;
      RECT 328.26 1875.745 351.33 1881.515 ;
      RECT 328.26 1889.635 351.33 1890.755 ;
      RECT 328.26 1892.755 351.33 1897.365 ;
      RECT 328.26 1899.365 351.33 1908.585 ;
      RECT 328.26 1910.585 351.33 1915.195 ;
      RECT 328.26 1917.195 351.33 1918.315 ;
      RECT 328.26 1926.435 351.33 1932.205 ;
      RECT 328.26 1934.205 351.33 1945.745 ;
      RECT 328.26 1947.745 351.33 1953.515 ;
      RECT 328.26 1961.635 351.33 1962.755 ;
      RECT 328.26 1964.755 351.33 1969.365 ;
      RECT 328.26 1971.365 351.33 1980.585 ;
      RECT 328.26 1982.585 351.33 1987.195 ;
      RECT 328.26 1989.195 351.33 1990.315 ;
      RECT 328.26 1998.435 351.33 2004.205 ;
      RECT 328.26 2006.205 351.33 2017.745 ;
      RECT 328.26 2019.745 351.33 2025.515 ;
      RECT 328.26 2033.635 351.33 2034.755 ;
      RECT 328.26 2036.755 351.33 2041.365 ;
      RECT 328.26 2043.365 351.33 2052.585 ;
      RECT 328.26 2054.585 351.33 2059.195 ;
      RECT 328.26 2061.195 351.33 2062.315 ;
      RECT 328.26 2070.435 351.33 2076.205 ;
      RECT 328.26 2078.205 351.33 2089.745 ;
      RECT 328.26 2091.745 351.33 2097.515 ;
      RECT 328.26 2105.635 351.33 2106.755 ;
      RECT 328.26 2108.755 351.33 2113.365 ;
      RECT 328.26 2115.365 351.33 2124.585 ;
      RECT 328.26 2126.585 351.33 2131.195 ;
      RECT 328.26 2133.195 351.33 2134.315 ;
      RECT 328.26 2142.435 351.33 2148.205 ;
      RECT 328.26 2150.205 351.33 2161.745 ;
      RECT 328.26 2163.745 351.33 2169.515 ;
      RECT 328.26 2177.635 351.33 2178.755 ;
      RECT 328.26 2180.755 351.33 2185.365 ;
      RECT 328.26 2187.365 351.33 2196.585 ;
      RECT 328.26 2198.585 351.33 2203.195 ;
      RECT 328.26 2205.195 351.33 2206.315 ;
      RECT 328.26 2214.435 351.33 2220.205 ;
      RECT 328.26 2222.205 351.33 2233.745 ;
      RECT 328.26 2235.745 351.33 2241.515 ;
      RECT 328.26 2249.635 351.33 2250.755 ;
      RECT 328.26 2252.755 351.33 2257.365 ;
      RECT 328.26 2259.365 351.33 2268.585 ;
      RECT 328.26 2270.585 351.33 2275.195 ;
      RECT 328.26 2277.195 351.33 2278.315 ;
      RECT 328.26 2286.435 351.33 2292.205 ;
      RECT 328.26 2294.205 351.33 2305.745 ;
      RECT 328.26 2307.745 351.33 2313.515 ;
      RECT 328.26 2321.635 351.33 2322.755 ;
      RECT 328.26 2324.755 351.33 2329.365 ;
      RECT 328.26 2331.365 351.33 2340.585 ;
      RECT 328.26 2342.585 351.33 2347.195 ;
      RECT 328.26 2349.195 351.33 2350.315 ;
      RECT 328.26 2358.435 351.33 2364.205 ;
      RECT 328.26 2366.205 351.33 2377.745 ;
      RECT 328.26 2379.745 351.33 2385.515 ;
      RECT 328.26 2393.635 351.33 2394.755 ;
      RECT 328.26 2396.755 351.33 2401.365 ;
      RECT 328.26 2403.365 351.33 2412.585 ;
      RECT 328.26 2414.585 351.33 2419.195 ;
      RECT 328.26 2421.195 351.33 2422.315 ;
      RECT 328.26 2430.435 351.33 2436.205 ;
      RECT 328.26 2438.205 351.33 2449.745 ;
      RECT 328.26 2451.745 351.33 2457.515 ;
      RECT 328.26 2465.635 351.33 2466.755 ;
      RECT 328.26 2468.755 351.33 2473.365 ;
      RECT 328.26 2475.365 351.33 2484.585 ;
      RECT 328.26 2486.585 351.33 2491.195 ;
      RECT 328.26 2493.195 351.33 2494.315 ;
      RECT 328.26 2502.435 351.33 2508.205 ;
      RECT 328.26 2510.205 351.33 2521.745 ;
      RECT 328.26 2523.745 351.33 2529.515 ;
      RECT 328.26 2537.635 351.33 2538.755 ;
      RECT 328.26 2540.755 351.33 2545.365 ;
      RECT 328.26 2547.365 351.33 2556.585 ;
      RECT 328.26 2558.585 351.33 2563.195 ;
      RECT 328.26 2565.195 351.33 2566.315 ;
      RECT 328.26 2574.435 351.33 2580.205 ;
      RECT 328.26 2582.205 351.33 2593.745 ;
      RECT 328.26 2595.745 351.33 2601.515 ;
      RECT 328.26 2609.635 351.33 2610.755 ;
      RECT 328.26 2612.755 351.33 2617.365 ;
      RECT 328.26 2619.365 351.33 2628.585 ;
      RECT 328.26 2630.585 351.33 2635.195 ;
      RECT 328.26 2637.195 351.33 2638.315 ;
      RECT 328.26 2646.435 351.33 2652.205 ;
      RECT 328.26 2654.205 351.33 2665.745 ;
      RECT 328.26 2667.745 351.33 2673.515 ;
      RECT 328.26 2681.635 351.33 2682.755 ;
      RECT 328.26 2684.755 351.33 2689.365 ;
      RECT 328.26 2691.365 351.33 2700.585 ;
      RECT 328.26 2702.585 351.33 2707.195 ;
      RECT 328.26 2709.195 351.33 2710.315 ;
      RECT 328.26 2718.435 351.33 2724.205 ;
      RECT 328.26 2726.205 351.33 2737.745 ;
      RECT 328.26 2739.745 351.33 2745.515 ;
      RECT 328.26 2753.635 351.33 2754.755 ;
      RECT 328.26 2756.755 351.33 2761.365 ;
      RECT 328.26 2763.365 351.33 2772.585 ;
      RECT 328.26 2774.585 351.33 2779.195 ;
      RECT 328.26 2781.195 351.33 2782.315 ;
      RECT 328.26 2790.435 351.33 2796.205 ;
      RECT 328.26 2798.205 351.33 2809.745 ;
      RECT 328.26 2811.745 351.33 2817.515 ;
      RECT 328.26 2825.635 351.33 2826.755 ;
      RECT 328.26 2828.755 351.33 2833.365 ;
      RECT 328.26 2835.365 351.33 2844.585 ;
      RECT 328.26 2846.585 351.33 2851.195 ;
      RECT 328.26 2853.195 351.33 2854.315 ;
      RECT 328.26 2862.435 351.33 2868.205 ;
      RECT 328.26 2870.205 351.33 2881.745 ;
      RECT 328.26 2883.745 351.33 2889.515 ;
      RECT 328.26 2897.635 351.33 2898.755 ;
      RECT 328.26 2900.755 351.33 2905.365 ;
      RECT 328.26 2907.365 351.33 2916.585 ;
      RECT 328.26 2918.585 351.33 2923.195 ;
      RECT 328.26 2925.195 351.33 2926.315 ;
      RECT 328.26 2934.435 351.33 2940.205 ;
      RECT 328.26 2942.205 351.33 2953.745 ;
      RECT 328.26 2955.745 351.33 2961.515 ;
      RECT 328.26 2969.635 351.33 2970.755 ;
      RECT 328.26 2972.755 351.33 2977.365 ;
      RECT 328.26 2979.365 351.33 2988.585 ;
      RECT 328.26 2990.585 351.33 2995.195 ;
      RECT 328.26 2997.195 351.33 2998.315 ;
      RECT 328.26 3006.435 351.33 3012.205 ;
      RECT 328.26 3014.205 351.33 3025.745 ;
      RECT 328.26 3027.745 351.33 3033.515 ;
      RECT 328.26 3041.635 351.33 3042.755 ;
      RECT 328.26 3044.755 351.33 3049.365 ;
      RECT 328.26 3051.365 351.33 3060.585 ;
      RECT 328.26 3062.585 351.33 3067.195 ;
      RECT 328.26 3069.195 351.33 3070.315 ;
      RECT 328.26 3078.435 351.33 3084.205 ;
      RECT 328.26 3086.205 351.33 3097.745 ;
      RECT 328.26 3099.745 351.33 3105.515 ;
      RECT 328.26 3113.635 351.33 3114.755 ;
      RECT 328.26 3116.755 351.33 3121.365 ;
      RECT 328.26 3123.365 351.33 3132.585 ;
      RECT 328.26 3134.585 351.33 3139.195 ;
      RECT 328.26 3141.195 351.33 3142.315 ;
      RECT 328.26 3150.435 351.33 3156.205 ;
      RECT 328.26 3158.205 351.33 3169.745 ;
      RECT 328.26 3171.745 351.33 3177.515 ;
      RECT 328.26 3185.635 351.33 3186.755 ;
      RECT 328.26 3188.755 351.33 3193.365 ;
      RECT 328.26 3195.365 351.33 3204.585 ;
      RECT 328.26 3206.585 351.33 3211.195 ;
      RECT 328.26 3213.195 351.33 3214.315 ;
      RECT 328.26 3222.435 351.33 3228.205 ;
      RECT 328.26 3230.205 351.33 3241.745 ;
      RECT 328.26 3243.745 351.33 3249.515 ;
      RECT 328.26 3257.635 351.33 3258.755 ;
      RECT 328.26 3260.755 351.33 3265.365 ;
      RECT 328.26 3267.365 351.33 3276.585 ;
      RECT 328.26 3278.585 351.33 3283.195 ;
      RECT 328.26 3285.195 351.33 3286.315 ;
      RECT 328.26 3294.435 351.33 3300.205 ;
      RECT 328.26 3302.205 351.33 3313.745 ;
      RECT 328.26 3315.745 351.33 3321.515 ;
      RECT 328.26 3329.635 351.33 3330.755 ;
      RECT 328.26 3332.755 351.33 3337.365 ;
      RECT 328.26 3339.365 351.33 3348.585 ;
      RECT 328.26 3350.585 351.33 3355.195 ;
      RECT 328.26 3357.195 351.33 3358.315 ;
      RECT 328.26 3366.435 351.33 3372.205 ;
      RECT 328.26 3374.205 351.33 3385.745 ;
      RECT 328.26 3387.745 351.33 3393.515 ;
      RECT 328.26 3401.635 351.33 3402.755 ;
      RECT 328.26 3404.755 351.33 3409.365 ;
      RECT 328.26 3411.365 351.33 3420.585 ;
      RECT 328.26 3422.585 351.33 3427.195 ;
      RECT 328.26 3429.195 351.33 3430.315 ;
      RECT 328.26 3438.435 351.33 3444.205 ;
      RECT 328.26 3446.205 351.33 3457.745 ;
      RECT 328.26 3459.745 351.33 3465.515 ;
      RECT 328.26 3473.635 351.33 3474.755 ;
      RECT 328.26 3476.755 351.33 3481.365 ;
      RECT 328.26 3483.365 351.33 3492.585 ;
      RECT 328.26 3494.585 351.33 3499.195 ;
      RECT 328.26 3501.195 351.33 3502.315 ;
      RECT 328.26 3510.435 351.33 3516.205 ;
      RECT 328.26 3518.205 351.33 3529.745 ;
      RECT 328.26 3531.745 351.33 3537.515 ;
      RECT 328.26 3545.635 351.33 3546.755 ;
      RECT 328.26 3548.755 351.33 3553.365 ;
      RECT 328.26 3555.365 351.33 3564.585 ;
      RECT 328.26 3566.585 351.33 3571.195 ;
      RECT 328.26 3573.195 351.33 3574.315 ;
      RECT 328.26 3582.435 351.33 3588.205 ;
      RECT 328.26 3590.205 351.33 3601.745 ;
      RECT 328.26 3603.745 351.33 3609.515 ;
      RECT 328.26 3617.635 351.33 3618.755 ;
      RECT 328.26 3620.755 351.33 3625.365 ;
      RECT 328.26 3627.365 351.33 3636.585 ;
      RECT 328.26 3638.585 351.33 3643.195 ;
      RECT 328.26 3645.195 351.33 3646.315 ;
      RECT 328.26 3654.435 351.33 3660.205 ;
      RECT 328.26 3662.205 351.33 3673.745 ;
      RECT 328.26 3675.745 351.33 3681.515 ;
      RECT 328.26 3689.635 351.33 3690.755 ;
      RECT 328.26 3692.755 351.33 3697.365 ;
      RECT 328.26 3699.365 351.33 3708.585 ;
      RECT 328.26 3710.585 351.33 3715.195 ;
      RECT 328.26 3717.195 351.33 3718.315 ;
      RECT 328.26 3726.435 351.33 3732.205 ;
      RECT 328.26 3734.205 351.33 3745.745 ;
      RECT 328.26 3747.745 351.33 3753.515 ;
      RECT 328.26 3761.635 351.33 3762.755 ;
      RECT 328.26 3764.755 351.33 3769.365 ;
      RECT 328.26 3771.365 351.33 3780.585 ;
      RECT 328.26 3782.585 351.33 3787.195 ;
      RECT 328.26 3789.195 351.33 3790.315 ;
      RECT 328.26 3798.435 351.33 3804.205 ;
      RECT 328.26 3806.205 351.33 3817.745 ;
      RECT 328.26 3819.745 351.33 3825.515 ;
      RECT 328.26 3833.635 351.33 3834.755 ;
      RECT 328.26 3836.755 351.33 3841.365 ;
      RECT 328.26 3843.365 351.33 3852.585 ;
      RECT 328.26 3854.585 351.33 3859.195 ;
      RECT 328.26 3861.195 351.33 3862.315 ;
      RECT 328.26 3870.435 351.33 3876.205 ;
      RECT 328.26 3878.205 351.33 3889.745 ;
      RECT 328.26 3891.745 351.33 3897.515 ;
      RECT 328.26 3905.635 351.33 3906.755 ;
      RECT 328.26 3908.755 351.33 3913.365 ;
      RECT 328.26 3915.365 351.33 3924.585 ;
      RECT 328.26 3926.585 351.33 3931.195 ;
      RECT 328.26 3933.195 351.33 3934.315 ;
      RECT 328.26 3942.435 351.33 3948.205 ;
      RECT 328.26 3950.205 351.33 3961.745 ;
      RECT 328.26 3963.745 351.33 3969.515 ;
      RECT 328.26 3977.635 351.33 3978.755 ;
      RECT 328.26 3980.755 351.33 3985.365 ;
      RECT 328.26 3987.365 351.33 3996.585 ;
      RECT 328.26 3998.585 351.33 4003.195 ;
      RECT 328.26 4005.195 351.33 4006.315 ;
      RECT 328.26 4014.435 351.33 4020.205 ;
      RECT 328.26 4022.205 351.33 4033.745 ;
      RECT 328.26 4035.745 351.33 4041.515 ;
      RECT 328.26 4049.635 351.33 4050.755 ;
      RECT 328.26 4052.755 351.33 4057.365 ;
      RECT 328.26 4059.365 351.33 4068.585 ;
      RECT 328.26 4070.585 351.33 4075.195 ;
      RECT 328.26 4077.195 351.33 4078.315 ;
      RECT 328.26 4086.435 351.33 4092.205 ;
      RECT 328.26 4094.205 351.33 4105.745 ;
      RECT 328.26 4107.745 351.33 4113.515 ;
      RECT 328.26 4121.635 351.33 4122.755 ;
      RECT 328.26 4124.755 351.33 4129.365 ;
      RECT 328.26 4131.365 351.33 4140.585 ;
      RECT 328.26 4142.585 351.33 4147.195 ;
      RECT 328.26 4149.195 351.33 4150.315 ;
      RECT 328.26 4158.435 351.33 4164.205 ;
      RECT 328.26 4166.205 351.33 4177.745 ;
      RECT 328.26 4179.745 351.33 4185.515 ;
      RECT 328.26 4193.635 351.33 4194.755 ;
      RECT 328.26 4196.755 351.33 4201.365 ;
      RECT 328.26 4203.365 351.33 4212.585 ;
      RECT 328.26 4214.585 351.33 4219.195 ;
      RECT 328.26 4221.195 351.33 4222.315 ;
      RECT 328.26 4230.435 351.33 4236.205 ;
      RECT 328.26 4238.205 351.33 4249.745 ;
      RECT 328.26 4251.745 351.33 4257.515 ;
      RECT 328.26 4265.635 351.33 4266.755 ;
      RECT 328.26 4268.755 351.33 4273.365 ;
      RECT 328.26 4275.365 351.33 4284.585 ;
      RECT 328.26 4286.585 351.33 4291.195 ;
      RECT 328.26 4293.195 351.33 4294.315 ;
      RECT 328.26 4302.435 351.33 4308.205 ;
      RECT 328.26 4310.205 351.33 4321.745 ;
      RECT 328.26 4323.745 351.33 4329.515 ;
      RECT 328.26 4337.635 351.33 4338.755 ;
      RECT 328.26 4340.755 351.33 4345.365 ;
      RECT 328.26 4347.365 351.33 4356.585 ;
      RECT 328.26 4358.585 351.33 4363.195 ;
      RECT 328.26 4365.195 351.33 4366.315 ;
      RECT 328.26 4374.435 351.33 4380.205 ;
      RECT 328.26 4382.205 351.33 4393.745 ;
      RECT 328.26 4395.745 351.33 4401.515 ;
      RECT 328.26 4409.635 351.33 4410.755 ;
      RECT 328.26 4412.755 351.33 4417.365 ;
      RECT 328.26 4419.365 351.33 4428.585 ;
      RECT 328.26 4430.585 351.33 4435.195 ;
      RECT 328.26 4437.195 351.33 4438.315 ;
      RECT 328.26 4446.435 351.33 4452.205 ;
      RECT 328.26 4454.205 351.33 4465.745 ;
      RECT 328.26 4467.745 351.33 4473.515 ;
      RECT 328.26 4481.635 351.33 4482.755 ;
      RECT 328.26 4484.755 351.33 4489.365 ;
      RECT 328.26 4491.365 351.33 4500.585 ;
      RECT 328.26 4502.585 351.33 4507.195 ;
      RECT 328.26 4509.195 351.33 4510.315 ;
      RECT 328.26 4518.435 351.33 4524.205 ;
      RECT 328.26 4526.205 351.33 4537.745 ;
      RECT 328.26 4539.745 351.33 4545.515 ;
      RECT 328.26 4553.635 351.33 4554.755 ;
      RECT 328.26 4556.755 351.33 4561.365 ;
      RECT 328.26 4563.365 351.33 4572.585 ;
      RECT 328.26 4574.585 351.33 4579.195 ;
      RECT 328.26 4581.195 351.33 4582.315 ;
      RECT 328.26 4590.435 351.33 4596.205 ;
      RECT 328.26 4598.205 351.33 4609.745 ;
      RECT 328.26 4611.745 351.33 4617.515 ;
      RECT 328.26 4625.635 351.33 4626.755 ;
      RECT 328.26 4628.755 351.33 4633.365 ;
      RECT 328.26 4635.365 351.33 4644.585 ;
      RECT 328.26 4646.585 351.33 4651.195 ;
      RECT 328.26 4653.195 351.33 4654.315 ;
      RECT 328.26 4662.435 351.33 4668.205 ;
      RECT 328.26 4670.205 351.33 4681.745 ;
      RECT 328.26 4683.745 351.33 4689.515 ;
      RECT 328.26 4697.635 351.33 4698.755 ;
      RECT 328.26 4700.755 351.33 4705.365 ;
      RECT 328.26 4707.365 351.33 4716.585 ;
      RECT 328.26 4718.585 351.33 4723.195 ;
      RECT 328.26 4725.195 351.33 4726.315 ;
      RECT 328.26 4734.435 351.33 4740.205 ;
      RECT 328.26 4742.205 351.33 4753.745 ;
      RECT 328.26 4755.745 351.33 4761.515 ;
      RECT 328.26 4769.635 351.33 4770.755 ;
      RECT 328.26 4772.755 351.33 4777.365 ;
      RECT 328.26 4779.365 351.33 4788.585 ;
      RECT 328.26 4790.585 351.33 4795.195 ;
      RECT 328.26 4797.195 351.33 4798.315 ;
      RECT 328.26 4806.435 351.33 4812.205 ;
      RECT 328.26 4814.205 351.33 4825.745 ;
      RECT 328.26 4827.745 351.33 4833.515 ;
      RECT 328.26 4841.635 351.33 4842.755 ;
      RECT 328.26 4844.755 351.33 4849.365 ;
      RECT 328.26 4851.365 351.33 4860.585 ;
      RECT 328.26 4862.585 351.33 4867.195 ;
      RECT 328.26 4869.195 351.33 4870.315 ;
      RECT 328.26 4878.435 351.33 4884.205 ;
      RECT 328.26 4886.205 351.33 4897.745 ;
      RECT 328.26 4899.745 351.33 4905.515 ;
      RECT 328.26 4913.635 351.33 4914.755 ;
      RECT 328.26 4916.755 351.33 4921.365 ;
      RECT 328.26 4923.365 351.33 4932.585 ;
      RECT 328.26 4934.585 351.33 4939.195 ;
      RECT 328.26 4941.195 351.33 4942.315 ;
      RECT 328.26 4950.435 351.33 4956.205 ;
      RECT 328.26 4958.205 351.33 4969.745 ;
      RECT 328.26 4971.745 351.33 4977.515 ;
      RECT 328.26 4985.635 351.33 4986.755 ;
      RECT 328.26 4988.755 351.33 4993.365 ;
      RECT 328.26 4995.365 351.33 5004.585 ;
      RECT 328.26 5006.585 351.33 5011.195 ;
      RECT 328.26 5013.195 351.33 5014.315 ;
      RECT 328.26 5022.435 351.33 5028.205 ;
      RECT 328.26 5030.205 351.33 5041.745 ;
      RECT 328.26 5043.745 351.33 5049.515 ;
      RECT 328.26 5057.635 351.33 5058.755 ;
      RECT 328.26 5060.755 351.33 5065.365 ;
      RECT 328.26 5067.365 351.33 5076.585 ;
      RECT 328.26 5078.585 351.33 5083.195 ;
      RECT 328.26 5085.195 351.33 5086.315 ;
      RECT 328.26 5094.435 351.33 5100.205 ;
      RECT 328.26 5102.205 351.33 5113.745 ;
      RECT 328.26 5115.745 351.33 5121.515 ;
      RECT 328.26 5129.635 351.33 5130.755 ;
      RECT 328.26 5132.755 351.33 5137.365 ;
      RECT 328.26 5139.365 351.33 5148.585 ;
      RECT 328.26 5150.585 351.33 5155.195 ;
      RECT 328.26 5157.195 351.33 5158.315 ;
      RECT 328.26 5166.435 351.33 5172.205 ;
      RECT 328.26 5174.205 351.33 5185.745 ;
      RECT 328.26 5187.745 351.33 5193.515 ;
      RECT 328.26 5201.635 351.33 5202.755 ;
      RECT 328.26 5204.755 351.33 5209.365 ;
      RECT 328.26 5211.365 351.33 5220.585 ;
      RECT 328.26 5222.585 351.33 5227.195 ;
      RECT 328.26 5229.195 351.33 5230.315 ;
      RECT 328.26 5238.435 351.33 5244.205 ;
      RECT 328.26 5246.205 351.33 5257.745 ;
      RECT 328.26 5259.745 351.33 5265.515 ;
      RECT 328.26 5273.635 351.33 5274.755 ;
      RECT 328.26 5276.755 351.33 5281.365 ;
      RECT 328.26 5283.365 351.33 5292.585 ;
      RECT 328.26 5294.585 351.33 5299.195 ;
      RECT 328.26 5301.195 351.33 5302.315 ;
      RECT 328.26 5310.435 351.33 5316.205 ;
      RECT 328.26 5318.205 351.33 5329.745 ;
      RECT 328.26 5331.745 351.33 5337.515 ;
      RECT 328.26 5345.635 351.33 5346.755 ;
      RECT 328.26 5348.755 351.33 5353.365 ;
      RECT 328.26 5355.365 351.33 5364.585 ;
      RECT 328.26 5366.585 351.33 5371.195 ;
      RECT 328.26 5373.195 351.33 5374.315 ;
      RECT 328.26 5382.435 351.33 5388.205 ;
      RECT 328.26 5390.205 351.33 5401.745 ;
      RECT 328.26 5403.745 351.33 5409.515 ;
      RECT 328.26 5417.635 351.33 5418.755 ;
      RECT 328.26 5420.755 351.33 5425.365 ;
      RECT 328.26 5427.365 351.33 5436.585 ;
      RECT 328.26 5438.585 351.33 5443.195 ;
      RECT 328.26 5445.195 351.33 5446.315 ;
      RECT 328.26 5454.435 351.33 5460.205 ;
      RECT 328.26 5462.205 351.33 5473.745 ;
      RECT 328.26 5475.745 351.33 5481.515 ;
      RECT 328.26 5489.635 351.33 5490.755 ;
      RECT 328.26 5492.755 351.33 5497.365 ;
      RECT 328.26 5499.365 351.33 5508.585 ;
      RECT 328.26 5510.585 351.33 5515.195 ;
      RECT 328.26 5517.195 351.33 5518.315 ;
      RECT 328.26 5526.435 351.33 5532.205 ;
      RECT 328.26 5534.205 351.33 5545.745 ;
      RECT 328.26 5547.745 351.33 5553.515 ;
      RECT 328.26 5561.635 351.33 5562.755 ;
      RECT 328.26 5564.755 351.33 5569.365 ;
      RECT 328.26 5571.365 351.33 5580.585 ;
      RECT 328.26 5582.585 351.33 5587.195 ;
      RECT 328.26 5589.195 351.33 5590.315 ;
      RECT 328.26 5598.435 351.33 5604.205 ;
      RECT 328.26 5606.205 351.33 5617.745 ;
      RECT 328.26 5619.745 351.33 5625.515 ;
      RECT 328.26 5633.635 351.33 5634.755 ;
      RECT 328.26 5636.755 351.33 5641.365 ;
      RECT 328.26 5643.365 351.33 5652.585 ;
      RECT 328.26 5654.585 351.33 5659.195 ;
      RECT 328.26 5661.195 351.33 5662.315 ;
      RECT 328.26 5670.435 351.33 5676.205 ;
      RECT 328.26 5678.205 351.33 5689.745 ;
      RECT 328.26 5691.745 351.33 5697.515 ;
      RECT 328.26 5705.635 351.33 5706.755 ;
      RECT 328.26 5708.755 351.33 5713.365 ;
      RECT 328.26 5715.365 351.33 5724.585 ;
      RECT 328.26 5726.585 351.33 5731.195 ;
      RECT 328.26 5733.195 351.33 5734.315 ;
      RECT 328.26 5742.435 351.33 5748.205 ;
      RECT 328.26 5750.205 351.33 5761.745 ;
      RECT 328.26 5763.745 351.33 5769.515 ;
      RECT 328.26 5777.635 351.33 5778.755 ;
      RECT 328.26 5780.755 351.33 5785.365 ;
      RECT 328.26 5787.365 351.33 5796.585 ;
      RECT 328.26 5798.585 351.33 5803.195 ;
      RECT 328.26 5805.195 351.33 5806.315 ;
      RECT 328.26 5814.435 351.33 5820.205 ;
      RECT 328.26 5822.205 351.33 5833.745 ;
      RECT 328.26 5835.745 351.33 5841.515 ;
      RECT 328.26 5849.635 351.33 5850.755 ;
      RECT 328.26 5852.755 351.33 5857.365 ;
      RECT 328.26 5859.365 351.33 5868.585 ;
      RECT 328.26 5870.585 351.33 5875.195 ;
      RECT 328.26 5877.195 351.33 5878.315 ;
      RECT 328.26 5886.435 351.33 5892.205 ;
      RECT 328.26 5894.205 351.33 5905.745 ;
      RECT 328.26 5907.745 351.33 5913.515 ;
      RECT 328.26 5921.635 351.33 5922.755 ;
      RECT 328.26 5924.755 351.33 5929.365 ;
      RECT 328.26 5931.365 351.33 5940.585 ;
      RECT 328.26 5942.585 351.33 5947.195 ;
      RECT 328.26 5949.195 351.33 5950.315 ;
      RECT 328.26 5958.435 351.33 5964.205 ;
      RECT 328.26 5966.205 351.33 5977.745 ;
      RECT 328.26 5979.745 351.33 5985.515 ;
      RECT 328.26 5993.635 351.33 5994.755 ;
      RECT 328.26 5996.755 351.33 6001.365 ;
      RECT 328.26 6003.365 351.33 6012.585 ;
      RECT 328.26 6014.585 351.33 6019.195 ;
      RECT 328.26 6021.195 351.33 6022.315 ;
      RECT 328.26 6030.435 351.33 6036.205 ;
      RECT 328.26 6038.205 351.33 6049.745 ;
      RECT 328.26 6051.745 351.33 6057.515 ;
      RECT 328.26 6065.635 351.33 6066.755 ;
      RECT 328.26 6068.755 351.33 6073.365 ;
      RECT 328.26 6075.365 351.33 6084.585 ;
      RECT 328.26 6086.585 351.33 6091.195 ;
      RECT 328.26 6093.195 351.33 6094.315 ;
      RECT 328.26 6102.435 351.33 6108.205 ;
      RECT 328.26 6110.205 351.33 6121.745 ;
      RECT 328.26 6123.745 351.33 6129.515 ;
      RECT 328.26 6137.635 351.33 6138.755 ;
      RECT 328.26 6140.755 351.33 6145.365 ;
      RECT 328.26 6147.365 351.33 6156.585 ;
      RECT 328.26 6158.585 351.33 6163.195 ;
      RECT 328.26 6165.195 351.33 6166.315 ;
      RECT 328.26 6174.435 351.33 6180.205 ;
      RECT 328.26 6182.205 351.33 6193.745 ;
      RECT 328.26 6195.745 351.33 6201.515 ;
      RECT 328.26 6209.635 351.33 6210.755 ;
      RECT 328.26 6212.755 351.33 6217.365 ;
      RECT 328.26 6219.365 351.33 6228.585 ;
      RECT 328.26 6230.585 351.33 6235.195 ;
      RECT 328.26 6237.195 351.33 6238.315 ;
      RECT 328.26 6246.435 351.33 6252.205 ;
      RECT 328.26 6254.205 351.33 6265.745 ;
      RECT 328.26 6267.745 351.33 6273.515 ;
      RECT 328.26 6281.635 351.33 6282.755 ;
      RECT 328.26 6284.755 351.33 6289.365 ;
      RECT 328.26 6291.365 351.33 6300.585 ;
      RECT 328.26 6302.585 351.33 6307.195 ;
      RECT 328.26 6309.195 351.33 6310.315 ;
      RECT 328.26 6318.435 351.33 6324.205 ;
      RECT 328.26 6326.205 351.33 6337.745 ;
      RECT 328.26 6339.745 351.33 6345.515 ;
      RECT 328.26 6353.635 351.33 6354.755 ;
      RECT 328.26 6356.755 351.33 6361.365 ;
      RECT 328.26 6363.365 351.33 6372.585 ;
      RECT 328.26 6374.585 351.33 6379.195 ;
      RECT 328.26 6381.195 351.33 6382.315 ;
      RECT 328.26 6390.435 351.33 6396.205 ;
      RECT 328.26 6398.205 351.33 6409.745 ;
      RECT 328.26 6411.745 351.33 6417.515 ;
      RECT 328.26 6425.635 351.33 6426.755 ;
      RECT 328.26 6428.755 351.33 6433.365 ;
      RECT 328.26 6435.365 351.33 6444.585 ;
      RECT 328.26 6446.585 351.33 6451.195 ;
      RECT 328.26 6453.195 351.33 6454.315 ;
      RECT 328.26 6462.435 351.33 6468.205 ;
      RECT 328.26 6470.205 351.33 6481.745 ;
      RECT 328.26 6483.745 351.33 6489.515 ;
      RECT 328.26 6497.635 351.33 6498.755 ;
      RECT 328.26 6500.755 351.33 6505.365 ;
      RECT 328.26 6507.365 351.33 6516.585 ;
      RECT 328.26 6518.585 351.33 6523.195 ;
      RECT 328.26 6525.195 351.33 6526.315 ;
      RECT 328.26 6534.435 351.33 6540.205 ;
      RECT 328.26 6542.205 351.33 6553.745 ;
      RECT 328.26 6555.745 351.33 6561.515 ;
      RECT 328.26 6569.635 351.33 6570.755 ;
      RECT 328.26 6572.755 351.33 6577.365 ;
      RECT 328.26 6579.365 351.33 6588.585 ;
      RECT 328.26 6590.585 351.33 6595.195 ;
      RECT 328.26 6597.195 351.33 6598.315 ;
      RECT 328.26 6606.435 351.33 6612.205 ;
      RECT 328.26 6614.205 351.33 6625.745 ;
      RECT 328.26 6627.745 351.33 6633.515 ;
      RECT 328.26 6641.635 351.33 6642.755 ;
      RECT 328.26 6644.755 351.33 6649.365 ;
      RECT 328.26 6651.365 351.33 6660.585 ;
      RECT 328.26 6662.585 351.33 6667.195 ;
      RECT 328.26 6669.195 351.33 6670.315 ;
      RECT 328.26 6678.435 351.33 6684.205 ;
      RECT 328.26 6686.205 351.33 6697.745 ;
      RECT 328.26 6699.745 351.33 6705.515 ;
      RECT 328.26 6713.635 351.33 6714.755 ;
      RECT 328.26 6716.755 351.33 6721.365 ;
      RECT 328.26 6723.365 351.33 6732.585 ;
      RECT 328.26 6734.585 351.33 6739.195 ;
      RECT 328.26 6741.195 351.33 6742.315 ;
      RECT 328.26 6750.435 351.33 6756.205 ;
      RECT 328.26 6758.205 351.33 6769.745 ;
      RECT 328.26 6771.745 351.33 6777.515 ;
      RECT 328.26 6785.635 351.33 6786.755 ;
      RECT 328.26 6788.755 351.33 6793.365 ;
      RECT 328.26 6795.365 351.33 6804.585 ;
      RECT 328.26 6806.585 351.33 6811.195 ;
      RECT 328.26 6813.195 351.33 6814.315 ;
      RECT 328.26 6822.435 351.33 6828.205 ;
      RECT 328.26 6830.205 351.33 6841.745 ;
      RECT 328.26 6843.745 351.33 6849.515 ;
      RECT 328.26 6857.635 351.33 6858.755 ;
      RECT 328.26 6860.755 351.33 6865.365 ;
      RECT 328.26 6867.365 351.33 6876.585 ;
      RECT 328.26 6878.585 351.33 6883.195 ;
      RECT 328.26 6885.195 351.33 6886.315 ;
      RECT 328.26 6894.435 351.33 6900.205 ;
      RECT 328.26 6902.205 351.33 6913.745 ;
      RECT 328.26 6915.745 351.33 6921.515 ;
      RECT 328.26 6929.635 351.33 6930.755 ;
      RECT 328.26 6932.755 351.33 6937.365 ;
      RECT 328.26 6939.365 351.33 6948.585 ;
      RECT 328.26 6950.585 351.33 6955.195 ;
      RECT 328.26 6957.195 351.33 6958.315 ;
      RECT 328.26 6966.435 351.33 6972.205 ;
      RECT 328.26 6974.205 351.33 6985.745 ;
      RECT 328.26 6987.745 351.33 6993.515 ;
      RECT 328.26 7001.635 351.33 7002.755 ;
      RECT 328.26 7004.755 351.33 7009.365 ;
      RECT 328.26 7011.365 351.33 7020.585 ;
      RECT 328.26 7022.585 351.33 7027.195 ;
      RECT 328.26 7029.195 351.33 7030.315 ;
      RECT 328.26 7038.435 351.33 7044.205 ;
      RECT 328.26 7046.205 351.33 7057.745 ;
      RECT 328.26 7059.745 351.33 7065.515 ;
      RECT 328.26 7073.635 351.33 7074.755 ;
      RECT 328.26 7076.755 351.33 7081.365 ;
      RECT 328.26 7083.365 351.33 7092.585 ;
      RECT 328.26 7094.585 351.33 7099.195 ;
      RECT 328.26 7101.195 351.33 7102.315 ;
      RECT 328.26 7110.435 351.33 7116.205 ;
      RECT 328.26 7118.205 351.33 7129.745 ;
      RECT 328.26 7131.745 351.33 7137.515 ;
      RECT 328.26 7145.635 351.33 7146.755 ;
      RECT 328.26 7148.755 351.33 7153.365 ;
      RECT 328.26 7155.365 351.33 7164.585 ;
      RECT 328.26 7166.585 351.33 7171.195 ;
      RECT 328.26 7173.195 351.33 7174.315 ;
      RECT 328.26 7182.435 351.33 7188.205 ;
      RECT 328.26 7190.205 351.33 7201.745 ;
      RECT 328.26 7203.745 351.33 7209.515 ;
      RECT 328.26 7217.635 351.33 7218.755 ;
      RECT 328.26 7220.755 351.33 7225.365 ;
      RECT 328.26 7227.365 351.33 7236.585 ;
      RECT 328.26 7238.585 351.33 7243.195 ;
      RECT 328.26 7245.195 351.33 7246.315 ;
      RECT 328.26 7254.435 351.33 7260.205 ;
      RECT 328.26 7262.205 351.33 7273.745 ;
      RECT 328.26 7275.745 351.33 7281.515 ;
      RECT 328.26 7289.635 351.33 7290.755 ;
      RECT 328.26 7292.755 351.33 7297.365 ;
      RECT 328.26 7299.365 351.33 7308.585 ;
      RECT 328.26 7310.585 351.33 7315.195 ;
      RECT 328.26 7317.195 351.33 7318.315 ;
      RECT 328.26 7326.435 351.33 7332.205 ;
      RECT 328.26 7334.205 351.33 7345.745 ;
      RECT 328.26 7347.745 351.33 7353.515 ;
      RECT 328.26 7361.635 351.33 7362.755 ;
      RECT 328.26 7364.755 351.33 7369.365 ;
      RECT 328.26 7371.365 351.33 7380.585 ;
      RECT 328.26 7382.585 351.33 7387.195 ;
      RECT 328.26 7389.195 351.33 7390.315 ;
      RECT 328.26 7398.435 351.33 7404.205 ;
      RECT 328.26 7406.205 351.33 7417.745 ;
      RECT 328.26 7419.745 351.33 7425.515 ;
      RECT 328.26 7433.635 351.33 7434.755 ;
      RECT 328.26 7436.755 351.33 7441.365 ;
      RECT 328.26 7443.365 351.33 7452.585 ;
      RECT 328.26 7454.585 351.33 7459.195 ;
      RECT 328.26 7461.195 351.33 7462.315 ;
      RECT 328.26 7470.435 351.33 7476.205 ;
      RECT 328.26 7478.205 351.33 7489.745 ;
      RECT 328.26 7491.745 351.33 7497.515 ;
      RECT 328.26 7505.635 351.33 7506.755 ;
      RECT 328.26 7508.755 351.33 7513.365 ;
      RECT 328.26 7515.365 351.33 7524.585 ;
      RECT 328.26 7526.585 351.33 7531.195 ;
      RECT 328.26 7533.195 351.33 7534.315 ;
      RECT 328.26 7542.435 351.33 7548.205 ;
      RECT 328.26 7550.205 351.33 7561.745 ;
      RECT 328.26 7563.745 351.33 7569.515 ;
      RECT 328.26 7577.635 351.33 7578.755 ;
      RECT 328.26 7580.755 351.33 7585.365 ;
      RECT 328.26 7587.365 351.33 7596.585 ;
      RECT 328.26 7598.585 351.33 7603.195 ;
      RECT 328.26 7605.195 351.33 7606.315 ;
      RECT 328.26 7614.435 351.33 7620.205 ;
      RECT 328.26 7622.205 351.33 7633.745 ;
      RECT 328.26 7635.745 351.33 7641.515 ;
      RECT 328.26 7649.635 351.33 7650.755 ;
      RECT 328.26 7652.755 351.33 7657.365 ;
      RECT 328.26 7659.365 351.33 7668.585 ;
      RECT 328.26 7670.585 351.33 7675.195 ;
      RECT 328.26 7677.195 351.33 7678.315 ;
      RECT 328.26 7686.435 351.33 7692.205 ;
      RECT 328.26 7694.205 351.33 7705.745 ;
      RECT 328.26 7707.745 351.33 7713.515 ;
      RECT 328.26 7721.635 351.33 7722.755 ;
      RECT 328.26 7724.755 351.33 7729.365 ;
      RECT 328.26 7731.365 351.33 7740.585 ;
      RECT 328.26 7742.585 351.33 7747.195 ;
      RECT 328.26 7749.195 351.33 7750.315 ;
      RECT 328.26 7758.435 351.33 7764.205 ;
      RECT 328.26 7766.205 351.33 7777.745 ;
      RECT 328.26 7779.745 351.33 7785.515 ;
      RECT 328.26 7793.635 351.33 7794.755 ;
      RECT 328.26 7796.755 351.33 7801.365 ;
      RECT 328.26 7803.365 351.33 7812.585 ;
      RECT 328.26 7814.585 351.33 7819.195 ;
      RECT 328.26 7821.195 351.33 7822.315 ;
      RECT 328.26 7830.435 351.33 7836.205 ;
      RECT 328.26 7838.205 351.33 7849.745 ;
      RECT 328.26 7851.745 351.33 7857.515 ;
      RECT 328.26 7865.635 351.33 7866.755 ;
      RECT 328.26 7868.755 351.33 7873.365 ;
      RECT 328.26 7875.365 351.33 7884.585 ;
      RECT 328.26 7886.585 351.33 7891.195 ;
      RECT 328.26 7893.195 351.33 7894.315 ;
      RECT 328.26 7902.435 351.33 7908.205 ;
      RECT 328.26 7910.205 351.33 7921.745 ;
      RECT 328.26 7923.745 351.33 7929.515 ;
      RECT 328.26 7937.635 351.33 7938.755 ;
      RECT 328.26 7940.755 351.33 7945.365 ;
      RECT 328.26 7947.365 351.33 7956.585 ;
      RECT 328.26 7958.585 351.33 7963.195 ;
      RECT 328.26 7965.195 351.33 7966.315 ;
      RECT 328.26 7974.435 351.33 7980.205 ;
      RECT 328.26 7982.205 351.33 7993.745 ;
      RECT 328.26 7995.745 351.33 8001.515 ;
      RECT 328.26 8009.635 351.33 8010.755 ;
      RECT 328.26 8012.755 351.33 8017.365 ;
      RECT 328.26 8019.365 351.33 8028.585 ;
      RECT 328.26 8030.585 351.33 8035.195 ;
      RECT 328.26 8037.195 351.33 8038.315 ;
      RECT 328.26 8046.435 351.33 8052.205 ;
      RECT 328.26 8054.205 351.33 8065.745 ;
      RECT 328.26 8067.745 351.33 8073.515 ;
      RECT 328.26 8081.635 351.33 8082.755 ;
      RECT 328.26 8084.755 351.33 8089.365 ;
      RECT 328.26 8091.365 351.33 8100.585 ;
      RECT 328.26 8102.585 351.33 8107.195 ;
      RECT 328.26 8109.195 351.33 8110.315 ;
      RECT 328.26 8118.435 351.33 8124.205 ;
      RECT 328.26 8126.205 351.33 8137.745 ;
      RECT 328.26 8139.745 351.33 8145.515 ;
      RECT 328.26 8153.635 351.33 8154.755 ;
      RECT 328.26 8156.755 351.33 8161.365 ;
      RECT 328.26 8163.365 351.33 8172.585 ;
      RECT 328.26 8174.585 351.33 8179.195 ;
      RECT 328.26 8181.195 351.33 8182.315 ;
      RECT 328.26 8190.435 351.33 8196.205 ;
      RECT 328.26 8198.205 351.33 8209.745 ;
      RECT 328.26 8211.745 351.33 8217.515 ;
      RECT 328.26 8225.635 351.33 8226.755 ;
      RECT 328.26 8228.755 351.33 8233.365 ;
      RECT 328.26 8235.365 351.33 8244.585 ;
      RECT 328.26 8246.585 351.33 8251.195 ;
      RECT 328.26 8253.195 351.33 8254.315 ;
      RECT 328.26 8262.435 351.33 8268.205 ;
      RECT 328.26 8270.205 351.33 8281.745 ;
      RECT 328.26 8283.745 351.33 8289.515 ;
      RECT 328.26 8297.635 351.33 8298.755 ;
      RECT 328.26 8300.755 351.33 8305.365 ;
      RECT 328.26 8307.365 351.33 8316.585 ;
      RECT 328.26 8318.585 351.33 8323.195 ;
      RECT 328.26 8325.195 351.33 8326.315 ;
      RECT 328.26 8334.435 351.33 8340.205 ;
      RECT 328.26 8342.205 351.33 8353.745 ;
      RECT 328.26 8355.745 351.33 8361.515 ;
      RECT 328.26 8369.635 351.33 8370.755 ;
      RECT 328.26 8372.755 351.33 8377.365 ;
      RECT 328.26 8379.365 351.33 8388.585 ;
      RECT 328.26 8390.585 351.33 8395.195 ;
      RECT 328.26 8397.195 351.33 8398.315 ;
      RECT 328.26 8406.435 351.33 8412.205 ;
      RECT 328.26 8414.205 351.33 8425.745 ;
      RECT 328.26 8427.745 351.33 8433.515 ;
      RECT 328.26 8441.635 351.33 8442.755 ;
      RECT 328.26 8444.755 351.33 8449.365 ;
      RECT 328.26 8451.365 351.33 8460.585 ;
      RECT 328.26 8462.585 351.33 8467.195 ;
      RECT 328.26 8469.195 351.33 8470.315 ;
      RECT 328.26 8478.435 351.33 8484.205 ;
      RECT 328.26 8486.205 351.33 8497.745 ;
      RECT 328.26 8499.745 351.33 8505.515 ;
      RECT 328.26 8513.635 351.33 8514.755 ;
      RECT 328.26 8516.755 351.33 8521.365 ;
      RECT 328.26 8523.365 351.33 8532.585 ;
      RECT 328.26 8534.585 351.33 8539.195 ;
      RECT 328.26 8541.195 351.33 8542.315 ;
      RECT 328.26 8550.435 351.33 8556.205 ;
      RECT 328.26 8558.205 351.33 8569.745 ;
      RECT 328.26 8571.745 351.33 8577.515 ;
      RECT 328.26 8585.635 351.33 8586.755 ;
      RECT 328.26 8588.755 351.33 8593.365 ;
      RECT 328.26 8595.365 351.33 8599.975 ;
    LAYER TOP_M SPACING 0.46 ;
      RECT 18488.23 551.045 18490.46 551.585 ;
      RECT 18488.23 187.44 18488.73 551.585 ;
      RECT 18488.23 547.925 18490.46 548.465 ;
      RECT 18488.23 541.315 18490.46 541.855 ;
      RECT 18488.23 523.41 18490.46 535.245 ;
      RECT 18488.23 514.995 18490.46 520.83 ;
      RECT 18488.23 510.175 18490.46 511.535 ;
      RECT 18488.23 507.175 18490.46 507.715 ;
      RECT 18488.23 324.005 18490.46 504.715 ;
      RECT 18488.23 307.005 18490.46 308.515 ;
      RECT 18488.23 290.005 18490.46 291.515 ;
      RECT 18488.23 228.005 18490.46 229.515 ;
      RECT 18488.23 211.005 18490.46 212.515 ;
      RECT 18488.23 194.005 18490.46 195.515 ;
      RECT 18488.23 187.44 18490.46 190.545 ;
      RECT 18488.23 586.245 18490.46 590.345 ;
      RECT 18488.23 553.605 18488.73 590.345 ;
      RECT 18488.23 578.475 18490.46 579.015 ;
      RECT 18488.23 564.935 18490.46 565.475 ;
      RECT 18488.23 553.605 18490.46 557.705 ;
      RECT 18488.23 623.045 18490.46 623.585 ;
      RECT 18488.23 592.365 18488.73 623.585 ;
      RECT 18488.23 619.925 18490.46 620.465 ;
      RECT 18488.23 613.315 18490.46 613.855 ;
      RECT 18488.23 602.095 18490.46 602.635 ;
      RECT 18488.23 595.485 18490.46 596.025 ;
      RECT 18488.23 592.365 18490.46 592.905 ;
      RECT 18488.23 658.245 18490.46 662.345 ;
      RECT 18488.23 625.605 18488.73 662.345 ;
      RECT 18488.23 650.475 18490.46 651.015 ;
      RECT 18488.23 636.935 18490.46 637.475 ;
      RECT 18488.23 625.605 18490.46 629.705 ;
      RECT 18488.23 695.045 18490.46 695.585 ;
      RECT 18488.23 664.365 18488.73 695.585 ;
      RECT 18488.23 691.925 18490.46 692.465 ;
      RECT 18488.23 685.315 18490.46 685.855 ;
      RECT 18488.23 674.095 18490.46 674.635 ;
      RECT 18488.23 667.485 18490.46 668.025 ;
      RECT 18488.23 664.365 18490.46 664.905 ;
      RECT 18488.23 730.245 18490.46 734.345 ;
      RECT 18488.23 697.605 18488.73 734.345 ;
      RECT 18488.23 722.475 18490.46 723.015 ;
      RECT 18488.23 708.935 18490.46 709.475 ;
      RECT 18488.23 697.605 18490.46 701.705 ;
      RECT 18488.23 767.045 18490.46 767.585 ;
      RECT 18488.23 736.365 18488.73 767.585 ;
      RECT 18488.23 763.925 18490.46 764.465 ;
      RECT 18488.23 757.315 18490.46 757.855 ;
      RECT 18488.23 746.095 18490.46 746.635 ;
      RECT 18488.23 739.485 18490.46 740.025 ;
      RECT 18488.23 736.365 18490.46 736.905 ;
      RECT 18488.23 802.245 18490.46 806.345 ;
      RECT 18488.23 769.605 18488.73 806.345 ;
      RECT 18488.23 794.475 18490.46 795.015 ;
      RECT 18488.23 780.935 18490.46 781.475 ;
      RECT 18488.23 769.605 18490.46 773.705 ;
      RECT 18488.23 839.045 18490.46 839.585 ;
      RECT 18488.23 808.365 18488.73 839.585 ;
      RECT 18488.23 835.925 18490.46 836.465 ;
      RECT 18488.23 829.315 18490.46 829.855 ;
      RECT 18488.23 818.095 18490.46 818.635 ;
      RECT 18488.23 811.485 18490.46 812.025 ;
      RECT 18488.23 808.365 18490.46 808.905 ;
      RECT 18488.23 874.245 18490.46 878.345 ;
      RECT 18488.23 841.605 18488.73 878.345 ;
      RECT 18488.23 866.475 18490.46 867.015 ;
      RECT 18488.23 852.935 18490.46 853.475 ;
      RECT 18488.23 841.605 18490.46 845.705 ;
      RECT 18488.23 911.045 18490.46 911.585 ;
      RECT 18488.23 880.365 18488.73 911.585 ;
      RECT 18488.23 907.925 18490.46 908.465 ;
      RECT 18488.23 901.315 18490.46 901.855 ;
      RECT 18488.23 890.095 18490.46 890.635 ;
      RECT 18488.23 883.485 18490.46 884.025 ;
      RECT 18488.23 880.365 18490.46 880.905 ;
      RECT 18488.23 946.245 18490.46 950.345 ;
      RECT 18488.23 913.605 18488.73 950.345 ;
      RECT 18488.23 938.475 18490.46 939.015 ;
      RECT 18488.23 924.935 18490.46 925.475 ;
      RECT 18488.23 913.605 18490.46 917.705 ;
      RECT 18488.23 983.045 18490.46 983.585 ;
      RECT 18488.23 952.365 18488.73 983.585 ;
      RECT 18488.23 979.925 18490.46 980.465 ;
      RECT 18488.23 973.315 18490.46 973.855 ;
      RECT 18488.23 962.095 18490.46 962.635 ;
      RECT 18488.23 955.485 18490.46 956.025 ;
      RECT 18488.23 952.365 18490.46 952.905 ;
      RECT 18488.23 1018.245 18490.46 1022.345 ;
      RECT 18488.23 985.605 18488.73 1022.345 ;
      RECT 18488.23 1010.475 18490.46 1011.015 ;
      RECT 18488.23 996.935 18490.46 997.475 ;
      RECT 18488.23 985.605 18490.46 989.705 ;
      RECT 18488.23 1055.045 18490.46 1055.585 ;
      RECT 18488.23 1024.365 18488.73 1055.585 ;
      RECT 18488.23 1051.925 18490.46 1052.465 ;
      RECT 18488.23 1045.315 18490.46 1045.855 ;
      RECT 18488.23 1034.095 18490.46 1034.635 ;
      RECT 18488.23 1027.485 18490.46 1028.025 ;
      RECT 18488.23 1024.365 18490.46 1024.905 ;
      RECT 18488.23 1090.245 18490.46 1094.345 ;
      RECT 18488.23 1057.605 18488.73 1094.345 ;
      RECT 18488.23 1082.475 18490.46 1083.015 ;
      RECT 18488.23 1068.935 18490.46 1069.475 ;
      RECT 18488.23 1057.605 18490.46 1061.705 ;
      RECT 18488.23 1127.045 18490.46 1127.585 ;
      RECT 18488.23 1096.365 18488.73 1127.585 ;
      RECT 18488.23 1123.925 18490.46 1124.465 ;
      RECT 18488.23 1117.315 18490.46 1117.855 ;
      RECT 18488.23 1106.095 18490.46 1106.635 ;
      RECT 18488.23 1099.485 18490.46 1100.025 ;
      RECT 18488.23 1096.365 18490.46 1096.905 ;
      RECT 18488.23 1162.245 18490.46 1166.345 ;
      RECT 18488.23 1129.605 18488.73 1166.345 ;
      RECT 18488.23 1154.475 18490.46 1155.015 ;
      RECT 18488.23 1140.935 18490.46 1141.475 ;
      RECT 18488.23 1129.605 18490.46 1133.705 ;
      RECT 18488.23 1199.045 18490.46 1199.585 ;
      RECT 18488.23 1168.365 18488.73 1199.585 ;
      RECT 18488.23 1195.925 18490.46 1196.465 ;
      RECT 18488.23 1189.315 18490.46 1189.855 ;
      RECT 18488.23 1178.095 18490.46 1178.635 ;
      RECT 18488.23 1171.485 18490.46 1172.025 ;
      RECT 18488.23 1168.365 18490.46 1168.905 ;
      RECT 18488.23 1234.245 18490.46 1238.345 ;
      RECT 18488.23 1201.605 18488.73 1238.345 ;
      RECT 18488.23 1226.475 18490.46 1227.015 ;
      RECT 18488.23 1212.935 18490.46 1213.475 ;
      RECT 18488.23 1201.605 18490.46 1205.705 ;
      RECT 18488.23 1271.045 18490.46 1271.585 ;
      RECT 18488.23 1240.365 18488.73 1271.585 ;
      RECT 18488.23 1267.925 18490.46 1268.465 ;
      RECT 18488.23 1261.315 18490.46 1261.855 ;
      RECT 18488.23 1250.095 18490.46 1250.635 ;
      RECT 18488.23 1243.485 18490.46 1244.025 ;
      RECT 18488.23 1240.365 18490.46 1240.905 ;
      RECT 18488.23 1306.245 18490.46 1310.345 ;
      RECT 18488.23 1273.605 18488.73 1310.345 ;
      RECT 18488.23 1298.475 18490.46 1299.015 ;
      RECT 18488.23 1284.935 18490.46 1285.475 ;
      RECT 18488.23 1273.605 18490.46 1277.705 ;
      RECT 18488.23 1343.045 18490.46 1343.585 ;
      RECT 18488.23 1312.365 18488.73 1343.585 ;
      RECT 18488.23 1339.925 18490.46 1340.465 ;
      RECT 18488.23 1333.315 18490.46 1333.855 ;
      RECT 18488.23 1322.095 18490.46 1322.635 ;
      RECT 18488.23 1315.485 18490.46 1316.025 ;
      RECT 18488.23 1312.365 18490.46 1312.905 ;
      RECT 18488.23 1378.245 18490.46 1382.345 ;
      RECT 18488.23 1345.605 18488.73 1382.345 ;
      RECT 18488.23 1370.475 18490.46 1371.015 ;
      RECT 18488.23 1356.935 18490.46 1357.475 ;
      RECT 18488.23 1345.605 18490.46 1349.705 ;
      RECT 18488.23 1415.045 18490.46 1415.585 ;
      RECT 18488.23 1384.365 18488.73 1415.585 ;
      RECT 18488.23 1411.925 18490.46 1412.465 ;
      RECT 18488.23 1405.315 18490.46 1405.855 ;
      RECT 18488.23 1394.095 18490.46 1394.635 ;
      RECT 18488.23 1387.485 18490.46 1388.025 ;
      RECT 18488.23 1384.365 18490.46 1384.905 ;
      RECT 18488.23 1450.245 18490.46 1454.345 ;
      RECT 18488.23 1417.605 18488.73 1454.345 ;
      RECT 18488.23 1442.475 18490.46 1443.015 ;
      RECT 18488.23 1428.935 18490.46 1429.475 ;
      RECT 18488.23 1417.605 18490.46 1421.705 ;
      RECT 18488.23 1487.045 18490.46 1487.585 ;
      RECT 18488.23 1456.365 18488.73 1487.585 ;
      RECT 18488.23 1483.925 18490.46 1484.465 ;
      RECT 18488.23 1477.315 18490.46 1477.855 ;
      RECT 18488.23 1466.095 18490.46 1466.635 ;
      RECT 18488.23 1459.485 18490.46 1460.025 ;
      RECT 18488.23 1456.365 18490.46 1456.905 ;
      RECT 18488.23 1522.245 18490.46 1526.345 ;
      RECT 18488.23 1489.605 18488.73 1526.345 ;
      RECT 18488.23 1514.475 18490.46 1515.015 ;
      RECT 18488.23 1500.935 18490.46 1501.475 ;
      RECT 18488.23 1489.605 18490.46 1493.705 ;
      RECT 18488.23 1559.045 18490.46 1559.585 ;
      RECT 18488.23 1528.365 18488.73 1559.585 ;
      RECT 18488.23 1555.925 18490.46 1556.465 ;
      RECT 18488.23 1549.315 18490.46 1549.855 ;
      RECT 18488.23 1538.095 18490.46 1538.635 ;
      RECT 18488.23 1531.485 18490.46 1532.025 ;
      RECT 18488.23 1528.365 18490.46 1528.905 ;
      RECT 2313.83 8584.365 18488.73 8610.835 ;
      RECT 2313.83 189.17 18488.23 8610.835 ;
      RECT 18375.79 187.44 18488.23 8610.835 ;
      RECT 2313.83 8545.605 18488.73 8582.345 ;
      RECT 2313.83 8512.365 18488.73 8543.585 ;
      RECT 2313.83 8473.605 18488.73 8510.345 ;
      RECT 2313.83 8440.365 18488.73 8471.585 ;
      RECT 2313.83 8401.605 18488.73 8438.345 ;
      RECT 2313.83 8368.365 18488.73 8399.585 ;
      RECT 2313.83 8329.605 18488.73 8366.345 ;
      RECT 2313.83 8296.365 18488.73 8327.585 ;
      RECT 2313.83 8257.605 18488.73 8294.345 ;
      RECT 2313.83 8224.365 18488.73 8255.585 ;
      RECT 2313.83 8185.605 18488.73 8222.345 ;
      RECT 2313.83 8152.365 18488.73 8183.585 ;
      RECT 2313.83 8113.605 18488.73 8150.345 ;
      RECT 2313.83 8080.365 18488.73 8111.585 ;
      RECT 2313.83 8041.605 18488.73 8078.345 ;
      RECT 2313.83 8008.365 18488.73 8039.585 ;
      RECT 2313.83 7969.605 18488.73 8006.345 ;
      RECT 2313.83 7936.365 18488.73 7967.585 ;
      RECT 2313.83 7897.605 18488.73 7934.345 ;
      RECT 2313.83 7864.365 18488.73 7895.585 ;
      RECT 2313.83 7825.605 18488.73 7862.345 ;
      RECT 2313.83 7792.365 18488.73 7823.585 ;
      RECT 2313.83 7753.605 18488.73 7790.345 ;
      RECT 2313.83 7720.365 18488.73 7751.585 ;
      RECT 2313.83 7681.605 18488.73 7718.345 ;
      RECT 2313.83 7648.365 18488.73 7679.585 ;
      RECT 2313.83 7609.605 18488.73 7646.345 ;
      RECT 2313.83 7576.365 18488.73 7607.585 ;
      RECT 2313.83 7537.605 18488.73 7574.345 ;
      RECT 2313.83 7504.365 18488.73 7535.585 ;
      RECT 2313.83 7465.605 18488.73 7502.345 ;
      RECT 2313.83 7432.365 18488.73 7463.585 ;
      RECT 2313.83 7393.605 18488.73 7430.345 ;
      RECT 2313.83 7360.365 18488.73 7391.585 ;
      RECT 2313.83 7321.605 18488.73 7358.345 ;
      RECT 2313.83 7288.365 18488.73 7319.585 ;
      RECT 2313.83 7249.605 18488.73 7286.345 ;
      RECT 2313.83 7216.365 18488.73 7247.585 ;
      RECT 2313.83 7177.605 18488.73 7214.345 ;
      RECT 2313.83 7144.365 18488.73 7175.585 ;
      RECT 2313.83 7105.605 18488.73 7142.345 ;
      RECT 2313.83 7072.365 18488.73 7103.585 ;
      RECT 2313.83 7033.605 18488.73 7070.345 ;
      RECT 2313.83 7000.365 18488.73 7031.585 ;
      RECT 2313.83 6961.605 18488.73 6998.345 ;
      RECT 2313.83 6928.365 18488.73 6959.585 ;
      RECT 2313.83 6889.605 18488.73 6926.345 ;
      RECT 2313.83 6856.365 18488.73 6887.585 ;
      RECT 2313.83 6817.605 18488.73 6854.345 ;
      RECT 2313.83 6784.365 18488.73 6815.585 ;
      RECT 2313.83 6745.605 18488.73 6782.345 ;
      RECT 2313.83 6712.365 18488.73 6743.585 ;
      RECT 2313.83 6673.605 18488.73 6710.345 ;
      RECT 2313.83 6640.365 18488.73 6671.585 ;
      RECT 2313.83 6601.605 18488.73 6638.345 ;
      RECT 2313.83 6568.365 18488.73 6599.585 ;
      RECT 2313.83 6529.605 18488.73 6566.345 ;
      RECT 2313.83 6496.365 18488.73 6527.585 ;
      RECT 2313.83 6457.605 18488.73 6494.345 ;
      RECT 2313.83 6424.365 18488.73 6455.585 ;
      RECT 2313.83 6385.605 18488.73 6422.345 ;
      RECT 2313.83 6352.365 18488.73 6383.585 ;
      RECT 2313.83 6313.605 18488.73 6350.345 ;
      RECT 2313.83 6280.365 18488.73 6311.585 ;
      RECT 2313.83 6241.605 18488.73 6278.345 ;
      RECT 2313.83 6208.365 18488.73 6239.585 ;
      RECT 2313.83 6169.605 18488.73 6206.345 ;
      RECT 2313.83 6136.365 18488.73 6167.585 ;
      RECT 2313.83 6097.605 18488.73 6134.345 ;
      RECT 2313.83 6064.365 18488.73 6095.585 ;
      RECT 2313.83 6025.605 18488.73 6062.345 ;
      RECT 2313.83 5992.365 18488.73 6023.585 ;
      RECT 2313.83 5953.605 18488.73 5990.345 ;
      RECT 2313.83 5920.365 18488.73 5951.585 ;
      RECT 2313.83 5881.605 18488.73 5918.345 ;
      RECT 2313.83 5848.365 18488.73 5879.585 ;
      RECT 2313.83 5809.605 18488.73 5846.345 ;
      RECT 2313.83 5776.365 18488.73 5807.585 ;
      RECT 2313.83 5737.605 18488.73 5774.345 ;
      RECT 2313.83 5704.365 18488.73 5735.585 ;
      RECT 2313.83 5665.605 18488.73 5702.345 ;
      RECT 2313.83 5632.365 18488.73 5663.585 ;
      RECT 2313.83 5593.605 18488.73 5630.345 ;
      RECT 2313.83 5560.365 18488.73 5591.585 ;
      RECT 2313.83 5521.605 18488.73 5558.345 ;
      RECT 2313.83 5488.365 18488.73 5519.585 ;
      RECT 2313.83 5449.605 18488.73 5486.345 ;
      RECT 2313.83 5416.365 18488.73 5447.585 ;
      RECT 2313.83 5377.605 18488.73 5414.345 ;
      RECT 2313.83 5344.365 18488.73 5375.585 ;
      RECT 2313.83 5305.605 18488.73 5342.345 ;
      RECT 2313.83 5272.365 18488.73 5303.585 ;
      RECT 2313.83 5233.605 18488.73 5270.345 ;
      RECT 2313.83 5200.365 18488.73 5231.585 ;
      RECT 2313.83 5161.605 18488.73 5198.345 ;
      RECT 2313.83 5128.365 18488.73 5159.585 ;
      RECT 2313.83 5089.605 18488.73 5126.345 ;
      RECT 2313.83 5056.365 18488.73 5087.585 ;
      RECT 2313.83 5017.605 18488.73 5054.345 ;
      RECT 2313.83 4984.365 18488.73 5015.585 ;
      RECT 2313.83 4945.605 18488.73 4982.345 ;
      RECT 2313.83 4912.365 18488.73 4943.585 ;
      RECT 2313.83 4873.605 18488.73 4910.345 ;
      RECT 2313.83 4840.365 18488.73 4871.585 ;
      RECT 2313.83 4801.605 18488.73 4838.345 ;
      RECT 2313.83 4768.365 18488.73 4799.585 ;
      RECT 2313.83 4729.605 18488.73 4766.345 ;
      RECT 2313.83 4696.365 18488.73 4727.585 ;
      RECT 2313.83 4657.605 18488.73 4694.345 ;
      RECT 2313.83 4624.365 18488.73 4655.585 ;
      RECT 2313.83 4585.605 18488.73 4622.345 ;
      RECT 2313.83 4552.365 18488.73 4583.585 ;
      RECT 2313.83 4513.605 18488.73 4550.345 ;
      RECT 2313.83 4480.365 18488.73 4511.585 ;
      RECT 2313.83 4441.605 18488.73 4478.345 ;
      RECT 2313.83 4408.365 18488.73 4439.585 ;
      RECT 2313.83 4369.605 18488.73 4406.345 ;
      RECT 2313.83 4336.365 18488.73 4367.585 ;
      RECT 2313.83 4297.605 18488.73 4334.345 ;
      RECT 2313.83 4264.365 18488.73 4295.585 ;
      RECT 2313.83 4225.605 18488.73 4262.345 ;
      RECT 2313.83 4192.365 18488.73 4223.585 ;
      RECT 2313.83 4153.605 18488.73 4190.345 ;
      RECT 2313.83 4120.365 18488.73 4151.585 ;
      RECT 2313.83 4081.605 18488.73 4118.345 ;
      RECT 2313.83 4048.365 18488.73 4079.585 ;
      RECT 2313.83 4009.605 18488.73 4046.345 ;
      RECT 2313.83 3976.365 18488.73 4007.585 ;
      RECT 2313.83 3937.605 18488.73 3974.345 ;
      RECT 2313.83 3904.365 18488.73 3935.585 ;
      RECT 2313.83 3865.605 18488.73 3902.345 ;
      RECT 2313.83 3832.365 18488.73 3863.585 ;
      RECT 2313.83 3793.605 18488.73 3830.345 ;
      RECT 2313.83 3760.365 18488.73 3791.585 ;
      RECT 2313.83 3721.605 18488.73 3758.345 ;
      RECT 2313.83 3688.365 18488.73 3719.585 ;
      RECT 2313.83 3649.605 18488.73 3686.345 ;
      RECT 2313.83 3616.365 18488.73 3647.585 ;
      RECT 2313.83 3577.605 18488.73 3614.345 ;
      RECT 2313.83 3544.365 18488.73 3575.585 ;
      RECT 2313.83 3505.605 18488.73 3542.345 ;
      RECT 2313.83 3472.365 18488.73 3503.585 ;
      RECT 2313.83 3433.605 18488.73 3470.345 ;
      RECT 2313.83 3400.365 18488.73 3431.585 ;
      RECT 2313.83 3361.605 18488.73 3398.345 ;
      RECT 2313.83 3328.365 18488.73 3359.585 ;
      RECT 2313.83 3289.605 18488.73 3326.345 ;
      RECT 2313.83 3256.365 18488.73 3287.585 ;
      RECT 2313.83 3217.605 18488.73 3254.345 ;
      RECT 2313.83 3184.365 18488.73 3215.585 ;
      RECT 2313.83 3145.605 18488.73 3182.345 ;
      RECT 2313.83 3112.365 18488.73 3143.585 ;
      RECT 2313.83 3073.605 18488.73 3110.345 ;
      RECT 2313.83 3040.365 18488.73 3071.585 ;
      RECT 2313.83 3001.605 18488.73 3038.345 ;
      RECT 2313.83 2968.365 18488.73 2999.585 ;
      RECT 2313.83 2929.605 18488.73 2966.345 ;
      RECT 2313.83 2896.365 18488.73 2927.585 ;
      RECT 2313.83 2857.605 18488.73 2894.345 ;
      RECT 2313.83 2824.365 18488.73 2855.585 ;
      RECT 2313.83 2785.605 18488.73 2822.345 ;
      RECT 2313.83 2752.365 18488.73 2783.585 ;
      RECT 2313.83 2713.605 18488.73 2750.345 ;
      RECT 2313.83 2680.365 18488.73 2711.585 ;
      RECT 2313.83 2641.605 18488.73 2678.345 ;
      RECT 2313.83 2608.365 18488.73 2639.585 ;
      RECT 2313.83 2569.605 18488.73 2606.345 ;
      RECT 2313.83 2536.365 18488.73 2567.585 ;
      RECT 2313.83 2497.605 18488.73 2534.345 ;
      RECT 2313.83 2464.365 18488.73 2495.585 ;
      RECT 2313.83 2425.605 18488.73 2462.345 ;
      RECT 2313.83 2392.365 18488.73 2423.585 ;
      RECT 2313.83 2353.605 18488.73 2390.345 ;
      RECT 2313.83 2320.365 18488.73 2351.585 ;
      RECT 2313.83 2281.605 18488.73 2318.345 ;
      RECT 2313.83 2248.365 18488.73 2279.585 ;
      RECT 2313.83 2209.605 18488.73 2246.345 ;
      RECT 2313.83 2176.365 18488.73 2207.585 ;
      RECT 2313.83 2137.605 18488.73 2174.345 ;
      RECT 2313.83 2104.365 18488.73 2135.585 ;
      RECT 2313.83 2065.605 18488.73 2102.345 ;
      RECT 2313.83 2032.365 18488.73 2063.585 ;
      RECT 2313.83 1993.605 18488.73 2030.345 ;
      RECT 2313.83 1960.365 18488.73 1991.585 ;
      RECT 2313.83 1921.605 18488.73 1958.345 ;
      RECT 2313.83 1888.365 18488.73 1919.585 ;
      RECT 2313.83 1849.605 18488.73 1886.345 ;
      RECT 2313.83 1816.365 18488.73 1847.585 ;
      RECT 2313.83 1777.605 18488.73 1814.345 ;
      RECT 2313.83 1744.365 18488.73 1775.585 ;
      RECT 2313.83 1705.605 18488.73 1742.345 ;
      RECT 2313.83 1672.365 18488.73 1703.585 ;
      RECT 2313.83 1633.605 18488.73 1670.345 ;
      RECT 2313.83 1600.365 18488.73 1631.585 ;
      RECT 2313.83 1561.605 18488.73 1598.345 ;
      RECT 18358.81 187.44 18361.33 8610.835 ;
      RECT 18343.29 187.44 18344.35 8610.835 ;
      RECT 18312.77 187.44 18313.83 8610.835 ;
      RECT 18295.79 187.44 18298.31 8610.835 ;
      RECT 18278.81 187.44 18281.33 8610.835 ;
      RECT 18263.29 187.44 18264.35 8610.835 ;
      RECT 18232.77 187.44 18233.83 8610.835 ;
      RECT 18215.79 187.44 18218.31 8610.835 ;
      RECT 18198.81 187.44 18201.33 8610.835 ;
      RECT 18183.29 187.44 18184.35 8610.835 ;
      RECT 18152.77 187.44 18153.83 8610.835 ;
      RECT 18135.79 187.44 18138.31 8610.835 ;
      RECT 18118.81 187.44 18121.33 8610.835 ;
      RECT 18103.29 187.44 18104.35 8610.835 ;
      RECT 18072.77 187.44 18073.83 8610.835 ;
      RECT 18055.79 187.44 18058.31 8610.835 ;
      RECT 18038.81 187.44 18041.33 8610.835 ;
      RECT 18023.29 187.44 18024.35 8610.835 ;
      RECT 17992.77 187.44 17993.83 8610.835 ;
      RECT 17975.79 187.44 17978.31 8610.835 ;
      RECT 17958.81 187.44 17961.33 8610.835 ;
      RECT 17943.29 187.44 17944.35 8610.835 ;
      RECT 17912.77 187.44 17913.83 8610.835 ;
      RECT 17895.79 187.44 17898.31 8610.835 ;
      RECT 17878.81 187.44 17881.33 8610.835 ;
      RECT 17863.29 187.44 17864.35 8610.835 ;
      RECT 17832.77 187.44 17833.83 8610.835 ;
      RECT 17815.79 187.44 17818.31 8610.835 ;
      RECT 17798.81 187.44 17801.33 8610.835 ;
      RECT 17783.29 187.44 17784.35 8610.835 ;
      RECT 17752.77 187.44 17753.83 8610.835 ;
      RECT 17735.79 187.44 17738.31 8610.835 ;
      RECT 17718.81 187.44 17721.33 8610.835 ;
      RECT 17703.29 187.44 17704.35 8610.835 ;
      RECT 17672.77 187.44 17673.83 8610.835 ;
      RECT 17655.79 187.44 17658.31 8610.835 ;
      RECT 17638.81 187.44 17641.33 8610.835 ;
      RECT 17623.29 187.44 17624.35 8610.835 ;
      RECT 17592.77 187.44 17593.83 8610.835 ;
      RECT 17575.79 187.44 17578.31 8610.835 ;
      RECT 17558.81 187.44 17561.33 8610.835 ;
      RECT 17543.29 187.44 17544.35 8610.835 ;
      RECT 17512.77 187.44 17513.83 8610.835 ;
      RECT 17495.79 187.44 17498.31 8610.835 ;
      RECT 17478.81 187.44 17481.33 8610.835 ;
      RECT 17463.29 187.44 17464.35 8610.835 ;
      RECT 17432.77 187.44 17433.83 8610.835 ;
      RECT 17415.79 187.44 17418.31 8610.835 ;
      RECT 17398.81 187.44 17401.33 8610.835 ;
      RECT 17383.29 187.44 17384.35 8610.835 ;
      RECT 17352.77 187.44 17353.83 8610.835 ;
      RECT 17335.79 187.44 17338.31 8610.835 ;
      RECT 17318.81 187.44 17321.33 8610.835 ;
      RECT 17303.29 187.44 17304.35 8610.835 ;
      RECT 17272.77 187.44 17273.83 8610.835 ;
      RECT 17255.79 187.44 17258.31 8610.835 ;
      RECT 17238.81 187.44 17241.33 8610.835 ;
      RECT 17223.29 187.44 17224.35 8610.835 ;
      RECT 17192.77 187.44 17193.83 8610.835 ;
      RECT 17175.79 187.44 17178.31 8610.835 ;
      RECT 17158.81 187.44 17161.33 8610.835 ;
      RECT 17143.29 187.44 17144.35 8610.835 ;
      RECT 17112.77 187.44 17113.83 8610.835 ;
      RECT 17095.79 187.44 17098.31 8610.835 ;
      RECT 17078.81 187.44 17081.33 8610.835 ;
      RECT 17063.29 187.44 17064.35 8610.835 ;
      RECT 17032.77 187.44 17033.83 8610.835 ;
      RECT 17015.79 187.44 17018.31 8610.835 ;
      RECT 16998.81 187.44 17001.33 8610.835 ;
      RECT 16983.29 187.44 16984.35 8610.835 ;
      RECT 16952.77 187.44 16953.83 8610.835 ;
      RECT 16935.79 187.44 16938.31 8610.835 ;
      RECT 16918.81 187.44 16921.33 8610.835 ;
      RECT 16903.29 187.44 16904.35 8610.835 ;
      RECT 16872.77 187.44 16873.83 8610.835 ;
      RECT 16855.79 187.44 16858.31 8610.835 ;
      RECT 16838.81 187.44 16841.33 8610.835 ;
      RECT 16823.29 187.44 16824.35 8610.835 ;
      RECT 16792.77 187.44 16793.83 8610.835 ;
      RECT 16775.79 187.44 16778.31 8610.835 ;
      RECT 16758.81 187.44 16761.33 8610.835 ;
      RECT 16743.29 187.44 16744.35 8610.835 ;
      RECT 16712.77 187.44 16713.83 8610.835 ;
      RECT 16695.79 187.44 16698.31 8610.835 ;
      RECT 16678.81 187.44 16681.33 8610.835 ;
      RECT 16663.29 187.44 16664.35 8610.835 ;
      RECT 16632.77 187.44 16633.83 8610.835 ;
      RECT 16615.79 187.44 16618.31 8610.835 ;
      RECT 16598.81 187.44 16601.33 8610.835 ;
      RECT 16583.29 187.44 16584.35 8610.835 ;
      RECT 16552.77 187.44 16553.83 8610.835 ;
      RECT 16535.79 187.44 16538.31 8610.835 ;
      RECT 16518.81 187.44 16521.33 8610.835 ;
      RECT 16503.29 187.44 16504.35 8610.835 ;
      RECT 16472.77 187.44 16473.83 8610.835 ;
      RECT 16455.79 187.44 16458.31 8610.835 ;
      RECT 16438.81 187.44 16441.33 8610.835 ;
      RECT 16423.29 187.44 16424.35 8610.835 ;
      RECT 16392.77 187.44 16393.83 8610.835 ;
      RECT 16375.79 187.44 16378.31 8610.835 ;
      RECT 16358.81 187.44 16361.33 8610.835 ;
      RECT 16343.29 187.44 16344.35 8610.835 ;
      RECT 16312.77 187.44 16313.83 8610.835 ;
      RECT 16295.79 187.44 16298.31 8610.835 ;
      RECT 16278.81 187.44 16281.33 8610.835 ;
      RECT 16263.29 187.44 16264.35 8610.835 ;
      RECT 16232.77 187.44 16233.83 8610.835 ;
      RECT 16215.79 187.44 16218.31 8610.835 ;
      RECT 16198.81 187.44 16201.33 8610.835 ;
      RECT 16183.29 187.44 16184.35 8610.835 ;
      RECT 16152.77 187.44 16153.83 8610.835 ;
      RECT 16135.79 187.44 16138.31 8610.835 ;
      RECT 16118.81 187.44 16121.33 8610.835 ;
      RECT 16103.29 187.44 16104.35 8610.835 ;
      RECT 16072.77 187.44 16073.83 8610.835 ;
      RECT 16055.79 187.44 16058.31 8610.835 ;
      RECT 16038.81 187.44 16041.33 8610.835 ;
      RECT 16023.29 187.44 16024.35 8610.835 ;
      RECT 15992.77 187.44 15993.83 8610.835 ;
      RECT 15975.79 187.44 15978.31 8610.835 ;
      RECT 15958.81 187.44 15961.33 8610.835 ;
      RECT 15943.29 187.44 15944.35 8610.835 ;
      RECT 15912.77 187.44 15913.83 8610.835 ;
      RECT 15895.79 187.44 15898.31 8610.835 ;
      RECT 15878.81 187.44 15881.33 8610.835 ;
      RECT 15863.29 187.44 15864.35 8610.835 ;
      RECT 15832.77 187.44 15833.83 8610.835 ;
      RECT 15815.79 187.44 15818.31 8610.835 ;
      RECT 15798.81 187.44 15801.33 8610.835 ;
      RECT 15783.29 187.44 15784.35 8610.835 ;
      RECT 15752.77 187.44 15753.83 8610.835 ;
      RECT 15735.79 187.44 15738.31 8610.835 ;
      RECT 15718.81 187.44 15721.33 8610.835 ;
      RECT 15703.29 187.44 15704.35 8610.835 ;
      RECT 15672.77 187.44 15673.83 8610.835 ;
      RECT 15655.79 187.44 15658.31 8610.835 ;
      RECT 15638.81 187.44 15641.33 8610.835 ;
      RECT 15623.29 187.44 15624.35 8610.835 ;
      RECT 15592.77 187.44 15593.83 8610.835 ;
      RECT 15575.79 187.44 15578.31 8610.835 ;
      RECT 15558.81 187.44 15561.33 8610.835 ;
      RECT 15543.29 187.44 15544.35 8610.835 ;
      RECT 15512.77 187.44 15513.83 8610.835 ;
      RECT 15495.79 187.44 15498.31 8610.835 ;
      RECT 15478.81 187.44 15481.33 8610.835 ;
      RECT 15463.29 187.44 15464.35 8610.835 ;
      RECT 15432.77 187.44 15433.83 8610.835 ;
      RECT 15415.79 187.44 15418.31 8610.835 ;
      RECT 15398.81 187.44 15401.33 8610.835 ;
      RECT 15383.29 187.44 15384.35 8610.835 ;
      RECT 15352.77 187.44 15353.83 8610.835 ;
      RECT 15335.79 187.44 15338.31 8610.835 ;
      RECT 15318.81 187.44 15321.33 8610.835 ;
      RECT 15303.29 187.44 15304.35 8610.835 ;
      RECT 15272.77 187.44 15273.83 8610.835 ;
      RECT 15255.79 187.44 15258.31 8610.835 ;
      RECT 15238.81 187.44 15241.33 8610.835 ;
      RECT 15223.29 187.44 15224.35 8610.835 ;
      RECT 15192.77 187.44 15193.83 8610.835 ;
      RECT 15175.79 187.44 15178.31 8610.835 ;
      RECT 15158.81 187.44 15161.33 8610.835 ;
      RECT 15143.29 187.44 15144.35 8610.835 ;
      RECT 15112.77 187.44 15113.83 8610.835 ;
      RECT 15095.79 187.44 15098.31 8610.835 ;
      RECT 15078.81 187.44 15081.33 8610.835 ;
      RECT 15063.29 187.44 15064.35 8610.835 ;
      RECT 15032.77 187.44 15033.83 8610.835 ;
      RECT 15015.79 187.44 15018.31 8610.835 ;
      RECT 14998.81 187.44 15001.33 8610.835 ;
      RECT 14983.29 187.44 14984.35 8610.835 ;
      RECT 14952.77 187.44 14953.83 8610.835 ;
      RECT 14935.79 187.44 14938.31 8610.835 ;
      RECT 14918.81 187.44 14921.33 8610.835 ;
      RECT 14903.29 187.44 14904.35 8610.835 ;
      RECT 14872.77 187.44 14873.83 8610.835 ;
      RECT 14855.79 187.44 14858.31 8610.835 ;
      RECT 14838.81 187.44 14841.33 8610.835 ;
      RECT 14823.29 187.44 14824.35 8610.835 ;
      RECT 14792.77 187.44 14793.83 8610.835 ;
      RECT 14775.79 187.44 14778.31 8610.835 ;
      RECT 14758.81 187.44 14761.33 8610.835 ;
      RECT 14743.29 187.44 14744.35 8610.835 ;
      RECT 14712.77 187.44 14713.83 8610.835 ;
      RECT 14695.79 187.44 14698.31 8610.835 ;
      RECT 14678.81 187.44 14681.33 8610.835 ;
      RECT 14663.29 187.44 14664.35 8610.835 ;
      RECT 14632.77 187.44 14633.83 8610.835 ;
      RECT 14615.79 187.44 14618.31 8610.835 ;
      RECT 14598.81 187.44 14601.33 8610.835 ;
      RECT 14583.29 187.44 14584.35 8610.835 ;
      RECT 14552.77 187.44 14553.83 8610.835 ;
      RECT 14535.79 187.44 14538.31 8610.835 ;
      RECT 14518.81 187.44 14521.33 8610.835 ;
      RECT 14503.29 187.44 14504.35 8610.835 ;
      RECT 14472.77 187.44 14473.83 8610.835 ;
      RECT 14455.79 187.44 14458.31 8610.835 ;
      RECT 14438.81 187.44 14441.33 8610.835 ;
      RECT 14423.29 187.44 14424.35 8610.835 ;
      RECT 14392.77 187.44 14393.83 8610.835 ;
      RECT 14375.79 187.44 14378.31 8610.835 ;
      RECT 14358.81 187.44 14361.33 8610.835 ;
      RECT 14343.29 187.44 14344.35 8610.835 ;
      RECT 14312.77 187.44 14313.83 8610.835 ;
      RECT 14295.79 187.44 14298.31 8610.835 ;
      RECT 14278.81 187.44 14281.33 8610.835 ;
      RECT 14263.29 187.44 14264.35 8610.835 ;
      RECT 14232.77 187.44 14233.83 8610.835 ;
      RECT 14215.79 187.44 14218.31 8610.835 ;
      RECT 14198.81 187.44 14201.33 8610.835 ;
      RECT 14183.29 187.44 14184.35 8610.835 ;
      RECT 14152.77 187.44 14153.83 8610.835 ;
      RECT 14135.79 187.44 14138.31 8610.835 ;
      RECT 14118.81 187.44 14121.33 8610.835 ;
      RECT 14103.29 187.44 14104.35 8610.835 ;
      RECT 14072.77 187.44 14073.83 8610.835 ;
      RECT 14055.79 187.44 14058.31 8610.835 ;
      RECT 14038.81 187.44 14041.33 8610.835 ;
      RECT 14023.29 187.44 14024.35 8610.835 ;
      RECT 13992.77 187.44 13993.83 8610.835 ;
      RECT 13975.79 187.44 13978.31 8610.835 ;
      RECT 13958.81 187.44 13961.33 8610.835 ;
      RECT 13943.29 187.44 13944.35 8610.835 ;
      RECT 13912.77 187.44 13913.83 8610.835 ;
      RECT 13895.79 187.44 13898.31 8610.835 ;
      RECT 13878.81 187.44 13881.33 8610.835 ;
      RECT 13863.29 187.44 13864.35 8610.835 ;
      RECT 13832.77 187.44 13833.83 8610.835 ;
      RECT 13815.79 187.44 13818.31 8610.835 ;
      RECT 13798.81 187.44 13801.33 8610.835 ;
      RECT 13783.29 187.44 13784.35 8610.835 ;
      RECT 13752.77 187.44 13753.83 8610.835 ;
      RECT 13735.79 187.44 13738.31 8610.835 ;
      RECT 13718.81 187.44 13721.33 8610.835 ;
      RECT 13703.29 187.44 13704.35 8610.835 ;
      RECT 13672.77 187.44 13673.83 8610.835 ;
      RECT 13655.79 187.44 13658.31 8610.835 ;
      RECT 13638.81 187.44 13641.33 8610.835 ;
      RECT 13623.29 187.44 13624.35 8610.835 ;
      RECT 13592.77 187.44 13593.83 8610.835 ;
      RECT 13575.79 187.44 13578.31 8610.835 ;
      RECT 13558.81 187.44 13561.33 8610.835 ;
      RECT 13543.29 187.44 13544.35 8610.835 ;
      RECT 13512.77 187.44 13513.83 8610.835 ;
      RECT 13495.79 187.44 13498.31 8610.835 ;
      RECT 13478.81 187.44 13481.33 8610.835 ;
      RECT 13463.29 187.44 13464.35 8610.835 ;
      RECT 13432.77 187.44 13433.83 8610.835 ;
      RECT 13415.79 187.44 13418.31 8610.835 ;
      RECT 13398.81 187.44 13401.33 8610.835 ;
      RECT 13383.29 187.44 13384.35 8610.835 ;
      RECT 13352.77 187.44 13353.83 8610.835 ;
      RECT 13335.79 187.44 13338.31 8610.835 ;
      RECT 13318.81 187.44 13321.33 8610.835 ;
      RECT 13303.29 187.44 13304.35 8610.835 ;
      RECT 13272.77 187.44 13273.83 8610.835 ;
      RECT 13255.79 187.44 13258.31 8610.835 ;
      RECT 13238.81 187.44 13241.33 8610.835 ;
      RECT 13223.29 187.44 13224.35 8610.835 ;
      RECT 13192.77 187.44 13193.83 8610.835 ;
      RECT 13175.79 187.44 13178.31 8610.835 ;
      RECT 13158.81 187.44 13161.33 8610.835 ;
      RECT 13143.29 187.44 13144.35 8610.835 ;
      RECT 13112.77 187.44 13113.83 8610.835 ;
      RECT 13095.79 187.44 13098.31 8610.835 ;
      RECT 13078.81 187.44 13081.33 8610.835 ;
      RECT 13063.29 187.44 13064.35 8610.835 ;
      RECT 13032.77 187.44 13033.83 8610.835 ;
      RECT 13015.79 187.44 13018.31 8610.835 ;
      RECT 12998.81 187.44 13001.33 8610.835 ;
      RECT 12983.29 187.44 12984.35 8610.835 ;
      RECT 12952.77 187.44 12953.83 8610.835 ;
      RECT 12935.79 187.44 12938.31 8610.835 ;
      RECT 12918.81 187.44 12921.33 8610.835 ;
      RECT 12903.29 187.44 12904.35 8610.835 ;
      RECT 12872.77 187.44 12873.83 8610.835 ;
      RECT 12855.79 187.44 12858.31 8610.835 ;
      RECT 12838.81 187.44 12841.33 8610.835 ;
      RECT 12823.29 187.44 12824.35 8610.835 ;
      RECT 12792.77 187.44 12793.83 8610.835 ;
      RECT 12775.79 187.44 12778.31 8610.835 ;
      RECT 12758.81 187.44 12761.33 8610.835 ;
      RECT 12743.29 187.44 12744.35 8610.835 ;
      RECT 12712.77 187.44 12713.83 8610.835 ;
      RECT 12695.79 187.44 12698.31 8610.835 ;
      RECT 12678.81 187.44 12681.33 8610.835 ;
      RECT 12663.29 187.44 12664.35 8610.835 ;
      RECT 12632.77 187.44 12633.83 8610.835 ;
      RECT 12615.79 187.44 12618.31 8610.835 ;
      RECT 12598.81 187.44 12601.33 8610.835 ;
      RECT 12583.29 187.44 12584.35 8610.835 ;
      RECT 12552.77 187.44 12553.83 8610.835 ;
      RECT 12535.79 187.44 12538.31 8610.835 ;
      RECT 12518.81 187.44 12521.33 8610.835 ;
      RECT 12503.29 187.44 12504.35 8610.835 ;
      RECT 12472.77 187.44 12473.83 8610.835 ;
      RECT 12455.79 187.44 12458.31 8610.835 ;
      RECT 12438.81 187.44 12441.33 8610.835 ;
      RECT 12423.29 187.44 12424.35 8610.835 ;
      RECT 12392.77 187.44 12393.83 8610.835 ;
      RECT 12375.79 187.44 12378.31 8610.835 ;
      RECT 12358.81 187.44 12361.33 8610.835 ;
      RECT 12343.29 187.44 12344.35 8610.835 ;
      RECT 12312.77 187.44 12313.83 8610.835 ;
      RECT 12295.79 187.44 12298.31 8610.835 ;
      RECT 12278.81 187.44 12281.33 8610.835 ;
      RECT 12263.29 187.44 12264.35 8610.835 ;
      RECT 12232.77 187.44 12233.83 8610.835 ;
      RECT 12215.79 187.44 12218.31 8610.835 ;
      RECT 12198.81 187.44 12201.33 8610.835 ;
      RECT 12183.29 187.44 12184.35 8610.835 ;
      RECT 12152.77 187.44 12153.83 8610.835 ;
      RECT 12135.79 187.44 12138.31 8610.835 ;
      RECT 12118.81 187.44 12121.33 8610.835 ;
      RECT 12103.29 187.44 12104.35 8610.835 ;
      RECT 12072.77 187.44 12073.83 8610.835 ;
      RECT 12055.79 187.44 12058.31 8610.835 ;
      RECT 12038.81 187.44 12041.33 8610.835 ;
      RECT 12023.29 187.44 12024.35 8610.835 ;
      RECT 11992.77 187.44 11993.83 8610.835 ;
      RECT 11975.79 187.44 11978.31 8610.835 ;
      RECT 11958.81 187.44 11961.33 8610.835 ;
      RECT 11943.29 187.44 11944.35 8610.835 ;
      RECT 11912.77 187.44 11913.83 8610.835 ;
      RECT 11895.79 187.44 11898.31 8610.835 ;
      RECT 11878.81 187.44 11881.33 8610.835 ;
      RECT 11863.29 187.44 11864.35 8610.835 ;
      RECT 11832.77 187.44 11833.83 8610.835 ;
      RECT 11815.79 187.44 11818.31 8610.835 ;
      RECT 11798.81 187.44 11801.33 8610.835 ;
      RECT 11783.29 187.44 11784.35 8610.835 ;
      RECT 11752.77 187.44 11753.83 8610.835 ;
      RECT 11735.79 187.44 11738.31 8610.835 ;
      RECT 11718.81 187.44 11721.33 8610.835 ;
      RECT 11703.29 187.44 11704.35 8610.835 ;
      RECT 11672.77 187.44 11673.83 8610.835 ;
      RECT 11655.79 187.44 11658.31 8610.835 ;
      RECT 11638.81 187.44 11641.33 8610.835 ;
      RECT 11623.29 187.44 11624.35 8610.835 ;
      RECT 11592.77 187.44 11593.83 8610.835 ;
      RECT 11575.79 187.44 11578.31 8610.835 ;
      RECT 11558.81 187.44 11561.33 8610.835 ;
      RECT 11543.29 187.44 11544.35 8610.835 ;
      RECT 11512.77 187.44 11513.83 8610.835 ;
      RECT 11495.79 187.44 11498.31 8610.835 ;
      RECT 11478.81 187.44 11481.33 8610.835 ;
      RECT 11463.29 187.44 11464.35 8610.835 ;
      RECT 11432.77 187.44 11433.83 8610.835 ;
      RECT 11415.79 187.44 11418.31 8610.835 ;
      RECT 11398.81 187.44 11401.33 8610.835 ;
      RECT 11383.29 187.44 11384.35 8610.835 ;
      RECT 11352.77 187.44 11353.83 8610.835 ;
      RECT 11335.79 187.44 11338.31 8610.835 ;
      RECT 11318.81 187.44 11321.33 8610.835 ;
      RECT 11303.29 187.44 11304.35 8610.835 ;
      RECT 11272.77 187.44 11273.83 8610.835 ;
      RECT 11255.79 187.44 11258.31 8610.835 ;
      RECT 11238.81 187.44 11241.33 8610.835 ;
      RECT 11223.29 187.44 11224.35 8610.835 ;
      RECT 11192.77 187.44 11193.83 8610.835 ;
      RECT 11175.79 187.44 11178.31 8610.835 ;
      RECT 11158.81 187.44 11161.33 8610.835 ;
      RECT 11143.29 187.44 11144.35 8610.835 ;
      RECT 11112.77 187.44 11113.83 8610.835 ;
      RECT 11095.79 187.44 11098.31 8610.835 ;
      RECT 11078.81 187.44 11081.33 8610.835 ;
      RECT 11063.29 187.44 11064.35 8610.835 ;
      RECT 11032.77 187.44 11033.83 8610.835 ;
      RECT 11015.79 187.44 11018.31 8610.835 ;
      RECT 10998.81 187.44 11001.33 8610.835 ;
      RECT 10983.29 187.44 10984.35 8610.835 ;
      RECT 10952.77 187.44 10953.83 8610.835 ;
      RECT 10935.79 187.44 10938.31 8610.835 ;
      RECT 10918.81 187.44 10921.33 8610.835 ;
      RECT 10903.29 187.44 10904.35 8610.835 ;
      RECT 10872.77 187.44 10873.83 8610.835 ;
      RECT 10855.79 187.44 10858.31 8610.835 ;
      RECT 10838.81 187.44 10841.33 8610.835 ;
      RECT 10823.29 187.44 10824.35 8610.835 ;
      RECT 10792.77 187.44 10793.83 8610.835 ;
      RECT 10775.79 187.44 10778.31 8610.835 ;
      RECT 10758.81 187.44 10761.33 8610.835 ;
      RECT 10743.29 187.44 10744.35 8610.835 ;
      RECT 10712.77 187.44 10713.83 8610.835 ;
      RECT 10695.79 187.44 10698.31 8610.835 ;
      RECT 10678.81 187.44 10681.33 8610.835 ;
      RECT 10663.29 187.44 10664.35 8610.835 ;
      RECT 10632.77 187.44 10633.83 8610.835 ;
      RECT 10615.79 187.44 10618.31 8610.835 ;
      RECT 10598.81 187.44 10601.33 8610.835 ;
      RECT 10583.29 187.44 10584.35 8610.835 ;
      RECT 10552.77 187.44 10553.83 8610.835 ;
      RECT 10535.79 187.44 10538.31 8610.835 ;
      RECT 10518.81 187.44 10521.33 8610.835 ;
      RECT 10503.29 187.44 10504.35 8610.835 ;
      RECT 10472.77 187.44 10473.83 8610.835 ;
      RECT 10455.79 187.44 10458.31 8610.835 ;
      RECT 10438.81 187.44 10441.33 8610.835 ;
      RECT 10423.29 187.44 10424.35 8610.835 ;
      RECT 10392.77 187.44 10393.83 8610.835 ;
      RECT 10375.79 187.44 10378.31 8610.835 ;
      RECT 10358.81 187.44 10361.33 8610.835 ;
      RECT 10343.29 187.44 10344.35 8610.835 ;
      RECT 10312.77 187.44 10313.83 8610.835 ;
      RECT 10295.79 187.44 10298.31 8610.835 ;
      RECT 10278.81 187.44 10281.33 8610.835 ;
      RECT 10263.29 187.44 10264.35 8610.835 ;
      RECT 10232.77 187.44 10233.83 8610.835 ;
      RECT 10215.79 187.44 10218.31 8610.835 ;
      RECT 10198.81 187.44 10201.33 8610.835 ;
      RECT 10183.29 187.44 10184.35 8610.835 ;
      RECT 10152.77 187.44 10153.83 8610.835 ;
      RECT 10135.79 187.44 10138.31 8610.835 ;
      RECT 10118.81 187.44 10121.33 8610.835 ;
      RECT 10103.29 187.44 10104.35 8610.835 ;
      RECT 10072.77 187.44 10073.83 8610.835 ;
      RECT 10055.79 187.44 10058.31 8610.835 ;
      RECT 10038.81 187.44 10041.33 8610.835 ;
      RECT 10023.29 187.44 10024.35 8610.835 ;
      RECT 9992.77 187.44 9993.83 8610.835 ;
      RECT 9975.79 187.44 9978.31 8610.835 ;
      RECT 9958.81 187.44 9961.33 8610.835 ;
      RECT 9943.29 187.44 9944.35 8610.835 ;
      RECT 9912.77 187.44 9913.83 8610.835 ;
      RECT 9895.79 187.44 9898.31 8610.835 ;
      RECT 9878.81 187.44 9881.33 8610.835 ;
      RECT 9863.29 187.44 9864.35 8610.835 ;
      RECT 9832.77 187.44 9833.83 8610.835 ;
      RECT 9815.79 187.44 9818.31 8610.835 ;
      RECT 9798.81 187.44 9801.33 8610.835 ;
      RECT 9783.29 187.44 9784.35 8610.835 ;
      RECT 9752.77 187.44 9753.83 8610.835 ;
      RECT 9735.79 187.44 9738.31 8610.835 ;
      RECT 9718.81 187.44 9721.33 8610.835 ;
      RECT 9703.29 187.44 9704.35 8610.835 ;
      RECT 9672.77 187.44 9673.83 8610.835 ;
      RECT 9655.79 187.44 9658.31 8610.835 ;
      RECT 9638.81 187.44 9641.33 8610.835 ;
      RECT 9623.29 187.44 9624.35 8610.835 ;
      RECT 9592.77 187.44 9593.83 8610.835 ;
      RECT 9575.79 187.44 9578.31 8610.835 ;
      RECT 9558.81 187.44 9561.33 8610.835 ;
      RECT 9543.29 187.44 9544.35 8610.835 ;
      RECT 9512.77 187.44 9513.83 8610.835 ;
      RECT 9495.79 187.44 9498.31 8610.835 ;
      RECT 9478.81 187.44 9481.33 8610.835 ;
      RECT 9463.29 187.44 9464.35 8610.835 ;
      RECT 9432.77 187.44 9433.83 8610.835 ;
      RECT 9415.79 187.44 9418.31 8610.835 ;
      RECT 9398.81 187.44 9401.33 8610.835 ;
      RECT 9383.29 187.44 9384.35 8610.835 ;
      RECT 9352.77 187.44 9353.83 8610.835 ;
      RECT 9335.79 187.44 9338.31 8610.835 ;
      RECT 9318.81 187.44 9321.33 8610.835 ;
      RECT 9303.29 187.44 9304.35 8610.835 ;
      RECT 9272.77 187.44 9273.83 8610.835 ;
      RECT 9255.79 187.44 9258.31 8610.835 ;
      RECT 9238.81 187.44 9241.33 8610.835 ;
      RECT 9223.29 187.44 9224.35 8610.835 ;
      RECT 9192.77 187.44 9193.83 8610.835 ;
      RECT 9175.79 187.44 9178.31 8610.835 ;
      RECT 9158.81 187.44 9161.33 8610.835 ;
      RECT 9143.29 187.44 9144.35 8610.835 ;
      RECT 9112.77 187.44 9113.83 8610.835 ;
      RECT 9095.79 187.44 9098.31 8610.835 ;
      RECT 9078.81 187.44 9081.33 8610.835 ;
      RECT 9063.29 187.44 9064.35 8610.835 ;
      RECT 9032.77 187.44 9033.83 8610.835 ;
      RECT 9015.79 187.44 9018.31 8610.835 ;
      RECT 8998.81 187.44 9001.33 8610.835 ;
      RECT 8983.29 187.44 8984.35 8610.835 ;
      RECT 8952.77 187.44 8953.83 8610.835 ;
      RECT 8935.79 187.44 8938.31 8610.835 ;
      RECT 8918.81 187.44 8921.33 8610.835 ;
      RECT 8903.29 187.44 8904.35 8610.835 ;
      RECT 8872.77 187.44 8873.83 8610.835 ;
      RECT 8855.79 187.44 8858.31 8610.835 ;
      RECT 8838.81 187.44 8841.33 8610.835 ;
      RECT 8823.29 187.44 8824.35 8610.835 ;
      RECT 8792.77 187.44 8793.83 8610.835 ;
      RECT 8775.79 187.44 8778.31 8610.835 ;
      RECT 8758.81 187.44 8761.33 8610.835 ;
      RECT 8743.29 187.44 8744.35 8610.835 ;
      RECT 8712.77 187.44 8713.83 8610.835 ;
      RECT 8695.79 187.44 8698.31 8610.835 ;
      RECT 8678.81 187.44 8681.33 8610.835 ;
      RECT 8663.29 187.44 8664.35 8610.835 ;
      RECT 8632.77 187.44 8633.83 8610.835 ;
      RECT 8615.79 187.44 8618.31 8610.835 ;
      RECT 8598.81 187.44 8601.33 8610.835 ;
      RECT 8583.29 187.44 8584.35 8610.835 ;
      RECT 8552.77 187.44 8553.83 8610.835 ;
      RECT 8535.79 187.44 8538.31 8610.835 ;
      RECT 8518.81 187.44 8521.33 8610.835 ;
      RECT 8503.29 187.44 8504.35 8610.835 ;
      RECT 8472.77 187.44 8473.83 8610.835 ;
      RECT 8455.79 187.44 8458.31 8610.835 ;
      RECT 8438.81 187.44 8441.33 8610.835 ;
      RECT 8423.29 187.44 8424.35 8610.835 ;
      RECT 8392.77 187.44 8393.83 8610.835 ;
      RECT 8375.79 187.44 8378.31 8610.835 ;
      RECT 8358.81 187.44 8361.33 8610.835 ;
      RECT 8343.29 187.44 8344.35 8610.835 ;
      RECT 8312.77 187.44 8313.83 8610.835 ;
      RECT 8295.79 187.44 8298.31 8610.835 ;
      RECT 8278.81 187.44 8281.33 8610.835 ;
      RECT 8263.29 187.44 8264.35 8610.835 ;
      RECT 8232.77 187.44 8233.83 8610.835 ;
      RECT 8215.79 187.44 8218.31 8610.835 ;
      RECT 8198.81 187.44 8201.33 8610.835 ;
      RECT 8183.29 187.44 8184.35 8610.835 ;
      RECT 8152.77 187.44 8153.83 8610.835 ;
      RECT 8135.79 187.44 8138.31 8610.835 ;
      RECT 8118.81 187.44 8121.33 8610.835 ;
      RECT 8103.29 187.44 8104.35 8610.835 ;
      RECT 8072.77 187.44 8073.83 8610.835 ;
      RECT 8055.79 187.44 8058.31 8610.835 ;
      RECT 8038.81 187.44 8041.33 8610.835 ;
      RECT 8023.29 187.44 8024.35 8610.835 ;
      RECT 7992.77 187.44 7993.83 8610.835 ;
      RECT 7975.79 187.44 7978.31 8610.835 ;
      RECT 7958.81 187.44 7961.33 8610.835 ;
      RECT 7943.29 187.44 7944.35 8610.835 ;
      RECT 7912.77 187.44 7913.83 8610.835 ;
      RECT 7895.79 187.44 7898.31 8610.835 ;
      RECT 7878.81 187.44 7881.33 8610.835 ;
      RECT 7863.29 187.44 7864.35 8610.835 ;
      RECT 7832.77 187.44 7833.83 8610.835 ;
      RECT 7815.79 187.44 7818.31 8610.835 ;
      RECT 7798.81 187.44 7801.33 8610.835 ;
      RECT 7783.29 187.44 7784.35 8610.835 ;
      RECT 7752.77 187.44 7753.83 8610.835 ;
      RECT 7735.79 187.44 7738.31 8610.835 ;
      RECT 7718.81 187.44 7721.33 8610.835 ;
      RECT 7703.29 187.44 7704.35 8610.835 ;
      RECT 7672.77 187.44 7673.83 8610.835 ;
      RECT 7655.79 187.44 7658.31 8610.835 ;
      RECT 7638.81 187.44 7641.33 8610.835 ;
      RECT 7623.29 187.44 7624.35 8610.835 ;
      RECT 7592.77 187.44 7593.83 8610.835 ;
      RECT 7575.79 187.44 7578.31 8610.835 ;
      RECT 7558.81 187.44 7561.33 8610.835 ;
      RECT 7543.29 187.44 7544.35 8610.835 ;
      RECT 7512.77 187.44 7513.83 8610.835 ;
      RECT 7495.79 187.44 7498.31 8610.835 ;
      RECT 7478.81 187.44 7481.33 8610.835 ;
      RECT 7463.29 187.44 7464.35 8610.835 ;
      RECT 7432.77 187.44 7433.83 8610.835 ;
      RECT 7415.79 187.44 7418.31 8610.835 ;
      RECT 7398.81 187.44 7401.33 8610.835 ;
      RECT 7383.29 187.44 7384.35 8610.835 ;
      RECT 7352.77 187.44 7353.83 8610.835 ;
      RECT 7335.79 187.44 7338.31 8610.835 ;
      RECT 7318.81 187.44 7321.33 8610.835 ;
      RECT 7303.29 187.44 7304.35 8610.835 ;
      RECT 7272.77 187.44 7273.83 8610.835 ;
      RECT 7255.79 187.44 7258.31 8610.835 ;
      RECT 7238.81 187.44 7241.33 8610.835 ;
      RECT 7223.29 187.44 7224.35 8610.835 ;
      RECT 7192.77 187.44 7193.83 8610.835 ;
      RECT 7175.79 187.44 7178.31 8610.835 ;
      RECT 7158.81 187.44 7161.33 8610.835 ;
      RECT 7143.29 187.44 7144.35 8610.835 ;
      RECT 7112.77 187.44 7113.83 8610.835 ;
      RECT 7095.79 187.44 7098.31 8610.835 ;
      RECT 7078.81 187.44 7081.33 8610.835 ;
      RECT 7063.29 187.44 7064.35 8610.835 ;
      RECT 7032.77 187.44 7033.83 8610.835 ;
      RECT 7015.79 187.44 7018.31 8610.835 ;
      RECT 6998.81 187.44 7001.33 8610.835 ;
      RECT 6983.29 187.44 6984.35 8610.835 ;
      RECT 6952.77 187.44 6953.83 8610.835 ;
      RECT 6935.79 187.44 6938.31 8610.835 ;
      RECT 6918.81 187.44 6921.33 8610.835 ;
      RECT 6903.29 187.44 6904.35 8610.835 ;
      RECT 6872.77 187.44 6873.83 8610.835 ;
      RECT 6855.79 187.44 6858.31 8610.835 ;
      RECT 6838.81 187.44 6841.33 8610.835 ;
      RECT 6823.29 187.44 6824.35 8610.835 ;
      RECT 6792.77 187.44 6793.83 8610.835 ;
      RECT 6775.79 187.44 6778.31 8610.835 ;
      RECT 6758.81 187.44 6761.33 8610.835 ;
      RECT 6743.29 187.44 6744.35 8610.835 ;
      RECT 6712.77 187.44 6713.83 8610.835 ;
      RECT 6695.79 187.44 6698.31 8610.835 ;
      RECT 6678.81 187.44 6681.33 8610.835 ;
      RECT 6663.29 187.44 6664.35 8610.835 ;
      RECT 6632.77 187.44 6633.83 8610.835 ;
      RECT 6615.79 187.44 6618.31 8610.835 ;
      RECT 6598.81 187.44 6601.33 8610.835 ;
      RECT 6583.29 187.44 6584.35 8610.835 ;
      RECT 6552.77 187.44 6553.83 8610.835 ;
      RECT 6535.79 187.44 6538.31 8610.835 ;
      RECT 6518.81 187.44 6521.33 8610.835 ;
      RECT 6503.29 187.44 6504.35 8610.835 ;
      RECT 6472.77 187.44 6473.83 8610.835 ;
      RECT 6455.79 187.44 6458.31 8610.835 ;
      RECT 6438.81 187.44 6441.33 8610.835 ;
      RECT 6423.29 187.44 6424.35 8610.835 ;
      RECT 6392.77 187.44 6393.83 8610.835 ;
      RECT 6375.79 187.44 6378.31 8610.835 ;
      RECT 6358.81 187.44 6361.33 8610.835 ;
      RECT 6343.29 187.44 6344.35 8610.835 ;
      RECT 6312.77 187.44 6313.83 8610.835 ;
      RECT 6295.79 187.44 6298.31 8610.835 ;
      RECT 6278.81 187.44 6281.33 8610.835 ;
      RECT 6263.29 187.44 6264.35 8610.835 ;
      RECT 6232.77 187.44 6233.83 8610.835 ;
      RECT 6215.79 187.44 6218.31 8610.835 ;
      RECT 6198.81 187.44 6201.33 8610.835 ;
      RECT 6183.29 187.44 6184.35 8610.835 ;
      RECT 6152.77 187.44 6153.83 8610.835 ;
      RECT 6135.79 187.44 6138.31 8610.835 ;
      RECT 6118.81 187.44 6121.33 8610.835 ;
      RECT 6103.29 187.44 6104.35 8610.835 ;
      RECT 6072.77 187.44 6073.83 8610.835 ;
      RECT 6055.79 187.44 6058.31 8610.835 ;
      RECT 6038.81 187.44 6041.33 8610.835 ;
      RECT 6023.29 187.44 6024.35 8610.835 ;
      RECT 5992.77 187.44 5993.83 8610.835 ;
      RECT 5975.79 187.44 5978.31 8610.835 ;
      RECT 5958.81 187.44 5961.33 8610.835 ;
      RECT 5943.29 187.44 5944.35 8610.835 ;
      RECT 5912.77 187.44 5913.83 8610.835 ;
      RECT 5895.79 187.44 5898.31 8610.835 ;
      RECT 5878.81 187.44 5881.33 8610.835 ;
      RECT 5863.29 187.44 5864.35 8610.835 ;
      RECT 5832.77 187.44 5833.83 8610.835 ;
      RECT 5815.79 187.44 5818.31 8610.835 ;
      RECT 5798.81 187.44 5801.33 8610.835 ;
      RECT 5783.29 187.44 5784.35 8610.835 ;
      RECT 5752.77 187.44 5753.83 8610.835 ;
      RECT 5735.79 187.44 5738.31 8610.835 ;
      RECT 5718.81 187.44 5721.33 8610.835 ;
      RECT 5703.29 187.44 5704.35 8610.835 ;
      RECT 5672.77 187.44 5673.83 8610.835 ;
      RECT 5655.79 187.44 5658.31 8610.835 ;
      RECT 5638.81 187.44 5641.33 8610.835 ;
      RECT 5623.29 187.44 5624.35 8610.835 ;
      RECT 5592.77 187.44 5593.83 8610.835 ;
      RECT 5575.79 187.44 5578.31 8610.835 ;
      RECT 5558.81 187.44 5561.33 8610.835 ;
      RECT 5543.29 187.44 5544.35 8610.835 ;
      RECT 5512.77 187.44 5513.83 8610.835 ;
      RECT 5495.79 187.44 5498.31 8610.835 ;
      RECT 5478.81 187.44 5481.33 8610.835 ;
      RECT 5463.29 187.44 5464.35 8610.835 ;
      RECT 5432.77 187.44 5433.83 8610.835 ;
      RECT 5415.79 187.44 5418.31 8610.835 ;
      RECT 5398.81 187.44 5401.33 8610.835 ;
      RECT 5383.29 187.44 5384.35 8610.835 ;
      RECT 5352.77 187.44 5353.83 8610.835 ;
      RECT 5335.79 187.44 5338.31 8610.835 ;
      RECT 5318.81 187.44 5321.33 8610.835 ;
      RECT 5303.29 187.44 5304.35 8610.835 ;
      RECT 5272.77 187.44 5273.83 8610.835 ;
      RECT 5255.79 187.44 5258.31 8610.835 ;
      RECT 5238.81 187.44 5241.33 8610.835 ;
      RECT 5223.29 187.44 5224.35 8610.835 ;
      RECT 5192.77 187.44 5193.83 8610.835 ;
      RECT 5175.79 187.44 5178.31 8610.835 ;
      RECT 5158.81 187.44 5161.33 8610.835 ;
      RECT 5143.29 187.44 5144.35 8610.835 ;
      RECT 5112.77 187.44 5113.83 8610.835 ;
      RECT 5095.79 187.44 5098.31 8610.835 ;
      RECT 5078.81 187.44 5081.33 8610.835 ;
      RECT 5063.29 187.44 5064.35 8610.835 ;
      RECT 5032.77 187.44 5033.83 8610.835 ;
      RECT 5015.79 187.44 5018.31 8610.835 ;
      RECT 4998.81 187.44 5001.33 8610.835 ;
      RECT 4983.29 187.44 4984.35 8610.835 ;
      RECT 4952.77 187.44 4953.83 8610.835 ;
      RECT 4935.79 187.44 4938.31 8610.835 ;
      RECT 4918.81 187.44 4921.33 8610.835 ;
      RECT 4903.29 187.44 4904.35 8610.835 ;
      RECT 4872.77 187.44 4873.83 8610.835 ;
      RECT 4855.79 187.44 4858.31 8610.835 ;
      RECT 4838.81 187.44 4841.33 8610.835 ;
      RECT 4823.29 187.44 4824.35 8610.835 ;
      RECT 4792.77 187.44 4793.83 8610.835 ;
      RECT 4775.79 187.44 4778.31 8610.835 ;
      RECT 4758.81 187.44 4761.33 8610.835 ;
      RECT 4743.29 187.44 4744.35 8610.835 ;
      RECT 4712.77 187.44 4713.83 8610.835 ;
      RECT 4695.79 187.44 4698.31 8610.835 ;
      RECT 4678.81 187.44 4681.33 8610.835 ;
      RECT 4663.29 187.44 4664.35 8610.835 ;
      RECT 4632.77 187.44 4633.83 8610.835 ;
      RECT 4615.79 187.44 4618.31 8610.835 ;
      RECT 4598.81 187.44 4601.33 8610.835 ;
      RECT 4583.29 187.44 4584.35 8610.835 ;
      RECT 4552.77 187.44 4553.83 8610.835 ;
      RECT 4535.79 187.44 4538.31 8610.835 ;
      RECT 4518.81 187.44 4521.33 8610.835 ;
      RECT 4503.29 187.44 4504.35 8610.835 ;
      RECT 4472.77 187.44 4473.83 8610.835 ;
      RECT 4455.79 187.44 4458.31 8610.835 ;
      RECT 4438.81 187.44 4441.33 8610.835 ;
      RECT 4423.29 187.44 4424.35 8610.835 ;
      RECT 4392.77 187.44 4393.83 8610.835 ;
      RECT 4375.79 187.44 4378.31 8610.835 ;
      RECT 4358.81 187.44 4361.33 8610.835 ;
      RECT 4343.29 187.44 4344.35 8610.835 ;
      RECT 4312.77 187.44 4313.83 8610.835 ;
      RECT 4295.79 187.44 4298.31 8610.835 ;
      RECT 4278.81 187.44 4281.33 8610.835 ;
      RECT 4263.29 187.44 4264.35 8610.835 ;
      RECT 4232.77 187.44 4233.83 8610.835 ;
      RECT 4215.79 187.44 4218.31 8610.835 ;
      RECT 4198.81 187.44 4201.33 8610.835 ;
      RECT 4183.29 187.44 4184.35 8610.835 ;
      RECT 4152.77 187.44 4153.83 8610.835 ;
      RECT 4135.79 187.44 4138.31 8610.835 ;
      RECT 4118.81 187.44 4121.33 8610.835 ;
      RECT 4103.29 187.44 4104.35 8610.835 ;
      RECT 4072.77 187.44 4073.83 8610.835 ;
      RECT 4055.79 187.44 4058.31 8610.835 ;
      RECT 4038.81 187.44 4041.33 8610.835 ;
      RECT 4023.29 187.44 4024.35 8610.835 ;
      RECT 3992.77 187.44 3993.83 8610.835 ;
      RECT 3975.79 187.44 3978.31 8610.835 ;
      RECT 3958.81 187.44 3961.33 8610.835 ;
      RECT 3943.29 187.44 3944.35 8610.835 ;
      RECT 3912.77 187.44 3913.83 8610.835 ;
      RECT 3895.79 187.44 3898.31 8610.835 ;
      RECT 3878.81 187.44 3881.33 8610.835 ;
      RECT 3863.29 187.44 3864.35 8610.835 ;
      RECT 3832.77 187.44 3833.83 8610.835 ;
      RECT 3815.79 187.44 3818.31 8610.835 ;
      RECT 3798.81 187.44 3801.33 8610.835 ;
      RECT 3783.29 187.44 3784.35 8610.835 ;
      RECT 3752.77 187.44 3753.83 8610.835 ;
      RECT 3735.79 187.44 3738.31 8610.835 ;
      RECT 3718.81 187.44 3721.33 8610.835 ;
      RECT 3703.29 187.44 3704.35 8610.835 ;
      RECT 3672.77 187.44 3673.83 8610.835 ;
      RECT 3655.79 187.44 3658.31 8610.835 ;
      RECT 3638.81 187.44 3641.33 8610.835 ;
      RECT 3623.29 187.44 3624.35 8610.835 ;
      RECT 3592.77 187.44 3593.83 8610.835 ;
      RECT 3575.79 187.44 3578.31 8610.835 ;
      RECT 3558.81 187.44 3561.33 8610.835 ;
      RECT 3543.29 187.44 3544.35 8610.835 ;
      RECT 3512.77 187.44 3513.83 8610.835 ;
      RECT 3495.79 187.44 3498.31 8610.835 ;
      RECT 3478.81 187.44 3481.33 8610.835 ;
      RECT 3463.29 187.44 3464.35 8610.835 ;
      RECT 3432.77 187.44 3433.83 8610.835 ;
      RECT 3415.79 187.44 3418.31 8610.835 ;
      RECT 3398.81 187.44 3401.33 8610.835 ;
      RECT 3383.29 187.44 3384.35 8610.835 ;
      RECT 3352.77 187.44 3353.83 8610.835 ;
      RECT 3335.79 187.44 3338.31 8610.835 ;
      RECT 3318.81 187.44 3321.33 8610.835 ;
      RECT 3303.29 187.44 3304.35 8610.835 ;
      RECT 3272.77 187.44 3273.83 8610.835 ;
      RECT 3255.79 187.44 3258.31 8610.835 ;
      RECT 3238.81 187.44 3241.33 8610.835 ;
      RECT 3223.29 187.44 3224.35 8610.835 ;
      RECT 3192.77 187.44 3193.83 8610.835 ;
      RECT 3175.79 187.44 3178.31 8610.835 ;
      RECT 3158.81 187.44 3161.33 8610.835 ;
      RECT 3143.29 187.44 3144.35 8610.835 ;
      RECT 3112.77 187.44 3113.83 8610.835 ;
      RECT 3095.79 187.44 3098.31 8610.835 ;
      RECT 3078.81 187.44 3081.33 8610.835 ;
      RECT 3063.29 187.44 3064.35 8610.835 ;
      RECT 3032.77 187.44 3033.83 8610.835 ;
      RECT 3015.79 187.44 3018.31 8610.835 ;
      RECT 2998.81 187.44 3001.33 8610.835 ;
      RECT 2983.29 187.44 2984.35 8610.835 ;
      RECT 2952.77 187.44 2953.83 8610.835 ;
      RECT 2935.79 187.44 2938.31 8610.835 ;
      RECT 2918.81 187.44 2921.33 8610.835 ;
      RECT 2903.29 187.44 2904.35 8610.835 ;
      RECT 2872.77 187.44 2873.83 8610.835 ;
      RECT 2855.79 187.44 2858.31 8610.835 ;
      RECT 2838.81 187.44 2841.33 8610.835 ;
      RECT 2823.29 187.44 2824.35 8610.835 ;
      RECT 2792.77 187.44 2793.83 8610.835 ;
      RECT 2775.79 187.44 2778.31 8610.835 ;
      RECT 2758.81 187.44 2761.33 8610.835 ;
      RECT 2743.29 187.44 2744.35 8610.835 ;
      RECT 2712.77 187.44 2713.83 8610.835 ;
      RECT 2695.79 187.44 2698.31 8610.835 ;
      RECT 2678.81 187.44 2681.33 8610.835 ;
      RECT 2663.29 187.44 2664.35 8610.835 ;
      RECT 2632.77 187.44 2633.83 8610.835 ;
      RECT 2615.79 187.44 2618.31 8610.835 ;
      RECT 2598.81 187.44 2601.33 8610.835 ;
      RECT 2583.29 187.44 2584.35 8610.835 ;
      RECT 2552.77 187.44 2553.83 8610.835 ;
      RECT 2535.79 187.44 2538.31 8610.835 ;
      RECT 2518.81 187.44 2521.33 8610.835 ;
      RECT 2503.29 187.44 2504.35 8610.835 ;
      RECT 2472.77 187.44 2473.83 8610.835 ;
      RECT 2455.79 187.44 2458.31 8610.835 ;
      RECT 2438.81 187.44 2441.33 8610.835 ;
      RECT 2423.29 187.44 2424.35 8610.835 ;
      RECT 2392.77 187.44 2393.83 8610.835 ;
      RECT 2375.79 187.44 2378.31 8610.835 ;
      RECT 2358.81 187.44 2361.33 8610.835 ;
      RECT 2343.29 187.44 2344.35 8610.835 ;
      RECT 326.66 8600.705 2313.83 8610.835 ;
      RECT 2312.77 187.44 2313.83 8610.835 ;
      RECT 328.39 189.17 2313.83 8610.835 ;
      RECT 326.66 8594.095 2313.83 8594.635 ;
      RECT 326.66 8587.485 2313.83 8588.025 ;
      RECT 326.66 8578.245 2313.83 8584.905 ;
      RECT 326.66 8570.475 2313.83 8571.015 ;
      RECT 326.66 8556.935 2313.83 8557.475 ;
      RECT 326.66 8543.045 2313.83 8549.705 ;
      RECT 326.66 8539.925 2313.83 8540.465 ;
      RECT 326.66 8533.315 2313.83 8533.855 ;
      RECT 326.66 8522.095 2313.83 8522.635 ;
      RECT 326.66 8515.485 2313.83 8516.025 ;
      RECT 326.66 8506.245 2313.83 8512.905 ;
      RECT 326.66 8498.475 2313.83 8499.015 ;
      RECT 326.66 8484.935 2313.83 8485.475 ;
      RECT 326.66 8471.045 2313.83 8477.705 ;
      RECT 326.66 8467.925 2313.83 8468.465 ;
      RECT 326.66 8461.315 2313.83 8461.855 ;
      RECT 326.66 8450.095 2313.83 8450.635 ;
      RECT 326.66 8443.485 2313.83 8444.025 ;
      RECT 326.66 8434.245 2313.83 8440.905 ;
      RECT 326.66 8426.475 2313.83 8427.015 ;
      RECT 326.66 8412.935 2313.83 8413.475 ;
      RECT 326.66 8399.045 2313.83 8405.705 ;
      RECT 326.66 8395.925 2313.83 8396.465 ;
      RECT 326.66 8389.315 2313.83 8389.855 ;
      RECT 326.66 8378.095 2313.83 8378.635 ;
      RECT 326.66 8371.485 2313.83 8372.025 ;
      RECT 326.66 8362.245 2313.83 8368.905 ;
      RECT 326.66 8354.475 2313.83 8355.015 ;
      RECT 326.66 8340.935 2313.83 8341.475 ;
      RECT 326.66 8327.045 2313.83 8333.705 ;
      RECT 326.66 8323.925 2313.83 8324.465 ;
      RECT 326.66 8317.315 2313.83 8317.855 ;
      RECT 326.66 8306.095 2313.83 8306.635 ;
      RECT 326.66 8299.485 2313.83 8300.025 ;
      RECT 326.66 8290.245 2313.83 8296.905 ;
      RECT 326.66 8282.475 2313.83 8283.015 ;
      RECT 326.66 8268.935 2313.83 8269.475 ;
      RECT 326.66 8255.045 2313.83 8261.705 ;
      RECT 326.66 8251.925 2313.83 8252.465 ;
      RECT 326.66 8245.315 2313.83 8245.855 ;
      RECT 326.66 8234.095 2313.83 8234.635 ;
      RECT 326.66 8227.485 2313.83 8228.025 ;
      RECT 326.66 8218.245 2313.83 8224.905 ;
      RECT 326.66 8210.475 2313.83 8211.015 ;
      RECT 326.66 8196.935 2313.83 8197.475 ;
      RECT 326.66 8183.045 2313.83 8189.705 ;
      RECT 326.66 8179.925 2313.83 8180.465 ;
      RECT 326.66 8173.315 2313.83 8173.855 ;
      RECT 326.66 8162.095 2313.83 8162.635 ;
      RECT 326.66 8155.485 2313.83 8156.025 ;
      RECT 326.66 8146.245 2313.83 8152.905 ;
      RECT 326.66 8138.475 2313.83 8139.015 ;
      RECT 326.66 8124.935 2313.83 8125.475 ;
      RECT 326.66 8111.045 2313.83 8117.705 ;
      RECT 326.66 8107.925 2313.83 8108.465 ;
      RECT 326.66 8101.315 2313.83 8101.855 ;
      RECT 326.66 8090.095 2313.83 8090.635 ;
      RECT 326.66 8083.485 2313.83 8084.025 ;
      RECT 326.66 8074.245 2313.83 8080.905 ;
      RECT 326.66 8066.475 2313.83 8067.015 ;
      RECT 326.66 8052.935 2313.83 8053.475 ;
      RECT 326.66 8039.045 2313.83 8045.705 ;
      RECT 326.66 8035.925 2313.83 8036.465 ;
      RECT 326.66 8029.315 2313.83 8029.855 ;
      RECT 326.66 8018.095 2313.83 8018.635 ;
      RECT 326.66 8011.485 2313.83 8012.025 ;
      RECT 326.66 8002.245 2313.83 8008.905 ;
      RECT 326.66 7994.475 2313.83 7995.015 ;
      RECT 326.66 7980.935 2313.83 7981.475 ;
      RECT 326.66 7967.045 2313.83 7973.705 ;
      RECT 326.66 7963.925 2313.83 7964.465 ;
      RECT 326.66 7957.315 2313.83 7957.855 ;
      RECT 326.66 7946.095 2313.83 7946.635 ;
      RECT 326.66 7939.485 2313.83 7940.025 ;
      RECT 326.66 7930.245 2313.83 7936.905 ;
      RECT 326.66 7922.475 2313.83 7923.015 ;
      RECT 326.66 7908.935 2313.83 7909.475 ;
      RECT 326.66 7895.045 2313.83 7901.705 ;
      RECT 326.66 7891.925 2313.83 7892.465 ;
      RECT 326.66 7885.315 2313.83 7885.855 ;
      RECT 326.66 7874.095 2313.83 7874.635 ;
      RECT 326.66 7867.485 2313.83 7868.025 ;
      RECT 326.66 7858.245 2313.83 7864.905 ;
      RECT 326.66 7850.475 2313.83 7851.015 ;
      RECT 326.66 7836.935 2313.83 7837.475 ;
      RECT 326.66 7823.045 2313.83 7829.705 ;
      RECT 326.66 7819.925 2313.83 7820.465 ;
      RECT 326.66 7813.315 2313.83 7813.855 ;
      RECT 326.66 7802.095 2313.83 7802.635 ;
      RECT 326.66 7795.485 2313.83 7796.025 ;
      RECT 326.66 7786.245 2313.83 7792.905 ;
      RECT 326.66 7778.475 2313.83 7779.015 ;
      RECT 326.66 7764.935 2313.83 7765.475 ;
      RECT 326.66 7751.045 2313.83 7757.705 ;
      RECT 326.66 7747.925 2313.83 7748.465 ;
      RECT 326.66 7741.315 2313.83 7741.855 ;
      RECT 326.66 7730.095 2313.83 7730.635 ;
      RECT 326.66 7723.485 2313.83 7724.025 ;
      RECT 326.66 7714.245 2313.83 7720.905 ;
      RECT 326.66 7706.475 2313.83 7707.015 ;
      RECT 326.66 7692.935 2313.83 7693.475 ;
      RECT 326.66 7679.045 2313.83 7685.705 ;
      RECT 326.66 7675.925 2313.83 7676.465 ;
      RECT 326.66 7669.315 2313.83 7669.855 ;
      RECT 326.66 7658.095 2313.83 7658.635 ;
      RECT 326.66 7651.485 2313.83 7652.025 ;
      RECT 326.66 7642.245 2313.83 7648.905 ;
      RECT 326.66 7634.475 2313.83 7635.015 ;
      RECT 326.66 7620.935 2313.83 7621.475 ;
      RECT 326.66 7607.045 2313.83 7613.705 ;
      RECT 326.66 7603.925 2313.83 7604.465 ;
      RECT 326.66 7597.315 2313.83 7597.855 ;
      RECT 326.66 7586.095 2313.83 7586.635 ;
      RECT 326.66 7579.485 2313.83 7580.025 ;
      RECT 326.66 7570.245 2313.83 7576.905 ;
      RECT 326.66 7562.475 2313.83 7563.015 ;
      RECT 326.66 7548.935 2313.83 7549.475 ;
      RECT 326.66 7535.045 2313.83 7541.705 ;
      RECT 326.66 7531.925 2313.83 7532.465 ;
      RECT 326.66 7525.315 2313.83 7525.855 ;
      RECT 326.66 7514.095 2313.83 7514.635 ;
      RECT 326.66 7507.485 2313.83 7508.025 ;
      RECT 326.66 7498.245 2313.83 7504.905 ;
      RECT 326.66 7490.475 2313.83 7491.015 ;
      RECT 326.66 7476.935 2313.83 7477.475 ;
      RECT 326.66 7463.045 2313.83 7469.705 ;
      RECT 326.66 7459.925 2313.83 7460.465 ;
      RECT 326.66 7453.315 2313.83 7453.855 ;
      RECT 326.66 7442.095 2313.83 7442.635 ;
      RECT 326.66 7435.485 2313.83 7436.025 ;
      RECT 326.66 7426.245 2313.83 7432.905 ;
      RECT 326.66 7418.475 2313.83 7419.015 ;
      RECT 326.66 7404.935 2313.83 7405.475 ;
      RECT 326.66 7391.045 2313.83 7397.705 ;
      RECT 326.66 7387.925 2313.83 7388.465 ;
      RECT 326.66 7381.315 2313.83 7381.855 ;
      RECT 326.66 7370.095 2313.83 7370.635 ;
      RECT 326.66 7363.485 2313.83 7364.025 ;
      RECT 326.66 7354.245 2313.83 7360.905 ;
      RECT 326.66 7346.475 2313.83 7347.015 ;
      RECT 326.66 7332.935 2313.83 7333.475 ;
      RECT 326.66 7319.045 2313.83 7325.705 ;
      RECT 326.66 7315.925 2313.83 7316.465 ;
      RECT 326.66 7309.315 2313.83 7309.855 ;
      RECT 326.66 7298.095 2313.83 7298.635 ;
      RECT 326.66 7291.485 2313.83 7292.025 ;
      RECT 326.66 7282.245 2313.83 7288.905 ;
      RECT 326.66 7274.475 2313.83 7275.015 ;
      RECT 326.66 7260.935 2313.83 7261.475 ;
      RECT 326.66 7247.045 2313.83 7253.705 ;
      RECT 326.66 7243.925 2313.83 7244.465 ;
      RECT 326.66 7237.315 2313.83 7237.855 ;
      RECT 326.66 7226.095 2313.83 7226.635 ;
      RECT 326.66 7219.485 2313.83 7220.025 ;
      RECT 326.66 7210.245 2313.83 7216.905 ;
      RECT 326.66 7202.475 2313.83 7203.015 ;
      RECT 326.66 7188.935 2313.83 7189.475 ;
      RECT 326.66 7175.045 2313.83 7181.705 ;
      RECT 326.66 7171.925 2313.83 7172.465 ;
      RECT 326.66 7165.315 2313.83 7165.855 ;
      RECT 326.66 7154.095 2313.83 7154.635 ;
      RECT 326.66 7147.485 2313.83 7148.025 ;
      RECT 326.66 7138.245 2313.83 7144.905 ;
      RECT 326.66 7130.475 2313.83 7131.015 ;
      RECT 326.66 7116.935 2313.83 7117.475 ;
      RECT 326.66 7103.045 2313.83 7109.705 ;
      RECT 326.66 7099.925 2313.83 7100.465 ;
      RECT 326.66 7093.315 2313.83 7093.855 ;
      RECT 326.66 7082.095 2313.83 7082.635 ;
      RECT 326.66 7075.485 2313.83 7076.025 ;
      RECT 326.66 7066.245 2313.83 7072.905 ;
      RECT 326.66 7058.475 2313.83 7059.015 ;
      RECT 326.66 7044.935 2313.83 7045.475 ;
      RECT 326.66 7031.045 2313.83 7037.705 ;
      RECT 326.66 7027.925 2313.83 7028.465 ;
      RECT 326.66 7021.315 2313.83 7021.855 ;
      RECT 326.66 7010.095 2313.83 7010.635 ;
      RECT 326.66 7003.485 2313.83 7004.025 ;
      RECT 326.66 6994.245 2313.83 7000.905 ;
      RECT 326.66 6986.475 2313.83 6987.015 ;
      RECT 326.66 6972.935 2313.83 6973.475 ;
      RECT 326.66 6959.045 2313.83 6965.705 ;
      RECT 326.66 6955.925 2313.83 6956.465 ;
      RECT 326.66 6949.315 2313.83 6949.855 ;
      RECT 326.66 6938.095 2313.83 6938.635 ;
      RECT 326.66 6931.485 2313.83 6932.025 ;
      RECT 326.66 6922.245 2313.83 6928.905 ;
      RECT 326.66 6914.475 2313.83 6915.015 ;
      RECT 326.66 6900.935 2313.83 6901.475 ;
      RECT 326.66 6887.045 2313.83 6893.705 ;
      RECT 326.66 6883.925 2313.83 6884.465 ;
      RECT 326.66 6877.315 2313.83 6877.855 ;
      RECT 326.66 6866.095 2313.83 6866.635 ;
      RECT 326.66 6859.485 2313.83 6860.025 ;
      RECT 326.66 6850.245 2313.83 6856.905 ;
      RECT 326.66 6842.475 2313.83 6843.015 ;
      RECT 326.66 6828.935 2313.83 6829.475 ;
      RECT 326.66 6815.045 2313.83 6821.705 ;
      RECT 326.66 6811.925 2313.83 6812.465 ;
      RECT 326.66 6805.315 2313.83 6805.855 ;
      RECT 326.66 6794.095 2313.83 6794.635 ;
      RECT 326.66 6787.485 2313.83 6788.025 ;
      RECT 326.66 6778.245 2313.83 6784.905 ;
      RECT 326.66 6770.475 2313.83 6771.015 ;
      RECT 326.66 6756.935 2313.83 6757.475 ;
      RECT 326.66 6743.045 2313.83 6749.705 ;
      RECT 326.66 6739.925 2313.83 6740.465 ;
      RECT 326.66 6733.315 2313.83 6733.855 ;
      RECT 326.66 6722.095 2313.83 6722.635 ;
      RECT 326.66 6715.485 2313.83 6716.025 ;
      RECT 326.66 6706.245 2313.83 6712.905 ;
      RECT 326.66 6698.475 2313.83 6699.015 ;
      RECT 326.66 6684.935 2313.83 6685.475 ;
      RECT 326.66 6671.045 2313.83 6677.705 ;
      RECT 326.66 6667.925 2313.83 6668.465 ;
      RECT 326.66 6661.315 2313.83 6661.855 ;
      RECT 326.66 6650.095 2313.83 6650.635 ;
      RECT 326.66 6643.485 2313.83 6644.025 ;
      RECT 326.66 6634.245 2313.83 6640.905 ;
      RECT 326.66 6626.475 2313.83 6627.015 ;
      RECT 326.66 6612.935 2313.83 6613.475 ;
      RECT 326.66 6599.045 2313.83 6605.705 ;
      RECT 326.66 6595.925 2313.83 6596.465 ;
      RECT 326.66 6589.315 2313.83 6589.855 ;
      RECT 326.66 6578.095 2313.83 6578.635 ;
      RECT 326.66 6571.485 2313.83 6572.025 ;
      RECT 326.66 6562.245 2313.83 6568.905 ;
      RECT 326.66 6554.475 2313.83 6555.015 ;
      RECT 326.66 6540.935 2313.83 6541.475 ;
      RECT 326.66 6527.045 2313.83 6533.705 ;
      RECT 326.66 6523.925 2313.83 6524.465 ;
      RECT 326.66 6517.315 2313.83 6517.855 ;
      RECT 326.66 6506.095 2313.83 6506.635 ;
      RECT 326.66 6499.485 2313.83 6500.025 ;
      RECT 326.66 6490.245 2313.83 6496.905 ;
      RECT 326.66 6482.475 2313.83 6483.015 ;
      RECT 326.66 6468.935 2313.83 6469.475 ;
      RECT 326.66 6455.045 2313.83 6461.705 ;
      RECT 326.66 6451.925 2313.83 6452.465 ;
      RECT 326.66 6445.315 2313.83 6445.855 ;
      RECT 326.66 6434.095 2313.83 6434.635 ;
      RECT 326.66 6427.485 2313.83 6428.025 ;
      RECT 326.66 6418.245 2313.83 6424.905 ;
      RECT 326.66 6410.475 2313.83 6411.015 ;
      RECT 326.66 6396.935 2313.83 6397.475 ;
      RECT 326.66 6383.045 2313.83 6389.705 ;
      RECT 326.66 6379.925 2313.83 6380.465 ;
      RECT 326.66 6373.315 2313.83 6373.855 ;
      RECT 326.66 6362.095 2313.83 6362.635 ;
      RECT 326.66 6355.485 2313.83 6356.025 ;
      RECT 326.66 6346.245 2313.83 6352.905 ;
      RECT 326.66 6338.475 2313.83 6339.015 ;
      RECT 326.66 6324.935 2313.83 6325.475 ;
      RECT 326.66 6311.045 2313.83 6317.705 ;
      RECT 326.66 6307.925 2313.83 6308.465 ;
      RECT 326.66 6301.315 2313.83 6301.855 ;
      RECT 326.66 6290.095 2313.83 6290.635 ;
      RECT 326.66 6283.485 2313.83 6284.025 ;
      RECT 326.66 6274.245 2313.83 6280.905 ;
      RECT 326.66 6266.475 2313.83 6267.015 ;
      RECT 326.66 6252.935 2313.83 6253.475 ;
      RECT 326.66 6239.045 2313.83 6245.705 ;
      RECT 326.66 6235.925 2313.83 6236.465 ;
      RECT 326.66 6229.315 2313.83 6229.855 ;
      RECT 326.66 6218.095 2313.83 6218.635 ;
      RECT 326.66 6211.485 2313.83 6212.025 ;
      RECT 326.66 6202.245 2313.83 6208.905 ;
      RECT 326.66 6194.475 2313.83 6195.015 ;
      RECT 326.66 6180.935 2313.83 6181.475 ;
      RECT 326.66 6167.045 2313.83 6173.705 ;
      RECT 326.66 6163.925 2313.83 6164.465 ;
      RECT 326.66 6157.315 2313.83 6157.855 ;
      RECT 326.66 6146.095 2313.83 6146.635 ;
      RECT 326.66 6139.485 2313.83 6140.025 ;
      RECT 326.66 6130.245 2313.83 6136.905 ;
      RECT 326.66 6122.475 2313.83 6123.015 ;
      RECT 326.66 6108.935 2313.83 6109.475 ;
      RECT 326.66 6095.045 2313.83 6101.705 ;
      RECT 326.66 6091.925 2313.83 6092.465 ;
      RECT 326.66 6085.315 2313.83 6085.855 ;
      RECT 326.66 6074.095 2313.83 6074.635 ;
      RECT 326.66 6067.485 2313.83 6068.025 ;
      RECT 326.66 6058.245 2313.83 6064.905 ;
      RECT 326.66 6050.475 2313.83 6051.015 ;
      RECT 326.66 6036.935 2313.83 6037.475 ;
      RECT 326.66 6023.045 2313.83 6029.705 ;
      RECT 326.66 6019.925 2313.83 6020.465 ;
      RECT 326.66 6013.315 2313.83 6013.855 ;
      RECT 326.66 6002.095 2313.83 6002.635 ;
      RECT 326.66 5995.485 2313.83 5996.025 ;
      RECT 326.66 5986.245 2313.83 5992.905 ;
      RECT 326.66 5978.475 2313.83 5979.015 ;
      RECT 326.66 5964.935 2313.83 5965.475 ;
      RECT 326.66 5951.045 2313.83 5957.705 ;
      RECT 326.66 5947.925 2313.83 5948.465 ;
      RECT 326.66 5941.315 2313.83 5941.855 ;
      RECT 326.66 5930.095 2313.83 5930.635 ;
      RECT 326.66 5923.485 2313.83 5924.025 ;
      RECT 326.66 5914.245 2313.83 5920.905 ;
      RECT 326.66 5906.475 2313.83 5907.015 ;
      RECT 326.66 5892.935 2313.83 5893.475 ;
      RECT 326.66 5879.045 2313.83 5885.705 ;
      RECT 326.66 5875.925 2313.83 5876.465 ;
      RECT 326.66 5869.315 2313.83 5869.855 ;
      RECT 326.66 5858.095 2313.83 5858.635 ;
      RECT 326.66 5851.485 2313.83 5852.025 ;
      RECT 326.66 5842.245 2313.83 5848.905 ;
      RECT 326.66 5834.475 2313.83 5835.015 ;
      RECT 326.66 5820.935 2313.83 5821.475 ;
      RECT 326.66 5807.045 2313.83 5813.705 ;
      RECT 326.66 5803.925 2313.83 5804.465 ;
      RECT 326.66 5797.315 2313.83 5797.855 ;
      RECT 326.66 5786.095 2313.83 5786.635 ;
      RECT 326.66 5779.485 2313.83 5780.025 ;
      RECT 326.66 5770.245 2313.83 5776.905 ;
      RECT 326.66 5762.475 2313.83 5763.015 ;
      RECT 326.66 5748.935 2313.83 5749.475 ;
      RECT 326.66 5735.045 2313.83 5741.705 ;
      RECT 326.66 5731.925 2313.83 5732.465 ;
      RECT 326.66 5725.315 2313.83 5725.855 ;
      RECT 326.66 5714.095 2313.83 5714.635 ;
      RECT 326.66 5707.485 2313.83 5708.025 ;
      RECT 326.66 5698.245 2313.83 5704.905 ;
      RECT 326.66 5690.475 2313.83 5691.015 ;
      RECT 326.66 5676.935 2313.83 5677.475 ;
      RECT 326.66 5663.045 2313.83 5669.705 ;
      RECT 326.66 5659.925 2313.83 5660.465 ;
      RECT 326.66 5653.315 2313.83 5653.855 ;
      RECT 326.66 5642.095 2313.83 5642.635 ;
      RECT 326.66 5635.485 2313.83 5636.025 ;
      RECT 326.66 5626.245 2313.83 5632.905 ;
      RECT 326.66 5618.475 2313.83 5619.015 ;
      RECT 326.66 5604.935 2313.83 5605.475 ;
      RECT 326.66 5591.045 2313.83 5597.705 ;
      RECT 326.66 5587.925 2313.83 5588.465 ;
      RECT 326.66 5581.315 2313.83 5581.855 ;
      RECT 326.66 5570.095 2313.83 5570.635 ;
      RECT 326.66 5563.485 2313.83 5564.025 ;
      RECT 326.66 5554.245 2313.83 5560.905 ;
      RECT 326.66 5546.475 2313.83 5547.015 ;
      RECT 326.66 5532.935 2313.83 5533.475 ;
      RECT 326.66 5519.045 2313.83 5525.705 ;
      RECT 326.66 5515.925 2313.83 5516.465 ;
      RECT 326.66 5509.315 2313.83 5509.855 ;
      RECT 326.66 5498.095 2313.83 5498.635 ;
      RECT 326.66 5491.485 2313.83 5492.025 ;
      RECT 326.66 5482.245 2313.83 5488.905 ;
      RECT 326.66 5474.475 2313.83 5475.015 ;
      RECT 326.66 5460.935 2313.83 5461.475 ;
      RECT 326.66 5447.045 2313.83 5453.705 ;
      RECT 326.66 5443.925 2313.83 5444.465 ;
      RECT 326.66 5437.315 2313.83 5437.855 ;
      RECT 326.66 5426.095 2313.83 5426.635 ;
      RECT 326.66 5419.485 2313.83 5420.025 ;
      RECT 326.66 5410.245 2313.83 5416.905 ;
      RECT 326.66 5402.475 2313.83 5403.015 ;
      RECT 326.66 5388.935 2313.83 5389.475 ;
      RECT 326.66 5375.045 2313.83 5381.705 ;
      RECT 326.66 5371.925 2313.83 5372.465 ;
      RECT 326.66 5365.315 2313.83 5365.855 ;
      RECT 326.66 5354.095 2313.83 5354.635 ;
      RECT 326.66 5347.485 2313.83 5348.025 ;
      RECT 326.66 5338.245 2313.83 5344.905 ;
      RECT 326.66 5330.475 2313.83 5331.015 ;
      RECT 326.66 5316.935 2313.83 5317.475 ;
      RECT 326.66 5303.045 2313.83 5309.705 ;
      RECT 326.66 5299.925 2313.83 5300.465 ;
      RECT 326.66 5293.315 2313.83 5293.855 ;
      RECT 326.66 5282.095 2313.83 5282.635 ;
      RECT 326.66 5275.485 2313.83 5276.025 ;
      RECT 326.66 5266.245 2313.83 5272.905 ;
      RECT 326.66 5258.475 2313.83 5259.015 ;
      RECT 326.66 5244.935 2313.83 5245.475 ;
      RECT 326.66 5231.045 2313.83 5237.705 ;
      RECT 326.66 5227.925 2313.83 5228.465 ;
      RECT 326.66 5221.315 2313.83 5221.855 ;
      RECT 326.66 5210.095 2313.83 5210.635 ;
      RECT 326.66 5203.485 2313.83 5204.025 ;
      RECT 326.66 5194.245 2313.83 5200.905 ;
      RECT 326.66 5186.475 2313.83 5187.015 ;
      RECT 326.66 5172.935 2313.83 5173.475 ;
      RECT 326.66 5159.045 2313.83 5165.705 ;
      RECT 326.66 5155.925 2313.83 5156.465 ;
      RECT 326.66 5149.315 2313.83 5149.855 ;
      RECT 326.66 5138.095 2313.83 5138.635 ;
      RECT 326.66 5131.485 2313.83 5132.025 ;
      RECT 326.66 5122.245 2313.83 5128.905 ;
      RECT 326.66 5114.475 2313.83 5115.015 ;
      RECT 326.66 5100.935 2313.83 5101.475 ;
      RECT 326.66 5087.045 2313.83 5093.705 ;
      RECT 326.66 5083.925 2313.83 5084.465 ;
      RECT 326.66 5077.315 2313.83 5077.855 ;
      RECT 326.66 5066.095 2313.83 5066.635 ;
      RECT 326.66 5059.485 2313.83 5060.025 ;
      RECT 326.66 5050.245 2313.83 5056.905 ;
      RECT 326.66 5042.475 2313.83 5043.015 ;
      RECT 326.66 5028.935 2313.83 5029.475 ;
      RECT 326.66 5015.045 2313.83 5021.705 ;
      RECT 326.66 5011.925 2313.83 5012.465 ;
      RECT 326.66 5005.315 2313.83 5005.855 ;
      RECT 326.66 4994.095 2313.83 4994.635 ;
      RECT 326.66 4987.485 2313.83 4988.025 ;
      RECT 326.66 4978.245 2313.83 4984.905 ;
      RECT 326.66 4970.475 2313.83 4971.015 ;
      RECT 326.66 4956.935 2313.83 4957.475 ;
      RECT 326.66 4943.045 2313.83 4949.705 ;
      RECT 326.66 4939.925 2313.83 4940.465 ;
      RECT 326.66 4933.315 2313.83 4933.855 ;
      RECT 326.66 4922.095 2313.83 4922.635 ;
      RECT 326.66 4915.485 2313.83 4916.025 ;
      RECT 326.66 4906.245 2313.83 4912.905 ;
      RECT 326.66 4898.475 2313.83 4899.015 ;
      RECT 326.66 4884.935 2313.83 4885.475 ;
      RECT 326.66 4871.045 2313.83 4877.705 ;
      RECT 326.66 4867.925 2313.83 4868.465 ;
      RECT 326.66 4861.315 2313.83 4861.855 ;
      RECT 326.66 4850.095 2313.83 4850.635 ;
      RECT 326.66 4843.485 2313.83 4844.025 ;
      RECT 326.66 4834.245 2313.83 4840.905 ;
      RECT 326.66 4826.475 2313.83 4827.015 ;
      RECT 326.66 4812.935 2313.83 4813.475 ;
      RECT 326.66 4799.045 2313.83 4805.705 ;
      RECT 326.66 4795.925 2313.83 4796.465 ;
      RECT 326.66 4789.315 2313.83 4789.855 ;
      RECT 326.66 4778.095 2313.83 4778.635 ;
      RECT 326.66 4771.485 2313.83 4772.025 ;
      RECT 326.66 4762.245 2313.83 4768.905 ;
      RECT 326.66 4754.475 2313.83 4755.015 ;
      RECT 326.66 4740.935 2313.83 4741.475 ;
      RECT 326.66 4727.045 2313.83 4733.705 ;
      RECT 326.66 4723.925 2313.83 4724.465 ;
      RECT 326.66 4717.315 2313.83 4717.855 ;
      RECT 326.66 4706.095 2313.83 4706.635 ;
      RECT 326.66 4699.485 2313.83 4700.025 ;
      RECT 326.66 4690.245 2313.83 4696.905 ;
      RECT 326.66 4682.475 2313.83 4683.015 ;
      RECT 326.66 4668.935 2313.83 4669.475 ;
      RECT 326.66 4655.045 2313.83 4661.705 ;
      RECT 326.66 4651.925 2313.83 4652.465 ;
      RECT 326.66 4645.315 2313.83 4645.855 ;
      RECT 326.66 4634.095 2313.83 4634.635 ;
      RECT 326.66 4627.485 2313.83 4628.025 ;
      RECT 326.66 4618.245 2313.83 4624.905 ;
      RECT 326.66 4610.475 2313.83 4611.015 ;
      RECT 326.66 4596.935 2313.83 4597.475 ;
      RECT 326.66 4583.045 2313.83 4589.705 ;
      RECT 326.66 4579.925 2313.83 4580.465 ;
      RECT 326.66 4573.315 2313.83 4573.855 ;
      RECT 326.66 4562.095 2313.83 4562.635 ;
      RECT 326.66 4555.485 2313.83 4556.025 ;
      RECT 326.66 4546.245 2313.83 4552.905 ;
      RECT 326.66 4538.475 2313.83 4539.015 ;
      RECT 326.66 4524.935 2313.83 4525.475 ;
      RECT 326.66 4511.045 2313.83 4517.705 ;
      RECT 326.66 4507.925 2313.83 4508.465 ;
      RECT 326.66 4501.315 2313.83 4501.855 ;
      RECT 326.66 4490.095 2313.83 4490.635 ;
      RECT 326.66 4483.485 2313.83 4484.025 ;
      RECT 326.66 4474.245 2313.83 4480.905 ;
      RECT 326.66 4466.475 2313.83 4467.015 ;
      RECT 326.66 4452.935 2313.83 4453.475 ;
      RECT 326.66 4439.045 2313.83 4445.705 ;
      RECT 326.66 4435.925 2313.83 4436.465 ;
      RECT 326.66 4429.315 2313.83 4429.855 ;
      RECT 326.66 4418.095 2313.83 4418.635 ;
      RECT 326.66 4411.485 2313.83 4412.025 ;
      RECT 326.66 4402.245 2313.83 4408.905 ;
      RECT 326.66 4394.475 2313.83 4395.015 ;
      RECT 326.66 4380.935 2313.83 4381.475 ;
      RECT 326.66 4367.045 2313.83 4373.705 ;
      RECT 326.66 4363.925 2313.83 4364.465 ;
      RECT 326.66 4357.315 2313.83 4357.855 ;
      RECT 326.66 4346.095 2313.83 4346.635 ;
      RECT 326.66 4339.485 2313.83 4340.025 ;
      RECT 326.66 4330.245 2313.83 4336.905 ;
      RECT 326.66 4322.475 2313.83 4323.015 ;
      RECT 326.66 4308.935 2313.83 4309.475 ;
      RECT 326.66 4295.045 2313.83 4301.705 ;
      RECT 326.66 4291.925 2313.83 4292.465 ;
      RECT 326.66 4285.315 2313.83 4285.855 ;
      RECT 326.66 4274.095 2313.83 4274.635 ;
      RECT 326.66 4267.485 2313.83 4268.025 ;
      RECT 326.66 4258.245 2313.83 4264.905 ;
      RECT 326.66 4250.475 2313.83 4251.015 ;
      RECT 326.66 4236.935 2313.83 4237.475 ;
      RECT 326.66 4223.045 2313.83 4229.705 ;
      RECT 326.66 4219.925 2313.83 4220.465 ;
      RECT 326.66 4213.315 2313.83 4213.855 ;
      RECT 326.66 4202.095 2313.83 4202.635 ;
      RECT 326.66 4195.485 2313.83 4196.025 ;
      RECT 326.66 4186.245 2313.83 4192.905 ;
      RECT 326.66 4178.475 2313.83 4179.015 ;
      RECT 326.66 4164.935 2313.83 4165.475 ;
      RECT 326.66 4151.045 2313.83 4157.705 ;
      RECT 326.66 4147.925 2313.83 4148.465 ;
      RECT 326.66 4141.315 2313.83 4141.855 ;
      RECT 326.66 4130.095 2313.83 4130.635 ;
      RECT 326.66 4123.485 2313.83 4124.025 ;
      RECT 326.66 4114.245 2313.83 4120.905 ;
      RECT 326.66 4106.475 2313.83 4107.015 ;
      RECT 326.66 4092.935 2313.83 4093.475 ;
      RECT 326.66 4079.045 2313.83 4085.705 ;
      RECT 326.66 4075.925 2313.83 4076.465 ;
      RECT 326.66 4069.315 2313.83 4069.855 ;
      RECT 326.66 4058.095 2313.83 4058.635 ;
      RECT 326.66 4051.485 2313.83 4052.025 ;
      RECT 326.66 4042.245 2313.83 4048.905 ;
      RECT 326.66 4034.475 2313.83 4035.015 ;
      RECT 326.66 4020.935 2313.83 4021.475 ;
      RECT 326.66 4007.045 2313.83 4013.705 ;
      RECT 326.66 4003.925 2313.83 4004.465 ;
      RECT 326.66 3997.315 2313.83 3997.855 ;
      RECT 326.66 3986.095 2313.83 3986.635 ;
      RECT 326.66 3979.485 2313.83 3980.025 ;
      RECT 326.66 3970.245 2313.83 3976.905 ;
      RECT 326.66 3962.475 2313.83 3963.015 ;
      RECT 326.66 3948.935 2313.83 3949.475 ;
      RECT 326.66 3935.045 2313.83 3941.705 ;
      RECT 326.66 3931.925 2313.83 3932.465 ;
      RECT 326.66 3925.315 2313.83 3925.855 ;
      RECT 326.66 3914.095 2313.83 3914.635 ;
      RECT 326.66 3907.485 2313.83 3908.025 ;
      RECT 326.66 3898.245 2313.83 3904.905 ;
      RECT 326.66 3890.475 2313.83 3891.015 ;
      RECT 326.66 3876.935 2313.83 3877.475 ;
      RECT 326.66 3863.045 2313.83 3869.705 ;
      RECT 326.66 3859.925 2313.83 3860.465 ;
      RECT 326.66 3853.315 2313.83 3853.855 ;
      RECT 326.66 3842.095 2313.83 3842.635 ;
      RECT 326.66 3835.485 2313.83 3836.025 ;
      RECT 326.66 3826.245 2313.83 3832.905 ;
      RECT 326.66 3818.475 2313.83 3819.015 ;
      RECT 326.66 3804.935 2313.83 3805.475 ;
      RECT 326.66 3791.045 2313.83 3797.705 ;
      RECT 326.66 3787.925 2313.83 3788.465 ;
      RECT 326.66 3781.315 2313.83 3781.855 ;
      RECT 326.66 3770.095 2313.83 3770.635 ;
      RECT 326.66 3763.485 2313.83 3764.025 ;
      RECT 326.66 3754.245 2313.83 3760.905 ;
      RECT 326.66 3746.475 2313.83 3747.015 ;
      RECT 326.66 3732.935 2313.83 3733.475 ;
      RECT 326.66 3719.045 2313.83 3725.705 ;
      RECT 326.66 3715.925 2313.83 3716.465 ;
      RECT 326.66 3709.315 2313.83 3709.855 ;
      RECT 326.66 3698.095 2313.83 3698.635 ;
      RECT 326.66 3691.485 2313.83 3692.025 ;
      RECT 326.66 3682.245 2313.83 3688.905 ;
      RECT 326.66 3674.475 2313.83 3675.015 ;
      RECT 326.66 3660.935 2313.83 3661.475 ;
      RECT 326.66 3647.045 2313.83 3653.705 ;
      RECT 326.66 3643.925 2313.83 3644.465 ;
      RECT 326.66 3637.315 2313.83 3637.855 ;
      RECT 326.66 3626.095 2313.83 3626.635 ;
      RECT 326.66 3619.485 2313.83 3620.025 ;
      RECT 326.66 3610.245 2313.83 3616.905 ;
      RECT 326.66 3602.475 2313.83 3603.015 ;
      RECT 326.66 3588.935 2313.83 3589.475 ;
      RECT 326.66 3575.045 2313.83 3581.705 ;
      RECT 326.66 3571.925 2313.83 3572.465 ;
      RECT 326.66 3565.315 2313.83 3565.855 ;
      RECT 326.66 3554.095 2313.83 3554.635 ;
      RECT 326.66 3547.485 2313.83 3548.025 ;
      RECT 326.66 3538.245 2313.83 3544.905 ;
      RECT 326.66 3530.475 2313.83 3531.015 ;
      RECT 326.66 3516.935 2313.83 3517.475 ;
      RECT 326.66 3503.045 2313.83 3509.705 ;
      RECT 326.66 3499.925 2313.83 3500.465 ;
      RECT 326.66 3493.315 2313.83 3493.855 ;
      RECT 326.66 3482.095 2313.83 3482.635 ;
      RECT 326.66 3475.485 2313.83 3476.025 ;
      RECT 326.66 3466.245 2313.83 3472.905 ;
      RECT 326.66 3458.475 2313.83 3459.015 ;
      RECT 326.66 3444.935 2313.83 3445.475 ;
      RECT 326.66 3431.045 2313.83 3437.705 ;
      RECT 326.66 3427.925 2313.83 3428.465 ;
      RECT 326.66 3421.315 2313.83 3421.855 ;
      RECT 326.66 3410.095 2313.83 3410.635 ;
      RECT 326.66 3403.485 2313.83 3404.025 ;
      RECT 326.66 3394.245 2313.83 3400.905 ;
      RECT 326.66 3386.475 2313.83 3387.015 ;
      RECT 326.66 3372.935 2313.83 3373.475 ;
      RECT 326.66 3359.045 2313.83 3365.705 ;
      RECT 326.66 3355.925 2313.83 3356.465 ;
      RECT 326.66 3349.315 2313.83 3349.855 ;
      RECT 326.66 3338.095 2313.83 3338.635 ;
      RECT 326.66 3331.485 2313.83 3332.025 ;
      RECT 326.66 3322.245 2313.83 3328.905 ;
      RECT 326.66 3314.475 2313.83 3315.015 ;
      RECT 326.66 3300.935 2313.83 3301.475 ;
      RECT 326.66 3287.045 2313.83 3293.705 ;
      RECT 326.66 3283.925 2313.83 3284.465 ;
      RECT 326.66 3277.315 2313.83 3277.855 ;
      RECT 326.66 3266.095 2313.83 3266.635 ;
      RECT 326.66 3259.485 2313.83 3260.025 ;
      RECT 326.66 3250.245 2313.83 3256.905 ;
      RECT 326.66 3242.475 2313.83 3243.015 ;
      RECT 326.66 3228.935 2313.83 3229.475 ;
      RECT 326.66 3215.045 2313.83 3221.705 ;
      RECT 326.66 3211.925 2313.83 3212.465 ;
      RECT 326.66 3205.315 2313.83 3205.855 ;
      RECT 326.66 3194.095 2313.83 3194.635 ;
      RECT 326.66 3187.485 2313.83 3188.025 ;
      RECT 326.66 3178.245 2313.83 3184.905 ;
      RECT 326.66 3170.475 2313.83 3171.015 ;
      RECT 326.66 3156.935 2313.83 3157.475 ;
      RECT 326.66 3143.045 2313.83 3149.705 ;
      RECT 326.66 3139.925 2313.83 3140.465 ;
      RECT 326.66 3133.315 2313.83 3133.855 ;
      RECT 326.66 3122.095 2313.83 3122.635 ;
      RECT 326.66 3115.485 2313.83 3116.025 ;
      RECT 326.66 3106.245 2313.83 3112.905 ;
      RECT 326.66 3098.475 2313.83 3099.015 ;
      RECT 326.66 3084.935 2313.83 3085.475 ;
      RECT 326.66 3071.045 2313.83 3077.705 ;
      RECT 326.66 3067.925 2313.83 3068.465 ;
      RECT 326.66 3061.315 2313.83 3061.855 ;
      RECT 326.66 3050.095 2313.83 3050.635 ;
      RECT 326.66 3043.485 2313.83 3044.025 ;
      RECT 326.66 3034.245 2313.83 3040.905 ;
      RECT 326.66 3026.475 2313.83 3027.015 ;
      RECT 326.66 3012.935 2313.83 3013.475 ;
      RECT 326.66 2999.045 2313.83 3005.705 ;
      RECT 326.66 2995.925 2313.83 2996.465 ;
      RECT 326.66 2989.315 2313.83 2989.855 ;
      RECT 326.66 2978.095 2313.83 2978.635 ;
      RECT 326.66 2971.485 2313.83 2972.025 ;
      RECT 326.66 2962.245 2313.83 2968.905 ;
      RECT 326.66 2954.475 2313.83 2955.015 ;
      RECT 326.66 2940.935 2313.83 2941.475 ;
      RECT 326.66 2927.045 2313.83 2933.705 ;
      RECT 326.66 2923.925 2313.83 2924.465 ;
      RECT 326.66 2917.315 2313.83 2917.855 ;
      RECT 326.66 2906.095 2313.83 2906.635 ;
      RECT 326.66 2899.485 2313.83 2900.025 ;
      RECT 326.66 2890.245 2313.83 2896.905 ;
      RECT 326.66 2882.475 2313.83 2883.015 ;
      RECT 326.66 2868.935 2313.83 2869.475 ;
      RECT 326.66 2855.045 2313.83 2861.705 ;
      RECT 326.66 2851.925 2313.83 2852.465 ;
      RECT 326.66 2845.315 2313.83 2845.855 ;
      RECT 326.66 2834.095 2313.83 2834.635 ;
      RECT 326.66 2827.485 2313.83 2828.025 ;
      RECT 326.66 2818.245 2313.83 2824.905 ;
      RECT 326.66 2810.475 2313.83 2811.015 ;
      RECT 326.66 2796.935 2313.83 2797.475 ;
      RECT 326.66 2783.045 2313.83 2789.705 ;
      RECT 326.66 2779.925 2313.83 2780.465 ;
      RECT 326.66 2773.315 2313.83 2773.855 ;
      RECT 326.66 2762.095 2313.83 2762.635 ;
      RECT 326.66 2755.485 2313.83 2756.025 ;
      RECT 326.66 2746.245 2313.83 2752.905 ;
      RECT 326.66 2738.475 2313.83 2739.015 ;
      RECT 326.66 2724.935 2313.83 2725.475 ;
      RECT 326.66 2711.045 2313.83 2717.705 ;
      RECT 326.66 2707.925 2313.83 2708.465 ;
      RECT 326.66 2701.315 2313.83 2701.855 ;
      RECT 326.66 2690.095 2313.83 2690.635 ;
      RECT 326.66 2683.485 2313.83 2684.025 ;
      RECT 326.66 2674.245 2313.83 2680.905 ;
      RECT 326.66 2666.475 2313.83 2667.015 ;
      RECT 326.66 2652.935 2313.83 2653.475 ;
      RECT 326.66 2639.045 2313.83 2645.705 ;
      RECT 326.66 2635.925 2313.83 2636.465 ;
      RECT 326.66 2629.315 2313.83 2629.855 ;
      RECT 326.66 2618.095 2313.83 2618.635 ;
      RECT 326.66 2611.485 2313.83 2612.025 ;
      RECT 326.66 2602.245 2313.83 2608.905 ;
      RECT 326.66 2594.475 2313.83 2595.015 ;
      RECT 326.66 2580.935 2313.83 2581.475 ;
      RECT 326.66 2567.045 2313.83 2573.705 ;
      RECT 326.66 2563.925 2313.83 2564.465 ;
      RECT 326.66 2557.315 2313.83 2557.855 ;
      RECT 326.66 2546.095 2313.83 2546.635 ;
      RECT 326.66 2539.485 2313.83 2540.025 ;
      RECT 326.66 2530.245 2313.83 2536.905 ;
      RECT 326.66 2522.475 2313.83 2523.015 ;
      RECT 326.66 2508.935 2313.83 2509.475 ;
      RECT 326.66 2495.045 2313.83 2501.705 ;
      RECT 326.66 2491.925 2313.83 2492.465 ;
      RECT 326.66 2485.315 2313.83 2485.855 ;
      RECT 326.66 2474.095 2313.83 2474.635 ;
      RECT 326.66 2467.485 2313.83 2468.025 ;
      RECT 326.66 2458.245 2313.83 2464.905 ;
      RECT 326.66 2450.475 2313.83 2451.015 ;
      RECT 326.66 2436.935 2313.83 2437.475 ;
      RECT 326.66 2423.045 2313.83 2429.705 ;
      RECT 326.66 2419.925 2313.83 2420.465 ;
      RECT 326.66 2413.315 2313.83 2413.855 ;
      RECT 326.66 2402.095 2313.83 2402.635 ;
      RECT 326.66 2395.485 2313.83 2396.025 ;
      RECT 326.66 2386.245 2313.83 2392.905 ;
      RECT 326.66 2378.475 2313.83 2379.015 ;
      RECT 326.66 2364.935 2313.83 2365.475 ;
      RECT 326.66 2351.045 2313.83 2357.705 ;
      RECT 326.66 2347.925 2313.83 2348.465 ;
      RECT 326.66 2341.315 2313.83 2341.855 ;
      RECT 326.66 2330.095 2313.83 2330.635 ;
      RECT 326.66 2323.485 2313.83 2324.025 ;
      RECT 326.66 2314.245 2313.83 2320.905 ;
      RECT 326.66 2306.475 2313.83 2307.015 ;
      RECT 326.66 2292.935 2313.83 2293.475 ;
      RECT 326.66 2279.045 2313.83 2285.705 ;
      RECT 326.66 2275.925 2313.83 2276.465 ;
      RECT 326.66 2269.315 2313.83 2269.855 ;
      RECT 326.66 2258.095 2313.83 2258.635 ;
      RECT 326.66 2251.485 2313.83 2252.025 ;
      RECT 326.66 2242.245 2313.83 2248.905 ;
      RECT 326.66 2234.475 2313.83 2235.015 ;
      RECT 326.66 2220.935 2313.83 2221.475 ;
      RECT 326.66 2207.045 2313.83 2213.705 ;
      RECT 326.66 2203.925 2313.83 2204.465 ;
      RECT 326.66 2197.315 2313.83 2197.855 ;
      RECT 326.66 2186.095 2313.83 2186.635 ;
      RECT 326.66 2179.485 2313.83 2180.025 ;
      RECT 326.66 2170.245 2313.83 2176.905 ;
      RECT 326.66 2162.475 2313.83 2163.015 ;
      RECT 326.66 2148.935 2313.83 2149.475 ;
      RECT 326.66 2135.045 2313.83 2141.705 ;
      RECT 326.66 2131.925 2313.83 2132.465 ;
      RECT 326.66 2125.315 2313.83 2125.855 ;
      RECT 326.66 2114.095 2313.83 2114.635 ;
      RECT 326.66 2107.485 2313.83 2108.025 ;
      RECT 326.66 2098.245 2313.83 2104.905 ;
      RECT 326.66 2090.475 2313.83 2091.015 ;
      RECT 326.66 2076.935 2313.83 2077.475 ;
      RECT 326.66 2063.045 2313.83 2069.705 ;
      RECT 326.66 2059.925 2313.83 2060.465 ;
      RECT 326.66 2053.315 2313.83 2053.855 ;
      RECT 326.66 2042.095 2313.83 2042.635 ;
      RECT 326.66 2035.485 2313.83 2036.025 ;
      RECT 326.66 2026.245 2313.83 2032.905 ;
      RECT 326.66 2018.475 2313.83 2019.015 ;
      RECT 326.66 2004.935 2313.83 2005.475 ;
      RECT 326.66 1991.045 2313.83 1997.705 ;
      RECT 326.66 1987.925 2313.83 1988.465 ;
      RECT 326.66 1981.315 2313.83 1981.855 ;
      RECT 326.66 1970.095 2313.83 1970.635 ;
      RECT 326.66 1963.485 2313.83 1964.025 ;
      RECT 326.66 1954.245 2313.83 1960.905 ;
      RECT 326.66 1946.475 2313.83 1947.015 ;
      RECT 326.66 1932.935 2313.83 1933.475 ;
      RECT 326.66 1919.045 2313.83 1925.705 ;
      RECT 326.66 1915.925 2313.83 1916.465 ;
      RECT 326.66 1909.315 2313.83 1909.855 ;
      RECT 326.66 1898.095 2313.83 1898.635 ;
      RECT 326.66 1891.485 2313.83 1892.025 ;
      RECT 326.66 1882.245 2313.83 1888.905 ;
      RECT 326.66 1874.475 2313.83 1875.015 ;
      RECT 326.66 1860.935 2313.83 1861.475 ;
      RECT 326.66 1847.045 2313.83 1853.705 ;
      RECT 326.66 1843.925 2313.83 1844.465 ;
      RECT 326.66 1837.315 2313.83 1837.855 ;
      RECT 326.66 1826.095 2313.83 1826.635 ;
      RECT 326.66 1819.485 2313.83 1820.025 ;
      RECT 326.66 1810.245 2313.83 1816.905 ;
      RECT 326.66 1802.475 2313.83 1803.015 ;
      RECT 326.66 1788.935 2313.83 1789.475 ;
      RECT 326.66 1775.045 2313.83 1781.705 ;
      RECT 326.66 1771.925 2313.83 1772.465 ;
      RECT 326.66 1765.315 2313.83 1765.855 ;
      RECT 326.66 1754.095 2313.83 1754.635 ;
      RECT 326.66 1747.485 2313.83 1748.025 ;
      RECT 326.66 1738.245 2313.83 1744.905 ;
      RECT 326.66 1730.475 2313.83 1731.015 ;
      RECT 326.66 1716.935 2313.83 1717.475 ;
      RECT 326.66 1703.045 2313.83 1709.705 ;
      RECT 326.66 1699.925 2313.83 1700.465 ;
      RECT 326.66 1693.315 2313.83 1693.855 ;
      RECT 326.66 1682.095 2313.83 1682.635 ;
      RECT 326.66 1675.485 2313.83 1676.025 ;
      RECT 326.66 1666.245 2313.83 1672.905 ;
      RECT 326.66 1658.475 2313.83 1659.015 ;
      RECT 326.66 1644.935 2313.83 1645.475 ;
      RECT 326.66 1631.045 2313.83 1637.705 ;
      RECT 326.66 1627.925 2313.83 1628.465 ;
      RECT 326.66 1621.315 2313.83 1621.855 ;
      RECT 326.66 1610.095 2313.83 1610.635 ;
      RECT 326.66 1603.485 2313.83 1604.025 ;
      RECT 326.66 1594.245 2313.83 1600.905 ;
      RECT 326.66 1586.475 2313.83 1587.015 ;
      RECT 326.66 1572.935 2313.83 1573.475 ;
      RECT 326.66 1559.045 2313.83 1565.705 ;
      RECT 326.66 1555.925 2313.83 1556.465 ;
      RECT 326.66 1549.315 2313.83 1549.855 ;
      RECT 326.66 1538.095 2313.83 1538.635 ;
      RECT 326.66 1531.485 2313.83 1532.025 ;
      RECT 326.66 1522.245 2313.83 1528.905 ;
      RECT 326.66 1514.475 2313.83 1515.015 ;
      RECT 326.66 1500.935 2313.83 1501.475 ;
      RECT 326.66 1487.045 2313.83 1493.705 ;
      RECT 326.66 1483.925 2313.83 1484.465 ;
      RECT 326.66 1477.315 2313.83 1477.855 ;
      RECT 326.66 1466.095 2313.83 1466.635 ;
      RECT 326.66 1459.485 2313.83 1460.025 ;
      RECT 326.66 1450.245 2313.83 1456.905 ;
      RECT 326.66 1442.475 2313.83 1443.015 ;
      RECT 326.66 1428.935 2313.83 1429.475 ;
      RECT 326.66 1415.045 2313.83 1421.705 ;
      RECT 326.66 1411.925 2313.83 1412.465 ;
      RECT 326.66 1405.315 2313.83 1405.855 ;
      RECT 326.66 1394.095 2313.83 1394.635 ;
      RECT 326.66 1387.485 2313.83 1388.025 ;
      RECT 326.66 1378.245 2313.83 1384.905 ;
      RECT 326.66 1370.475 2313.83 1371.015 ;
      RECT 326.66 1356.935 2313.83 1357.475 ;
      RECT 326.66 1343.045 2313.83 1349.705 ;
      RECT 326.66 1339.925 2313.83 1340.465 ;
      RECT 326.66 1333.315 2313.83 1333.855 ;
      RECT 326.66 1322.095 2313.83 1322.635 ;
      RECT 326.66 1315.485 2313.83 1316.025 ;
      RECT 326.66 1306.245 2313.83 1312.905 ;
      RECT 326.66 1298.475 2313.83 1299.015 ;
      RECT 326.66 1284.935 2313.83 1285.475 ;
      RECT 326.66 1271.045 2313.83 1277.705 ;
      RECT 326.66 1267.925 2313.83 1268.465 ;
      RECT 326.66 1261.315 2313.83 1261.855 ;
      RECT 326.66 1250.095 2313.83 1250.635 ;
      RECT 326.66 1243.485 2313.83 1244.025 ;
      RECT 326.66 1234.245 2313.83 1240.905 ;
      RECT 326.66 1226.475 2313.83 1227.015 ;
      RECT 326.66 1212.935 2313.83 1213.475 ;
      RECT 326.66 1199.045 2313.83 1205.705 ;
      RECT 326.66 1195.925 2313.83 1196.465 ;
      RECT 326.66 1189.315 2313.83 1189.855 ;
      RECT 326.66 1178.095 2313.83 1178.635 ;
      RECT 326.66 1171.485 2313.83 1172.025 ;
      RECT 326.66 1162.245 2313.83 1168.905 ;
      RECT 326.66 1154.475 2313.83 1155.015 ;
      RECT 326.66 1140.935 2313.83 1141.475 ;
      RECT 326.66 1127.045 2313.83 1133.705 ;
      RECT 326.66 1123.925 2313.83 1124.465 ;
      RECT 326.66 1117.315 2313.83 1117.855 ;
      RECT 326.66 1106.095 2313.83 1106.635 ;
      RECT 326.66 1099.485 2313.83 1100.025 ;
      RECT 326.66 1090.245 2313.83 1096.905 ;
      RECT 326.66 1082.475 2313.83 1083.015 ;
      RECT 326.66 1068.935 2313.83 1069.475 ;
      RECT 326.66 1055.045 2313.83 1061.705 ;
      RECT 326.66 1051.925 2313.83 1052.465 ;
      RECT 326.66 1045.315 2313.83 1045.855 ;
      RECT 326.66 1034.095 2313.83 1034.635 ;
      RECT 326.66 1027.485 2313.83 1028.025 ;
      RECT 326.66 1018.245 2313.83 1024.905 ;
      RECT 326.66 1010.475 2313.83 1011.015 ;
      RECT 326.66 996.935 2313.83 997.475 ;
      RECT 326.66 983.045 2313.83 989.705 ;
      RECT 326.66 979.925 2313.83 980.465 ;
      RECT 326.66 973.315 2313.83 973.855 ;
      RECT 326.66 962.095 2313.83 962.635 ;
      RECT 326.66 955.485 2313.83 956.025 ;
      RECT 326.66 946.245 2313.83 952.905 ;
      RECT 326.66 938.475 2313.83 939.015 ;
      RECT 326.66 924.935 2313.83 925.475 ;
      RECT 326.66 911.045 2313.83 917.705 ;
      RECT 326.66 907.925 2313.83 908.465 ;
      RECT 326.66 901.315 2313.83 901.855 ;
      RECT 326.66 890.095 2313.83 890.635 ;
      RECT 326.66 883.485 2313.83 884.025 ;
      RECT 326.66 874.245 2313.83 880.905 ;
      RECT 326.66 866.475 2313.83 867.015 ;
      RECT 326.66 852.935 2313.83 853.475 ;
      RECT 326.66 839.045 2313.83 845.705 ;
      RECT 326.66 835.925 2313.83 836.465 ;
      RECT 326.66 829.315 2313.83 829.855 ;
      RECT 326.66 818.095 2313.83 818.635 ;
      RECT 326.66 811.485 2313.83 812.025 ;
      RECT 326.66 802.245 2313.83 808.905 ;
      RECT 326.66 794.475 2313.83 795.015 ;
      RECT 326.66 780.935 2313.83 781.475 ;
      RECT 326.66 767.045 2313.83 773.705 ;
      RECT 326.66 763.925 2313.83 764.465 ;
      RECT 326.66 757.315 2313.83 757.855 ;
      RECT 326.66 746.095 2313.83 746.635 ;
      RECT 326.66 739.485 2313.83 740.025 ;
      RECT 326.66 730.245 2313.83 736.905 ;
      RECT 326.66 722.475 2313.83 723.015 ;
      RECT 326.66 708.935 2313.83 709.475 ;
      RECT 326.66 695.045 2313.83 701.705 ;
      RECT 326.66 691.925 2313.83 692.465 ;
      RECT 326.66 685.315 2313.83 685.855 ;
      RECT 326.66 674.095 2313.83 674.635 ;
      RECT 326.66 667.485 2313.83 668.025 ;
      RECT 326.66 658.245 2313.83 664.905 ;
      RECT 326.66 650.475 2313.83 651.015 ;
      RECT 326.66 636.935 2313.83 637.475 ;
      RECT 326.66 623.045 2313.83 629.705 ;
      RECT 326.66 619.925 2313.83 620.465 ;
      RECT 326.66 613.315 2313.83 613.855 ;
      RECT 326.66 602.095 2313.83 602.635 ;
      RECT 326.66 595.485 2313.83 596.025 ;
      RECT 326.66 586.245 2313.83 592.905 ;
      RECT 326.66 578.475 2313.83 579.015 ;
      RECT 326.66 564.935 2313.83 565.475 ;
      RECT 326.66 551.045 2313.83 557.705 ;
      RECT 326.66 547.925 2313.83 548.465 ;
      RECT 326.66 541.315 2313.83 541.855 ;
      RECT 326.66 523.41 2313.83 535.245 ;
      RECT 326.66 514.995 2313.83 520.83 ;
      RECT 326.66 510.995 2313.83 511.535 ;
      RECT 326.66 324.005 2313.83 499.535 ;
      RECT 326.66 307.005 2313.83 308.515 ;
      RECT 326.66 290.005 2313.83 291.515 ;
      RECT 326.66 228.005 2313.83 229.515 ;
      RECT 326.66 211.005 2313.83 212.515 ;
      RECT 326.66 194.005 2313.83 195.515 ;
      RECT 326.66 187.44 458.31 190.545 ;
      RECT 2295.79 187.44 2298.31 8610.835 ;
      RECT 2278.81 187.44 2281.33 8610.835 ;
      RECT 2263.29 187.44 2264.35 8610.835 ;
      RECT 2232.77 187.44 2233.83 8610.835 ;
      RECT 2215.79 187.44 2218.31 8610.835 ;
      RECT 2198.81 187.44 2201.33 8610.835 ;
      RECT 2183.29 187.44 2184.35 8610.835 ;
      RECT 2152.77 187.44 2153.83 8610.835 ;
      RECT 2135.79 187.44 2138.31 8610.835 ;
      RECT 2118.81 187.44 2121.33 8610.835 ;
      RECT 2103.29 187.44 2104.35 8610.835 ;
      RECT 2072.77 187.44 2073.83 8610.835 ;
      RECT 2055.79 187.44 2058.31 8610.835 ;
      RECT 2038.81 187.44 2041.33 8610.835 ;
      RECT 2023.29 187.44 2024.35 8610.835 ;
      RECT 1992.77 187.44 1993.83 8610.835 ;
      RECT 1975.79 187.44 1978.31 8610.835 ;
      RECT 1958.81 187.44 1961.33 8610.835 ;
      RECT 1943.29 187.44 1944.35 8610.835 ;
      RECT 1912.77 187.44 1913.83 8610.835 ;
      RECT 1895.79 187.44 1898.31 8610.835 ;
      RECT 1878.81 187.44 1881.33 8610.835 ;
      RECT 1863.29 187.44 1864.35 8610.835 ;
      RECT 1832.77 187.44 1833.83 8610.835 ;
      RECT 1815.79 187.44 1818.31 8610.835 ;
      RECT 1798.81 187.44 1801.33 8610.835 ;
      RECT 1783.29 187.44 1784.35 8610.835 ;
      RECT 1752.77 187.44 1753.83 8610.835 ;
      RECT 1735.79 187.44 1738.31 8610.835 ;
      RECT 1718.81 187.44 1721.33 8610.835 ;
      RECT 1703.29 187.44 1704.35 8610.835 ;
      RECT 1672.77 187.44 1673.83 8610.835 ;
      RECT 1655.79 187.44 1658.31 8610.835 ;
      RECT 1638.81 187.44 1641.33 8610.835 ;
      RECT 1623.29 187.44 1624.35 8610.835 ;
      RECT 1592.77 187.44 1593.83 8610.835 ;
      RECT 1575.79 187.44 1578.31 8610.835 ;
      RECT 1558.81 187.44 1561.33 8610.835 ;
      RECT 1543.29 187.44 1544.35 8610.835 ;
      RECT 1512.77 187.44 1513.83 8610.835 ;
      RECT 1495.79 187.44 1498.31 8610.835 ;
      RECT 1478.81 187.44 1481.33 8610.835 ;
      RECT 1463.29 187.44 1464.35 8610.835 ;
      RECT 1432.77 187.44 1433.83 8610.835 ;
      RECT 1415.79 187.44 1418.31 8610.835 ;
      RECT 1398.81 187.44 1401.33 8610.835 ;
      RECT 1383.29 187.44 1384.35 8610.835 ;
      RECT 1352.77 187.44 1353.83 8610.835 ;
      RECT 1335.79 187.44 1338.31 8610.835 ;
      RECT 1318.81 187.44 1321.33 8610.835 ;
      RECT 1303.29 187.44 1304.35 8610.835 ;
      RECT 1272.77 187.44 1273.83 8610.835 ;
      RECT 1255.79 187.44 1258.31 8610.835 ;
      RECT 1238.81 187.44 1241.33 8610.835 ;
      RECT 1223.29 187.44 1224.35 8610.835 ;
      RECT 1192.77 187.44 1193.83 8610.835 ;
      RECT 1175.79 187.44 1178.31 8610.835 ;
      RECT 1158.81 187.44 1161.33 8610.835 ;
      RECT 1143.29 187.44 1144.35 8610.835 ;
      RECT 1112.77 187.44 1113.83 8610.835 ;
      RECT 1095.79 187.44 1098.31 8610.835 ;
      RECT 1078.81 187.44 1081.33 8610.835 ;
      RECT 1063.29 187.44 1064.35 8610.835 ;
      RECT 1032.77 187.44 1033.83 8610.835 ;
      RECT 1015.79 187.44 1018.31 8610.835 ;
      RECT 998.81 187.44 1001.33 8610.835 ;
      RECT 983.29 187.44 984.35 8610.835 ;
      RECT 952.77 187.44 953.83 8610.835 ;
      RECT 935.79 187.44 938.31 8610.835 ;
      RECT 918.81 187.44 921.33 8610.835 ;
      RECT 903.29 187.44 904.35 8610.835 ;
      RECT 872.77 187.44 873.83 8610.835 ;
      RECT 855.79 187.44 858.31 8610.835 ;
      RECT 838.81 187.44 841.33 8610.835 ;
      RECT 823.29 187.44 824.35 8610.835 ;
      RECT 792.77 187.44 793.83 8610.835 ;
      RECT 775.79 187.44 778.31 8610.835 ;
      RECT 758.81 187.44 761.33 8610.835 ;
      RECT 743.29 187.44 744.35 8610.835 ;
      RECT 712.77 187.44 713.83 8610.835 ;
      RECT 695.79 187.44 698.31 8610.835 ;
      RECT 678.81 187.44 681.33 8610.835 ;
      RECT 663.29 187.44 664.35 8610.835 ;
      RECT 632.77 187.44 633.83 8610.835 ;
      RECT 615.79 187.44 618.31 8610.835 ;
      RECT 598.81 187.44 601.33 8610.835 ;
      RECT 583.29 187.44 584.35 8610.835 ;
      RECT 552.77 187.44 553.83 8610.835 ;
      RECT 535.79 187.44 538.31 8610.835 ;
      RECT 518.81 187.44 521.33 8610.835 ;
      RECT 503.29 187.44 504.35 8610.835 ;
      RECT 472.77 187.44 473.83 8610.835 ;
      RECT 18488.73 1561.605 18490.46 1565.705 ;
      RECT 18488.73 1572.935 18490.46 1573.475 ;
      RECT 18488.73 1586.475 18490.46 1587.015 ;
      RECT 18488.73 1594.245 18490.46 1598.345 ;
      RECT 18488.73 1600.365 18490.46 1600.905 ;
      RECT 18488.73 1603.485 18490.46 1604.025 ;
      RECT 18488.73 1610.095 18490.46 1610.635 ;
      RECT 18488.73 1621.315 18490.46 1621.855 ;
      RECT 18488.73 1627.925 18490.46 1628.465 ;
      RECT 18488.73 1631.045 18490.46 1631.585 ;
      RECT 18488.73 1633.605 18490.46 1637.705 ;
      RECT 18488.73 1644.935 18490.46 1645.475 ;
      RECT 18488.73 1658.475 18490.46 1659.015 ;
      RECT 18488.73 1666.245 18490.46 1670.345 ;
      RECT 18488.73 1672.365 18490.46 1672.905 ;
      RECT 18488.73 1675.485 18490.46 1676.025 ;
      RECT 18488.73 1682.095 18490.46 1682.635 ;
      RECT 18488.73 1693.315 18490.46 1693.855 ;
      RECT 18488.73 1699.925 18490.46 1700.465 ;
      RECT 18488.73 1703.045 18490.46 1703.585 ;
      RECT 18488.73 1705.605 18490.46 1709.705 ;
      RECT 18488.73 1716.935 18490.46 1717.475 ;
      RECT 18488.73 1730.475 18490.46 1731.015 ;
      RECT 18488.73 1738.245 18490.46 1742.345 ;
      RECT 18488.73 1744.365 18490.46 1744.905 ;
      RECT 18488.73 1747.485 18490.46 1748.025 ;
      RECT 18488.73 1754.095 18490.46 1754.635 ;
      RECT 18488.73 1765.315 18490.46 1765.855 ;
      RECT 18488.73 1771.925 18490.46 1772.465 ;
      RECT 18488.73 1775.045 18490.46 1775.585 ;
      RECT 18488.73 1777.605 18490.46 1781.705 ;
      RECT 18488.73 1788.935 18490.46 1789.475 ;
      RECT 18488.73 1802.475 18490.46 1803.015 ;
      RECT 18488.73 1810.245 18490.46 1814.345 ;
      RECT 18488.73 1816.365 18490.46 1816.905 ;
      RECT 18488.73 1819.485 18490.46 1820.025 ;
      RECT 18488.73 1826.095 18490.46 1826.635 ;
      RECT 18488.73 1837.315 18490.46 1837.855 ;
      RECT 18488.73 1843.925 18490.46 1844.465 ;
      RECT 18488.73 1847.045 18490.46 1847.585 ;
      RECT 18488.73 1849.605 18490.46 1853.705 ;
      RECT 18488.73 1860.935 18490.46 1861.475 ;
      RECT 18488.73 1874.475 18490.46 1875.015 ;
      RECT 18488.73 1882.245 18490.46 1886.345 ;
      RECT 18488.73 1888.365 18490.46 1888.905 ;
      RECT 18488.73 1891.485 18490.46 1892.025 ;
      RECT 18488.73 1898.095 18490.46 1898.635 ;
      RECT 18488.73 1909.315 18490.46 1909.855 ;
      RECT 18488.73 1915.925 18490.46 1916.465 ;
      RECT 18488.73 1919.045 18490.46 1919.585 ;
      RECT 18488.73 1921.605 18490.46 1925.705 ;
      RECT 18488.73 1932.935 18490.46 1933.475 ;
      RECT 18488.73 1946.475 18490.46 1947.015 ;
      RECT 18488.73 1954.245 18490.46 1958.345 ;
      RECT 18488.73 1960.365 18490.46 1960.905 ;
      RECT 18488.73 1963.485 18490.46 1964.025 ;
      RECT 18488.73 1970.095 18490.46 1970.635 ;
      RECT 18488.73 1981.315 18490.46 1981.855 ;
      RECT 18488.73 1987.925 18490.46 1988.465 ;
      RECT 18488.73 1991.045 18490.46 1991.585 ;
      RECT 18488.73 1993.605 18490.46 1997.705 ;
      RECT 18488.73 2004.935 18490.46 2005.475 ;
      RECT 18488.73 2018.475 18490.46 2019.015 ;
      RECT 18488.73 2026.245 18490.46 2030.345 ;
      RECT 18488.73 2032.365 18490.46 2032.905 ;
      RECT 18488.73 2035.485 18490.46 2036.025 ;
      RECT 18488.73 2042.095 18490.46 2042.635 ;
      RECT 18488.73 2053.315 18490.46 2053.855 ;
      RECT 18488.73 2059.925 18490.46 2060.465 ;
      RECT 18488.73 2063.045 18490.46 2063.585 ;
      RECT 18488.73 2065.605 18490.46 2069.705 ;
      RECT 18488.73 2076.935 18490.46 2077.475 ;
      RECT 18488.73 2090.475 18490.46 2091.015 ;
      RECT 18488.73 2098.245 18490.46 2102.345 ;
      RECT 18488.73 2104.365 18490.46 2104.905 ;
      RECT 18488.73 2107.485 18490.46 2108.025 ;
      RECT 18488.73 2114.095 18490.46 2114.635 ;
      RECT 18488.73 2125.315 18490.46 2125.855 ;
      RECT 18488.73 2131.925 18490.46 2132.465 ;
      RECT 18488.73 2135.045 18490.46 2135.585 ;
      RECT 18488.73 2137.605 18490.46 2141.705 ;
      RECT 18488.73 2148.935 18490.46 2149.475 ;
      RECT 18488.73 2162.475 18490.46 2163.015 ;
      RECT 18488.73 2170.245 18490.46 2174.345 ;
      RECT 18488.73 2176.365 18490.46 2176.905 ;
      RECT 18488.73 2179.485 18490.46 2180.025 ;
      RECT 18488.73 2186.095 18490.46 2186.635 ;
      RECT 18488.73 2197.315 18490.46 2197.855 ;
      RECT 18488.73 2203.925 18490.46 2204.465 ;
      RECT 18488.73 2207.045 18490.46 2207.585 ;
      RECT 18488.73 2209.605 18490.46 2213.705 ;
      RECT 18488.73 2220.935 18490.46 2221.475 ;
      RECT 18488.73 2234.475 18490.46 2235.015 ;
      RECT 18488.73 2242.245 18490.46 2246.345 ;
      RECT 18488.73 2248.365 18490.46 2248.905 ;
      RECT 18488.73 2251.485 18490.46 2252.025 ;
      RECT 18488.73 2258.095 18490.46 2258.635 ;
      RECT 18488.73 2269.315 18490.46 2269.855 ;
      RECT 18488.73 2275.925 18490.46 2276.465 ;
      RECT 18488.73 2279.045 18490.46 2279.585 ;
      RECT 18488.73 2281.605 18490.46 2285.705 ;
      RECT 18488.73 2292.935 18490.46 2293.475 ;
      RECT 18488.73 2306.475 18490.46 2307.015 ;
      RECT 18488.73 2314.245 18490.46 2318.345 ;
      RECT 18488.73 2320.365 18490.46 2320.905 ;
      RECT 18488.73 2323.485 18490.46 2324.025 ;
      RECT 18488.73 2330.095 18490.46 2330.635 ;
      RECT 18488.73 2341.315 18490.46 2341.855 ;
      RECT 18488.73 2347.925 18490.46 2348.465 ;
      RECT 18488.73 2351.045 18490.46 2351.585 ;
      RECT 18488.73 2353.605 18490.46 2357.705 ;
      RECT 18488.73 2364.935 18490.46 2365.475 ;
      RECT 18488.73 2378.475 18490.46 2379.015 ;
      RECT 18488.73 2386.245 18490.46 2390.345 ;
      RECT 18488.73 2392.365 18490.46 2392.905 ;
      RECT 18488.73 2395.485 18490.46 2396.025 ;
      RECT 18488.73 2402.095 18490.46 2402.635 ;
      RECT 18488.73 2413.315 18490.46 2413.855 ;
      RECT 18488.73 2419.925 18490.46 2420.465 ;
      RECT 18488.73 2423.045 18490.46 2423.585 ;
      RECT 18488.73 2425.605 18490.46 2429.705 ;
      RECT 18488.73 2436.935 18490.46 2437.475 ;
      RECT 18488.73 2450.475 18490.46 2451.015 ;
      RECT 18488.73 2458.245 18490.46 2462.345 ;
      RECT 18488.73 2464.365 18490.46 2464.905 ;
      RECT 18488.73 2467.485 18490.46 2468.025 ;
      RECT 18488.73 2474.095 18490.46 2474.635 ;
      RECT 18488.73 2485.315 18490.46 2485.855 ;
      RECT 18488.73 2491.925 18490.46 2492.465 ;
      RECT 18488.73 2495.045 18490.46 2495.585 ;
      RECT 18488.73 2497.605 18490.46 2501.705 ;
      RECT 18488.73 2508.935 18490.46 2509.475 ;
      RECT 18488.73 2522.475 18490.46 2523.015 ;
      RECT 18488.73 2530.245 18490.46 2534.345 ;
      RECT 18488.73 2536.365 18490.46 2536.905 ;
      RECT 18488.73 2539.485 18490.46 2540.025 ;
      RECT 18488.73 2546.095 18490.46 2546.635 ;
      RECT 18488.73 2557.315 18490.46 2557.855 ;
      RECT 18488.73 2563.925 18490.46 2564.465 ;
      RECT 18488.73 2567.045 18490.46 2567.585 ;
      RECT 18488.73 2569.605 18490.46 2573.705 ;
      RECT 18488.73 2580.935 18490.46 2581.475 ;
      RECT 18488.73 2594.475 18490.46 2595.015 ;
      RECT 18488.73 2602.245 18490.46 2606.345 ;
      RECT 18488.73 2608.365 18490.46 2608.905 ;
      RECT 18488.73 2611.485 18490.46 2612.025 ;
      RECT 18488.73 2618.095 18490.46 2618.635 ;
      RECT 18488.73 2629.315 18490.46 2629.855 ;
      RECT 18488.73 2635.925 18490.46 2636.465 ;
      RECT 18488.73 2639.045 18490.46 2639.585 ;
      RECT 18488.73 2641.605 18490.46 2645.705 ;
      RECT 18488.73 2652.935 18490.46 2653.475 ;
      RECT 18488.73 2666.475 18490.46 2667.015 ;
      RECT 18488.73 2674.245 18490.46 2678.345 ;
      RECT 18488.73 2680.365 18490.46 2680.905 ;
      RECT 18488.73 2683.485 18490.46 2684.025 ;
      RECT 18488.73 2690.095 18490.46 2690.635 ;
      RECT 18488.73 2701.315 18490.46 2701.855 ;
      RECT 18488.73 2707.925 18490.46 2708.465 ;
      RECT 18488.73 2711.045 18490.46 2711.585 ;
      RECT 18488.73 2713.605 18490.46 2717.705 ;
      RECT 18488.73 2724.935 18490.46 2725.475 ;
      RECT 18488.73 2738.475 18490.46 2739.015 ;
      RECT 18488.73 2746.245 18490.46 2750.345 ;
      RECT 18488.73 2752.365 18490.46 2752.905 ;
      RECT 18488.73 2755.485 18490.46 2756.025 ;
      RECT 18488.73 2762.095 18490.46 2762.635 ;
      RECT 18488.73 2773.315 18490.46 2773.855 ;
      RECT 18488.73 2779.925 18490.46 2780.465 ;
      RECT 18488.73 2783.045 18490.46 2783.585 ;
      RECT 18488.73 2785.605 18490.46 2789.705 ;
      RECT 18488.73 2796.935 18490.46 2797.475 ;
      RECT 18488.73 2810.475 18490.46 2811.015 ;
      RECT 18488.73 2818.245 18490.46 2822.345 ;
      RECT 18488.73 2824.365 18490.46 2824.905 ;
      RECT 18488.73 2827.485 18490.46 2828.025 ;
      RECT 18488.73 2834.095 18490.46 2834.635 ;
      RECT 18488.73 2845.315 18490.46 2845.855 ;
      RECT 18488.73 2851.925 18490.46 2852.465 ;
      RECT 18488.73 2855.045 18490.46 2855.585 ;
      RECT 18488.73 2857.605 18490.46 2861.705 ;
      RECT 18488.73 2868.935 18490.46 2869.475 ;
      RECT 18488.73 2882.475 18490.46 2883.015 ;
      RECT 18488.73 2890.245 18490.46 2894.345 ;
      RECT 18488.73 2896.365 18490.46 2896.905 ;
      RECT 18488.73 2899.485 18490.46 2900.025 ;
      RECT 18488.73 2906.095 18490.46 2906.635 ;
      RECT 18488.73 2917.315 18490.46 2917.855 ;
      RECT 18488.73 2923.925 18490.46 2924.465 ;
      RECT 18488.73 2927.045 18490.46 2927.585 ;
      RECT 18488.73 2929.605 18490.46 2933.705 ;
      RECT 18488.73 2940.935 18490.46 2941.475 ;
      RECT 18488.73 2954.475 18490.46 2955.015 ;
      RECT 18488.73 2962.245 18490.46 2966.345 ;
      RECT 18488.73 2968.365 18490.46 2968.905 ;
      RECT 18488.73 2971.485 18490.46 2972.025 ;
      RECT 18488.73 2978.095 18490.46 2978.635 ;
      RECT 18488.73 2989.315 18490.46 2989.855 ;
      RECT 18488.73 2995.925 18490.46 2996.465 ;
      RECT 18488.73 2999.045 18490.46 2999.585 ;
      RECT 18488.73 3001.605 18490.46 3005.705 ;
      RECT 18488.73 3012.935 18490.46 3013.475 ;
      RECT 18488.73 3026.475 18490.46 3027.015 ;
      RECT 18488.73 3034.245 18490.46 3038.345 ;
      RECT 18488.73 3040.365 18490.46 3040.905 ;
      RECT 18488.73 3043.485 18490.46 3044.025 ;
      RECT 18488.73 3050.095 18490.46 3050.635 ;
      RECT 18488.73 3061.315 18490.46 3061.855 ;
      RECT 18488.73 3067.925 18490.46 3068.465 ;
      RECT 18488.73 3071.045 18490.46 3071.585 ;
      RECT 18488.73 3073.605 18490.46 3077.705 ;
      RECT 18488.73 3084.935 18490.46 3085.475 ;
      RECT 18488.73 3098.475 18490.46 3099.015 ;
      RECT 18488.73 3106.245 18490.46 3110.345 ;
      RECT 18488.73 3112.365 18490.46 3112.905 ;
      RECT 18488.73 3115.485 18490.46 3116.025 ;
      RECT 18488.73 3122.095 18490.46 3122.635 ;
      RECT 18488.73 3133.315 18490.46 3133.855 ;
      RECT 18488.73 3139.925 18490.46 3140.465 ;
      RECT 18488.73 3143.045 18490.46 3143.585 ;
      RECT 18488.73 3145.605 18490.46 3149.705 ;
      RECT 18488.73 3156.935 18490.46 3157.475 ;
      RECT 18488.73 3170.475 18490.46 3171.015 ;
      RECT 18488.73 3178.245 18490.46 3182.345 ;
      RECT 18488.73 3184.365 18490.46 3184.905 ;
      RECT 18488.73 3187.485 18490.46 3188.025 ;
      RECT 18488.73 3194.095 18490.46 3194.635 ;
      RECT 18488.73 3205.315 18490.46 3205.855 ;
      RECT 18488.73 3211.925 18490.46 3212.465 ;
      RECT 18488.73 3215.045 18490.46 3215.585 ;
      RECT 18488.73 3217.605 18490.46 3221.705 ;
      RECT 18488.73 3228.935 18490.46 3229.475 ;
      RECT 18488.73 3242.475 18490.46 3243.015 ;
      RECT 18488.73 3250.245 18490.46 3254.345 ;
      RECT 18488.73 3256.365 18490.46 3256.905 ;
      RECT 18488.73 3259.485 18490.46 3260.025 ;
      RECT 18488.73 3266.095 18490.46 3266.635 ;
      RECT 18488.73 3277.315 18490.46 3277.855 ;
      RECT 18488.73 3283.925 18490.46 3284.465 ;
      RECT 18488.73 3287.045 18490.46 3287.585 ;
      RECT 18488.73 3289.605 18490.46 3293.705 ;
      RECT 18488.73 3300.935 18490.46 3301.475 ;
      RECT 18488.73 3314.475 18490.46 3315.015 ;
      RECT 18488.73 3322.245 18490.46 3326.345 ;
      RECT 18488.73 3328.365 18490.46 3328.905 ;
      RECT 18488.73 3331.485 18490.46 3332.025 ;
      RECT 18488.73 3338.095 18490.46 3338.635 ;
      RECT 18488.73 3349.315 18490.46 3349.855 ;
      RECT 18488.73 3355.925 18490.46 3356.465 ;
      RECT 18488.73 3359.045 18490.46 3359.585 ;
      RECT 18488.73 3361.605 18490.46 3365.705 ;
      RECT 18488.73 3372.935 18490.46 3373.475 ;
      RECT 18488.73 3386.475 18490.46 3387.015 ;
      RECT 18488.73 3394.245 18490.46 3398.345 ;
      RECT 18488.73 3400.365 18490.46 3400.905 ;
      RECT 18488.73 3403.485 18490.46 3404.025 ;
      RECT 18488.73 3410.095 18490.46 3410.635 ;
      RECT 18488.73 3421.315 18490.46 3421.855 ;
      RECT 18488.73 3427.925 18490.46 3428.465 ;
      RECT 18488.73 3431.045 18490.46 3431.585 ;
      RECT 18488.73 3433.605 18490.46 3437.705 ;
      RECT 18488.73 3444.935 18490.46 3445.475 ;
      RECT 18488.73 3458.475 18490.46 3459.015 ;
      RECT 18488.73 3466.245 18490.46 3470.345 ;
      RECT 18488.73 3472.365 18490.46 3472.905 ;
      RECT 18488.73 3475.485 18490.46 3476.025 ;
      RECT 18488.73 3482.095 18490.46 3482.635 ;
      RECT 18488.73 3493.315 18490.46 3493.855 ;
      RECT 18488.73 3499.925 18490.46 3500.465 ;
      RECT 18488.73 3503.045 18490.46 3503.585 ;
      RECT 18488.73 3505.605 18490.46 3509.705 ;
      RECT 18488.73 3516.935 18490.46 3517.475 ;
      RECT 18488.73 3530.475 18490.46 3531.015 ;
      RECT 18488.73 3538.245 18490.46 3542.345 ;
      RECT 18488.73 3544.365 18490.46 3544.905 ;
      RECT 18488.73 3547.485 18490.46 3548.025 ;
      RECT 18488.73 3554.095 18490.46 3554.635 ;
      RECT 18488.73 3565.315 18490.46 3565.855 ;
      RECT 18488.73 3571.925 18490.46 3572.465 ;
      RECT 18488.73 3575.045 18490.46 3575.585 ;
      RECT 18488.73 3577.605 18490.46 3581.705 ;
      RECT 18488.73 3588.935 18490.46 3589.475 ;
      RECT 18488.73 3602.475 18490.46 3603.015 ;
      RECT 18488.73 3610.245 18490.46 3614.345 ;
      RECT 18488.73 3616.365 18490.46 3616.905 ;
      RECT 18488.73 3619.485 18490.46 3620.025 ;
      RECT 18488.73 3626.095 18490.46 3626.635 ;
      RECT 18488.73 3637.315 18490.46 3637.855 ;
      RECT 18488.73 3643.925 18490.46 3644.465 ;
      RECT 18488.73 3647.045 18490.46 3647.585 ;
      RECT 18488.73 3649.605 18490.46 3653.705 ;
      RECT 18488.73 3660.935 18490.46 3661.475 ;
      RECT 18488.73 3674.475 18490.46 3675.015 ;
      RECT 18488.73 3682.245 18490.46 3686.345 ;
      RECT 18488.73 3688.365 18490.46 3688.905 ;
      RECT 18488.73 3691.485 18490.46 3692.025 ;
      RECT 18488.73 3698.095 18490.46 3698.635 ;
      RECT 18488.73 3709.315 18490.46 3709.855 ;
      RECT 18488.73 3715.925 18490.46 3716.465 ;
      RECT 18488.73 3719.045 18490.46 3719.585 ;
      RECT 18488.73 3721.605 18490.46 3725.705 ;
      RECT 18488.73 3732.935 18490.46 3733.475 ;
      RECT 18488.73 3746.475 18490.46 3747.015 ;
      RECT 18488.73 3754.245 18490.46 3758.345 ;
      RECT 18488.73 3760.365 18490.46 3760.905 ;
      RECT 18488.73 3763.485 18490.46 3764.025 ;
      RECT 18488.73 3770.095 18490.46 3770.635 ;
      RECT 18488.73 3781.315 18490.46 3781.855 ;
      RECT 18488.73 3787.925 18490.46 3788.465 ;
      RECT 18488.73 3791.045 18490.46 3791.585 ;
      RECT 18488.73 3793.605 18490.46 3797.705 ;
      RECT 18488.73 3804.935 18490.46 3805.475 ;
      RECT 18488.73 3818.475 18490.46 3819.015 ;
      RECT 18488.73 3826.245 18490.46 3830.345 ;
      RECT 18488.73 3832.365 18490.46 3832.905 ;
      RECT 18488.73 3835.485 18490.46 3836.025 ;
      RECT 18488.73 3842.095 18490.46 3842.635 ;
      RECT 18488.73 3853.315 18490.46 3853.855 ;
      RECT 18488.73 3859.925 18490.46 3860.465 ;
      RECT 18488.73 3863.045 18490.46 3863.585 ;
      RECT 18488.73 3865.605 18490.46 3869.705 ;
      RECT 18488.73 3876.935 18490.46 3877.475 ;
      RECT 18488.73 3890.475 18490.46 3891.015 ;
      RECT 18488.73 3898.245 18490.46 3902.345 ;
      RECT 18488.73 3904.365 18490.46 3904.905 ;
      RECT 18488.73 3907.485 18490.46 3908.025 ;
      RECT 18488.73 3914.095 18490.46 3914.635 ;
      RECT 18488.73 3925.315 18490.46 3925.855 ;
      RECT 18488.73 3931.925 18490.46 3932.465 ;
      RECT 18488.73 3935.045 18490.46 3935.585 ;
      RECT 18488.73 3937.605 18490.46 3941.705 ;
      RECT 18488.73 3948.935 18490.46 3949.475 ;
      RECT 18488.73 3962.475 18490.46 3963.015 ;
      RECT 18488.73 3970.245 18490.46 3974.345 ;
      RECT 18488.73 3976.365 18490.46 3976.905 ;
      RECT 18488.73 3979.485 18490.46 3980.025 ;
      RECT 18488.73 3986.095 18490.46 3986.635 ;
      RECT 18488.73 3997.315 18490.46 3997.855 ;
      RECT 18488.73 4003.925 18490.46 4004.465 ;
      RECT 18488.73 4007.045 18490.46 4007.585 ;
      RECT 18488.73 4009.605 18490.46 4013.705 ;
      RECT 18488.73 4020.935 18490.46 4021.475 ;
      RECT 18488.73 4034.475 18490.46 4035.015 ;
      RECT 18488.73 4042.245 18490.46 4046.345 ;
      RECT 18488.73 4048.365 18490.46 4048.905 ;
      RECT 18488.73 4051.485 18490.46 4052.025 ;
      RECT 18488.73 4058.095 18490.46 4058.635 ;
      RECT 18488.73 4069.315 18490.46 4069.855 ;
      RECT 18488.73 4075.925 18490.46 4076.465 ;
      RECT 18488.73 4079.045 18490.46 4079.585 ;
      RECT 18488.73 4081.605 18490.46 4085.705 ;
      RECT 18488.73 4092.935 18490.46 4093.475 ;
      RECT 18488.73 4106.475 18490.46 4107.015 ;
      RECT 18488.73 4114.245 18490.46 4118.345 ;
      RECT 18488.73 4120.365 18490.46 4120.905 ;
      RECT 18488.73 4123.485 18490.46 4124.025 ;
      RECT 18488.73 4130.095 18490.46 4130.635 ;
      RECT 18488.73 4141.315 18490.46 4141.855 ;
      RECT 18488.73 4147.925 18490.46 4148.465 ;
      RECT 18488.73 4151.045 18490.46 4151.585 ;
      RECT 18488.73 4153.605 18490.46 4157.705 ;
      RECT 18488.73 4164.935 18490.46 4165.475 ;
      RECT 18488.73 4178.475 18490.46 4179.015 ;
      RECT 18488.73 4186.245 18490.46 4190.345 ;
      RECT 18488.73 4192.365 18490.46 4192.905 ;
      RECT 18488.73 4195.485 18490.46 4196.025 ;
      RECT 18488.73 4202.095 18490.46 4202.635 ;
      RECT 18488.73 4213.315 18490.46 4213.855 ;
      RECT 18488.73 4219.925 18490.46 4220.465 ;
      RECT 18488.73 4223.045 18490.46 4223.585 ;
      RECT 18488.73 4225.605 18490.46 4229.705 ;
      RECT 18488.73 4236.935 18490.46 4237.475 ;
      RECT 18488.73 4250.475 18490.46 4251.015 ;
      RECT 18488.73 4258.245 18490.46 4262.345 ;
      RECT 18488.73 4264.365 18490.46 4264.905 ;
      RECT 18488.73 4267.485 18490.46 4268.025 ;
      RECT 18488.73 4274.095 18490.46 4274.635 ;
      RECT 18488.73 4285.315 18490.46 4285.855 ;
      RECT 18488.73 4291.925 18490.46 4292.465 ;
      RECT 18488.73 4295.045 18490.46 4295.585 ;
      RECT 18488.73 4297.605 18490.46 4301.705 ;
      RECT 18488.73 4308.935 18490.46 4309.475 ;
      RECT 18488.73 4322.475 18490.46 4323.015 ;
      RECT 18488.73 4330.245 18490.46 4334.345 ;
      RECT 18488.73 4336.365 18490.46 4336.905 ;
      RECT 18488.73 4339.485 18490.46 4340.025 ;
      RECT 18488.73 4346.095 18490.46 4346.635 ;
      RECT 18488.73 4357.315 18490.46 4357.855 ;
      RECT 18488.73 4363.925 18490.46 4364.465 ;
      RECT 18488.73 4367.045 18490.46 4367.585 ;
      RECT 18488.73 4369.605 18490.46 4373.705 ;
      RECT 18488.73 4380.935 18490.46 4381.475 ;
      RECT 18488.73 4394.475 18490.46 4395.015 ;
      RECT 18488.73 4402.245 18490.46 4406.345 ;
      RECT 18488.73 4408.365 18490.46 4408.905 ;
      RECT 18488.73 4411.485 18490.46 4412.025 ;
      RECT 18488.73 4418.095 18490.46 4418.635 ;
      RECT 18488.73 4429.315 18490.46 4429.855 ;
      RECT 18488.73 4435.925 18490.46 4436.465 ;
      RECT 18488.73 4439.045 18490.46 4439.585 ;
      RECT 18488.73 4441.605 18490.46 4445.705 ;
      RECT 18488.73 4452.935 18490.46 4453.475 ;
      RECT 18488.73 4466.475 18490.46 4467.015 ;
      RECT 18488.73 4474.245 18490.46 4478.345 ;
      RECT 18488.73 4480.365 18490.46 4480.905 ;
      RECT 18488.73 4483.485 18490.46 4484.025 ;
      RECT 18488.73 4490.095 18490.46 4490.635 ;
      RECT 18488.73 4501.315 18490.46 4501.855 ;
      RECT 18488.73 4507.925 18490.46 4508.465 ;
      RECT 18488.73 4511.045 18490.46 4511.585 ;
      RECT 18488.73 4513.605 18490.46 4517.705 ;
      RECT 18488.73 4524.935 18490.46 4525.475 ;
      RECT 18488.73 4538.475 18490.46 4539.015 ;
      RECT 18488.73 4546.245 18490.46 4550.345 ;
      RECT 18488.73 4552.365 18490.46 4552.905 ;
      RECT 18488.73 4555.485 18490.46 4556.025 ;
      RECT 18488.73 4562.095 18490.46 4562.635 ;
      RECT 18488.73 4573.315 18490.46 4573.855 ;
      RECT 18488.73 4579.925 18490.46 4580.465 ;
      RECT 18488.73 4583.045 18490.46 4583.585 ;
      RECT 18488.73 4585.605 18490.46 4589.705 ;
      RECT 18488.73 4596.935 18490.46 4597.475 ;
      RECT 18488.73 4610.475 18490.46 4611.015 ;
      RECT 18488.73 4618.245 18490.46 4622.345 ;
      RECT 18488.73 4624.365 18490.46 4624.905 ;
      RECT 18488.73 4627.485 18490.46 4628.025 ;
      RECT 18488.73 4634.095 18490.46 4634.635 ;
      RECT 18488.73 4645.315 18490.46 4645.855 ;
      RECT 18488.73 4651.925 18490.46 4652.465 ;
      RECT 18488.73 4655.045 18490.46 4655.585 ;
      RECT 18488.73 4657.605 18490.46 4661.705 ;
      RECT 18488.73 4668.935 18490.46 4669.475 ;
      RECT 18488.73 4682.475 18490.46 4683.015 ;
      RECT 18488.73 4690.245 18490.46 4694.345 ;
      RECT 18488.73 4696.365 18490.46 4696.905 ;
      RECT 18488.73 4699.485 18490.46 4700.025 ;
      RECT 18488.73 4706.095 18490.46 4706.635 ;
      RECT 18488.73 4717.315 18490.46 4717.855 ;
      RECT 18488.73 4723.925 18490.46 4724.465 ;
      RECT 18488.73 4727.045 18490.46 4727.585 ;
      RECT 18488.73 4729.605 18490.46 4733.705 ;
      RECT 18488.73 4740.935 18490.46 4741.475 ;
      RECT 18488.73 4754.475 18490.46 4755.015 ;
      RECT 18488.73 4762.245 18490.46 4766.345 ;
      RECT 18488.73 4768.365 18490.46 4768.905 ;
      RECT 18488.73 4771.485 18490.46 4772.025 ;
      RECT 18488.73 4778.095 18490.46 4778.635 ;
      RECT 18488.73 4789.315 18490.46 4789.855 ;
      RECT 18488.73 4795.925 18490.46 4796.465 ;
      RECT 18488.73 4799.045 18490.46 4799.585 ;
      RECT 18488.73 4801.605 18490.46 4805.705 ;
      RECT 18488.73 4812.935 18490.46 4813.475 ;
      RECT 18488.73 4826.475 18490.46 4827.015 ;
      RECT 18488.73 4834.245 18490.46 4838.345 ;
      RECT 18488.73 4840.365 18490.46 4840.905 ;
      RECT 18488.73 4843.485 18490.46 4844.025 ;
      RECT 18488.73 4850.095 18490.46 4850.635 ;
      RECT 18488.73 4861.315 18490.46 4861.855 ;
      RECT 18488.73 4867.925 18490.46 4868.465 ;
      RECT 18488.73 4871.045 18490.46 4871.585 ;
      RECT 18488.73 4873.605 18490.46 4877.705 ;
      RECT 18488.73 4884.935 18490.46 4885.475 ;
      RECT 18488.73 4898.475 18490.46 4899.015 ;
      RECT 18488.73 4906.245 18490.46 4910.345 ;
      RECT 18488.73 4912.365 18490.46 4912.905 ;
      RECT 18488.73 4915.485 18490.46 4916.025 ;
      RECT 18488.73 4922.095 18490.46 4922.635 ;
      RECT 18488.73 4933.315 18490.46 4933.855 ;
      RECT 18488.73 4939.925 18490.46 4940.465 ;
      RECT 18488.73 4943.045 18490.46 4943.585 ;
      RECT 18488.73 4945.605 18490.46 4949.705 ;
      RECT 18488.73 4956.935 18490.46 4957.475 ;
      RECT 18488.73 4970.475 18490.46 4971.015 ;
      RECT 18488.73 4978.245 18490.46 4982.345 ;
      RECT 18488.73 4984.365 18490.46 4984.905 ;
      RECT 18488.73 4987.485 18490.46 4988.025 ;
      RECT 18488.73 4994.095 18490.46 4994.635 ;
      RECT 18488.73 5005.315 18490.46 5005.855 ;
      RECT 18488.73 5011.925 18490.46 5012.465 ;
      RECT 18488.73 5015.045 18490.46 5015.585 ;
      RECT 18488.73 5017.605 18490.46 5021.705 ;
      RECT 18488.73 5028.935 18490.46 5029.475 ;
      RECT 18488.73 5042.475 18490.46 5043.015 ;
      RECT 18488.73 5050.245 18490.46 5054.345 ;
      RECT 18488.73 5056.365 18490.46 5056.905 ;
      RECT 18488.73 5059.485 18490.46 5060.025 ;
      RECT 18488.73 5066.095 18490.46 5066.635 ;
      RECT 18488.73 5077.315 18490.46 5077.855 ;
      RECT 18488.73 5083.925 18490.46 5084.465 ;
      RECT 18488.73 5087.045 18490.46 5087.585 ;
      RECT 18488.73 5089.605 18490.46 5093.705 ;
      RECT 18488.73 5100.935 18490.46 5101.475 ;
      RECT 18488.73 5114.475 18490.46 5115.015 ;
      RECT 18488.73 5122.245 18490.46 5126.345 ;
      RECT 18488.73 5128.365 18490.46 5128.905 ;
      RECT 18488.73 5131.485 18490.46 5132.025 ;
      RECT 18488.73 5138.095 18490.46 5138.635 ;
      RECT 18488.73 5149.315 18490.46 5149.855 ;
      RECT 18488.73 5155.925 18490.46 5156.465 ;
      RECT 18488.73 5159.045 18490.46 5159.585 ;
      RECT 18488.73 5161.605 18490.46 5165.705 ;
      RECT 18488.73 5172.935 18490.46 5173.475 ;
      RECT 18488.73 5186.475 18490.46 5187.015 ;
      RECT 18488.73 5194.245 18490.46 5198.345 ;
      RECT 18488.73 5200.365 18490.46 5200.905 ;
      RECT 18488.73 5203.485 18490.46 5204.025 ;
      RECT 18488.73 5210.095 18490.46 5210.635 ;
      RECT 18488.73 5221.315 18490.46 5221.855 ;
      RECT 18488.73 5227.925 18490.46 5228.465 ;
      RECT 18488.73 5231.045 18490.46 5231.585 ;
      RECT 18488.73 5233.605 18490.46 5237.705 ;
      RECT 18488.73 5244.935 18490.46 5245.475 ;
      RECT 18488.73 5258.475 18490.46 5259.015 ;
      RECT 18488.73 5266.245 18490.46 5270.345 ;
      RECT 18488.73 5272.365 18490.46 5272.905 ;
      RECT 18488.73 5275.485 18490.46 5276.025 ;
      RECT 18488.73 5282.095 18490.46 5282.635 ;
      RECT 18488.73 5293.315 18490.46 5293.855 ;
      RECT 18488.73 5299.925 18490.46 5300.465 ;
      RECT 18488.73 5303.045 18490.46 5303.585 ;
      RECT 18488.73 5305.605 18490.46 5309.705 ;
      RECT 18488.73 5316.935 18490.46 5317.475 ;
      RECT 18488.73 5330.475 18490.46 5331.015 ;
      RECT 18488.73 5338.245 18490.46 5342.345 ;
      RECT 18488.73 5344.365 18490.46 5344.905 ;
      RECT 18488.73 5347.485 18490.46 5348.025 ;
      RECT 18488.73 5354.095 18490.46 5354.635 ;
      RECT 18488.73 5365.315 18490.46 5365.855 ;
      RECT 18488.73 5371.925 18490.46 5372.465 ;
      RECT 18488.73 5375.045 18490.46 5375.585 ;
      RECT 18488.73 5377.605 18490.46 5381.705 ;
      RECT 18488.73 5388.935 18490.46 5389.475 ;
      RECT 18488.73 5402.475 18490.46 5403.015 ;
      RECT 18488.73 5410.245 18490.46 5414.345 ;
      RECT 18488.73 5416.365 18490.46 5416.905 ;
      RECT 18488.73 5419.485 18490.46 5420.025 ;
      RECT 18488.73 5426.095 18490.46 5426.635 ;
      RECT 18488.73 5437.315 18490.46 5437.855 ;
      RECT 18488.73 5443.925 18490.46 5444.465 ;
      RECT 18488.73 5447.045 18490.46 5447.585 ;
      RECT 18488.73 5449.605 18490.46 5453.705 ;
      RECT 18488.73 5460.935 18490.46 5461.475 ;
      RECT 18488.73 5474.475 18490.46 5475.015 ;
      RECT 18488.73 5482.245 18490.46 5486.345 ;
      RECT 18488.73 5488.365 18490.46 5488.905 ;
      RECT 18488.73 5491.485 18490.46 5492.025 ;
      RECT 18488.73 5498.095 18490.46 5498.635 ;
      RECT 18488.73 5509.315 18490.46 5509.855 ;
      RECT 18488.73 5515.925 18490.46 5516.465 ;
      RECT 18488.73 5519.045 18490.46 5519.585 ;
      RECT 18488.73 5521.605 18490.46 5525.705 ;
      RECT 18488.73 5532.935 18490.46 5533.475 ;
      RECT 18488.73 5546.475 18490.46 5547.015 ;
      RECT 18488.73 5554.245 18490.46 5558.345 ;
      RECT 18488.73 5560.365 18490.46 5560.905 ;
      RECT 18488.73 5563.485 18490.46 5564.025 ;
      RECT 18488.73 5570.095 18490.46 5570.635 ;
      RECT 18488.73 5581.315 18490.46 5581.855 ;
      RECT 18488.73 5587.925 18490.46 5588.465 ;
      RECT 18488.73 5591.045 18490.46 5591.585 ;
      RECT 18488.73 5593.605 18490.46 5597.705 ;
      RECT 18488.73 5604.935 18490.46 5605.475 ;
      RECT 18488.73 5618.475 18490.46 5619.015 ;
      RECT 18488.73 5626.245 18490.46 5630.345 ;
      RECT 18488.73 5632.365 18490.46 5632.905 ;
      RECT 18488.73 5635.485 18490.46 5636.025 ;
      RECT 18488.73 5642.095 18490.46 5642.635 ;
      RECT 18488.73 5653.315 18490.46 5653.855 ;
      RECT 18488.73 5659.925 18490.46 5660.465 ;
      RECT 18488.73 5663.045 18490.46 5663.585 ;
      RECT 18488.73 5665.605 18490.46 5669.705 ;
      RECT 18488.73 5676.935 18490.46 5677.475 ;
      RECT 18488.73 5690.475 18490.46 5691.015 ;
      RECT 18488.73 5698.245 18490.46 5702.345 ;
      RECT 18488.73 5704.365 18490.46 5704.905 ;
      RECT 18488.73 5707.485 18490.46 5708.025 ;
      RECT 18488.73 5714.095 18490.46 5714.635 ;
      RECT 18488.73 5725.315 18490.46 5725.855 ;
      RECT 18488.73 5731.925 18490.46 5732.465 ;
      RECT 18488.73 5735.045 18490.46 5735.585 ;
      RECT 18488.73 5737.605 18490.46 5741.705 ;
      RECT 18488.73 5748.935 18490.46 5749.475 ;
      RECT 18488.73 5762.475 18490.46 5763.015 ;
      RECT 18488.73 5770.245 18490.46 5774.345 ;
      RECT 18488.73 5776.365 18490.46 5776.905 ;
      RECT 18488.73 5779.485 18490.46 5780.025 ;
      RECT 18488.73 5786.095 18490.46 5786.635 ;
      RECT 18488.73 5797.315 18490.46 5797.855 ;
      RECT 18488.73 5803.925 18490.46 5804.465 ;
      RECT 18488.73 5807.045 18490.46 5807.585 ;
      RECT 18488.73 5809.605 18490.46 5813.705 ;
      RECT 18488.73 5820.935 18490.46 5821.475 ;
      RECT 18488.73 5834.475 18490.46 5835.015 ;
      RECT 18488.73 5842.245 18490.46 5846.345 ;
      RECT 18488.73 5848.365 18490.46 5848.905 ;
      RECT 18488.73 5851.485 18490.46 5852.025 ;
      RECT 18488.73 5858.095 18490.46 5858.635 ;
      RECT 18488.73 5869.315 18490.46 5869.855 ;
      RECT 18488.73 5875.925 18490.46 5876.465 ;
      RECT 18488.73 5879.045 18490.46 5879.585 ;
      RECT 18488.73 5881.605 18490.46 5885.705 ;
      RECT 18488.73 5892.935 18490.46 5893.475 ;
      RECT 18488.73 5906.475 18490.46 5907.015 ;
      RECT 18488.73 5914.245 18490.46 5918.345 ;
      RECT 18488.73 5920.365 18490.46 5920.905 ;
      RECT 18488.73 5923.485 18490.46 5924.025 ;
      RECT 18488.73 5930.095 18490.46 5930.635 ;
      RECT 18488.73 5941.315 18490.46 5941.855 ;
      RECT 18488.73 5947.925 18490.46 5948.465 ;
      RECT 18488.73 5951.045 18490.46 5951.585 ;
      RECT 18488.73 5953.605 18490.46 5957.705 ;
      RECT 18488.73 5964.935 18490.46 5965.475 ;
      RECT 18488.73 5978.475 18490.46 5979.015 ;
      RECT 18488.73 5986.245 18490.46 5990.345 ;
      RECT 18488.73 5992.365 18490.46 5992.905 ;
      RECT 18488.73 5995.485 18490.46 5996.025 ;
      RECT 18488.73 6002.095 18490.46 6002.635 ;
      RECT 18488.73 6013.315 18490.46 6013.855 ;
      RECT 18488.73 6019.925 18490.46 6020.465 ;
      RECT 18488.73 6023.045 18490.46 6023.585 ;
      RECT 18488.73 6025.605 18490.46 6029.705 ;
      RECT 18488.73 6036.935 18490.46 6037.475 ;
      RECT 18488.73 6050.475 18490.46 6051.015 ;
      RECT 18488.73 6058.245 18490.46 6062.345 ;
      RECT 18488.73 6064.365 18490.46 6064.905 ;
      RECT 18488.73 6067.485 18490.46 6068.025 ;
      RECT 18488.73 6074.095 18490.46 6074.635 ;
      RECT 18488.73 6085.315 18490.46 6085.855 ;
      RECT 18488.73 6091.925 18490.46 6092.465 ;
      RECT 18488.73 6095.045 18490.46 6095.585 ;
      RECT 18488.73 6097.605 18490.46 6101.705 ;
      RECT 18488.73 6108.935 18490.46 6109.475 ;
      RECT 18488.73 6122.475 18490.46 6123.015 ;
      RECT 18488.73 6130.245 18490.46 6134.345 ;
      RECT 18488.73 6136.365 18490.46 6136.905 ;
      RECT 18488.73 6139.485 18490.46 6140.025 ;
      RECT 18488.73 6146.095 18490.46 6146.635 ;
      RECT 18488.73 6157.315 18490.46 6157.855 ;
      RECT 18488.73 6163.925 18490.46 6164.465 ;
      RECT 18488.73 6167.045 18490.46 6167.585 ;
      RECT 18488.73 6169.605 18490.46 6173.705 ;
      RECT 18488.73 6180.935 18490.46 6181.475 ;
      RECT 18488.73 6194.475 18490.46 6195.015 ;
      RECT 18488.73 6202.245 18490.46 6206.345 ;
      RECT 18488.73 6208.365 18490.46 6208.905 ;
      RECT 18488.73 6211.485 18490.46 6212.025 ;
      RECT 18488.73 6218.095 18490.46 6218.635 ;
      RECT 18488.73 6229.315 18490.46 6229.855 ;
      RECT 18488.73 6235.925 18490.46 6236.465 ;
      RECT 18488.73 6239.045 18490.46 6239.585 ;
      RECT 18488.73 6241.605 18490.46 6245.705 ;
      RECT 18488.73 6252.935 18490.46 6253.475 ;
      RECT 18488.73 6266.475 18490.46 6267.015 ;
      RECT 18488.73 6274.245 18490.46 6278.345 ;
      RECT 18488.73 6280.365 18490.46 6280.905 ;
      RECT 18488.73 6283.485 18490.46 6284.025 ;
      RECT 18488.73 6290.095 18490.46 6290.635 ;
      RECT 18488.73 6301.315 18490.46 6301.855 ;
      RECT 18488.73 6307.925 18490.46 6308.465 ;
      RECT 18488.73 6311.045 18490.46 6311.585 ;
      RECT 18488.73 6313.605 18490.46 6317.705 ;
      RECT 18488.73 6324.935 18490.46 6325.475 ;
      RECT 18488.73 6338.475 18490.46 6339.015 ;
      RECT 18488.73 6346.245 18490.46 6350.345 ;
      RECT 18488.73 6352.365 18490.46 6352.905 ;
      RECT 18488.73 6355.485 18490.46 6356.025 ;
      RECT 18488.73 6362.095 18490.46 6362.635 ;
      RECT 18488.73 6373.315 18490.46 6373.855 ;
      RECT 18488.73 6379.925 18490.46 6380.465 ;
      RECT 18488.73 6383.045 18490.46 6383.585 ;
      RECT 18488.73 6385.605 18490.46 6389.705 ;
      RECT 18488.73 6396.935 18490.46 6397.475 ;
      RECT 18488.73 6410.475 18490.46 6411.015 ;
      RECT 18488.73 6418.245 18490.46 6422.345 ;
      RECT 18488.73 6424.365 18490.46 6424.905 ;
      RECT 18488.73 6427.485 18490.46 6428.025 ;
      RECT 18488.73 6434.095 18490.46 6434.635 ;
      RECT 18488.73 6445.315 18490.46 6445.855 ;
      RECT 18488.73 6451.925 18490.46 6452.465 ;
      RECT 18488.73 6455.045 18490.46 6455.585 ;
      RECT 18488.73 6457.605 18490.46 6461.705 ;
      RECT 18488.73 6468.935 18490.46 6469.475 ;
      RECT 18488.73 6482.475 18490.46 6483.015 ;
      RECT 18488.73 6490.245 18490.46 6494.345 ;
      RECT 18488.73 6496.365 18490.46 6496.905 ;
      RECT 18488.73 6499.485 18490.46 6500.025 ;
      RECT 18488.73 6506.095 18490.46 6506.635 ;
      RECT 18488.73 6517.315 18490.46 6517.855 ;
      RECT 18488.73 6523.925 18490.46 6524.465 ;
      RECT 18488.73 6527.045 18490.46 6527.585 ;
      RECT 18488.73 6529.605 18490.46 6533.705 ;
      RECT 18488.73 6540.935 18490.46 6541.475 ;
      RECT 18488.73 6554.475 18490.46 6555.015 ;
      RECT 18488.73 6562.245 18490.46 6566.345 ;
      RECT 18488.73 6568.365 18490.46 6568.905 ;
      RECT 18488.73 6571.485 18490.46 6572.025 ;
      RECT 18488.73 6578.095 18490.46 6578.635 ;
      RECT 18488.73 6589.315 18490.46 6589.855 ;
      RECT 18488.73 6595.925 18490.46 6596.465 ;
      RECT 18488.73 6599.045 18490.46 6599.585 ;
      RECT 18488.73 6601.605 18490.46 6605.705 ;
      RECT 18488.73 6612.935 18490.46 6613.475 ;
      RECT 18488.73 6626.475 18490.46 6627.015 ;
      RECT 18488.73 6634.245 18490.46 6638.345 ;
      RECT 18488.73 6640.365 18490.46 6640.905 ;
      RECT 18488.73 6643.485 18490.46 6644.025 ;
      RECT 18488.73 6650.095 18490.46 6650.635 ;
      RECT 18488.73 6661.315 18490.46 6661.855 ;
      RECT 18488.73 6667.925 18490.46 6668.465 ;
      RECT 18488.73 6671.045 18490.46 6671.585 ;
      RECT 18488.73 6673.605 18490.46 6677.705 ;
      RECT 18488.73 6684.935 18490.46 6685.475 ;
      RECT 18488.73 6698.475 18490.46 6699.015 ;
      RECT 18488.73 6706.245 18490.46 6710.345 ;
      RECT 18488.73 6712.365 18490.46 6712.905 ;
      RECT 18488.73 6715.485 18490.46 6716.025 ;
      RECT 18488.73 6722.095 18490.46 6722.635 ;
      RECT 18488.73 6733.315 18490.46 6733.855 ;
      RECT 18488.73 6739.925 18490.46 6740.465 ;
      RECT 18488.73 6743.045 18490.46 6743.585 ;
      RECT 18488.73 6745.605 18490.46 6749.705 ;
      RECT 18488.73 6756.935 18490.46 6757.475 ;
      RECT 18488.73 6770.475 18490.46 6771.015 ;
      RECT 18488.73 6778.245 18490.46 6782.345 ;
      RECT 18488.73 6784.365 18490.46 6784.905 ;
      RECT 18488.73 6787.485 18490.46 6788.025 ;
      RECT 18488.73 6794.095 18490.46 6794.635 ;
      RECT 18488.73 6805.315 18490.46 6805.855 ;
      RECT 18488.73 6811.925 18490.46 6812.465 ;
      RECT 18488.73 6815.045 18490.46 6815.585 ;
      RECT 18488.73 6817.605 18490.46 6821.705 ;
      RECT 18488.73 6828.935 18490.46 6829.475 ;
      RECT 18488.73 6842.475 18490.46 6843.015 ;
      RECT 18488.73 6850.245 18490.46 6854.345 ;
      RECT 18488.73 6856.365 18490.46 6856.905 ;
      RECT 18488.73 6859.485 18490.46 6860.025 ;
      RECT 18488.73 6866.095 18490.46 6866.635 ;
      RECT 18488.73 6877.315 18490.46 6877.855 ;
      RECT 18488.73 6883.925 18490.46 6884.465 ;
      RECT 18488.73 6887.045 18490.46 6887.585 ;
      RECT 18488.73 6889.605 18490.46 6893.705 ;
      RECT 18488.73 6900.935 18490.46 6901.475 ;
      RECT 18488.73 6914.475 18490.46 6915.015 ;
      RECT 18488.73 6922.245 18490.46 6926.345 ;
      RECT 18488.73 6928.365 18490.46 6928.905 ;
      RECT 18488.73 6931.485 18490.46 6932.025 ;
      RECT 18488.73 6938.095 18490.46 6938.635 ;
      RECT 18488.73 6949.315 18490.46 6949.855 ;
      RECT 18488.73 6955.925 18490.46 6956.465 ;
      RECT 18488.73 6959.045 18490.46 6959.585 ;
      RECT 18488.73 6961.605 18490.46 6965.705 ;
      RECT 18488.73 6972.935 18490.46 6973.475 ;
      RECT 18488.73 6986.475 18490.46 6987.015 ;
      RECT 18488.73 6994.245 18490.46 6998.345 ;
      RECT 18488.73 7000.365 18490.46 7000.905 ;
      RECT 18488.73 7003.485 18490.46 7004.025 ;
      RECT 18488.73 7010.095 18490.46 7010.635 ;
      RECT 18488.73 7021.315 18490.46 7021.855 ;
      RECT 18488.73 7027.925 18490.46 7028.465 ;
      RECT 18488.73 7031.045 18490.46 7031.585 ;
      RECT 18488.73 7033.605 18490.46 7037.705 ;
      RECT 18488.73 7044.935 18490.46 7045.475 ;
      RECT 18488.73 7058.475 18490.46 7059.015 ;
      RECT 18488.73 7066.245 18490.46 7070.345 ;
      RECT 18488.73 7072.365 18490.46 7072.905 ;
      RECT 18488.73 7075.485 18490.46 7076.025 ;
      RECT 18488.73 7082.095 18490.46 7082.635 ;
      RECT 18488.73 7093.315 18490.46 7093.855 ;
      RECT 18488.73 7099.925 18490.46 7100.465 ;
      RECT 18488.73 7103.045 18490.46 7103.585 ;
      RECT 18488.73 7105.605 18490.46 7109.705 ;
      RECT 18488.73 7116.935 18490.46 7117.475 ;
      RECT 18488.73 7130.475 18490.46 7131.015 ;
      RECT 18488.73 7138.245 18490.46 7142.345 ;
      RECT 18488.73 7144.365 18490.46 7144.905 ;
      RECT 18488.73 7147.485 18490.46 7148.025 ;
      RECT 18488.73 7154.095 18490.46 7154.635 ;
      RECT 18488.73 7165.315 18490.46 7165.855 ;
      RECT 18488.73 7171.925 18490.46 7172.465 ;
      RECT 18488.73 7175.045 18490.46 7175.585 ;
      RECT 18488.73 7177.605 18490.46 7181.705 ;
      RECT 18488.73 7188.935 18490.46 7189.475 ;
      RECT 18488.73 7202.475 18490.46 7203.015 ;
      RECT 18488.73 7210.245 18490.46 7214.345 ;
      RECT 18488.73 7216.365 18490.46 7216.905 ;
      RECT 18488.73 7219.485 18490.46 7220.025 ;
      RECT 18488.73 7226.095 18490.46 7226.635 ;
      RECT 18488.73 7237.315 18490.46 7237.855 ;
      RECT 18488.73 7243.925 18490.46 7244.465 ;
      RECT 18488.73 7247.045 18490.46 7247.585 ;
      RECT 18488.73 7249.605 18490.46 7253.705 ;
      RECT 18488.73 7260.935 18490.46 7261.475 ;
      RECT 18488.73 7274.475 18490.46 7275.015 ;
      RECT 18488.73 7282.245 18490.46 7286.345 ;
      RECT 18488.73 7288.365 18490.46 7288.905 ;
      RECT 18488.73 7291.485 18490.46 7292.025 ;
      RECT 18488.73 7298.095 18490.46 7298.635 ;
      RECT 18488.73 7309.315 18490.46 7309.855 ;
      RECT 18488.73 7315.925 18490.46 7316.465 ;
      RECT 18488.73 7319.045 18490.46 7319.585 ;
      RECT 18488.73 7321.605 18490.46 7325.705 ;
      RECT 18488.73 7332.935 18490.46 7333.475 ;
      RECT 18488.73 7346.475 18490.46 7347.015 ;
      RECT 18488.73 7354.245 18490.46 7358.345 ;
      RECT 18488.73 7360.365 18490.46 7360.905 ;
      RECT 18488.73 7363.485 18490.46 7364.025 ;
      RECT 18488.73 7370.095 18490.46 7370.635 ;
      RECT 18488.73 7381.315 18490.46 7381.855 ;
      RECT 18488.73 7387.925 18490.46 7388.465 ;
      RECT 18488.73 7391.045 18490.46 7391.585 ;
      RECT 18488.73 7393.605 18490.46 7397.705 ;
      RECT 18488.73 7404.935 18490.46 7405.475 ;
      RECT 18488.73 7418.475 18490.46 7419.015 ;
      RECT 18488.73 7426.245 18490.46 7430.345 ;
      RECT 18488.73 7432.365 18490.46 7432.905 ;
      RECT 18488.73 7435.485 18490.46 7436.025 ;
      RECT 18488.73 7442.095 18490.46 7442.635 ;
      RECT 18488.73 7453.315 18490.46 7453.855 ;
      RECT 18488.73 7459.925 18490.46 7460.465 ;
      RECT 18488.73 7463.045 18490.46 7463.585 ;
      RECT 18488.73 7465.605 18490.46 7469.705 ;
      RECT 18488.73 7476.935 18490.46 7477.475 ;
      RECT 18488.73 7490.475 18490.46 7491.015 ;
      RECT 18488.73 7498.245 18490.46 7502.345 ;
      RECT 18488.73 7504.365 18490.46 7504.905 ;
      RECT 18488.73 7507.485 18490.46 7508.025 ;
      RECT 18488.73 7514.095 18490.46 7514.635 ;
      RECT 18488.73 7525.315 18490.46 7525.855 ;
      RECT 18488.73 7531.925 18490.46 7532.465 ;
      RECT 18488.73 7535.045 18490.46 7535.585 ;
      RECT 18488.73 7537.605 18490.46 7541.705 ;
      RECT 18488.73 7548.935 18490.46 7549.475 ;
      RECT 18488.73 7562.475 18490.46 7563.015 ;
      RECT 18488.73 7570.245 18490.46 7574.345 ;
      RECT 18488.73 7576.365 18490.46 7576.905 ;
      RECT 18488.73 7579.485 18490.46 7580.025 ;
      RECT 18488.73 7586.095 18490.46 7586.635 ;
      RECT 18488.73 7597.315 18490.46 7597.855 ;
      RECT 18488.73 7603.925 18490.46 7604.465 ;
      RECT 18488.73 7607.045 18490.46 7607.585 ;
      RECT 18488.73 7609.605 18490.46 7613.705 ;
      RECT 18488.73 7620.935 18490.46 7621.475 ;
      RECT 18488.73 7634.475 18490.46 7635.015 ;
      RECT 18488.73 7642.245 18490.46 7646.345 ;
      RECT 18488.73 7648.365 18490.46 7648.905 ;
      RECT 18488.73 7651.485 18490.46 7652.025 ;
      RECT 18488.73 7658.095 18490.46 7658.635 ;
      RECT 18488.73 7669.315 18490.46 7669.855 ;
      RECT 18488.73 7675.925 18490.46 7676.465 ;
      RECT 18488.73 7679.045 18490.46 7679.585 ;
      RECT 18488.73 7681.605 18490.46 7685.705 ;
      RECT 18488.73 7692.935 18490.46 7693.475 ;
      RECT 18488.73 7706.475 18490.46 7707.015 ;
      RECT 18488.73 7714.245 18490.46 7718.345 ;
      RECT 18488.73 7720.365 18490.46 7720.905 ;
      RECT 18488.73 7723.485 18490.46 7724.025 ;
      RECT 18488.73 7730.095 18490.46 7730.635 ;
      RECT 18488.73 7741.315 18490.46 7741.855 ;
      RECT 18488.73 7747.925 18490.46 7748.465 ;
      RECT 18488.73 7751.045 18490.46 7751.585 ;
      RECT 18488.73 7753.605 18490.46 7757.705 ;
      RECT 18488.73 7764.935 18490.46 7765.475 ;
      RECT 18488.73 7778.475 18490.46 7779.015 ;
      RECT 18488.73 7786.245 18490.46 7790.345 ;
      RECT 18488.73 7792.365 18490.46 7792.905 ;
      RECT 18488.73 7795.485 18490.46 7796.025 ;
      RECT 18488.73 7802.095 18490.46 7802.635 ;
      RECT 18488.73 7813.315 18490.46 7813.855 ;
      RECT 18488.73 7819.925 18490.46 7820.465 ;
      RECT 18488.73 7823.045 18490.46 7823.585 ;
      RECT 18488.73 7825.605 18490.46 7829.705 ;
      RECT 18488.73 7836.935 18490.46 7837.475 ;
      RECT 18488.73 7850.475 18490.46 7851.015 ;
      RECT 18488.73 7858.245 18490.46 7862.345 ;
      RECT 18488.73 7864.365 18490.46 7864.905 ;
      RECT 18488.73 7867.485 18490.46 7868.025 ;
      RECT 18488.73 7874.095 18490.46 7874.635 ;
      RECT 18488.73 7885.315 18490.46 7885.855 ;
      RECT 18488.73 7891.925 18490.46 7892.465 ;
      RECT 18488.73 7895.045 18490.46 7895.585 ;
      RECT 18488.73 7897.605 18490.46 7901.705 ;
      RECT 18488.73 7908.935 18490.46 7909.475 ;
      RECT 18488.73 7922.475 18490.46 7923.015 ;
      RECT 18488.73 7930.245 18490.46 7934.345 ;
      RECT 18488.73 7936.365 18490.46 7936.905 ;
      RECT 18488.73 7939.485 18490.46 7940.025 ;
      RECT 18488.73 7946.095 18490.46 7946.635 ;
      RECT 18488.73 7957.315 18490.46 7957.855 ;
      RECT 18488.73 7963.925 18490.46 7964.465 ;
      RECT 18488.73 7967.045 18490.46 7967.585 ;
      RECT 18488.73 7969.605 18490.46 7973.705 ;
      RECT 18488.73 7980.935 18490.46 7981.475 ;
      RECT 18488.73 7994.475 18490.46 7995.015 ;
      RECT 18488.73 8002.245 18490.46 8006.345 ;
      RECT 18488.73 8008.365 18490.46 8008.905 ;
      RECT 18488.73 8011.485 18490.46 8012.025 ;
      RECT 18488.73 8018.095 18490.46 8018.635 ;
      RECT 18488.73 8029.315 18490.46 8029.855 ;
      RECT 18488.73 8035.925 18490.46 8036.465 ;
      RECT 18488.73 8039.045 18490.46 8039.585 ;
      RECT 18488.73 8041.605 18490.46 8045.705 ;
      RECT 18488.73 8052.935 18490.46 8053.475 ;
      RECT 18488.73 8066.475 18490.46 8067.015 ;
      RECT 18488.73 8074.245 18490.46 8078.345 ;
      RECT 18488.73 8080.365 18490.46 8080.905 ;
      RECT 18488.73 8083.485 18490.46 8084.025 ;
      RECT 18488.73 8090.095 18490.46 8090.635 ;
      RECT 18488.73 8101.315 18490.46 8101.855 ;
      RECT 18488.73 8107.925 18490.46 8108.465 ;
      RECT 18488.73 8111.045 18490.46 8111.585 ;
      RECT 18488.73 8113.605 18490.46 8117.705 ;
      RECT 18488.73 8124.935 18490.46 8125.475 ;
      RECT 18488.73 8138.475 18490.46 8139.015 ;
      RECT 18488.73 8146.245 18490.46 8150.345 ;
      RECT 18488.73 8152.365 18490.46 8152.905 ;
      RECT 18488.73 8155.485 18490.46 8156.025 ;
      RECT 18488.73 8162.095 18490.46 8162.635 ;
      RECT 18488.73 8173.315 18490.46 8173.855 ;
      RECT 18488.73 8179.925 18490.46 8180.465 ;
      RECT 18488.73 8183.045 18490.46 8183.585 ;
      RECT 18488.73 8185.605 18490.46 8189.705 ;
      RECT 18488.73 8196.935 18490.46 8197.475 ;
      RECT 18488.73 8210.475 18490.46 8211.015 ;
      RECT 18488.73 8218.245 18490.46 8222.345 ;
      RECT 18488.73 8224.365 18490.46 8224.905 ;
      RECT 18488.73 8227.485 18490.46 8228.025 ;
      RECT 18488.73 8234.095 18490.46 8234.635 ;
      RECT 18488.73 8245.315 18490.46 8245.855 ;
      RECT 18488.73 8251.925 18490.46 8252.465 ;
      RECT 18488.73 8255.045 18490.46 8255.585 ;
      RECT 18488.73 8257.605 18490.46 8261.705 ;
      RECT 18488.73 8268.935 18490.46 8269.475 ;
      RECT 18488.73 8282.475 18490.46 8283.015 ;
      RECT 18488.73 8290.245 18490.46 8294.345 ;
      RECT 18488.73 8296.365 18490.46 8296.905 ;
      RECT 18488.73 8299.485 18490.46 8300.025 ;
      RECT 18488.73 8306.095 18490.46 8306.635 ;
      RECT 18488.73 8317.315 18490.46 8317.855 ;
      RECT 18488.73 8323.925 18490.46 8324.465 ;
      RECT 18488.73 8327.045 18490.46 8327.585 ;
      RECT 18488.73 8329.605 18490.46 8333.705 ;
      RECT 18488.73 8340.935 18490.46 8341.475 ;
      RECT 18488.73 8354.475 18490.46 8355.015 ;
      RECT 18488.73 8362.245 18490.46 8366.345 ;
      RECT 18488.73 8368.365 18490.46 8368.905 ;
      RECT 18488.73 8371.485 18490.46 8372.025 ;
      RECT 18488.73 8378.095 18490.46 8378.635 ;
      RECT 18488.73 8389.315 18490.46 8389.855 ;
      RECT 18488.73 8395.925 18490.46 8396.465 ;
      RECT 18488.73 8399.045 18490.46 8399.585 ;
      RECT 18488.73 8401.605 18490.46 8405.705 ;
      RECT 18488.73 8412.935 18490.46 8413.475 ;
      RECT 18488.73 8426.475 18490.46 8427.015 ;
      RECT 18488.73 8434.245 18490.46 8438.345 ;
      RECT 18488.73 8440.365 18490.46 8440.905 ;
      RECT 18488.73 8443.485 18490.46 8444.025 ;
      RECT 18488.73 8450.095 18490.46 8450.635 ;
      RECT 18488.73 8461.315 18490.46 8461.855 ;
      RECT 18488.73 8467.925 18490.46 8468.465 ;
      RECT 18488.73 8471.045 18490.46 8471.585 ;
      RECT 18488.73 8473.605 18490.46 8477.705 ;
      RECT 18488.73 8484.935 18490.46 8485.475 ;
      RECT 18488.73 8498.475 18490.46 8499.015 ;
      RECT 18488.73 8506.245 18490.46 8510.345 ;
      RECT 18488.73 8512.365 18490.46 8512.905 ;
      RECT 18488.73 8515.485 18490.46 8516.025 ;
      RECT 18488.73 8522.095 18490.46 8522.635 ;
      RECT 18488.73 8533.315 18490.46 8533.855 ;
      RECT 18488.73 8539.925 18490.46 8540.465 ;
      RECT 18488.73 8543.045 18490.46 8543.585 ;
      RECT 18488.73 8545.605 18490.46 8549.705 ;
      RECT 18488.73 8556.935 18490.46 8557.475 ;
      RECT 18488.73 8570.475 18490.46 8571.015 ;
      RECT 18488.73 8578.245 18490.46 8582.345 ;
      RECT 18488.73 8584.365 18490.46 8584.905 ;
      RECT 18488.73 8587.485 18490.46 8588.025 ;
      RECT 18488.73 8594.095 18490.46 8594.635 ;
      RECT 18488.73 8600.705 18490.46 8610.835 ;
  END
  PROPERTY CatenaDesignType "asic" ;
END matrix_dac

END LIBRARY
