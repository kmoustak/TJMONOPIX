VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO Pulldown_pol_IO_lowcap_EN
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN Pulldown_pol_IO_lowcap_EN 0 0 ;
  SIZE 100 BY 120 ;
  SYMMETRY X Y R90 ;
  PIN PAD
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 4 4 96 96 ;
        RECT 33.245 4 67.155 99.65 ;
    END
  END PAD
  PIN OEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7.75 117 10.75 120 ;
    END
  END OEN
  PIN SUB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
        RECT 0 4 100 8 ;
      LAYER M3 ;
        RECT 0 4 100 8 ;
      LAYER V4 ;
        RECT 0.35 6.59 0.61 6.85 ;
        RECT 0.35 5.83 0.61 6.09 ;
        RECT 0.35 5.07 0.61 5.33 ;
        RECT 1.11 6.59 1.37 6.85 ;
        RECT 1.11 5.83 1.37 6.09 ;
        RECT 1.11 5.07 1.37 5.33 ;
        RECT 1.87 6.59 2.13 6.85 ;
        RECT 1.87 5.83 2.13 6.09 ;
        RECT 1.87 5.07 2.13 5.33 ;
        RECT 2.63 6.59 2.89 6.85 ;
        RECT 2.63 5.83 2.89 6.09 ;
        RECT 2.63 5.07 2.89 5.33 ;
        RECT 3.39 6.59 3.65 6.85 ;
        RECT 3.39 5.83 3.65 6.09 ;
        RECT 3.39 5.07 3.65 5.33 ;
        RECT 96.35 6.59 96.61 6.85 ;
        RECT 96.35 5.83 96.61 6.09 ;
        RECT 96.35 5.07 96.61 5.33 ;
        RECT 97.11 6.59 97.37 6.85 ;
        RECT 97.11 5.83 97.37 6.09 ;
        RECT 97.11 5.07 97.37 5.33 ;
        RECT 97.87 6.59 98.13 6.85 ;
        RECT 97.87 5.83 98.13 6.09 ;
        RECT 97.87 5.07 98.13 5.33 ;
        RECT 98.63 6.59 98.89 6.85 ;
        RECT 98.63 5.83 98.89 6.09 ;
        RECT 98.63 5.07 98.89 5.33 ;
        RECT 99.39 6.59 99.65 6.85 ;
        RECT 99.39 5.83 99.65 6.09 ;
        RECT 99.39 5.07 99.65 5.33 ;
    END
  END SUB
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
        RECT 0 66 100 96 ;
      LAYER M3 ;
        RECT 0 66 100 96 ;
      LAYER V4 ;
        RECT 0.35 91.2 0.61 91.46 ;
        RECT 0.35 90.44 0.61 90.7 ;
        RECT 0.35 89.68 0.61 89.94 ;
        RECT 0.35 88.92 0.61 89.18 ;
        RECT 0.35 88.16 0.61 88.42 ;
        RECT 0.35 87.4 0.61 87.66 ;
        RECT 0.35 86.64 0.61 86.9 ;
        RECT 0.35 85.88 0.61 86.14 ;
        RECT 0.35 85.12 0.61 85.38 ;
        RECT 0.35 84.36 0.61 84.62 ;
        RECT 0.35 83.6 0.61 83.86 ;
        RECT 0.35 82.84 0.61 83.1 ;
        RECT 0.35 82.08 0.61 82.34 ;
        RECT 0.35 81.32 0.61 81.58 ;
        RECT 0.35 80.56 0.61 80.82 ;
        RECT 0.35 79.8 0.61 80.06 ;
        RECT 0.35 79.04 0.61 79.3 ;
        RECT 0.35 78.28 0.61 78.54 ;
        RECT 0.35 77.52 0.61 77.78 ;
        RECT 0.35 76.76 0.61 77.02 ;
        RECT 0.35 76 0.61 76.26 ;
        RECT 0.35 75.24 0.61 75.5 ;
        RECT 0.35 74.48 0.61 74.74 ;
        RECT 0.35 73.72 0.61 73.98 ;
        RECT 0.35 72.96 0.61 73.22 ;
        RECT 0.35 72.2 0.61 72.46 ;
        RECT 0.35 71.44 0.61 71.7 ;
        RECT 0.35 70.68 0.61 70.94 ;
        RECT 0.35 69.92 0.61 70.18 ;
        RECT 0.35 69.16 0.61 69.42 ;
        RECT 1.11 91.2 1.37 91.46 ;
        RECT 1.11 90.44 1.37 90.7 ;
        RECT 1.11 89.68 1.37 89.94 ;
        RECT 1.11 88.92 1.37 89.18 ;
        RECT 1.11 88.16 1.37 88.42 ;
        RECT 1.11 87.4 1.37 87.66 ;
        RECT 1.11 86.64 1.37 86.9 ;
        RECT 1.11 85.88 1.37 86.14 ;
        RECT 1.11 85.12 1.37 85.38 ;
        RECT 1.11 84.36 1.37 84.62 ;
        RECT 1.11 83.6 1.37 83.86 ;
        RECT 1.11 82.84 1.37 83.1 ;
        RECT 1.11 82.08 1.37 82.34 ;
        RECT 1.11 81.32 1.37 81.58 ;
        RECT 1.11 80.56 1.37 80.82 ;
        RECT 1.11 79.8 1.37 80.06 ;
        RECT 1.11 79.04 1.37 79.3 ;
        RECT 1.11 78.28 1.37 78.54 ;
        RECT 1.11 77.52 1.37 77.78 ;
        RECT 1.11 76.76 1.37 77.02 ;
        RECT 1.11 76 1.37 76.26 ;
        RECT 1.11 75.24 1.37 75.5 ;
        RECT 1.11 74.48 1.37 74.74 ;
        RECT 1.11 73.72 1.37 73.98 ;
        RECT 1.11 72.96 1.37 73.22 ;
        RECT 1.11 72.2 1.37 72.46 ;
        RECT 1.11 71.44 1.37 71.7 ;
        RECT 1.11 70.68 1.37 70.94 ;
        RECT 1.11 69.92 1.37 70.18 ;
        RECT 1.11 69.16 1.37 69.42 ;
        RECT 1.87 91.2 2.13 91.46 ;
        RECT 1.87 90.44 2.13 90.7 ;
        RECT 1.87 89.68 2.13 89.94 ;
        RECT 1.87 88.92 2.13 89.18 ;
        RECT 1.87 88.16 2.13 88.42 ;
        RECT 1.87 87.4 2.13 87.66 ;
        RECT 1.87 86.64 2.13 86.9 ;
        RECT 1.87 85.88 2.13 86.14 ;
        RECT 1.87 85.12 2.13 85.38 ;
        RECT 1.87 84.36 2.13 84.62 ;
        RECT 1.87 83.6 2.13 83.86 ;
        RECT 1.87 82.84 2.13 83.1 ;
        RECT 1.87 82.08 2.13 82.34 ;
        RECT 1.87 81.32 2.13 81.58 ;
        RECT 1.87 80.56 2.13 80.82 ;
        RECT 1.87 79.8 2.13 80.06 ;
        RECT 1.87 79.04 2.13 79.3 ;
        RECT 1.87 78.28 2.13 78.54 ;
        RECT 1.87 77.52 2.13 77.78 ;
        RECT 1.87 76.76 2.13 77.02 ;
        RECT 1.87 76 2.13 76.26 ;
        RECT 1.87 75.24 2.13 75.5 ;
        RECT 1.87 74.48 2.13 74.74 ;
        RECT 1.87 73.72 2.13 73.98 ;
        RECT 1.87 72.96 2.13 73.22 ;
        RECT 1.87 72.2 2.13 72.46 ;
        RECT 1.87 71.44 2.13 71.7 ;
        RECT 1.87 70.68 2.13 70.94 ;
        RECT 1.87 69.92 2.13 70.18 ;
        RECT 1.87 69.16 2.13 69.42 ;
        RECT 2.63 91.2 2.89 91.46 ;
        RECT 2.63 90.44 2.89 90.7 ;
        RECT 2.63 89.68 2.89 89.94 ;
        RECT 2.63 88.92 2.89 89.18 ;
        RECT 2.63 88.16 2.89 88.42 ;
        RECT 2.63 87.4 2.89 87.66 ;
        RECT 2.63 86.64 2.89 86.9 ;
        RECT 2.63 85.88 2.89 86.14 ;
        RECT 2.63 85.12 2.89 85.38 ;
        RECT 2.63 84.36 2.89 84.62 ;
        RECT 2.63 83.6 2.89 83.86 ;
        RECT 2.63 82.84 2.89 83.1 ;
        RECT 2.63 82.08 2.89 82.34 ;
        RECT 2.63 81.32 2.89 81.58 ;
        RECT 2.63 80.56 2.89 80.82 ;
        RECT 2.63 79.8 2.89 80.06 ;
        RECT 2.63 79.04 2.89 79.3 ;
        RECT 2.63 78.28 2.89 78.54 ;
        RECT 2.63 77.52 2.89 77.78 ;
        RECT 2.63 76.76 2.89 77.02 ;
        RECT 2.63 76 2.89 76.26 ;
        RECT 2.63 75.24 2.89 75.5 ;
        RECT 2.63 74.48 2.89 74.74 ;
        RECT 2.63 73.72 2.89 73.98 ;
        RECT 2.63 72.96 2.89 73.22 ;
        RECT 2.63 72.2 2.89 72.46 ;
        RECT 2.63 71.44 2.89 71.7 ;
        RECT 2.63 70.68 2.89 70.94 ;
        RECT 2.63 69.92 2.89 70.18 ;
        RECT 2.63 69.16 2.89 69.42 ;
        RECT 3.39 91.2 3.65 91.46 ;
        RECT 3.39 90.44 3.65 90.7 ;
        RECT 3.39 89.68 3.65 89.94 ;
        RECT 3.39 88.92 3.65 89.18 ;
        RECT 3.39 88.16 3.65 88.42 ;
        RECT 3.39 87.4 3.65 87.66 ;
        RECT 3.39 86.64 3.65 86.9 ;
        RECT 3.39 85.88 3.65 86.14 ;
        RECT 3.39 85.12 3.65 85.38 ;
        RECT 3.39 84.36 3.65 84.62 ;
        RECT 3.39 83.6 3.65 83.86 ;
        RECT 3.39 82.84 3.65 83.1 ;
        RECT 3.39 82.08 3.65 82.34 ;
        RECT 3.39 81.32 3.65 81.58 ;
        RECT 3.39 80.56 3.65 80.82 ;
        RECT 3.39 79.8 3.65 80.06 ;
        RECT 3.39 79.04 3.65 79.3 ;
        RECT 3.39 78.28 3.65 78.54 ;
        RECT 3.39 77.52 3.65 77.78 ;
        RECT 3.39 76.76 3.65 77.02 ;
        RECT 3.39 76 3.65 76.26 ;
        RECT 3.39 75.24 3.65 75.5 ;
        RECT 3.39 74.48 3.65 74.74 ;
        RECT 3.39 73.72 3.65 73.98 ;
        RECT 3.39 72.96 3.65 73.22 ;
        RECT 3.39 72.2 3.65 72.46 ;
        RECT 3.39 71.44 3.65 71.7 ;
        RECT 3.39 70.68 3.65 70.94 ;
        RECT 3.39 69.92 3.65 70.18 ;
        RECT 3.39 69.16 3.65 69.42 ;
        RECT 96.35 91.2 96.61 91.46 ;
        RECT 96.35 90.44 96.61 90.7 ;
        RECT 96.35 89.68 96.61 89.94 ;
        RECT 96.35 88.92 96.61 89.18 ;
        RECT 96.35 88.16 96.61 88.42 ;
        RECT 96.35 87.4 96.61 87.66 ;
        RECT 96.35 86.64 96.61 86.9 ;
        RECT 96.35 85.88 96.61 86.14 ;
        RECT 96.35 85.12 96.61 85.38 ;
        RECT 96.35 84.36 96.61 84.62 ;
        RECT 96.35 83.6 96.61 83.86 ;
        RECT 96.35 82.84 96.61 83.1 ;
        RECT 96.35 82.08 96.61 82.34 ;
        RECT 96.35 81.32 96.61 81.58 ;
        RECT 96.35 80.56 96.61 80.82 ;
        RECT 96.35 79.8 96.61 80.06 ;
        RECT 96.35 79.04 96.61 79.3 ;
        RECT 96.35 78.28 96.61 78.54 ;
        RECT 96.35 77.52 96.61 77.78 ;
        RECT 96.35 76.76 96.61 77.02 ;
        RECT 96.35 76 96.61 76.26 ;
        RECT 96.35 75.24 96.61 75.5 ;
        RECT 96.35 74.48 96.61 74.74 ;
        RECT 96.35 73.72 96.61 73.98 ;
        RECT 96.35 72.96 96.61 73.22 ;
        RECT 96.35 72.2 96.61 72.46 ;
        RECT 96.35 71.44 96.61 71.7 ;
        RECT 96.35 70.68 96.61 70.94 ;
        RECT 96.35 69.92 96.61 70.18 ;
        RECT 96.35 69.16 96.61 69.42 ;
        RECT 97.11 91.2 97.37 91.46 ;
        RECT 97.11 90.44 97.37 90.7 ;
        RECT 97.11 89.68 97.37 89.94 ;
        RECT 97.11 88.92 97.37 89.18 ;
        RECT 97.11 88.16 97.37 88.42 ;
        RECT 97.11 87.4 97.37 87.66 ;
        RECT 97.11 86.64 97.37 86.9 ;
        RECT 97.11 85.88 97.37 86.14 ;
        RECT 97.11 85.12 97.37 85.38 ;
        RECT 97.11 84.36 97.37 84.62 ;
        RECT 97.11 83.6 97.37 83.86 ;
        RECT 97.11 82.84 97.37 83.1 ;
        RECT 97.11 82.08 97.37 82.34 ;
        RECT 97.11 81.32 97.37 81.58 ;
        RECT 97.11 80.56 97.37 80.82 ;
        RECT 97.11 79.8 97.37 80.06 ;
        RECT 97.11 79.04 97.37 79.3 ;
        RECT 97.11 78.28 97.37 78.54 ;
        RECT 97.11 77.52 97.37 77.78 ;
        RECT 97.11 76.76 97.37 77.02 ;
        RECT 97.11 76 97.37 76.26 ;
        RECT 97.11 75.24 97.37 75.5 ;
        RECT 97.11 74.48 97.37 74.74 ;
        RECT 97.11 73.72 97.37 73.98 ;
        RECT 97.11 72.96 97.37 73.22 ;
        RECT 97.11 72.2 97.37 72.46 ;
        RECT 97.11 71.44 97.37 71.7 ;
        RECT 97.11 70.68 97.37 70.94 ;
        RECT 97.11 69.92 97.37 70.18 ;
        RECT 97.11 69.16 97.37 69.42 ;
        RECT 97.87 91.2 98.13 91.46 ;
        RECT 97.87 90.44 98.13 90.7 ;
        RECT 97.87 89.68 98.13 89.94 ;
        RECT 97.87 88.92 98.13 89.18 ;
        RECT 97.87 88.16 98.13 88.42 ;
        RECT 97.87 87.4 98.13 87.66 ;
        RECT 97.87 86.64 98.13 86.9 ;
        RECT 97.87 85.88 98.13 86.14 ;
        RECT 97.87 85.12 98.13 85.38 ;
        RECT 97.87 84.36 98.13 84.62 ;
        RECT 97.87 83.6 98.13 83.86 ;
        RECT 97.87 82.84 98.13 83.1 ;
        RECT 97.87 82.08 98.13 82.34 ;
        RECT 97.87 81.32 98.13 81.58 ;
        RECT 97.87 80.56 98.13 80.82 ;
        RECT 97.87 79.8 98.13 80.06 ;
        RECT 97.87 79.04 98.13 79.3 ;
        RECT 97.87 78.28 98.13 78.54 ;
        RECT 97.87 77.52 98.13 77.78 ;
        RECT 97.87 76.76 98.13 77.02 ;
        RECT 97.87 76 98.13 76.26 ;
        RECT 97.87 75.24 98.13 75.5 ;
        RECT 97.87 74.48 98.13 74.74 ;
        RECT 97.87 73.72 98.13 73.98 ;
        RECT 97.87 72.96 98.13 73.22 ;
        RECT 97.87 72.2 98.13 72.46 ;
        RECT 97.87 71.44 98.13 71.7 ;
        RECT 97.87 70.68 98.13 70.94 ;
        RECT 97.87 69.92 98.13 70.18 ;
        RECT 97.87 69.16 98.13 69.42 ;
        RECT 98.63 91.2 98.89 91.46 ;
        RECT 98.63 90.44 98.89 90.7 ;
        RECT 98.63 89.68 98.89 89.94 ;
        RECT 98.63 88.92 98.89 89.18 ;
        RECT 98.63 88.16 98.89 88.42 ;
        RECT 98.63 87.4 98.89 87.66 ;
        RECT 98.63 86.64 98.89 86.9 ;
        RECT 98.63 85.88 98.89 86.14 ;
        RECT 98.63 85.12 98.89 85.38 ;
        RECT 98.63 84.36 98.89 84.62 ;
        RECT 98.63 83.6 98.89 83.86 ;
        RECT 98.63 82.84 98.89 83.1 ;
        RECT 98.63 82.08 98.89 82.34 ;
        RECT 98.63 81.32 98.89 81.58 ;
        RECT 98.63 80.56 98.89 80.82 ;
        RECT 98.63 79.8 98.89 80.06 ;
        RECT 98.63 79.04 98.89 79.3 ;
        RECT 98.63 78.28 98.89 78.54 ;
        RECT 98.63 77.52 98.89 77.78 ;
        RECT 98.63 76.76 98.89 77.02 ;
        RECT 98.63 76 98.89 76.26 ;
        RECT 98.63 75.24 98.89 75.5 ;
        RECT 98.63 74.48 98.89 74.74 ;
        RECT 98.63 73.72 98.89 73.98 ;
        RECT 98.63 72.96 98.89 73.22 ;
        RECT 98.63 72.2 98.89 72.46 ;
        RECT 98.63 71.44 98.89 71.7 ;
        RECT 98.63 70.68 98.89 70.94 ;
        RECT 98.63 69.92 98.89 70.18 ;
        RECT 98.63 69.16 98.89 69.42 ;
        RECT 99.39 91.2 99.65 91.46 ;
        RECT 99.39 90.44 99.65 90.7 ;
        RECT 99.39 89.68 99.65 89.94 ;
        RECT 99.39 88.92 99.65 89.18 ;
        RECT 99.39 88.16 99.65 88.42 ;
        RECT 99.39 87.4 99.65 87.66 ;
        RECT 99.39 86.64 99.65 86.9 ;
        RECT 99.39 85.88 99.65 86.14 ;
        RECT 99.39 85.12 99.65 85.38 ;
        RECT 99.39 84.36 99.65 84.62 ;
        RECT 99.39 83.6 99.65 83.86 ;
        RECT 99.39 82.84 99.65 83.1 ;
        RECT 99.39 82.08 99.65 82.34 ;
        RECT 99.39 81.32 99.65 81.58 ;
        RECT 99.39 80.56 99.65 80.82 ;
        RECT 99.39 79.8 99.65 80.06 ;
        RECT 99.39 79.04 99.65 79.3 ;
        RECT 99.39 78.28 99.65 78.54 ;
        RECT 99.39 77.52 99.65 77.78 ;
        RECT 99.39 76.76 99.65 77.02 ;
        RECT 99.39 76 99.65 76.26 ;
        RECT 99.39 75.24 99.65 75.5 ;
        RECT 99.39 74.48 99.65 74.74 ;
        RECT 99.39 73.72 99.65 73.98 ;
        RECT 99.39 72.96 99.65 73.22 ;
        RECT 99.39 72.2 99.65 72.46 ;
        RECT 99.39 71.44 99.65 71.7 ;
        RECT 99.39 70.68 99.65 70.94 ;
        RECT 99.39 69.92 99.65 70.18 ;
        RECT 99.39 69.16 99.65 69.42 ;
    END
  END DVSS
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
        RECT 0 34 100 64 ;
      LAYER M3 ;
        RECT 0 34 100 64 ;
      LAYER V4 ;
        RECT 0.35 58.725 0.61 58.985 ;
        RECT 0.35 57.965 0.61 58.225 ;
        RECT 0.35 57.205 0.61 57.465 ;
        RECT 0.35 56.445 0.61 56.705 ;
        RECT 0.35 55.685 0.61 55.945 ;
        RECT 0.35 54.925 0.61 55.185 ;
        RECT 0.35 54.165 0.61 54.425 ;
        RECT 0.35 53.405 0.61 53.665 ;
        RECT 0.35 52.645 0.61 52.905 ;
        RECT 0.35 51.885 0.61 52.145 ;
        RECT 0.35 51.125 0.61 51.385 ;
        RECT 0.35 50.365 0.61 50.625 ;
        RECT 0.35 49.605 0.61 49.865 ;
        RECT 0.35 48.845 0.61 49.105 ;
        RECT 0.35 48.085 0.61 48.345 ;
        RECT 0.35 47.325 0.61 47.585 ;
        RECT 0.35 46.565 0.61 46.825 ;
        RECT 0.35 45.805 0.61 46.065 ;
        RECT 0.35 45.045 0.61 45.305 ;
        RECT 0.35 44.285 0.61 44.545 ;
        RECT 0.35 43.525 0.61 43.785 ;
        RECT 0.35 42.765 0.61 43.025 ;
        RECT 0.35 42.005 0.61 42.265 ;
        RECT 0.35 41.245 0.61 41.505 ;
        RECT 0.35 40.485 0.61 40.745 ;
        RECT 0.35 39.725 0.61 39.985 ;
        RECT 0.35 38.965 0.61 39.225 ;
        RECT 0.35 38.205 0.61 38.465 ;
        RECT 0.35 37.445 0.61 37.705 ;
        RECT 0.35 36.685 0.61 36.945 ;
        RECT 1.11 58.725 1.37 58.985 ;
        RECT 1.11 57.965 1.37 58.225 ;
        RECT 1.11 57.205 1.37 57.465 ;
        RECT 1.11 56.445 1.37 56.705 ;
        RECT 1.11 55.685 1.37 55.945 ;
        RECT 1.11 54.925 1.37 55.185 ;
        RECT 1.11 54.165 1.37 54.425 ;
        RECT 1.11 53.405 1.37 53.665 ;
        RECT 1.11 52.645 1.37 52.905 ;
        RECT 1.11 51.885 1.37 52.145 ;
        RECT 1.11 51.125 1.37 51.385 ;
        RECT 1.11 50.365 1.37 50.625 ;
        RECT 1.11 49.605 1.37 49.865 ;
        RECT 1.11 48.845 1.37 49.105 ;
        RECT 1.11 48.085 1.37 48.345 ;
        RECT 1.11 47.325 1.37 47.585 ;
        RECT 1.11 46.565 1.37 46.825 ;
        RECT 1.11 45.805 1.37 46.065 ;
        RECT 1.11 45.045 1.37 45.305 ;
        RECT 1.11 44.285 1.37 44.545 ;
        RECT 1.11 43.525 1.37 43.785 ;
        RECT 1.11 42.765 1.37 43.025 ;
        RECT 1.11 42.005 1.37 42.265 ;
        RECT 1.11 41.245 1.37 41.505 ;
        RECT 1.11 40.485 1.37 40.745 ;
        RECT 1.11 39.725 1.37 39.985 ;
        RECT 1.11 38.965 1.37 39.225 ;
        RECT 1.11 38.205 1.37 38.465 ;
        RECT 1.11 37.445 1.37 37.705 ;
        RECT 1.11 36.685 1.37 36.945 ;
        RECT 1.87 58.725 2.13 58.985 ;
        RECT 1.87 57.965 2.13 58.225 ;
        RECT 1.87 57.205 2.13 57.465 ;
        RECT 1.87 56.445 2.13 56.705 ;
        RECT 1.87 55.685 2.13 55.945 ;
        RECT 1.87 54.925 2.13 55.185 ;
        RECT 1.87 54.165 2.13 54.425 ;
        RECT 1.87 53.405 2.13 53.665 ;
        RECT 1.87 52.645 2.13 52.905 ;
        RECT 1.87 51.885 2.13 52.145 ;
        RECT 1.87 51.125 2.13 51.385 ;
        RECT 1.87 50.365 2.13 50.625 ;
        RECT 1.87 49.605 2.13 49.865 ;
        RECT 1.87 48.845 2.13 49.105 ;
        RECT 1.87 48.085 2.13 48.345 ;
        RECT 1.87 47.325 2.13 47.585 ;
        RECT 1.87 46.565 2.13 46.825 ;
        RECT 1.87 45.805 2.13 46.065 ;
        RECT 1.87 45.045 2.13 45.305 ;
        RECT 1.87 44.285 2.13 44.545 ;
        RECT 1.87 43.525 2.13 43.785 ;
        RECT 1.87 42.765 2.13 43.025 ;
        RECT 1.87 42.005 2.13 42.265 ;
        RECT 1.87 41.245 2.13 41.505 ;
        RECT 1.87 40.485 2.13 40.745 ;
        RECT 1.87 39.725 2.13 39.985 ;
        RECT 1.87 38.965 2.13 39.225 ;
        RECT 1.87 38.205 2.13 38.465 ;
        RECT 1.87 37.445 2.13 37.705 ;
        RECT 1.87 36.685 2.13 36.945 ;
        RECT 2.63 58.725 2.89 58.985 ;
        RECT 2.63 57.965 2.89 58.225 ;
        RECT 2.63 57.205 2.89 57.465 ;
        RECT 2.63 56.445 2.89 56.705 ;
        RECT 2.63 55.685 2.89 55.945 ;
        RECT 2.63 54.925 2.89 55.185 ;
        RECT 2.63 54.165 2.89 54.425 ;
        RECT 2.63 53.405 2.89 53.665 ;
        RECT 2.63 52.645 2.89 52.905 ;
        RECT 2.63 51.885 2.89 52.145 ;
        RECT 2.63 51.125 2.89 51.385 ;
        RECT 2.63 50.365 2.89 50.625 ;
        RECT 2.63 49.605 2.89 49.865 ;
        RECT 2.63 48.845 2.89 49.105 ;
        RECT 2.63 48.085 2.89 48.345 ;
        RECT 2.63 47.325 2.89 47.585 ;
        RECT 2.63 46.565 2.89 46.825 ;
        RECT 2.63 45.805 2.89 46.065 ;
        RECT 2.63 45.045 2.89 45.305 ;
        RECT 2.63 44.285 2.89 44.545 ;
        RECT 2.63 43.525 2.89 43.785 ;
        RECT 2.63 42.765 2.89 43.025 ;
        RECT 2.63 42.005 2.89 42.265 ;
        RECT 2.63 41.245 2.89 41.505 ;
        RECT 2.63 40.485 2.89 40.745 ;
        RECT 2.63 39.725 2.89 39.985 ;
        RECT 2.63 38.965 2.89 39.225 ;
        RECT 2.63 38.205 2.89 38.465 ;
        RECT 2.63 37.445 2.89 37.705 ;
        RECT 2.63 36.685 2.89 36.945 ;
        RECT 3.39 58.725 3.65 58.985 ;
        RECT 3.39 57.965 3.65 58.225 ;
        RECT 3.39 57.205 3.65 57.465 ;
        RECT 3.39 56.445 3.65 56.705 ;
        RECT 3.39 55.685 3.65 55.945 ;
        RECT 3.39 54.925 3.65 55.185 ;
        RECT 3.39 54.165 3.65 54.425 ;
        RECT 3.39 53.405 3.65 53.665 ;
        RECT 3.39 52.645 3.65 52.905 ;
        RECT 3.39 51.885 3.65 52.145 ;
        RECT 3.39 51.125 3.65 51.385 ;
        RECT 3.39 50.365 3.65 50.625 ;
        RECT 3.39 49.605 3.65 49.865 ;
        RECT 3.39 48.845 3.65 49.105 ;
        RECT 3.39 48.085 3.65 48.345 ;
        RECT 3.39 47.325 3.65 47.585 ;
        RECT 3.39 46.565 3.65 46.825 ;
        RECT 3.39 45.805 3.65 46.065 ;
        RECT 3.39 45.045 3.65 45.305 ;
        RECT 3.39 44.285 3.65 44.545 ;
        RECT 3.39 43.525 3.65 43.785 ;
        RECT 3.39 42.765 3.65 43.025 ;
        RECT 3.39 42.005 3.65 42.265 ;
        RECT 3.39 41.245 3.65 41.505 ;
        RECT 3.39 40.485 3.65 40.745 ;
        RECT 3.39 39.725 3.65 39.985 ;
        RECT 3.39 38.965 3.65 39.225 ;
        RECT 3.39 38.205 3.65 38.465 ;
        RECT 3.39 37.445 3.65 37.705 ;
        RECT 3.39 36.685 3.65 36.945 ;
        RECT 96.35 58.725 96.61 58.985 ;
        RECT 96.35 57.965 96.61 58.225 ;
        RECT 96.35 57.205 96.61 57.465 ;
        RECT 96.35 56.445 96.61 56.705 ;
        RECT 96.35 55.685 96.61 55.945 ;
        RECT 96.35 54.925 96.61 55.185 ;
        RECT 96.35 54.165 96.61 54.425 ;
        RECT 96.35 53.405 96.61 53.665 ;
        RECT 96.35 52.645 96.61 52.905 ;
        RECT 96.35 51.885 96.61 52.145 ;
        RECT 96.35 51.125 96.61 51.385 ;
        RECT 96.35 50.365 96.61 50.625 ;
        RECT 96.35 49.605 96.61 49.865 ;
        RECT 96.35 48.845 96.61 49.105 ;
        RECT 96.35 48.085 96.61 48.345 ;
        RECT 96.35 47.325 96.61 47.585 ;
        RECT 96.35 46.565 96.61 46.825 ;
        RECT 96.35 45.805 96.61 46.065 ;
        RECT 96.35 45.045 96.61 45.305 ;
        RECT 96.35 44.285 96.61 44.545 ;
        RECT 96.35 43.525 96.61 43.785 ;
        RECT 96.35 42.765 96.61 43.025 ;
        RECT 96.35 42.005 96.61 42.265 ;
        RECT 96.35 41.245 96.61 41.505 ;
        RECT 96.35 40.485 96.61 40.745 ;
        RECT 96.35 39.725 96.61 39.985 ;
        RECT 96.35 38.965 96.61 39.225 ;
        RECT 96.35 38.205 96.61 38.465 ;
        RECT 96.35 37.445 96.61 37.705 ;
        RECT 96.35 36.685 96.61 36.945 ;
        RECT 97.11 58.725 97.37 58.985 ;
        RECT 97.11 57.965 97.37 58.225 ;
        RECT 97.11 57.205 97.37 57.465 ;
        RECT 97.11 56.445 97.37 56.705 ;
        RECT 97.11 55.685 97.37 55.945 ;
        RECT 97.11 54.925 97.37 55.185 ;
        RECT 97.11 54.165 97.37 54.425 ;
        RECT 97.11 53.405 97.37 53.665 ;
        RECT 97.11 52.645 97.37 52.905 ;
        RECT 97.11 51.885 97.37 52.145 ;
        RECT 97.11 51.125 97.37 51.385 ;
        RECT 97.11 50.365 97.37 50.625 ;
        RECT 97.11 49.605 97.37 49.865 ;
        RECT 97.11 48.845 97.37 49.105 ;
        RECT 97.11 48.085 97.37 48.345 ;
        RECT 97.11 47.325 97.37 47.585 ;
        RECT 97.11 46.565 97.37 46.825 ;
        RECT 97.11 45.805 97.37 46.065 ;
        RECT 97.11 45.045 97.37 45.305 ;
        RECT 97.11 44.285 97.37 44.545 ;
        RECT 97.11 43.525 97.37 43.785 ;
        RECT 97.11 42.765 97.37 43.025 ;
        RECT 97.11 42.005 97.37 42.265 ;
        RECT 97.11 41.245 97.37 41.505 ;
        RECT 97.11 40.485 97.37 40.745 ;
        RECT 97.11 39.725 97.37 39.985 ;
        RECT 97.11 38.965 97.37 39.225 ;
        RECT 97.11 38.205 97.37 38.465 ;
        RECT 97.11 37.445 97.37 37.705 ;
        RECT 97.11 36.685 97.37 36.945 ;
        RECT 97.87 58.725 98.13 58.985 ;
        RECT 97.87 57.965 98.13 58.225 ;
        RECT 97.87 57.205 98.13 57.465 ;
        RECT 97.87 56.445 98.13 56.705 ;
        RECT 97.87 55.685 98.13 55.945 ;
        RECT 97.87 54.925 98.13 55.185 ;
        RECT 97.87 54.165 98.13 54.425 ;
        RECT 97.87 53.405 98.13 53.665 ;
        RECT 97.87 52.645 98.13 52.905 ;
        RECT 97.87 51.885 98.13 52.145 ;
        RECT 97.87 51.125 98.13 51.385 ;
        RECT 97.87 50.365 98.13 50.625 ;
        RECT 97.87 49.605 98.13 49.865 ;
        RECT 97.87 48.845 98.13 49.105 ;
        RECT 97.87 48.085 98.13 48.345 ;
        RECT 97.87 47.325 98.13 47.585 ;
        RECT 97.87 46.565 98.13 46.825 ;
        RECT 97.87 45.805 98.13 46.065 ;
        RECT 97.87 45.045 98.13 45.305 ;
        RECT 97.87 44.285 98.13 44.545 ;
        RECT 97.87 43.525 98.13 43.785 ;
        RECT 97.87 42.765 98.13 43.025 ;
        RECT 97.87 42.005 98.13 42.265 ;
        RECT 97.87 41.245 98.13 41.505 ;
        RECT 97.87 40.485 98.13 40.745 ;
        RECT 97.87 39.725 98.13 39.985 ;
        RECT 97.87 38.965 98.13 39.225 ;
        RECT 97.87 38.205 98.13 38.465 ;
        RECT 97.87 37.445 98.13 37.705 ;
        RECT 97.87 36.685 98.13 36.945 ;
        RECT 98.63 58.725 98.89 58.985 ;
        RECT 98.63 57.965 98.89 58.225 ;
        RECT 98.63 57.205 98.89 57.465 ;
        RECT 98.63 56.445 98.89 56.705 ;
        RECT 98.63 55.685 98.89 55.945 ;
        RECT 98.63 54.925 98.89 55.185 ;
        RECT 98.63 54.165 98.89 54.425 ;
        RECT 98.63 53.405 98.89 53.665 ;
        RECT 98.63 52.645 98.89 52.905 ;
        RECT 98.63 51.885 98.89 52.145 ;
        RECT 98.63 51.125 98.89 51.385 ;
        RECT 98.63 50.365 98.89 50.625 ;
        RECT 98.63 49.605 98.89 49.865 ;
        RECT 98.63 48.845 98.89 49.105 ;
        RECT 98.63 48.085 98.89 48.345 ;
        RECT 98.63 47.325 98.89 47.585 ;
        RECT 98.63 46.565 98.89 46.825 ;
        RECT 98.63 45.805 98.89 46.065 ;
        RECT 98.63 45.045 98.89 45.305 ;
        RECT 98.63 44.285 98.89 44.545 ;
        RECT 98.63 43.525 98.89 43.785 ;
        RECT 98.63 42.765 98.89 43.025 ;
        RECT 98.63 42.005 98.89 42.265 ;
        RECT 98.63 41.245 98.89 41.505 ;
        RECT 98.63 40.485 98.89 40.745 ;
        RECT 98.63 39.725 98.89 39.985 ;
        RECT 98.63 38.965 98.89 39.225 ;
        RECT 98.63 38.205 98.89 38.465 ;
        RECT 98.63 37.445 98.89 37.705 ;
        RECT 98.63 36.685 98.89 36.945 ;
        RECT 99.39 58.725 99.65 58.985 ;
        RECT 99.39 57.965 99.65 58.225 ;
        RECT 99.39 57.205 99.65 57.465 ;
        RECT 99.39 56.445 99.65 56.705 ;
        RECT 99.39 55.685 99.65 55.945 ;
        RECT 99.39 54.925 99.65 55.185 ;
        RECT 99.39 54.165 99.65 54.425 ;
        RECT 99.39 53.405 99.65 53.665 ;
        RECT 99.39 52.645 99.65 52.905 ;
        RECT 99.39 51.885 99.65 52.145 ;
        RECT 99.39 51.125 99.65 51.385 ;
        RECT 99.39 50.365 99.65 50.625 ;
        RECT 99.39 49.605 99.65 49.865 ;
        RECT 99.39 48.845 99.65 49.105 ;
        RECT 99.39 48.085 99.65 48.345 ;
        RECT 99.39 47.325 99.65 47.585 ;
        RECT 99.39 46.565 99.65 46.825 ;
        RECT 99.39 45.805 99.65 46.065 ;
        RECT 99.39 45.045 99.65 45.305 ;
        RECT 99.39 44.285 99.65 44.545 ;
        RECT 99.39 43.525 99.65 43.785 ;
        RECT 99.39 42.765 99.65 43.025 ;
        RECT 99.39 42.005 99.65 42.265 ;
        RECT 99.39 41.245 99.65 41.505 ;
        RECT 99.39 40.485 99.65 40.745 ;
        RECT 99.39 39.725 99.65 39.985 ;
        RECT 99.39 38.965 99.65 39.225 ;
        RECT 99.39 38.205 99.65 38.465 ;
        RECT 99.39 37.445 99.65 37.705 ;
        RECT 99.39 36.685 99.65 36.945 ;
    END
  END DVDD
  PIN AVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
        RECT 0 22 100 32 ;
      LAYER M3 ;
        RECT 0 22 100 32 ;
      LAYER V4 ;
        RECT 0.35 30.215 0.61 30.475 ;
        RECT 0.35 29.455 0.61 29.715 ;
        RECT 0.35 28.695 0.61 28.955 ;
        RECT 0.35 27.935 0.61 28.195 ;
        RECT 0.35 27.175 0.61 27.435 ;
        RECT 0.35 26.415 0.61 26.675 ;
        RECT 0.35 25.655 0.61 25.915 ;
        RECT 0.35 24.895 0.61 25.155 ;
        RECT 0.35 24.135 0.61 24.395 ;
        RECT 0.35 23.375 0.61 23.635 ;
        RECT 1.11 30.215 1.37 30.475 ;
        RECT 1.11 29.455 1.37 29.715 ;
        RECT 1.11 28.695 1.37 28.955 ;
        RECT 1.11 27.935 1.37 28.195 ;
        RECT 1.11 27.175 1.37 27.435 ;
        RECT 1.11 26.415 1.37 26.675 ;
        RECT 1.11 25.655 1.37 25.915 ;
        RECT 1.11 24.895 1.37 25.155 ;
        RECT 1.11 24.135 1.37 24.395 ;
        RECT 1.11 23.375 1.37 23.635 ;
        RECT 1.87 30.215 2.13 30.475 ;
        RECT 1.87 29.455 2.13 29.715 ;
        RECT 1.87 28.695 2.13 28.955 ;
        RECT 1.87 27.935 2.13 28.195 ;
        RECT 1.87 27.175 2.13 27.435 ;
        RECT 1.87 26.415 2.13 26.675 ;
        RECT 1.87 25.655 2.13 25.915 ;
        RECT 1.87 24.895 2.13 25.155 ;
        RECT 1.87 24.135 2.13 24.395 ;
        RECT 1.87 23.375 2.13 23.635 ;
        RECT 2.63 30.215 2.89 30.475 ;
        RECT 2.63 29.455 2.89 29.715 ;
        RECT 2.63 28.695 2.89 28.955 ;
        RECT 2.63 27.935 2.89 28.195 ;
        RECT 2.63 27.175 2.89 27.435 ;
        RECT 2.63 26.415 2.89 26.675 ;
        RECT 2.63 25.655 2.89 25.915 ;
        RECT 2.63 24.895 2.89 25.155 ;
        RECT 2.63 24.135 2.89 24.395 ;
        RECT 2.63 23.375 2.89 23.635 ;
        RECT 3.39 30.215 3.65 30.475 ;
        RECT 3.39 29.455 3.65 29.715 ;
        RECT 3.39 28.695 3.65 28.955 ;
        RECT 3.39 27.935 3.65 28.195 ;
        RECT 3.39 27.175 3.65 27.435 ;
        RECT 3.39 26.415 3.65 26.675 ;
        RECT 3.39 25.655 3.65 25.915 ;
        RECT 3.39 24.895 3.65 25.155 ;
        RECT 3.39 24.135 3.65 24.395 ;
        RECT 3.39 23.375 3.65 23.635 ;
        RECT 96.35 30.215 96.61 30.475 ;
        RECT 96.35 29.455 96.61 29.715 ;
        RECT 96.35 28.695 96.61 28.955 ;
        RECT 96.35 27.935 96.61 28.195 ;
        RECT 96.35 27.175 96.61 27.435 ;
        RECT 96.35 26.415 96.61 26.675 ;
        RECT 96.35 25.655 96.61 25.915 ;
        RECT 96.35 24.895 96.61 25.155 ;
        RECT 96.35 24.135 96.61 24.395 ;
        RECT 96.35 23.375 96.61 23.635 ;
        RECT 97.11 30.215 97.37 30.475 ;
        RECT 97.11 29.455 97.37 29.715 ;
        RECT 97.11 28.695 97.37 28.955 ;
        RECT 97.11 27.935 97.37 28.195 ;
        RECT 97.11 27.175 97.37 27.435 ;
        RECT 97.11 26.415 97.37 26.675 ;
        RECT 97.11 25.655 97.37 25.915 ;
        RECT 97.11 24.895 97.37 25.155 ;
        RECT 97.11 24.135 97.37 24.395 ;
        RECT 97.11 23.375 97.37 23.635 ;
        RECT 97.87 30.215 98.13 30.475 ;
        RECT 97.87 29.455 98.13 29.715 ;
        RECT 97.87 28.695 98.13 28.955 ;
        RECT 97.87 27.935 98.13 28.195 ;
        RECT 97.87 27.175 98.13 27.435 ;
        RECT 97.87 26.415 98.13 26.675 ;
        RECT 97.87 25.655 98.13 25.915 ;
        RECT 97.87 24.895 98.13 25.155 ;
        RECT 97.87 24.135 98.13 24.395 ;
        RECT 97.87 23.375 98.13 23.635 ;
        RECT 98.63 30.215 98.89 30.475 ;
        RECT 98.63 29.455 98.89 29.715 ;
        RECT 98.63 28.695 98.89 28.955 ;
        RECT 98.63 27.935 98.89 28.195 ;
        RECT 98.63 27.175 98.89 27.435 ;
        RECT 98.63 26.415 98.89 26.675 ;
        RECT 98.63 25.655 98.89 25.915 ;
        RECT 98.63 24.895 98.89 25.155 ;
        RECT 98.63 24.135 98.89 24.395 ;
        RECT 98.63 23.375 98.89 23.635 ;
        RECT 99.39 30.215 99.65 30.475 ;
        RECT 99.39 29.455 99.65 29.715 ;
        RECT 99.39 28.695 99.65 28.955 ;
        RECT 99.39 27.935 99.65 28.195 ;
        RECT 99.39 27.175 99.65 27.435 ;
        RECT 99.39 26.415 99.65 26.675 ;
        RECT 99.39 25.655 99.65 25.915 ;
        RECT 99.39 24.895 99.65 25.155 ;
        RECT 99.39 24.135 99.65 24.395 ;
        RECT 99.39 23.375 99.65 23.635 ;
    END
  END AVSS
  PIN AVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
        RECT 0 10 100 20 ;
      LAYER M3 ;
        RECT 0 10 100 20 ;
      LAYER V4 ;
        RECT 0.35 18.24 0.61 18.5 ;
        RECT 0.35 17.48 0.61 17.74 ;
        RECT 0.35 16.72 0.61 16.98 ;
        RECT 0.35 15.96 0.61 16.22 ;
        RECT 0.35 15.2 0.61 15.46 ;
        RECT 0.35 14.44 0.61 14.7 ;
        RECT 0.35 13.68 0.61 13.94 ;
        RECT 0.35 12.92 0.61 13.18 ;
        RECT 0.35 12.16 0.61 12.42 ;
        RECT 0.35 11.4 0.61 11.66 ;
        RECT 1.11 18.24 1.37 18.5 ;
        RECT 1.11 17.48 1.37 17.74 ;
        RECT 1.11 16.72 1.37 16.98 ;
        RECT 1.11 15.96 1.37 16.22 ;
        RECT 1.11 15.2 1.37 15.46 ;
        RECT 1.11 14.44 1.37 14.7 ;
        RECT 1.11 13.68 1.37 13.94 ;
        RECT 1.11 12.92 1.37 13.18 ;
        RECT 1.11 12.16 1.37 12.42 ;
        RECT 1.11 11.4 1.37 11.66 ;
        RECT 1.87 18.24 2.13 18.5 ;
        RECT 1.87 17.48 2.13 17.74 ;
        RECT 1.87 16.72 2.13 16.98 ;
        RECT 1.87 15.96 2.13 16.22 ;
        RECT 1.87 15.2 2.13 15.46 ;
        RECT 1.87 14.44 2.13 14.7 ;
        RECT 1.87 13.68 2.13 13.94 ;
        RECT 1.87 12.92 2.13 13.18 ;
        RECT 1.87 12.16 2.13 12.42 ;
        RECT 1.87 11.4 2.13 11.66 ;
        RECT 2.63 18.24 2.89 18.5 ;
        RECT 2.63 17.48 2.89 17.74 ;
        RECT 2.63 16.72 2.89 16.98 ;
        RECT 2.63 15.96 2.89 16.22 ;
        RECT 2.63 15.2 2.89 15.46 ;
        RECT 2.63 14.44 2.89 14.7 ;
        RECT 2.63 13.68 2.89 13.94 ;
        RECT 2.63 12.92 2.89 13.18 ;
        RECT 2.63 12.16 2.89 12.42 ;
        RECT 2.63 11.4 2.89 11.66 ;
        RECT 3.39 18.24 3.65 18.5 ;
        RECT 3.39 17.48 3.65 17.74 ;
        RECT 3.39 16.72 3.65 16.98 ;
        RECT 3.39 15.96 3.65 16.22 ;
        RECT 3.39 15.2 3.65 15.46 ;
        RECT 3.39 14.44 3.65 14.7 ;
        RECT 3.39 13.68 3.65 13.94 ;
        RECT 3.39 12.92 3.65 13.18 ;
        RECT 3.39 12.16 3.65 12.42 ;
        RECT 3.39 11.4 3.65 11.66 ;
        RECT 96.35 18.24 96.61 18.5 ;
        RECT 96.35 17.48 96.61 17.74 ;
        RECT 96.35 16.72 96.61 16.98 ;
        RECT 96.35 15.96 96.61 16.22 ;
        RECT 96.35 15.2 96.61 15.46 ;
        RECT 96.35 14.44 96.61 14.7 ;
        RECT 96.35 13.68 96.61 13.94 ;
        RECT 96.35 12.92 96.61 13.18 ;
        RECT 96.35 12.16 96.61 12.42 ;
        RECT 96.35 11.4 96.61 11.66 ;
        RECT 97.11 18.24 97.37 18.5 ;
        RECT 97.11 17.48 97.37 17.74 ;
        RECT 97.11 16.72 97.37 16.98 ;
        RECT 97.11 15.96 97.37 16.22 ;
        RECT 97.11 15.2 97.37 15.46 ;
        RECT 97.11 14.44 97.37 14.7 ;
        RECT 97.11 13.68 97.37 13.94 ;
        RECT 97.11 12.92 97.37 13.18 ;
        RECT 97.11 12.16 97.37 12.42 ;
        RECT 97.11 11.4 97.37 11.66 ;
        RECT 97.87 18.24 98.13 18.5 ;
        RECT 97.87 17.48 98.13 17.74 ;
        RECT 97.87 16.72 98.13 16.98 ;
        RECT 97.87 15.96 98.13 16.22 ;
        RECT 97.87 15.2 98.13 15.46 ;
        RECT 97.87 14.44 98.13 14.7 ;
        RECT 97.87 13.68 98.13 13.94 ;
        RECT 97.87 12.92 98.13 13.18 ;
        RECT 97.87 12.16 98.13 12.42 ;
        RECT 97.87 11.4 98.13 11.66 ;
        RECT 98.63 18.24 98.89 18.5 ;
        RECT 98.63 17.48 98.89 17.74 ;
        RECT 98.63 16.72 98.89 16.98 ;
        RECT 98.63 15.96 98.89 16.22 ;
        RECT 98.63 15.2 98.89 15.46 ;
        RECT 98.63 14.44 98.89 14.7 ;
        RECT 98.63 13.68 98.89 13.94 ;
        RECT 98.63 12.92 98.89 13.18 ;
        RECT 98.63 12.16 98.89 12.42 ;
        RECT 98.63 11.4 98.89 11.66 ;
        RECT 99.39 18.24 99.65 18.5 ;
        RECT 99.39 17.48 99.65 17.74 ;
        RECT 99.39 16.72 99.65 16.98 ;
        RECT 99.39 15.96 99.65 16.22 ;
        RECT 99.39 15.2 99.65 15.46 ;
        RECT 99.39 14.44 99.65 14.7 ;
        RECT 99.39 13.68 99.65 13.94 ;
        RECT 99.39 12.92 99.65 13.18 ;
        RECT 99.39 12.16 99.65 12.42 ;
        RECT 99.39 11.4 99.65 11.66 ;
    END
  END AVDD
  PIN DOUT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12.955 117 15.955 120 ;
    END
  END DOUT
  PIN CIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 84.56 117 87.56 120 ;
    END
  END CIN
  OBS
    LAYER M1 ;
      RECT 76.895 72.415 95.64 74.845 ;
      RECT 88.955 31.9 95.64 74.845 ;
      RECT 67.965 72.415 95.64 74.775 ;
      RECT 57.89 72.415 95.64 73.605 ;
      RECT 60.695 72.185 78.635 73.605 ;
      RECT 57.89 60.325 58.85 73.605 ;
      RECT 17 69.53 58.85 70.72 ;
      RECT 44.545 67.1 49.815 70.72 ;
      RECT 28.565 69.1 38.235 70.72 ;
      RECT 38.005 61.95 38.235 70.72 ;
      RECT 17.29 61.95 17.52 70.72 ;
      RECT 36.565 61.95 36.795 70.72 ;
      RECT 30.005 61.95 30.235 70.72 ;
      RECT 28.565 61.95 28.795 70.72 ;
      RECT 44.545 67.1 55.14 67.33 ;
      RECT 54.91 61.95 55.14 67.33 ;
      RECT 53.43 61.95 53.66 67.33 ;
      RECT 51.95 61.95 52.18 67.33 ;
      RECT 50.47 61.95 50.7 67.33 ;
      RECT 48.99 61.95 49.22 70.72 ;
      RECT 47.51 61.95 47.74 70.72 ;
      RECT 46.03 61.95 46.26 70.72 ;
      RECT 44.55 61.95 44.78 70.72 ;
      RECT 57.89 60.325 75.83 60.555 ;
      RECT 64.14 31.9 95.64 39.91 ;
      RECT 10.195 28.97 90.08 30.33 ;
      RECT 88.71 9.56 90.08 30.33 ;
      RECT 10.195 9.56 11.565 30.33 ;
      RECT 10.195 9.56 90.08 10.92 ;
      RECT 12.37 26.895 36.15 27.175 ;
      RECT 12.37 26.92 87.905 27.15 ;
      RECT 12.375 23.595 12.605 27.175 ;
      RECT 12.355 23.595 36.135 23.875 ;
      RECT 12.355 23.62 87.905 23.85 ;
      RECT 72.89 78.115 85.24 79.525 ;
      RECT 85.01 78.075 85.24 79.525 ;
      RECT 64.335 18.745 84.995 19.025 ;
      RECT 15.375 18.75 84.995 18.98 ;
      RECT 15.375 15.45 15.605 18.98 ;
      RECT 64.335 15.415 84.995 15.695 ;
      RECT 15.375 15.45 84.995 15.68 ;
      RECT 32.885 43.35 33.115 52.74 ;
      RECT 31.445 43.35 31.675 52.74 ;
      RECT 30.005 43.35 30.235 52.74 ;
      RECT 28.565 43.35 28.795 52.74 ;
      RECT 24.885 43.35 25.115 52.74 ;
      RECT 23.445 43.35 23.675 52.74 ;
      RECT 22.005 43.35 22.235 52.74 ;
      RECT 20.565 43.35 20.795 52.74 ;
      RECT 17.29 43.35 17.52 52.74 ;
      RECT 78.59 43.35 78.82 50.845 ;
      RECT 77.11 43.35 77.34 50.845 ;
      RECT 75.63 43.35 75.86 50.845 ;
      RECT 74.15 43.35 74.38 50.845 ;
      RECT 72.67 43.35 72.9 50.845 ;
      RECT 71.19 43.35 71.42 50.845 ;
      RECT 69.71 43.35 69.94 50.845 ;
      RECT 68.23 43.35 68.46 50.845 ;
      RECT 66.75 43.35 66.98 50.845 ;
      RECT 65.27 43.35 65.5 50.845 ;
      RECT 63.79 43.35 64.02 50.845 ;
      RECT 62.31 43.35 62.54 50.845 ;
      RECT 60.83 43.35 61.06 50.845 ;
      RECT 59.35 43.35 59.58 50.845 ;
      RECT 57.87 43.35 58.1 50.845 ;
      RECT 56.39 43.35 56.62 50.845 ;
      RECT 54.91 43.35 55.14 50.845 ;
      RECT 53.43 43.35 53.66 50.845 ;
      RECT 51.95 43.35 52.18 50.845 ;
      RECT 50.47 43.35 50.7 50.845 ;
      RECT 48.99 43.35 49.22 50.845 ;
      RECT 47.51 43.35 47.74 50.845 ;
      RECT 46.03 43.35 46.26 50.845 ;
      RECT 44.55 43.35 44.78 50.845 ;
      RECT 44.55 43.35 78.82 45.695 ;
      RECT 28.565 43.35 33.115 45.59 ;
      RECT 20.565 43.35 25.115 45.59 ;
      RECT 16.775 43.35 84.55 44.285 ;
      RECT 77.505 61.655 77.735 65.035 ;
      RECT 75.825 61.655 76.055 65.035 ;
      RECT 74.145 61.655 74.375 65.035 ;
      RECT 72.465 61.655 72.695 65.035 ;
      RECT 70.785 61.655 71.015 65.035 ;
      RECT 79.59 64.505 79.99 64.905 ;
      RECT 77.48 62.33 77.76 64.79 ;
      RECT 75.8 62.33 76.08 64.79 ;
      RECT 74.12 62.33 74.4 64.79 ;
      RECT 72.44 62.33 72.72 64.79 ;
      RECT 70.76 62.33 71.04 64.79 ;
      RECT 78.46 64.505 79.99 64.765 ;
      RECT 78.46 61.655 78.79 64.765 ;
      RECT 80.97 61.655 81.21 64.145 ;
      RECT 78.46 61.655 78.86 63.525 ;
      RECT 77.505 61.655 82.23 63.255 ;
      RECT 70.785 61.655 82.23 61.885 ;
      RECT 78.23 67.375 82.23 70.355 ;
      RECT 80.91 67.115 81.31 70.355 ;
      RECT 79.05 67.115 79.45 70.355 ;
      RECT 78.67 66.225 81.75 66.655 ;
      RECT 81.47 64.575 81.75 66.655 ;
      RECT 80.23 64.575 82.03 64.975 ;
      RECT 80.23 63.885 80.47 64.975 ;
      RECT 79.03 63.885 80.47 64.125 ;
      RECT 70.37 61.195 80.895 61.425 ;
      RECT 79.995 61.145 80.895 61.425 ;
      RECT 79.995 70.585 80.895 70.865 ;
      RECT 76.25 70.585 80.895 70.815 ;
      RECT 76.25 70.13 77.31 70.815 ;
      RECT 76.665 62.115 76.895 69.895 ;
      RECT 78.78 65.095 79.37 65.615 ;
      RECT 69.945 65.265 79.37 65.495 ;
      RECT 74.985 62.115 75.215 65.495 ;
      RECT 73.305 62.115 73.535 65.495 ;
      RECT 71.625 62.115 71.855 65.495 ;
      RECT 69.945 62.115 70.175 65.495 ;
      RECT 22.725 61.44 22.955 68.82 ;
      RECT 21.285 61.44 21.515 68.82 ;
      RECT 21.285 61.44 26.565 61.67 ;
      RECT 26.285 52.97 26.565 61.67 ;
      RECT 21.285 52.97 33.835 53.2 ;
      RECT 33.605 45.36 33.835 53.2 ;
      RECT 32.165 45.82 32.395 53.2 ;
      RECT 30.725 45.82 30.955 53.2 ;
      RECT 29.285 45.82 29.515 53.2 ;
      RECT 25.605 45.82 25.835 53.2 ;
      RECT 24.165 45.82 24.395 53.2 ;
      RECT 22.725 45.82 22.955 53.2 ;
      RECT 21.285 45.82 21.515 53.2 ;
      RECT 41.605 45.36 41.835 52.74 ;
      RECT 40.165 45.36 40.395 52.74 ;
      RECT 38.725 45.36 38.955 52.74 ;
      RECT 37.285 45.36 37.515 52.74 ;
      RECT 41.605 51.535 78.395 51.765 ;
      RECT 33.605 45.36 41.835 45.59 ;
      RECT 45.29 51.075 78.08 51.305 ;
      RECT 77.85 45.925 78.08 51.305 ;
      RECT 76.37 45.925 76.6 51.305 ;
      RECT 74.89 45.925 75.12 51.305 ;
      RECT 73.41 45.925 73.64 51.305 ;
      RECT 71.93 45.925 72.16 51.305 ;
      RECT 70.45 45.925 70.68 51.305 ;
      RECT 68.97 45.925 69.2 51.305 ;
      RECT 67.49 45.925 67.72 51.305 ;
      RECT 66.01 45.925 66.24 51.305 ;
      RECT 64.53 45.925 64.76 51.305 ;
      RECT 63.05 45.925 63.28 51.305 ;
      RECT 61.57 45.925 61.8 51.305 ;
      RECT 60.09 45.925 60.32 51.305 ;
      RECT 58.61 45.925 58.84 51.305 ;
      RECT 57.13 45.925 57.36 51.305 ;
      RECT 55.65 45.925 55.88 51.305 ;
      RECT 54.17 45.925 54.4 51.305 ;
      RECT 52.69 45.925 52.92 51.305 ;
      RECT 51.21 45.925 51.44 51.305 ;
      RECT 49.73 45.925 49.96 51.305 ;
      RECT 48.25 45.925 48.48 51.305 ;
      RECT 46.77 45.925 47 51.305 ;
      RECT 45.29 45.925 45.52 51.305 ;
      RECT 77.825 46.115 78.105 50.655 ;
      RECT 76.345 46.115 76.625 50.655 ;
      RECT 74.865 46.115 75.145 50.655 ;
      RECT 73.385 46.115 73.665 50.655 ;
      RECT 71.905 46.115 72.185 50.655 ;
      RECT 70.425 46.115 70.705 50.655 ;
      RECT 68.945 46.115 69.225 50.655 ;
      RECT 67.465 46.115 67.745 50.655 ;
      RECT 65.985 46.115 66.265 50.655 ;
      RECT 64.505 46.115 64.785 50.655 ;
      RECT 63.025 46.115 63.305 50.655 ;
      RECT 61.545 46.115 61.825 50.655 ;
      RECT 60.065 46.115 60.345 50.655 ;
      RECT 58.585 46.115 58.865 50.655 ;
      RECT 57.105 46.115 57.385 50.655 ;
      RECT 55.625 46.115 55.905 50.655 ;
      RECT 54.145 46.115 54.425 50.655 ;
      RECT 52.665 46.115 52.945 50.655 ;
      RECT 51.185 46.115 51.465 50.655 ;
      RECT 49.705 46.115 49.985 50.655 ;
      RECT 48.225 46.115 48.505 50.655 ;
      RECT 46.745 46.115 47.025 50.655 ;
      RECT 45.265 46.115 45.545 50.655 ;
      RECT 77.505 65.975 77.735 69.895 ;
      RECT 77.48 66.98 77.76 69.44 ;
      RECT 75.825 65.975 76.055 69.895 ;
      RECT 75.8 66.98 76.08 69.44 ;
      RECT 61.365 70.125 74.555 70.355 ;
      RECT 74.325 66.475 74.555 70.355 ;
      RECT 74.25 70.025 74.63 70.305 ;
      RECT 72.81 70.025 73.19 70.355 ;
      RECT 71.37 70.025 71.75 70.355 ;
      RECT 69.93 70.025 70.31 70.355 ;
      RECT 68.49 70.025 68.87 70.355 ;
      RECT 67.05 70.025 67.43 70.355 ;
      RECT 65.61 70.025 65.99 70.355 ;
      RECT 64.17 70.025 64.55 70.355 ;
      RECT 62.73 70.025 63.11 70.355 ;
      RECT 61.29 70.025 61.67 70.305 ;
      RECT 72.885 66.475 73.115 70.355 ;
      RECT 71.445 66.475 71.675 70.355 ;
      RECT 70.005 66.475 70.235 70.355 ;
      RECT 68.565 66.475 68.795 70.355 ;
      RECT 67.125 66.475 67.355 70.355 ;
      RECT 65.685 66.475 65.915 70.355 ;
      RECT 64.245 66.475 64.475 70.355 ;
      RECT 62.805 66.475 63.035 70.355 ;
      RECT 61.365 61.72 61.595 70.355 ;
      RECT 67.125 61.72 67.355 65.1 ;
      RECT 65.685 61.72 65.915 65.1 ;
      RECT 64.245 61.72 64.475 65.1 ;
      RECT 62.805 61.72 63.035 65.1 ;
      RECT 67.05 61.72 67.43 62 ;
      RECT 65.61 61.72 65.99 62 ;
      RECT 64.17 61.72 64.55 62 ;
      RECT 62.73 61.72 63.11 62 ;
      RECT 61.29 61.72 61.67 62 ;
      RECT 61.29 61.72 67.43 61.95 ;
      RECT 60.375 70.585 74.13 70.84 ;
      RECT 60.375 61.115 60.655 70.84 ;
      RECT 59.425 63.485 60.655 64.385 ;
      RECT 67.83 63.65 69.61 63.88 ;
      RECT 67.83 61.115 68.11 63.88 ;
      RECT 61.79 61.115 66.93 61.49 ;
      RECT 60.375 61.115 68.11 61.395 ;
      RECT 73.605 65.775 73.835 69.895 ;
      RECT 72.165 65.775 72.395 69.895 ;
      RECT 70.725 65.775 70.955 69.895 ;
      RECT 69.285 65.775 69.515 69.895 ;
      RECT 67.845 65.775 68.075 69.895 ;
      RECT 66.405 62.18 66.635 69.895 ;
      RECT 64.965 62.18 65.195 69.895 ;
      RECT 63.525 62.18 63.755 69.895 ;
      RECT 62.085 62.18 62.315 69.895 ;
      RECT 73.58 66.98 73.86 69.44 ;
      RECT 72.14 66.98 72.42 69.44 ;
      RECT 70.7 66.98 70.98 69.44 ;
      RECT 69.26 66.98 69.54 69.44 ;
      RECT 67.82 66.98 68.1 69.44 ;
      RECT 66.38 66.98 66.66 69.44 ;
      RECT 64.94 66.98 65.22 69.44 ;
      RECT 63.5 66.98 63.78 69.44 ;
      RECT 62.06 66.98 62.34 69.44 ;
      RECT 62.085 65.775 73.835 66.245 ;
      RECT 62.085 65.33 66.635 66.245 ;
      RECT 66.38 62.42 66.66 64.88 ;
      RECT 64.94 62.42 65.22 64.88 ;
      RECT 63.5 62.42 63.78 64.88 ;
      RECT 62.06 62.42 62.34 64.88 ;
      RECT 69.105 62.135 69.335 63.24 ;
      RECT 69.08 62.305 69.36 63.205 ;
      RECT 68.905 64.115 69.135 65.035 ;
      RECT 68.88 64.125 69.16 65.025 ;
      RECT 7.75 75.1 56.855 75.38 ;
      RECT 56.575 74.48 56.855 75.38 ;
      RECT 55.65 61.49 55.88 66.87 ;
      RECT 54.17 61.49 54.4 66.87 ;
      RECT 52.69 61.49 52.92 66.87 ;
      RECT 51.21 61.49 51.44 66.87 ;
      RECT 49.73 61.49 49.96 66.87 ;
      RECT 48.25 61.49 48.48 66.87 ;
      RECT 46.77 61.49 47 66.87 ;
      RECT 45.29 61.49 45.52 66.87 ;
      RECT 55.625 62.14 55.905 66.68 ;
      RECT 54.145 62.14 54.425 66.68 ;
      RECT 52.665 62.14 52.945 66.68 ;
      RECT 51.185 62.14 51.465 66.68 ;
      RECT 49.705 62.14 49.985 66.68 ;
      RECT 48.225 62.14 48.505 66.68 ;
      RECT 46.745 62.14 47.025 66.68 ;
      RECT 45.265 62.14 45.545 66.68 ;
      RECT 45.29 61.49 55.88 61.72 ;
      RECT 20.565 69.05 27.93 69.28 ;
      RECT 27.7 61.49 27.93 69.28 ;
      RECT 22.005 61.9 22.235 69.28 ;
      RECT 20.565 61.9 20.795 69.28 ;
      RECT 38.725 61.49 38.955 68.87 ;
      RECT 37.285 61.49 37.515 68.87 ;
      RECT 30.725 61.49 30.955 68.87 ;
      RECT 29.285 61.49 29.515 68.87 ;
      RECT 27.7 61.49 43.8 61.72 ;
      RECT 43.57 61.03 43.8 61.72 ;
      RECT 35.825 52.97 36.055 61.72 ;
      RECT 43.57 61.03 55.455 61.26 ;
      RECT 35.825 52.97 41.115 53.2 ;
      RECT 40.885 45.82 41.115 53.2 ;
      RECT 39.445 45.82 39.675 53.2 ;
      RECT 38.005 45.82 38.235 53.2 ;
      RECT 36.565 45.82 36.795 53.2 ;
      RECT 36.99 60.98 38.53 61.26 ;
      RECT 38.25 53.43 38.53 61.26 ;
      RECT 36.99 53.43 41.41 53.66 ;
      RECT 28.99 61.03 30.53 61.26 ;
      RECT 30.3 53.43 30.53 61.26 ;
      RECT 30.3 59.43 32.74 60.24 ;
      RECT 29.505 55.44 30.925 56.76 ;
      RECT 28.99 53.43 33.41 53.66 ;
      RECT 18.13 61.95 18.59 66.87 ;
      RECT 18.36 45.82 18.59 66.87 ;
      RECT 18.36 60.98 22.53 61.21 ;
      RECT 18.36 53.43 25.41 53.66 ;
      RECT 18.13 45.82 18.59 52.74 ;
      RECT 17.1 61.31 17.935 61.65 ;
      RECT 17.1 53.04 17.38 61.65 ;
      RECT 15.61 59.6 17.38 60.41 ;
      RECT 17.095 57.58 17.38 58.48 ;
      RECT 7.77 53.38 10.75 54.7 ;
      RECT 7.77 53.605 17.38 54.415 ;
      RECT 17.1 53.04 17.935 53.38 ;
      RECT 5.135 4.5 95.14 7.49 ;
      RECT 13.14 24.385 87.14 26.385 ;
      RECT 79.865 76.375 85.24 77.785 ;
      RECT 16.14 16.215 84.14 18.215 ;
      RECT 78.37 54.215 81.055 59.495 ;
      RECT 24.275 80.77 76.155 82.775 ;
      RECT 24.275 85.205 76.155 87.21 ;
      RECT 45.91 54.215 46.2 59.495 ;
      RECT 10.195 37.46 36.075 40.54 ;
      RECT 14.35 76.375 14.58 79.445 ;
    LAYER M2 SPACING 0.28 ;
      RECT 56.395 98.41 56.715 99.64 ;
      RECT 43.715 98.41 44.035 99.64 ;
    LAYER M2 ;
      RECT 84.56 65.115 87.56 116.58 ;
      RECT 81.47 65.115 87.56 66.015 ;
      RECT 68.88 62.375 69.16 65.025 ;
      RECT 70.76 62.33 77.76 64.79 ;
      RECT 70.76 62.33 79.315 63.255 ;
      RECT 69.08 62.305 69.36 63.205 ;
      RECT 68.88 62.375 79.315 63.175 ;
      RECT 60.375 70.025 74.63 71.585 ;
      RECT 60.375 70.025 79.15 70.305 ;
      RECT 78.35 67.615 79.15 70.305 ;
      RECT 60.375 61.695 61.67 71.585 ;
      RECT 67.05 61.695 67.43 62 ;
      RECT 65.61 61.695 65.99 62 ;
      RECT 64.17 61.695 64.55 62 ;
      RECT 62.73 61.695 63.11 62 ;
      RECT 60.375 61.695 67.43 61.975 ;
      RECT 44.455 16.215 55.975 82.78 ;
      RECT 44.455 45.885 78.915 50.885 ;
      RECT 38.03 16.215 62.03 39.91 ;
      RECT 62.06 66.72 77.76 69.7 ;
      RECT 62.06 62.42 66.66 69.7 ;
      RECT 57.77 72.415 58.85 73.605 ;
      RECT 57.77 72.535 64.46 73.435 ;
      RECT 56.575 63.795 56.855 75.38 ;
      RECT 59.425 63.485 59.705 64.385 ;
      RECT 56.575 63.795 59.705 64.075 ;
      RECT 38.2 57.63 38.58 58.43 ;
      RECT 17.045 57.63 17.425 58.43 ;
      RECT 17.045 57.63 38.58 57.91 ;
      RECT 12.14 9.56 36.14 44.285 ;
      RECT 10.195 37.46 36.14 40.54 ;
      RECT 12.955 55.445 15.955 116.58 ;
      RECT 14.185 55.44 30.925 56.76 ;
      RECT 5.28 4.505 95 7.485 ;
      RECT 64.14 14.34 88.14 39.91 ;
      RECT 58.785 43.365 84.545 44.265 ;
      RECT 79.865 54.215 81.055 77.785 ;
      RECT 72.89 78.115 78.865 79.525 ;
      RECT 68.015 72.365 77.135 74.825 ;
      RECT 56.715 98.41 65.585 99.64 ;
      RECT 34.815 98.41 43.715 99.64 ;
      RECT 19.15 69.675 42.31 70.575 ;
      RECT 7.75 53.33 10.75 116.58 ;
    LAYER M3 ;
      RECT 33.165 98.41 67.235 99.64 ;
    LAYER M4 ;
      RECT 33.165 98.41 67.235 99.64 ;
    LAYER M5 ;
      RECT 4 4 96 96 ;
      RECT 33.165 98.41 67.235 99.64 ;
  END
END Pulldown_pol_IO_lowcap_EN

END LIBRARY
