//Verilog HDL for "pALPIDEfs_V2_BLOCKS_CAM", "PAD_DVSS" "functional"
`timescale 1ns / 1ps

module PAD_DVSS ( AVDD, AVSS/*, DVDD, DVSS, SUB*/ );

//  inout DVDD;
  inout AVSS;
//  inout SUB;
//  inout DVSS;
  inout AVDD;
  
endmodule
