VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO MONOPIX_TOP
  CLASS BLOCK ;
  ORIGIN -998.1 -1046.435 ;
  FOREIGN MONOPIX_TOP 998.1 1046.435 ;
  SIZE 18163.8 BY 8953.565 ;
  SYMMETRY X Y R90 ;
  PIN INJ_ROW[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8948.585 1046.435 8948.865 1047.435 ;
    END
  END INJ_ROW[97]
  PIN Data_PMOS[869]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8946.905 1046.435 8947.185 1047.435 ;
    END
  END Data_PMOS[869]
  PIN Data_PMOS[866]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8945.225 1046.435 8945.505 1047.435 ;
    END
  END Data_PMOS[866]
  PIN Data_PMOS[875]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8943.545 1046.435 8943.825 1047.435 ;
    END
  END Data_PMOS[875]
  PIN INJ_IN[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8941.305 1046.435 8941.585 1047.435 ;
    END
  END INJ_IN[195]
  PIN BcidMtx[585]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8924.505 1046.435 8924.785 1047.435 ;
    END
  END BcidMtx[585]
  PIN Read_PMOS[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8923.385 1046.435 8923.665 1047.435 ;
    END
  END Read_PMOS[41]
  PIN BcidMtx[582]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8921.705 1046.435 8921.985 1047.435 ;
    END
  END BcidMtx[582]
  PIN Data_PMOS[870]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8918.345 1046.435 8918.625 1047.435 ;
    END
  END Data_PMOS[870]
  PIN Data_PMOS[871]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8917.225 1046.435 8917.505 1047.435 ;
    END
  END Data_PMOS[871]
  PIN Data_PMOS[872]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8915.545 1046.435 8915.825 1047.435 ;
    END
  END Data_PMOS[872]
  PIN Data_PMOS[878]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8913.865 1046.435 8914.145 1047.435 ;
    END
  END Data_PMOS[878]
  PIN MASKD[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8873.545 1046.435 8873.825 1047.435 ;
    END
  END MASKD[194]
  PIN DIG_MON_SEL[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8870.745 1046.435 8871.025 1047.435 ;
    END
  END DIG_MON_SEL[194]
  PIN DIG_MON_PMOS[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8867.945 1046.435 8868.225 1047.435 ;
    END
  END DIG_MON_PMOS[81]
  PIN Data_PMOS[858]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8865.705 1046.435 8865.985 1047.435 ;
    END
  END Data_PMOS[858]
  PIN Data_PMOS[859]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8864.025 1046.435 8864.305 1047.435 ;
    END
  END Data_PMOS[859]
  PIN Data_PMOS[854]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8861.785 1046.435 8862.065 1047.435 ;
    END
  END Data_PMOS[854]
  PIN Data_PMOS[846]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8852.265 1046.435 8852.545 1047.435 ;
    END
  END Data_PMOS[846]
  PIN Data_HV[1068]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18641.345 1046.435 18641.625 1047.435 ;
    END
  END Data_HV[1068]
  PIN BcidMtx[579]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8847.785 1046.435 8848.065 1047.435 ;
    END
  END BcidMtx[579]
  PIN BcidMtx[578]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8846.105 1046.435 8846.385 1047.435 ;
    END
  END BcidMtx[578]
  PIN INJ_IN[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8841.905 1046.435 8842.185 1047.435 ;
    END
  END INJ_IN[192]
  PIN Data_PMOS[849]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8839.665 1046.435 8839.945 1047.435 ;
    END
  END Data_PMOS[849]
  PIN Data_PMOS[844]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8812.505 1046.435 8812.785 1047.435 ;
    END
  END Data_PMOS[844]
  PIN Data_PMOS[841]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8810.825 1046.435 8811.105 1047.435 ;
    END
  END Data_PMOS[841]
  PIN MASKV[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8809.145 1046.435 8809.425 1047.435 ;
    END
  END MASKV[192]
  PIN DIG_MON_PMOS[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8806.905 1046.435 8807.185 1047.435 ;
    END
  END DIG_MON_PMOS[80]
  PIN DIG_MON_SEL[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8804.665 1046.435 8804.945 1047.435 ;
    END
  END DIG_MON_SEL[191]
  PIN MASKV[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8800.745 1046.435 8801.025 1047.435 ;
    END
  END MASKV[191]
  PIN Data_PMOS[827]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8799.625 1046.435 8799.905 1047.435 ;
    END
  END Data_PMOS[827]
  PIN Data_PMOS[824]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8785.065 1046.435 8785.345 1047.435 ;
    END
  END Data_PMOS[824]
  PIN Data_PMOS[826]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8782.825 1046.435 8783.105 1047.435 ;
    END
  END Data_PMOS[826]
  PIN INJ_IN[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8781.145 1046.435 8781.425 1047.435 ;
    END
  END INJ_IN[191]
  PIN BcidMtx[574]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8778.345 1046.435 8778.625 1047.435 ;
    END
  END BcidMtx[574]
  PIN Read_PMOS[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8776.665 1046.435 8776.945 1047.435 ;
    END
  END Read_PMOS[39]
  PIN BcidMtx[570]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8774.985 1046.435 8775.265 1047.435 ;
    END
  END BcidMtx[570]
  PIN Data_PMOS[821]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8733.545 1046.435 8733.825 1047.435 ;
    END
  END Data_PMOS[821]
  PIN Data_PMOS[829]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8731.865 1046.435 8732.145 1047.435 ;
    END
  END Data_PMOS[829]
  PIN Data_PMOS[830]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8730.185 1046.435 8730.465 1047.435 ;
    END
  END Data_PMOS[830]
  PIN Data_PMOS[836]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8728.505 1046.435 8728.785 1047.435 ;
    END
  END Data_PMOS[836]
  PIN MASKD[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8726.825 1046.435 8727.105 1047.435 ;
    END
  END MASKD[190]
  PIN DIG_MON_SEL[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8724.025 1046.435 8724.305 1047.435 ;
    END
  END DIG_MON_SEL[190]
  PIN DIG_MON_PMOS[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8721.225 1046.435 8721.505 1047.435 ;
    END
  END DIG_MON_PMOS[77]
  PIN Data_PMOS[816]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8710.585 1046.435 8710.865 1047.435 ;
    END
  END Data_PMOS[816]
  PIN Data_PMOS[817]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8708.905 1046.435 8709.185 1047.435 ;
    END
  END Data_PMOS[817]
  PIN Data_PMOS[818]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8707.225 1046.435 8707.505 1047.435 ;
    END
  END Data_PMOS[818]
  PIN Data_PMOS[804]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8705.545 1046.435 8705.825 1047.435 ;
    END
  END Data_PMOS[804]
  PIN BcidMtx[569]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8700.225 1046.435 8700.505 1047.435 ;
    END
  END BcidMtx[569]
  PIN Read_PMOS[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8672.505 1046.435 8672.785 1047.435 ;
    END
  END Read_PMOS[38]
  PIN INJ_IN[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8669.705 1046.435 8669.985 1047.435 ;
    END
  END INJ_IN[188]
  PIN Data_PMOS[800]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8668.025 1046.435 8668.305 1047.435 ;
    END
  END Data_PMOS[800]
  PIN Data_PMOS[808]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8666.345 1046.435 8666.625 1047.435 ;
    END
  END Data_PMOS[808]
  PIN Data_PMOS[814]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8665.225 1046.435 8665.505 1047.435 ;
    END
  END Data_PMOS[814]
  PIN Data_PMOS[798]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8663.545 1046.435 8663.825 1047.435 ;
    END
  END Data_PMOS[798]
  PIN MASKV[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8662.425 1046.435 8662.705 1047.435 ;
    END
  END MASKV[188]
  PIN MASKD[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8643.945 1046.435 8644.225 1047.435 ;
    END
  END MASKD[187]
  PIN INJ_ROW[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8641.705 1046.435 8641.985 1047.435 ;
    END
  END INJ_ROW[93]
  PIN MASKV[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18641.905 1046.435 18642.185 1047.435 ;
    END
  END MASKV[437]
  PIN Data_PMOS[789]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8639.465 1046.435 8639.745 1047.435 ;
    END
  END Data_PMOS[789]
  PIN Data_PMOS[790]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8637.785 1046.435 8638.065 1047.435 ;
    END
  END Data_PMOS[790]
  PIN Data_PMOS[784]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8636.105 1046.435 8636.385 1047.435 ;
    END
  END Data_PMOS[784]
  PIN INJ_IN[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8634.425 1046.435 8634.705 1047.435 ;
    END
  END INJ_IN[187]
  PIN BcidMtx[561]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8591.865 1046.435 8592.145 1047.435 ;
    END
  END BcidMtx[561]
  PIN BcidMtx[560]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8590.185 1046.435 8590.465 1047.435 ;
    END
  END BcidMtx[560]
  PIN BcidMtx[558]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8589.065 1046.435 8589.345 1047.435 ;
    END
  END BcidMtx[558]
  PIN Data_PMOS[779]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8586.265 1046.435 8586.545 1047.435 ;
    END
  END Data_PMOS[779]
  PIN Data_PMOS[792]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8585.145 1046.435 8585.425 1047.435 ;
    END
  END Data_PMOS[792]
  PIN Data_PMOS[788]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8582.905 1046.435 8583.185 1047.435 ;
    END
  END Data_PMOS[788]
  PIN Data_PMOS[777]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8581.785 1046.435 8582.065 1047.435 ;
    END
  END Data_PMOS[777]
  PIN MASKH[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8571.705 1046.435 8571.985 1047.435 ;
    END
  END MASKH[93]
  PIN DIG_MON_SEL[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8567.785 1046.435 8568.065 1047.435 ;
    END
  END DIG_MON_SEL[185]
  PIN DIG_MON_PMOS[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8565.545 1046.435 8565.825 1047.435 ;
    END
  END DIG_MON_PMOS[73]
  PIN Data_PMOS[774]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8561.345 1046.435 8561.625 1047.435 ;
    END
  END Data_PMOS[774]
  PIN Data_PMOS[761]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8559.105 1046.435 8559.385 1047.435 ;
    END
  END Data_PMOS[761]
  PIN Data_PMOS[776]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8532.505 1046.435 8532.785 1047.435 ;
    END
  END Data_PMOS[776]
  PIN Data_PMOS[763]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8531.385 1046.435 8531.665 1047.435 ;
    END
  END Data_PMOS[763]
  PIN BcidMtx[557]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8527.465 1046.435 8527.745 1047.435 ;
    END
  END BcidMtx[557]
  PIN FREEZE_PMOS[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8525.785 1046.435 8526.065 1047.435 ;
    END
  END FREEZE_PMOS[36]
  PIN BcidMtx[554]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8524.665 1046.435 8524.945 1047.435 ;
    END
  END BcidMtx[554]
  PIN INJ_IN[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8522.425 1046.435 8522.705 1047.435 ;
    END
  END INJ_IN[184]
  PIN Data_PMOS[765]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8520.185 1046.435 8520.465 1047.435 ;
    END
  END Data_PMOS[765]
  PIN Data_PMOS[760]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8505.625 1046.435 8505.905 1047.435 ;
    END
  END Data_PMOS[760]
  PIN Data_PMOS[757]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8503.945 1046.435 8504.225 1047.435 ;
    END
  END Data_PMOS[757]
  PIN Data_PMOS[773]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8502.825 1046.435 8503.105 1047.435 ;
    END
  END Data_PMOS[773]
  PIN MASKH[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8501.705 1046.435 8501.985 1047.435 ;
    END
  END MASKH[92]
  PIN DIG_MON_SEL[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8497.785 1046.435 8498.065 1047.435 ;
    END
  END DIG_MON_SEL[183]
  PIN DIG_MON_PMOS[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8495.545 1046.435 8495.825 1047.435 ;
    END
  END DIG_MON_PMOS[71]
  PIN Data_PMOS[743]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8452.985 1046.435 8453.265 1047.435 ;
    END
  END Data_PMOS[743]
  PIN Data_PMOS[740]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8451.305 1046.435 8451.585 1047.435 ;
    END
  END Data_PMOS[740]
  PIN Data_PMOS[755]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8450.185 1046.435 8450.465 1047.435 ;
    END
  END Data_PMOS[755]
  PIN Data_HV[1060]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18586.185 1046.435 18586.465 1047.435 ;
    END
  END Data_HV[1060]
  PIN nTOK_PMOS[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8446.265 1046.435 8446.545 1047.435 ;
    END
  END nTOK_PMOS[35]
  PIN BcidMtx[550]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8444.585 1046.435 8444.865 1047.435 ;
    END
  END BcidMtx[550]
  PIN Read_PMOS[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8442.905 1046.435 8443.185 1047.435 ;
    END
  END Read_PMOS[35]
  PIN INJ_IN[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8431.705 1046.435 8431.985 1047.435 ;
    END
  END INJ_IN[182]
  PIN Data_PMOS[737]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8430.025 1046.435 8430.305 1047.435 ;
    END
  END Data_PMOS[737]
  PIN Data_PMOS[739]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8427.785 1046.435 8428.065 1047.435 ;
    END
  END Data_PMOS[739]
  PIN Data_PMOS[736]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8426.105 1046.435 8426.385 1047.435 ;
    END
  END Data_PMOS[736]
  PIN Data_PMOS[752]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8424.985 1046.435 8425.265 1047.435 ;
    END
  END Data_PMOS[752]
  PIN MASKD[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12341.345 1046.435 12341.625 1047.435 ;
    END
  END MASKD[280]
  PIN DIG_MON_SEL[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12338.545 1046.435 12338.825 1047.435 ;
    END
  END DIG_MON_SEL[280]
  PIN MASKD[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13430.825 1046.435 13431.105 1047.435 ;
    END
  END MASKD[307]
  PIN MASKV[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13428.025 1046.435 13428.305 1047.435 ;
    END
  END MASKV[307]
  PIN Data_COMP[873]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13426.345 1046.435 13426.625 1047.435 ;
    END
  END Data_COMP[873]
  PIN Data_COMP[874]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13424.665 1046.435 13424.945 1047.435 ;
    END
  END Data_COMP[874]
  PIN Data_COMP[868]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13422.985 1046.435 13423.265 1047.435 ;
    END
  END Data_COMP[868]
  PIN INJ_IN[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13421.305 1046.435 13421.585 1047.435 ;
    END
  END INJ_IN[307]
  PIN BcidMtx[922]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13405.065 1046.435 13405.345 1047.435 ;
    END
  END BcidMtx[922]
  PIN Read_COMP[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13403.385 1046.435 13403.665 1047.435 ;
    END
  END Read_COMP[41]
  PIN BcidMtx[918]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13401.705 1046.435 13401.985 1047.435 ;
    END
  END BcidMtx[918]
  PIN Data_COMP[863]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13398.905 1046.435 13399.185 1047.435 ;
    END
  END Data_COMP[863]
  PIN Data_COMP[871]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13397.225 1046.435 13397.505 1047.435 ;
    END
  END Data_COMP[871]
  PIN Data_COMP[872]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13395.545 1046.435 13395.825 1047.435 ;
    END
  END Data_COMP[872]
  PIN Data_COMP[878]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13393.865 1046.435 13394.145 1047.435 ;
    END
  END Data_COMP[878]
  PIN MASKD[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13353.545 1046.435 13353.825 1047.435 ;
    END
  END MASKD[306]
  PIN DIG_MON_SEL[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13350.745 1046.435 13351.025 1047.435 ;
    END
  END DIG_MON_SEL[306]
  PIN DIG_MON_COMP[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13347.945 1046.435 13348.225 1047.435 ;
    END
  END DIG_MON_COMP[81]
  PIN Data_COMP[858]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13345.705 1046.435 13345.985 1047.435 ;
    END
  END Data_COMP[858]
  PIN Data_COMP[859]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13344.025 1046.435 13344.305 1047.435 ;
    END
  END Data_COMP[859]
  PIN Data_COMP[860]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13342.345 1046.435 13342.625 1047.435 ;
    END
  END Data_COMP[860]
  PIN Data_COMP[846]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13332.265 1046.435 13332.545 1047.435 ;
    END
  END Data_COMP[846]
  PIN BcidMtx[917]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13328.905 1046.435 13329.185 1047.435 ;
    END
  END BcidMtx[917]
  PIN FREEZE_COMP[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13327.225 1046.435 13327.505 1047.435 ;
    END
  END FREEZE_COMP[40]
  PIN BcidMtx[913]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13325.545 1046.435 13325.825 1047.435 ;
    END
  END BcidMtx[913]
  PIN Data_COMP[843]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13320.785 1046.435 13321.065 1047.435 ;
    END
  END Data_COMP[843]
  PIN Data_COMP[855]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13319.105 1046.435 13319.385 1047.435 ;
    END
  END Data_COMP[855]
  PIN Data_COMP[856]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13291.945 1046.435 13292.225 1047.435 ;
    END
  END Data_COMP[856]
  PIN Data_COMP[840]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13290.265 1046.435 13290.545 1047.435 ;
    END
  END Data_COMP[840]
  PIN MASKV[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13289.145 1046.435 13289.425 1047.435 ;
    END
  END MASKV[304]
  PIN MASKD[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13283.545 1046.435 13283.825 1047.435 ;
    END
  END MASKD[303]
  PIN MASKV[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13280.745 1046.435 13281.025 1047.435 ;
    END
  END MASKV[303]
  PIN Data_COMP[831]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13266.185 1046.435 13266.465 1047.435 ;
    END
  END Data_COMP[831]
  PIN Data_COMP[832]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13264.505 1046.435 13264.785 1047.435 ;
    END
  END Data_COMP[832]
  PIN Data_COMP[826]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13262.825 1046.435 13263.105 1047.435 ;
    END
  END Data_COMP[826]
  PIN nTOK_COMP[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13260.025 1046.435 13260.305 1047.435 ;
    END
  END nTOK_COMP[39]
  PIN BcidMtx[909]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13257.785 1046.435 13258.065 1047.435 ;
    END
  END BcidMtx[909]
  PIN BcidMtx[908]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13256.105 1046.435 13256.385 1047.435 ;
    END
  END BcidMtx[908]
  PIN INJ_IN[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13253.865 1046.435 13254.145 1047.435 ;
    END
  END INJ_IN[302]
  PIN Data_COMP[828]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13212.985 1046.435 13213.265 1047.435 ;
    END
  END Data_COMP[828]
  PIN Data_COMP[823]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13211.305 1046.435 13211.585 1047.435 ;
    END
  END Data_COMP[823]
  PIN Data_COMP[820]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13209.625 1046.435 13209.905 1047.435 ;
    END
  END Data_COMP[820]
  PIN MASKV[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13207.945 1046.435 13208.225 1047.435 ;
    END
  END MASKV[302]
  PIN DIG_MON_COMP[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13205.705 1046.435 13205.985 1047.435 ;
    END
  END DIG_MON_COMP[78]
  PIN DIG_MON_SEL[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13203.465 1046.435 13203.745 1047.435 ;
    END
  END DIG_MON_SEL[301]
  PIN MASKD[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13202.345 1046.435 13202.625 1047.435 ;
    END
  END MASKD[301]
  PIN MASKV[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13191.145 1046.435 13191.425 1047.435 ;
    END
  END MASKV[301]
  PIN Data_COMP[810]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13189.465 1046.435 13189.745 1047.435 ;
    END
  END Data_COMP[810]
  PIN Data_COMP[811]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13187.785 1046.435 13188.065 1047.435 ;
    END
  END Data_COMP[811]
  PIN Data_COMP[805]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13186.105 1046.435 13186.385 1047.435 ;
    END
  END Data_COMP[805]
  PIN nTOK_COMP[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13181.345 1046.435 13181.625 1047.435 ;
    END
  END nTOK_COMP[38]
  PIN BcidMtx[903]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13179.105 1046.435 13179.385 1047.435 ;
    END
  END BcidMtx[903]
  PIN BcidMtx[901]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13151.385 1046.435 13151.665 1047.435 ;
    END
  END BcidMtx[901]
  PIN Data_COMP[801]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13148.585 1046.435 13148.865 1047.435 ;
    END
  END Data_COMP[801]
  PIN Data_COMP[813]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13146.905 1046.435 13147.185 1047.435 ;
    END
  END Data_COMP[813]
  PIN Data_COMP[814]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13145.225 1046.435 13145.505 1047.435 ;
    END
  END Data_COMP[814]
  PIN Data_COMP[798]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13143.545 1046.435 13143.825 1047.435 ;
    END
  END Data_COMP[798]
  PIN MASKH[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13141.865 1046.435 13142.145 1047.435 ;
    END
  END MASKH[150]
  PIN MASKD[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13123.945 1046.435 13124.225 1047.435 ;
    END
  END MASKD[299]
  PIN INJ_ROW[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13121.705 1046.435 13121.985 1047.435 ;
    END
  END INJ_ROW[149]
  PIN nTOK_HV[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18608.585 1046.435 18608.865 1047.435 ;
    END
  END nTOK_HV[50]
  PIN Data_COMP[789]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13119.465 1046.435 13119.745 1047.435 ;
    END
  END Data_COMP[789]
  PIN Data_COMP[790]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13117.785 1046.435 13118.065 1047.435 ;
    END
  END Data_COMP[790]
  PIN Data_COMP[784]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13116.105 1046.435 13116.385 1047.435 ;
    END
  END Data_COMP[784]
  PIN nTOK_COMP[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13074.105 1046.435 13074.385 1047.435 ;
    END
  END nTOK_COMP[37]
  PIN BcidMtx[897]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13071.865 1046.435 13072.145 1047.435 ;
    END
  END BcidMtx[897]
  PIN BcidMtx[896]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13070.185 1046.435 13070.465 1047.435 ;
    END
  END BcidMtx[896]
  PIN INJ_IN[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13067.945 1046.435 13068.225 1047.435 ;
    END
  END INJ_IN[298]
  PIN Data_COMP[786]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13065.705 1046.435 13065.985 1047.435 ;
    END
  END Data_COMP[786]
  PIN Data_COMP[781]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13064.025 1046.435 13064.305 1047.435 ;
    END
  END Data_COMP[781]
  PIN Data_COMP[778]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13062.345 1046.435 13062.625 1047.435 ;
    END
  END Data_COMP[778]
  PIN MASKV[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13052.265 1046.435 13052.545 1047.435 ;
    END
  END MASKV[298]
  PIN DIG_MON_COMP[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13050.025 1046.435 13050.305 1047.435 ;
    END
  END DIG_MON_COMP[74]
  PIN MASKD[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13046.665 1046.435 13046.945 1047.435 ;
    END
  END MASKD[297]
  PIN Data_HV[1096]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18745.785 1046.435 18746.065 1047.435 ;
    END
  END Data_HV[1096]
  PIN MASKV[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13041.905 1046.435 13042.185 1047.435 ;
    END
  END MASKV[297]
  PIN Data_COMP[775]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13039.665 1046.435 13039.945 1047.435 ;
    END
  END Data_COMP[775]
  PIN Data_COMP[761]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13039.105 1046.435 13039.385 1047.435 ;
    END
  END Data_COMP[761]
  PIN Data_COMP[770]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13011.945 1046.435 13012.225 1047.435 ;
    END
  END Data_COMP[770]
  PIN INJ_IN[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13009.705 1046.435 13009.985 1047.435 ;
    END
  END INJ_IN[297]
  PIN BcidMtx[892]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13006.905 1046.435 13007.185 1047.435 ;
    END
  END BcidMtx[892]
  PIN Read_COMP[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13005.225 1046.435 13005.505 1047.435 ;
    END
  END Read_COMP[36]
  PIN BcidMtx[888]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13003.545 1046.435 13003.825 1047.435 ;
    END
  END BcidMtx[888]
  PIN Data_COMP[758]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13000.745 1046.435 13001.025 1047.435 ;
    END
  END Data_COMP[758]
  PIN Data_COMP[766]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12986.185 1046.435 12986.465 1047.435 ;
    END
  END Data_COMP[766]
  PIN Data_COMP[767]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12984.505 1046.435 12984.785 1047.435 ;
    END
  END Data_COMP[767]
  PIN Data_COMP[773]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12982.825 1046.435 12983.105 1047.435 ;
    END
  END Data_COMP[773]
  PIN MASKD[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12981.145 1046.435 12981.425 1047.435 ;
    END
  END MASKD[296]
  PIN DIG_MON_SEL[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12978.345 1046.435 12978.625 1047.435 ;
    END
  END DIG_MON_SEL[296]
  PIN DIG_MON_COMP[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12975.545 1046.435 12975.825 1047.435 ;
    END
  END DIG_MON_COMP[71]
  PIN Data_COMP[753]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12933.545 1046.435 12933.825 1047.435 ;
    END
  END Data_COMP[753]
  PIN Data_COMP[754]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12931.865 1046.435 12932.145 1047.435 ;
    END
  END Data_COMP[754]
  PIN Data_COMP[755]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12930.185 1046.435 12930.465 1047.435 ;
    END
  END Data_COMP[755]
  PIN Data_COMP[741]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12928.505 1046.435 12928.785 1047.435 ;
    END
  END Data_COMP[741]
  PIN BcidMtx[887]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12925.145 1046.435 12925.425 1047.435 ;
    END
  END BcidMtx[887]
  PIN FREEZE_COMP[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12923.465 1046.435 12923.745 1047.435 ;
    END
  END FREEZE_COMP[35]
  PIN BcidMtx[883]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12921.785 1046.435 12922.065 1047.435 ;
    END
  END BcidMtx[883]
  PIN Data_COMP[738]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12910.585 1046.435 12910.865 1047.435 ;
    END
  END Data_COMP[738]
  PIN Data_COMP[750]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12908.905 1046.435 12909.185 1047.435 ;
    END
  END Data_COMP[750]
  PIN Data_COMP[751]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12907.225 1046.435 12907.505 1047.435 ;
    END
  END Data_COMP[751]
  PIN Data_COMP[458]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11784.985 1046.435 11785.265 1047.435 ;
    END
  END Data_COMP[458]
  PIN DIG_MON_SEL[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12871.945 1046.435 12872.225 1047.435 ;
    END
  END DIG_MON_SEL[293]
  PIN DIG_MON_COMP[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12869.705 1046.435 12869.985 1047.435 ;
    END
  END DIG_MON_COMP[69]
  PIN Data_COMP[722]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12866.905 1046.435 12867.185 1047.435 ;
    END
  END Data_COMP[722]
  PIN Data_COMP[719]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12865.225 1046.435 12865.505 1047.435 ;
    END
  END Data_COMP[719]
  PIN Data_COMP[734]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12864.105 1046.435 12864.385 1047.435 ;
    END
  END Data_COMP[734]
  PIN INJ_IN[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12861.305 1046.435 12861.585 1047.435 ;
    END
  END INJ_IN[293]
  PIN BcidMtx[880]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12845.065 1046.435 12845.345 1047.435 ;
    END
  END BcidMtx[880]
  PIN BcidMtx[879]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12844.505 1046.435 12844.785 1047.435 ;
    END
  END BcidMtx[879]
  PIN BcidMtx[878]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12842.825 1046.435 12843.105 1047.435 ;
    END
  END BcidMtx[878]
  PIN Data_COMP[717]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12839.465 1046.435 12839.745 1047.435 ;
    END
  END Data_COMP[717]
  PIN Data_COMP[723]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12838.345 1046.435 12838.625 1047.435 ;
    END
  END Data_COMP[723]
  PIN Data_COMP[718]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12836.665 1046.435 12836.945 1047.435 ;
    END
  END Data_COMP[718]
  PIN Data_COMP[714]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12834.425 1046.435 12834.705 1047.435 ;
    END
  END Data_COMP[714]
  PIN MASKV[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12794.665 1046.435 12794.945 1047.435 ;
    END
  END MASKV[292]
  PIN DIG_MON_COMP[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12792.425 1046.435 12792.705 1047.435 ;
    END
  END DIG_MON_COMP[68]
  PIN DIG_MON_COMP[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12787.945 1046.435 12788.225 1047.435 ;
    END
  END DIG_MON_COMP[67]
  PIN MASKV[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12786.265 1046.435 12786.545 1047.435 ;
    END
  END MASKV[291]
  PIN Data_COMP[701]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12785.145 1046.435 12785.425 1047.435 ;
    END
  END Data_COMP[701]
  PIN Data_COMP[713]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12782.345 1046.435 12782.625 1047.435 ;
    END
  END Data_COMP[713]
  PIN Data_COMP[707]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12781.785 1046.435 12782.065 1047.435 ;
    END
  END Data_COMP[707]
  PIN INJ_IN[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12771.145 1046.435 12771.425 1047.435 ;
    END
  END INJ_IN[291]
  PIN FREEZE_COMP[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12767.225 1046.435 12767.505 1047.435 ;
    END
  END FREEZE_COMP[33]
  PIN BcidMtx[872]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12766.105 1046.435 12766.385 1047.435 ;
    END
  END BcidMtx[872]
  PIN BcidMtx[870]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12764.985 1046.435 12765.265 1047.435 ;
    END
  END BcidMtx[870]
  PIN Data_COMP[695]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12760.225 1046.435 12760.505 1047.435 ;
    END
  END Data_COMP[695]
  PIN Data_COMP[697]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12732.505 1046.435 12732.785 1047.435 ;
    END
  END Data_COMP[697]
  PIN Data_COMP[693]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12730.265 1046.435 12730.545 1047.435 ;
    END
  END Data_COMP[693]
  PIN MASKH[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12728.585 1046.435 12728.865 1047.435 ;
    END
  END MASKH[145]
  PIN MASKD[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12723.545 1046.435 12723.825 1047.435 ;
    END
  END MASKD[289]
  PIN MASKV[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12720.745 1046.435 12721.025 1047.435 ;
    END
  END MASKV[289]
  PIN Data_COMP[684]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12706.185 1046.435 12706.465 1047.435 ;
    END
  END Data_COMP[684]
  PIN Data_COMP[685]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12704.505 1046.435 12704.785 1047.435 ;
    END
  END Data_COMP[685]
  PIN Data_COMP[679]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12702.825 1046.435 12703.105 1047.435 ;
    END
  END Data_COMP[679]
  PIN nTOK_COMP[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12700.025 1046.435 12700.305 1047.435 ;
    END
  END nTOK_COMP[32]
  PIN BcidMtx[867]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12697.785 1046.435 12698.065 1047.435 ;
    END
  END BcidMtx[867]
  PIN BcidMtx[866]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12696.105 1046.435 12696.385 1047.435 ;
    END
  END BcidMtx[866]
  PIN BcidMtx[865]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12695.545 1046.435 12695.825 1047.435 ;
    END
  END BcidMtx[865]
  PIN Data_COMP[681]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12652.985 1046.435 12653.265 1047.435 ;
    END
  END Data_COMP[681]
  PIN Data_COMP[676]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12651.305 1046.435 12651.585 1047.435 ;
    END
  END Data_COMP[676]
  PIN Data_COMP[673]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12649.625 1046.435 12649.905 1047.435 ;
    END
  END Data_COMP[673]
  PIN MASKV[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12647.945 1046.435 12648.225 1047.435 ;
    END
  END MASKV[288]
  PIN DIG_MON_COMP[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12645.705 1046.435 12645.985 1047.435 ;
    END
  END DIG_MON_COMP[64]
  PIN DIG_MON_SEL[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12643.465 1046.435 12643.745 1047.435 ;
    END
  END DIG_MON_SEL[287]
  PIN INJ_ROW[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12631.705 1046.435 12631.985 1047.435 ;
    END
  END INJ_ROW[143]
  PIN BcidMtx[1322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18751.945 1046.435 18752.225 1047.435 ;
    END
  END BcidMtx[1322]
  PIN Data_COMP[670]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12628.905 1046.435 12629.185 1047.435 ;
    END
  END Data_COMP[670]
  PIN Data_COMP[671]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12627.225 1046.435 12627.505 1047.435 ;
    END
  END Data_COMP[671]
  PIN Data_COMP[657]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12625.545 1046.435 12625.825 1047.435 ;
    END
  END Data_COMP[657]
  PIN BcidMtx[863]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12620.225 1046.435 12620.505 1047.435 ;
    END
  END BcidMtx[863]
  PIN Read_COMP[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12592.505 1046.435 12592.785 1047.435 ;
    END
  END Read_COMP[31]
  PIN BcidMtx[858]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12590.825 1046.435 12591.105 1047.435 ;
    END
  END BcidMtx[858]
  PIN Data_COMP[653]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12588.025 1046.435 12588.305 1047.435 ;
    END
  END Data_COMP[653]
  PIN Data_COMP[661]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12586.345 1046.435 12586.625 1047.435 ;
    END
  END Data_COMP[661]
  PIN Data_COMP[662]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12584.665 1046.435 12584.945 1047.435 ;
    END
  END Data_COMP[662]
  PIN Data_COMP[668]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12582.985 1046.435 12583.265 1047.435 ;
    END
  END Data_COMP[668]
  PIN MASKD[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12581.305 1046.435 12581.585 1047.435 ;
    END
  END MASKD[286]
  PIN DIG_MON_SEL[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12565.625 1046.435 12565.905 1047.435 ;
    END
  END DIG_MON_SEL[286]
  PIN DIG_MON_COMP[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12562.825 1046.435 12563.105 1047.435 ;
    END
  END DIG_MON_COMP[61]
  PIN Data_COMP[648]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12560.585 1046.435 12560.865 1047.435 ;
    END
  END Data_COMP[648]
  PIN Data_COMP[649]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12558.905 1046.435 12559.185 1047.435 ;
    END
  END Data_COMP[649]
  PIN Data_COMP[650]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12557.225 1046.435 12557.505 1047.435 ;
    END
  END Data_COMP[650]
  PIN Data_COMP[637]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12556.105 1046.435 12556.385 1047.435 ;
    END
  END Data_COMP[637]
  PIN nTOK_COMP[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12514.105 1046.435 12514.385 1047.435 ;
    END
  END nTOK_COMP[30]
  PIN BcidMtx[855]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12511.865 1046.435 12512.145 1047.435 ;
    END
  END BcidMtx[855]
  PIN BcidMtx[854]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12510.185 1046.435 12510.465 1047.435 ;
    END
  END BcidMtx[854]
  PIN INJ_IN[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12507.945 1046.435 12508.225 1047.435 ;
    END
  END INJ_IN[284]
  PIN Data_COMP[639]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12505.705 1046.435 12505.985 1047.435 ;
    END
  END Data_COMP[639]
  PIN Data_COMP[634]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12504.025 1046.435 12504.305 1047.435 ;
    END
  END Data_COMP[634]
  PIN Data_COMP[631]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12502.345 1046.435 12502.625 1047.435 ;
    END
  END Data_COMP[631]
  PIN MASKV[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12492.265 1046.435 12492.545 1047.435 ;
    END
  END MASKV[284]
  PIN DIG_MON_COMP[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12490.025 1046.435 12490.305 1047.435 ;
    END
  END DIG_MON_COMP[60]
  PIN DIG_MON_SEL[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12487.785 1046.435 12488.065 1047.435 ;
    END
  END DIG_MON_SEL[283]
  PIN INJ_ROW[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12482.465 1046.435 12482.745 1047.435 ;
    END
  END INJ_ROW[141]
  PIN Data_COMP[617]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12480.785 1046.435 12481.065 1047.435 ;
    END
  END Data_COMP[617]
  PIN Data_HV[1095]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18748.585 1046.435 18748.865 1047.435 ;
    END
  END Data_HV[1095]
  PIN Data_COMP[629]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12452.505 1046.435 12452.785 1047.435 ;
    END
  END Data_COMP[629]
  PIN Data_COMP[615]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12450.825 1046.435 12451.105 1047.435 ;
    END
  END Data_COMP[615]
  PIN BcidMtx[851]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12447.465 1046.435 12447.745 1047.435 ;
    END
  END BcidMtx[851]
  PIN FREEZE_COMP[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12445.785 1046.435 12446.065 1047.435 ;
    END
  END FREEZE_COMP[29]
  PIN BcidMtx[847]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12444.105 1046.435 12444.385 1047.435 ;
    END
  END BcidMtx[847]
  PIN Data_COMP[612]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12441.305 1046.435 12441.585 1047.435 ;
    END
  END Data_COMP[612]
  PIN Data_COMP[624]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12426.745 1046.435 12427.025 1047.435 ;
    END
  END Data_COMP[624]
  PIN Data_COMP[625]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12425.065 1046.435 12425.345 1047.435 ;
    END
  END Data_COMP[625]
  PIN Data_COMP[609]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12423.385 1046.435 12423.665 1047.435 ;
    END
  END Data_COMP[609]
  PIN MASKH[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12421.705 1046.435 12421.985 1047.435 ;
    END
  END MASKH[141]
  PIN MASKD[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12416.665 1046.435 12416.945 1047.435 ;
    END
  END MASKD[281]
  PIN MASKV[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12413.865 1046.435 12414.145 1047.435 ;
    END
  END MASKV[281]
  PIN Data_COMP[600]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12372.425 1046.435 12372.705 1047.435 ;
    END
  END Data_COMP[600]
  PIN Data_COMP[601]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12370.745 1046.435 12371.025 1047.435 ;
    END
  END Data_COMP[601]
  PIN Data_COMP[602]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12369.625 1046.435 12369.905 1047.435 ;
    END
  END Data_COMP[602]
  PIN INJ_IN[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12367.385 1046.435 12367.665 1047.435 ;
    END
  END INJ_IN[281]
  PIN BcidMtx[844]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12364.585 1046.435 12364.865 1047.435 ;
    END
  END BcidMtx[844]
  PIN Read_COMP[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12362.905 1046.435 12363.185 1047.435 ;
    END
  END Read_COMP[28]
  PIN BcidMtx[840]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12361.225 1046.435 12361.505 1047.435 ;
    END
  END BcidMtx[840]
  PIN Data_COMP[590]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12350.025 1046.435 12350.305 1047.435 ;
    END
  END Data_COMP[590]
  PIN Data_COMP[598]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12348.345 1046.435 12348.625 1047.435 ;
    END
  END Data_COMP[598]
  PIN Data_COMP[599]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12346.665 1046.435 12346.945 1047.435 ;
    END
  END Data_COMP[599]
  PIN Data_COMP[605]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12344.985 1046.435 12345.265 1047.435 ;
    END
  END Data_COMP[605]
  PIN Data_COMP[294]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11225.545 1046.435 11225.825 1047.435 ;
    END
  END Data_COMP[294]
  PIN MASKH[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11221.905 1046.435 11222.185 1047.435 ;
    END
  END MASKH[126]
  PIN DIG_MON_SEL[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12311.945 1046.435 12312.225 1047.435 ;
    END
  END DIG_MON_SEL[279]
  PIN INJ_ROW[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12308.585 1046.435 12308.865 1047.435 ;
    END
  END INJ_ROW[139]
  PIN Data_COMP[575]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12306.905 1046.435 12307.185 1047.435 ;
    END
  END Data_COMP[575]
  PIN Data_COMP[572]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12305.225 1046.435 12305.505 1047.435 ;
    END
  END Data_COMP[572]
  PIN Data_COMP[581]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12303.545 1046.435 12303.825 1047.435 ;
    END
  END Data_COMP[581]
  PIN INJ_IN[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12301.305 1046.435 12301.585 1047.435 ;
    END
  END INJ_IN[279]
  PIN BcidMtx[838]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12285.065 1046.435 12285.345 1047.435 ;
    END
  END BcidMtx[838]
  PIN Read_COMP[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12283.385 1046.435 12283.665 1047.435 ;
    END
  END Read_COMP[27]
  PIN BcidMtx[834]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12281.705 1046.435 12281.985 1047.435 ;
    END
  END BcidMtx[834]
  PIN INJ_IN[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12280.585 1046.435 12280.865 1047.435 ;
    END
  END INJ_IN[278]
  PIN Data_COMP[576]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12278.345 1046.435 12278.625 1047.435 ;
    END
  END Data_COMP[576]
  PIN Data_COMP[571]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12276.665 1046.435 12276.945 1047.435 ;
    END
  END Data_COMP[571]
  PIN Data_COMP[568]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12274.985 1046.435 12275.265 1047.435 ;
    END
  END Data_COMP[568]
  PIN MASKV[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12234.665 1046.435 12234.945 1047.435 ;
    END
  END MASKV[278]
  PIN DIG_MON_COMP[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12232.425 1046.435 12232.705 1047.435 ;
    END
  END DIG_MON_COMP[54]
  PIN MASKD[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12229.065 1046.435 12229.345 1047.435 ;
    END
  END MASKD[277]
  PIN MASKV[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12226.265 1046.435 12226.545 1047.435 ;
    END
  END MASKV[277]
  PIN Data_COMP[554]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12225.145 1046.435 12225.425 1047.435 ;
    END
  END Data_COMP[554]
  PIN Data_COMP[559]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12222.905 1046.435 12223.185 1047.435 ;
    END
  END Data_COMP[559]
  PIN Data_COMP[553]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12221.225 1046.435 12221.505 1047.435 ;
    END
  END Data_COMP[553]
  PIN INJ_IN[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12211.145 1046.435 12211.425 1047.435 ;
    END
  END INJ_IN[277]
  PIN BcidMtx[831]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12207.785 1046.435 12208.065 1047.435 ;
    END
  END BcidMtx[831]
  PIN BcidMtx[830]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12206.105 1046.435 12206.385 1047.435 ;
    END
  END BcidMtx[830]
  PIN BcidMtx[828]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12204.985 1046.435 12205.265 1047.435 ;
    END
  END BcidMtx[828]
  PIN Data_COMP[555]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12199.665 1046.435 12199.945 1047.435 ;
    END
  END Data_COMP[555]
  PIN Data_COMP[550]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12172.505 1046.435 12172.785 1047.435 ;
    END
  END Data_COMP[550]
  PIN Data_COMP[557]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12171.385 1046.435 12171.665 1047.435 ;
    END
  END Data_COMP[557]
  PIN MASKV[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12169.145 1046.435 12169.425 1047.435 ;
    END
  END MASKV[276]
  PIN DIG_MON_COMP[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12166.905 1046.435 12167.185 1047.435 ;
    END
  END DIG_MON_COMP[52]
  PIN DIG_MON_SEL[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12165.225 1046.435 12165.505 1047.435 ;
    END
  END DIG_MON_SEL[276]
  PIN INJ_ROW[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12161.305 1046.435 12161.585 1047.435 ;
    END
  END INJ_ROW[137]
  PIN Data_COMP[533]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12159.625 1046.435 12159.905 1047.435 ;
    END
  END Data_COMP[533]
  PIN Data_COMP[544]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12145.625 1046.435 12145.905 1047.435 ;
    END
  END Data_COMP[544]
  PIN Data_COMP[532]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12142.825 1046.435 12143.105 1047.435 ;
    END
  END Data_COMP[532]
  PIN INJ_IN[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12141.145 1046.435 12141.425 1047.435 ;
    END
  END INJ_IN[275]
  PIN BcidMtx[827]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12138.905 1046.435 12139.185 1047.435 ;
    END
  END BcidMtx[827]
  PIN Read_COMP[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12136.665 1046.435 12136.945 1047.435 ;
    END
  END Read_COMP[25]
  PIN BcidMtx[822]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12134.985 1046.435 12135.265 1047.435 ;
    END
  END BcidMtx[822]
  PIN INJ_IN[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12133.865 1046.435 12134.145 1047.435 ;
    END
  END INJ_IN[274]
  PIN Data_COMP[535]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12091.865 1046.435 12092.145 1047.435 ;
    END
  END Data_COMP[535]
  PIN Data_COMP[536]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12090.185 1046.435 12090.465 1047.435 ;
    END
  END Data_COMP[536]
  PIN Data_COMP[526]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12089.625 1046.435 12089.905 1047.435 ;
    END
  END Data_COMP[526]
  PIN MASKD[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12086.825 1046.435 12087.105 1047.435 ;
    END
  END MASKD[274]
  PIN DIG_MON_SEL[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12084.025 1046.435 12084.305 1047.435 ;
    END
  END DIG_MON_SEL[274]
  PIN DIG_MON_SEL[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12083.465 1046.435 12083.745 1047.435 ;
    END
  END DIG_MON_SEL[273]
  PIN Data_COMP[522]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12070.585 1046.435 12070.865 1047.435 ;
    END
  END Data_COMP[522]
  PIN Data_COMP[523]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12068.905 1046.435 12069.185 1047.435 ;
    END
  END Data_COMP[523]
  PIN Data_COMP[509]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12068.345 1046.435 12068.625 1047.435 ;
    END
  END Data_COMP[509]
  PIN Data_HV[1057]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18611.385 1046.435 18611.665 1047.435 ;
    END
  END Data_HV[1057]
  PIN nTOK_COMP[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12061.345 1046.435 12061.625 1047.435 ;
    END
  END nTOK_COMP[24]
  PIN BcidMtx[821]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12060.225 1046.435 12060.505 1047.435 ;
    END
  END BcidMtx[821]
  PIN BcidMtx[817]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12031.385 1046.435 12031.665 1047.435 ;
    END
  END BcidMtx[817]
  PIN Data_COMP[507]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12028.585 1046.435 12028.865 1047.435 ;
    END
  END Data_COMP[507]
  PIN Data_COMP[513]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12027.465 1046.435 12027.745 1047.435 ;
    END
  END Data_COMP[513]
  PIN Data_COMP[520]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12025.225 1046.435 12025.505 1047.435 ;
    END
  END Data_COMP[520]
  PIN Data_COMP[504]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12023.545 1046.435 12023.825 1047.435 ;
    END
  END Data_COMP[504]
  PIN MASKV[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12022.425 1046.435 12022.705 1047.435 ;
    END
  END MASKV[272]
  PIN DIG_MON_SEL[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12005.625 1046.435 12005.905 1047.435 ;
    END
  END DIG_MON_SEL[272]
  PIN DIG_MON_COMP[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12002.825 1046.435 12003.105 1047.435 ;
    END
  END DIG_MON_COMP[47]
  PIN INJ_ROW[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12001.705 1046.435 12001.985 1047.435 ;
    END
  END INJ_ROW[135]
  PIN Data_COMP[502]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11998.905 1046.435 11999.185 1047.435 ;
    END
  END Data_COMP[502]
  PIN Data_COMP[503]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11997.225 1046.435 11997.505 1047.435 ;
    END
  END Data_COMP[503]
  PIN Data_COMP[497]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11996.665 1046.435 11996.945 1047.435 ;
    END
  END Data_COMP[497]
  PIN BcidMtx[1321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18751.385 1046.435 18751.665 1047.435 ;
    END
  END BcidMtx[1321]
  PIN BcidMtx[813]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11951.865 1046.435 11952.145 1047.435 ;
    END
  END BcidMtx[813]
  PIN FREEZE_COMP[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11951.305 1046.435 11951.585 1047.435 ;
    END
  END FREEZE_COMP[23]
  PIN INJ_IN[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11947.945 1046.435 11948.225 1047.435 ;
    END
  END INJ_IN[270]
  PIN Data_COMP[492]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11945.705 1046.435 11945.985 1047.435 ;
    END
  END Data_COMP[492]
  PIN Data_COMP[498]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11945.145 1046.435 11945.425 1047.435 ;
    END
  END Data_COMP[498]
  PIN Data_COMP[484]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11942.345 1046.435 11942.625 1047.435 ;
    END
  END Data_COMP[484]
  PIN MASKV[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11932.265 1046.435 11932.545 1047.435 ;
    END
  END MASKV[270]
  PIN MASKH[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11931.705 1046.435 11931.985 1047.435 ;
    END
  END MASKH[135]
  PIN DIG_MON_SEL[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11927.785 1046.435 11928.065 1047.435 ;
    END
  END DIG_MON_SEL[269]
  PIN INJ_ROW[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11922.465 1046.435 11922.745 1047.435 ;
    END
  END INJ_ROW[134]
  PIN MASKV[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11921.905 1046.435 11922.185 1047.435 ;
    END
  END MASKV[269]
  PIN Data_COMP[474]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11920.225 1046.435 11920.505 1047.435 ;
    END
  END Data_COMP[474]
  PIN Data_COMP[476]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11891.945 1046.435 11892.225 1047.435 ;
    END
  END Data_COMP[476]
  PIN Data_COMP[468]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11890.825 1046.435 11891.105 1047.435 ;
    END
  END Data_COMP[468]
  PIN BcidMtx[809]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11887.465 1046.435 11887.745 1047.435 ;
    END
  END BcidMtx[809]
  PIN BcidMtx[807]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11886.345 1046.435 11886.625 1047.435 ;
    END
  END BcidMtx[807]
  PIN BcidMtx[806]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11884.665 1046.435 11884.945 1047.435 ;
    END
  END BcidMtx[806]
  PIN BcidMtx[804]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11883.545 1046.435 11883.825 1047.435 ;
    END
  END BcidMtx[804]
  PIN Data_COMP[464]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11880.745 1046.435 11881.025 1047.435 ;
    END
  END Data_COMP[464]
  PIN Data_COMP[466]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11865.625 1046.435 11865.905 1047.435 ;
    END
  END Data_COMP[466]
  PIN Data_COMP[473]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11864.505 1046.435 11864.785 1047.435 ;
    END
  END Data_COMP[473]
  PIN Data_COMP[479]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11862.825 1046.435 11863.105 1047.435 ;
    END
  END Data_COMP[479]
  PIN DIG_MON_COMP[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11860.025 1046.435 11860.305 1047.435 ;
    END
  END DIG_MON_COMP[44]
  PIN DIG_MON_SEL[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11858.345 1046.435 11858.625 1047.435 ;
    END
  END DIG_MON_SEL[268]
  PIN DIG_MON_COMP[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11855.545 1046.435 11855.825 1047.435 ;
    END
  END DIG_MON_COMP[43]
  PIN Data_COMP[453]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11812.425 1046.435 11812.705 1047.435 ;
    END
  END Data_COMP[453]
  PIN Data_COMP[446]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11811.305 1046.435 11811.585 1047.435 ;
    END
  END Data_COMP[446]
  PIN Data_COMP[455]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11809.625 1046.435 11809.905 1047.435 ;
    END
  END Data_COMP[455]
  PIN nTOK_COMP[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11806.265 1046.435 11806.545 1047.435 ;
    END
  END nTOK_COMP[21]
  PIN BcidMtx[802]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11804.585 1046.435 11804.865 1047.435 ;
    END
  END BcidMtx[802]
  PIN BcidMtx[799]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11801.785 1046.435 11802.065 1047.435 ;
    END
  END BcidMtx[799]
  PIN INJ_IN[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11791.705 1046.435 11791.985 1047.435 ;
    END
  END INJ_IN[266]
  PIN Data_COMP[443]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11790.025 1046.435 11790.305 1047.435 ;
    END
  END Data_COMP[443]
  PIN Data_COMP[451]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11788.345 1046.435 11788.625 1047.435 ;
    END
  END Data_COMP[451]
  PIN Data_COMP[441]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11785.545 1046.435 11785.825 1047.435 ;
    END
  END Data_COMP[441]
  PIN BcidMtx[1262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17962.345 1046.435 17962.625 1047.435 ;
    END
  END BcidMtx[1262]
  PIN Data_HV[884]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17950.025 1046.435 17950.305 1047.435 ;
    END
  END Data_HV[884]
  PIN Data_HV[897]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17948.905 1046.435 17949.185 1047.435 ;
    END
  END Data_HV[897]
  PIN Data_HV[886]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17947.785 1046.435 17948.065 1047.435 ;
    END
  END Data_HV[886]
  PIN Data_HV[883]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17946.105 1046.435 17946.385 1047.435 ;
    END
  END Data_HV[883]
  PIN MASKH[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17941.905 1046.435 17942.185 1047.435 ;
    END
  END MASKH[210]
  PIN DIG_MON_HV[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17940.225 1046.435 17940.505 1047.435 ;
    END
  END DIG_MON_HV[84]
  PIN FREEZE_HV[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18193.065 1046.435 18193.345 1047.435 ;
    END
  END FREEZE_HV[45]
  PIN INJ_ROW[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 19028.585 1046.435 19028.865 1047.435 ;
    END
  END INJ_ROW[223]
  PIN Data_HV[1173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 19027.465 1046.435 19027.745 1047.435 ;
    END
  END Data_HV[1173]
  PIN Data_HV[1174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 19025.785 1046.435 19026.065 1047.435 ;
    END
  END Data_HV[1174]
  PIN Data_HV[1169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 19023.545 1046.435 19023.825 1047.435 ;
    END
  END Data_HV[1169]
  PIN Data_HV[1161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 19022.425 1046.435 19022.705 1047.435 ;
    END
  END Data_HV[1161]
  PIN BcidMtx[1343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 19005.625 1046.435 19005.905 1047.435 ;
    END
  END BcidMtx[1343]
  PIN BcidMtx[1340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 19002.825 1046.435 19003.105 1047.435 ;
    END
  END BcidMtx[1340]
  PIN BcidMtx[1338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 19001.705 1046.435 19001.985 1047.435 ;
    END
  END BcidMtx[1338]
  PIN Data_HV[1157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18998.905 1046.435 18999.185 1047.435 ;
    END
  END Data_HV[1157]
  PIN Data_HV[1159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18996.665 1046.435 18996.945 1047.435 ;
    END
  END Data_HV[1159]
  PIN Data_HV[1166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18995.545 1046.435 18995.825 1047.435 ;
    END
  END Data_HV[1166]
  PIN MASKH[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18954.105 1046.435 18954.385 1047.435 ;
    END
  END MASKH[223]
  PIN DIG_MON_HV[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18952.425 1046.435 18952.705 1047.435 ;
    END
  END DIG_MON_HV[110]
  PIN DIG_MON_SEL[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18950.745 1046.435 18951.025 1047.435 ;
    END
  END DIG_MON_SEL[446]
  PIN DIG_MON_HV[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18947.945 1046.435 18948.225 1047.435 ;
    END
  END DIG_MON_HV[109]
  PIN Data_HV[1146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18944.585 1046.435 18944.865 1047.435 ;
    END
  END Data_HV[1146]
  PIN Data_HV[1153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18944.025 1046.435 18944.305 1047.435 ;
    END
  END Data_HV[1153]
  PIN Data_HV[1141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18941.225 1046.435 18941.505 1047.435 ;
    END
  END Data_HV[1141]
  PIN nTOK_HV[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18930.025 1046.435 18930.305 1047.435 ;
    END
  END nTOK_HV[54]
  PIN BcidMtx[1336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18928.345 1046.435 18928.625 1047.435 ;
    END
  END BcidMtx[1336]
  PIN BcidMtx[1334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18926.105 1046.435 18926.385 1047.435 ;
    END
  END BcidMtx[1334]
  PIN INJ_IN[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18921.905 1046.435 18922.185 1047.435 ;
    END
  END INJ_IN[444]
  PIN Data_HV[1031]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18510.025 1046.435 18510.305 1047.435 ;
    END
  END Data_HV[1031]
  PIN FREEZE_HV[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18523.465 1046.435 18523.745 1047.435 ;
    END
  END FREEZE_HV[49]
  PIN Data_HV[1046]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18504.985 1046.435 18505.265 1047.435 ;
    END
  END Data_HV[1046]
  PIN Data_HV[1043]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18529.625 1046.435 18529.905 1047.435 ;
    END
  END Data_HV[1043]
  PIN Data_HV[1038]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18509.465 1046.435 18509.745 1047.435 ;
    END
  END Data_HV[1038]
  PIN Data_HV[1143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18919.665 1046.435 18919.945 1047.435 ;
    END
  END Data_HV[1143]
  PIN Data_HV[1149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18919.105 1046.435 18919.385 1047.435 ;
    END
  END Data_HV[1149]
  PIN Data_HV[1144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18918.545 1046.435 18918.825 1047.435 ;
    END
  END Data_HV[1144]
  PIN Data_HV[1053]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18601.305 1046.435 18601.585 1047.435 ;
    END
  END Data_HV[1053]
  PIN DIG_MON_HV[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18575.545 1046.435 18575.825 1047.435 ;
    END
  END DIG_MON_HV[99]
  PIN INJ_ROW[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18574.425 1046.435 18574.705 1047.435 ;
    END
  END INJ_ROW[217]
  PIN MASKV[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18573.865 1046.435 18574.145 1047.435 ;
    END
  END MASKV[435]
  PIN Data_HV[1047]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18533.545 1046.435 18533.825 1047.435 ;
    END
  END Data_HV[1047]
  PIN MASKD[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18501.345 1046.435 18501.625 1047.435 ;
    END
  END MASKD[434]
  PIN Read_HV[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18522.905 1046.435 18523.185 1047.435 ;
    END
  END Read_HV[49]
  PIN MASKV[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18502.465 1046.435 18502.745 1047.435 ;
    END
  END MASKV[434]
  PIN Data_HV[1036]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18529.065 1046.435 18529.345 1047.435 ;
    END
  END Data_HV[1036]
  PIN Data_HV[1044]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18508.905 1046.435 18509.185 1047.435 ;
    END
  END Data_HV[1044]
  PIN DIG_MON_HV[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18500.225 1046.435 18500.505 1047.435 ;
    END
  END DIG_MON_HV[98]
  PIN MASKH[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18501.905 1046.435 18502.185 1047.435 ;
    END
  END MASKH[217]
  PIN Data_HV[1035]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18528.505 1046.435 18528.785 1047.435 ;
    END
  END Data_HV[1035]
  PIN Data_HV[1039]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18508.345 1046.435 18508.625 1047.435 ;
    END
  END Data_HV[1039]
  PIN BcidMtx[1304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18522.345 1046.435 18522.625 1047.435 ;
    END
  END BcidMtx[1304]
  PIN Data_HV[1033]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18507.785 1046.435 18508.065 1047.435 ;
    END
  END Data_HV[1033]
  PIN DIG_MON_SEL[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18498.545 1046.435 18498.825 1047.435 ;
    END
  END DIG_MON_SEL[434]
  PIN BcidMtx[1303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18521.785 1046.435 18522.065 1047.435 ;
    END
  END BcidMtx[1303]
  PIN nTOK_HV[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18526.265 1046.435 18526.545 1047.435 ;
    END
  END nTOK_HV[49]
  PIN Data_HV[1045]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18507.225 1046.435 18507.505 1047.435 ;
    END
  END Data_HV[1045]
  PIN BcidMtx[1302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18521.225 1046.435 18521.505 1047.435 ;
    END
  END BcidMtx[1302]
  PIN BcidMtx[1307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18525.145 1046.435 18525.425 1047.435 ;
    END
  END BcidMtx[1307]
  PIN Data_HV[1040]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18506.665 1046.435 18506.945 1047.435 ;
    END
  END Data_HV[1040]
  PIN FREEZE_HV[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18753.065 1046.435 18753.345 1047.435 ;
    END
  END FREEZE_HV[52]
  PIN INJ_IN[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18511.705 1046.435 18511.985 1047.435 ;
    END
  END INJ_IN[434]
  PIN BcidMtx[1306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18524.585 1046.435 18524.865 1047.435 ;
    END
  END BcidMtx[1306]
  PIN Data_HV[1030]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18506.105 1046.435 18506.385 1047.435 ;
    END
  END Data_HV[1030]
  PIN Data_HV[1032]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18510.585 1046.435 18510.865 1047.435 ;
    END
  END Data_HV[1032]
  PIN BcidMtx[1305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18524.025 1046.435 18524.305 1047.435 ;
    END
  END BcidMtx[1305]
  PIN Data_HV[1029]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18505.545 1046.435 18505.825 1047.435 ;
    END
  END Data_HV[1029]
  PIN INJ_IN_MON_L
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1137.985 1046.435 1138.265 1047.435 ;
    END
  END INJ_IN_MON_L
  PIN INJ_IN_MON_R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 19032.505 1046.435 19032.785 1047.435 ;
    END
  END INJ_IN_MON_R
  PIN Data_COMP[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10666.105 1046.435 10666.385 1047.435 ;
    END
  END Data_COMP[148]
  PIN MASKV[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10662.465 1046.435 10662.745 1047.435 ;
    END
  END MASKV[238]
  PIN MASKD[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10661.345 1046.435 10661.625 1047.435 ;
    END
  END MASKD[238]
  PIN FREEZE_COMP[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10913.065 1046.435 10913.345 1047.435 ;
    END
  END FREEZE_COMP[10]
  PIN DIG_MON_COMP[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11749.705 1046.435 11749.985 1047.435 ;
    END
  END DIG_MON_COMP[41]
  PIN MASKV[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11748.025 1046.435 11748.305 1047.435 ;
    END
  END MASKV[265]
  PIN Data_COMP[439]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11745.785 1046.435 11746.065 1047.435 ;
    END
  END Data_COMP[439]
  PIN Data_COMP[440]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11744.105 1046.435 11744.385 1047.435 ;
    END
  END Data_COMP[440]
  PIN Data_COMP[427]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11742.985 1046.435 11743.265 1047.435 ;
    END
  END Data_COMP[427]
  PIN BcidMtx[797]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11725.625 1046.435 11725.905 1047.435 ;
    END
  END BcidMtx[797]
  PIN FREEZE_COMP[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11723.945 1046.435 11724.225 1047.435 ;
    END
  END FREEZE_COMP[20]
  PIN BcidMtx[794]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11722.825 1046.435 11723.105 1047.435 ;
    END
  END BcidMtx[794]
  PIN Data_COMP[423]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11719.465 1046.435 11719.745 1047.435 ;
    END
  END Data_COMP[423]
  PIN Data_COMP[435]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11717.785 1046.435 11718.065 1047.435 ;
    END
  END Data_COMP[435]
  PIN Data_COMP[424]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11716.665 1046.435 11716.945 1047.435 ;
    END
  END Data_COMP[424]
  PIN Data_COMP[420]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11714.425 1046.435 11714.705 1047.435 ;
    END
  END Data_COMP[420]
  PIN MASKH[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11674.105 1046.435 11674.385 1047.435 ;
    END
  END MASKH[132]
  PIN DIG_MON_COMP[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11672.425 1046.435 11672.705 1047.435 ;
    END
  END DIG_MON_COMP[40]
  PIN MASKD[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11669.065 1046.435 11669.345 1047.435 ;
    END
  END MASKD[263]
  PIN MASKV[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11666.265 1046.435 11666.545 1047.435 ;
    END
  END MASKV[263]
  PIN Data_COMP[407]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11665.145 1046.435 11665.425 1047.435 ;
    END
  END Data_COMP[407]
  PIN Data_COMP[412]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11662.905 1046.435 11663.185 1047.435 ;
    END
  END Data_COMP[412]
  PIN Data_COMP[406]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11661.225 1046.435 11661.505 1047.435 ;
    END
  END Data_COMP[406]
  PIN INJ_IN[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11651.145 1046.435 11651.425 1047.435 ;
    END
  END INJ_IN[263]
  PIN BcidMtx[789]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11647.785 1046.435 11648.065 1047.435 ;
    END
  END BcidMtx[789]
  PIN BcidMtx[788]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11646.105 1046.435 11646.385 1047.435 ;
    END
  END BcidMtx[788]
  PIN BcidMtx[786]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11644.985 1046.435 11645.265 1047.435 ;
    END
  END BcidMtx[786]
  PIN Data_COMP[408]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11639.665 1046.435 11639.945 1047.435 ;
    END
  END Data_COMP[408]
  PIN Data_COMP[403]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11612.505 1046.435 11612.785 1047.435 ;
    END
  END Data_COMP[403]
  PIN Data_COMP[410]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11611.385 1046.435 11611.665 1047.435 ;
    END
  END Data_COMP[410]
  PIN MASKV[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11609.145 1046.435 11609.425 1047.435 ;
    END
  END MASKV[262]
  PIN DIG_MON_COMP[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11606.905 1046.435 11607.185 1047.435 ;
    END
  END DIG_MON_COMP[38]
  PIN DIG_MON_SEL[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11605.225 1046.435 11605.505 1047.435 ;
    END
  END DIG_MON_SEL[262]
  PIN INJ_ROW[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11601.305 1046.435 11601.585 1047.435 ;
    END
  END INJ_ROW[130]
  PIN Data_COMP[386]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11599.625 1046.435 11599.905 1047.435 ;
    END
  END Data_COMP[386]
  PIN Data_COMP[397]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11585.625 1046.435 11585.905 1047.435 ;
    END
  END Data_COMP[397]
  PIN Data_COMP[392]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11583.385 1046.435 11583.665 1047.435 ;
    END
  END Data_COMP[392]
  PIN INJ_IN[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11581.145 1046.435 11581.425 1047.435 ;
    END
  END INJ_IN[261]
  PIN BcidMtx[785]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11578.905 1046.435 11579.185 1047.435 ;
    END
  END BcidMtx[785]
  PIN Read_COMP[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11576.665 1046.435 11576.945 1047.435 ;
    END
  END Read_COMP[18]
  PIN BcidMtx[780]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11574.985 1046.435 11575.265 1047.435 ;
    END
  END BcidMtx[780]
  PIN Data_COMP[381]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11534.105 1046.435 11534.385 1047.435 ;
    END
  END Data_COMP[381]
  PIN Data_COMP[388]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11531.865 1046.435 11532.145 1047.435 ;
    END
  END Data_COMP[388]
  PIN Data_COMP[389]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11530.185 1046.435 11530.465 1047.435 ;
    END
  END Data_COMP[389]
  PIN Data_COMP[378]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11529.065 1046.435 11529.345 1047.435 ;
    END
  END Data_COMP[378]
  PIN MASKD[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11526.825 1046.435 11527.105 1047.435 ;
    END
  END MASKD[260]
  PIN DIG_MON_SEL[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11524.025 1046.435 11524.305 1047.435 ;
    END
  END DIG_MON_SEL[260]
  PIN MASKD[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11522.345 1046.435 11522.625 1047.435 ;
    END
  END MASKD[259]
  PIN Data_COMP[375]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11510.585 1046.435 11510.865 1047.435 ;
    END
  END Data_COMP[375]
  PIN Data_COMP[376]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11508.905 1046.435 11509.185 1047.435 ;
    END
  END Data_COMP[376]
  PIN Data_COMP[370]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11507.785 1046.435 11508.065 1047.435 ;
    END
  END Data_COMP[370]
  PIN Data_COMP[363]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11505.545 1046.435 11505.825 1047.435 ;
    END
  END Data_COMP[363]
  PIN BcidMtx[779]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11500.225 1046.435 11500.505 1047.435 ;
    END
  END BcidMtx[779]
  PIN BcidMtx[777]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11499.105 1046.435 11499.385 1047.435 ;
    END
  END BcidMtx[777]
  PIN BcidMtx[774]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11470.825 1046.435 11471.105 1047.435 ;
    END
  END BcidMtx[774]
  PIN Data_COMP[359]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11468.025 1046.435 11468.305 1047.435 ;
    END
  END Data_COMP[359]
  PIN Data_COMP[372]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11466.905 1046.435 11467.185 1047.435 ;
    END
  END Data_COMP[372]
  PIN Data_COMP[368]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11464.665 1046.435 11464.945 1047.435 ;
    END
  END Data_COMP[368]
  PIN Data_COMP[374]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11462.985 1046.435 11463.265 1047.435 ;
    END
  END Data_COMP[374]
  PIN MASKH[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11461.865 1046.435 11462.145 1047.435 ;
    END
  END MASKH[129]
  PIN DIG_MON_SEL[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11445.625 1046.435 11445.905 1047.435 ;
    END
  END DIG_MON_SEL[258]
  PIN DIG_MON_COMP[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11442.825 1046.435 11443.105 1047.435 ;
    END
  END DIG_MON_COMP[33]
  PIN MASKV[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11441.145 1046.435 11441.425 1047.435 ;
    END
  END MASKV[257]
  PIN Data_COMP[355]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11438.905 1046.435 11439.185 1047.435 ;
    END
  END Data_COMP[355]
  PIN Data_COMP[356]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11437.225 1046.435 11437.505 1047.435 ;
    END
  END Data_COMP[356]
  PIN Data_COMP[343]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11436.105 1046.435 11436.385 1047.435 ;
    END
  END Data_COMP[343]
  PIN BcidMtx[773]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11392.985 1046.435 11393.265 1047.435 ;
    END
  END BcidMtx[773]
  PIN FREEZE_COMP[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11391.305 1046.435 11391.585 1047.435 ;
    END
  END FREEZE_COMP[16]
  PIN BcidMtx[770]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11390.185 1046.435 11390.465 1047.435 ;
    END
  END BcidMtx[770]
  PIN BcidMtx[768]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11389.065 1046.435 11389.345 1047.435 ;
    END
  END BcidMtx[768]
  PIN Data_COMP[338]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11386.265 1046.435 11386.545 1047.435 ;
    END
  END Data_COMP[338]
  PIN Data_COMP[351]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11385.145 1046.435 11385.425 1047.435 ;
    END
  END Data_COMP[351]
  PIN Data_COMP[347]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11382.905 1046.435 11383.185 1047.435 ;
    END
  END Data_COMP[347]
  PIN Data_COMP[353]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11381.225 1046.435 11381.505 1047.435 ;
    END
  END Data_COMP[353]
  PIN MASKH[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11371.705 1046.435 11371.985 1047.435 ;
    END
  END MASKH[128]
  PIN DIG_MON_SEL[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11368.345 1046.435 11368.625 1047.435 ;
    END
  END DIG_MON_SEL[256]
  PIN DIG_MON_COMP[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11365.545 1046.435 11365.825 1047.435 ;
    END
  END DIG_MON_COMP[31]
  PIN MASKV[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11361.905 1046.435 11362.185 1047.435 ;
    END
  END MASKV[255]
  PIN Data_COMP[334]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11359.665 1046.435 11359.945 1047.435 ;
    END
  END Data_COMP[334]
  PIN Data_COMP[335]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11332.505 1046.435 11332.785 1047.435 ;
    END
  END Data_COMP[335]
  PIN Data_COMP[322]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11331.385 1046.435 11331.665 1047.435 ;
    END
  END Data_COMP[322]
  PIN BcidMtx[767]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11327.465 1046.435 11327.745 1047.435 ;
    END
  END BcidMtx[767]
  PIN FREEZE_COMP[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11325.785 1046.435 11326.065 1047.435 ;
    END
  END FREEZE_COMP[15]
  PIN BcidMtx[764]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11324.665 1046.435 11324.945 1047.435 ;
    END
  END BcidMtx[764]
  PIN BcidMtx[1324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18779.665 1046.435 18779.945 1047.435 ;
    END
  END BcidMtx[1324]
  PIN Data_COMP[324]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11320.185 1046.435 11320.465 1047.435 ;
    END
  END Data_COMP[324]
  PIN Data_COMP[325]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11306.185 1046.435 11306.465 1047.435 ;
    END
  END Data_COMP[325]
  PIN Data_COMP[316]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11303.945 1046.435 11304.225 1047.435 ;
    END
  END Data_COMP[316]
  PIN MASKV[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11302.265 1046.435 11302.545 1047.435 ;
    END
  END MASKV[254]
  PIN DIG_MON_COMP[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11300.025 1046.435 11300.305 1047.435 ;
    END
  END DIG_MON_COMP[30]
  PIN DIG_MON_SEL[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11297.785 1046.435 11298.065 1047.435 ;
    END
  END DIG_MON_SEL[253]
  PIN INJ_ROW[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11294.425 1046.435 11294.705 1047.435 ;
    END
  END INJ_ROW[126]
  PIN Data_COMP[302]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11252.985 1046.435 11253.265 1047.435 ;
    END
  END Data_COMP[302]
  PIN Data_COMP[299]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11251.305 1046.435 11251.585 1047.435 ;
    END
  END Data_COMP[299]
  PIN Data_COMP[308]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11249.625 1046.435 11249.905 1047.435 ;
    END
  END Data_COMP[308]
  PIN INJ_IN[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11247.385 1046.435 11247.665 1047.435 ;
    END
  END INJ_IN[253]
  PIN BcidMtx[760]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11244.585 1046.435 11244.865 1047.435 ;
    END
  END BcidMtx[760]
  PIN Read_COMP[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11242.905 1046.435 11243.185 1047.435 ;
    END
  END Read_COMP[14]
  PIN BcidMtx[1323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18779.105 1046.435 18779.385 1047.435 ;
    END
  END BcidMtx[1323]
  PIN Data_COMP[297]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11230.585 1046.435 11230.865 1047.435 ;
    END
  END Data_COMP[297]
  PIN Data_COMP[309]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11228.905 1046.435 11229.185 1047.435 ;
    END
  END Data_COMP[309]
  PIN Data_COMP[310]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11227.225 1046.435 11227.505 1047.435 ;
    END
  END Data_COMP[310]
  PIN MASKH[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10101.905 1046.435 10102.185 1047.435 ;
    END
  END MASKH[112]
  PIN DIG_MON_SEL[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11191.945 1046.435 11192.225 1047.435 ;
    END
  END DIG_MON_SEL[251]
  PIN INJ_ROW[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11188.585 1046.435 11188.865 1047.435 ;
    END
  END INJ_ROW[125]
  PIN Data_COMP[281]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11186.905 1046.435 11187.185 1047.435 ;
    END
  END Data_COMP[281]
  PIN Data_COMP[278]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11185.225 1046.435 11185.505 1047.435 ;
    END
  END Data_COMP[278]
  PIN Data_COMP[287]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11183.545 1046.435 11183.825 1047.435 ;
    END
  END Data_COMP[287]
  PIN INJ_IN[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11181.305 1046.435 11181.585 1047.435 ;
    END
  END INJ_IN[251]
  PIN BcidMtx[754]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11165.065 1046.435 11165.345 1047.435 ;
    END
  END BcidMtx[754]
  PIN Read_COMP[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11163.385 1046.435 11163.665 1047.435 ;
    END
  END Read_COMP[13]
  PIN BcidMtx[750]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11161.705 1046.435 11161.985 1047.435 ;
    END
  END BcidMtx[750]
  PIN Data_COMP[275]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11158.905 1046.435 11159.185 1047.435 ;
    END
  END Data_COMP[275]
  PIN Data_COMP[283]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11157.225 1046.435 11157.505 1047.435 ;
    END
  END Data_COMP[283]
  PIN Data_COMP[284]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11155.545 1046.435 11155.825 1047.435 ;
    END
  END Data_COMP[284]
  PIN Data_COMP[290]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11153.865 1046.435 11154.145 1047.435 ;
    END
  END Data_COMP[290]
  PIN Data_HV[1070]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18612.505 1046.435 18612.785 1047.435 ;
    END
  END Data_HV[1070]
  PIN DIG_MON_COMP[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11112.425 1046.435 11112.705 1047.435 ;
    END
  END DIG_MON_COMP[26]
  PIN DIG_MON_SEL[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11110.745 1046.435 11111.025 1047.435 ;
    END
  END DIG_MON_SEL[250]
  PIN Data_COMP[270]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11105.705 1046.435 11105.985 1047.435 ;
    END
  END Data_COMP[270]
  PIN Data_COMP[264]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11104.585 1046.435 11104.865 1047.435 ;
    END
  END Data_COMP[264]
  PIN Data_COMP[257]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11103.465 1046.435 11103.745 1047.435 ;
    END
  END Data_COMP[257]
  PIN Data_COMP[266]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11101.785 1046.435 11102.065 1047.435 ;
    END
  END Data_COMP[266]
  PIN INJ_IN[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11091.145 1046.435 11091.425 1047.435 ;
    END
  END INJ_IN[249]
  PIN BcidMtx[749]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11088.905 1046.435 11089.185 1047.435 ;
    END
  END BcidMtx[749]
  PIN Read_COMP[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11086.665 1046.435 11086.945 1047.435 ;
    END
  END Read_COMP[12]
  PIN BcidMtx[744]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11084.985 1046.435 11085.265 1047.435 ;
    END
  END BcidMtx[744]
  PIN Data_COMP[255]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11080.785 1046.435 11081.065 1047.435 ;
    END
  END Data_COMP[255]
  PIN Data_COMP[262]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11078.545 1046.435 11078.825 1047.435 ;
    END
  END Data_COMP[262]
  PIN Data_COMP[263]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11051.385 1046.435 11051.665 1047.435 ;
    END
  END Data_COMP[263]
  PIN Data_COMP[252]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11050.265 1046.435 11050.545 1047.435 ;
    END
  END Data_COMP[252]
  PIN MASKD[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11048.025 1046.435 11048.305 1047.435 ;
    END
  END MASKD[248]
  PIN DIG_MON_SEL[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11045.225 1046.435 11045.505 1047.435 ;
    END
  END DIG_MON_SEL[248]
  PIN MASKD[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11043.545 1046.435 11043.825 1047.435 ;
    END
  END MASKD[247]
  PIN Data_COMP[249]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11040.185 1046.435 11040.465 1047.435 ;
    END
  END Data_COMP[249]
  PIN Data_COMP[250]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11025.625 1046.435 11025.905 1047.435 ;
    END
  END Data_COMP[250]
  PIN Data_COMP[244]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11024.505 1046.435 11024.785 1047.435 ;
    END
  END Data_COMP[244]
  PIN Data_COMP[237]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11022.265 1046.435 11022.545 1047.435 ;
    END
  END Data_COMP[237]
  PIN BcidMtx[743]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11018.905 1046.435 11019.185 1047.435 ;
    END
  END BcidMtx[743]
  PIN BcidMtx[741]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11017.785 1046.435 11018.065 1047.435 ;
    END
  END BcidMtx[741]
  PIN BcidMtx[739]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11015.545 1046.435 11015.825 1047.435 ;
    END
  END BcidMtx[739]
  PIN Data_COMP[234]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10974.105 1046.435 10974.385 1047.435 ;
    END
  END Data_COMP[234]
  PIN Data_COMP[240]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10972.985 1046.435 10973.265 1047.435 ;
    END
  END Data_COMP[240]
  PIN Data_COMP[247]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10970.745 1046.435 10971.025 1047.435 ;
    END
  END Data_COMP[247]
  PIN Data_COMP[231]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10969.065 1046.435 10969.345 1047.435 ;
    END
  END Data_COMP[231]
  PIN MASKV[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10967.945 1046.435 10968.225 1047.435 ;
    END
  END MASKV[246]
  PIN MASKD[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10962.345 1046.435 10962.625 1047.435 ;
    END
  END MASKD[245]
  PIN INJ_ROW[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10951.705 1046.435 10951.985 1047.435 ;
    END
  END INJ_ROW[122]
  PIN Data_COMP[222]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10949.465 1046.435 10949.745 1047.435 ;
    END
  END Data_COMP[222]
  PIN Data_COMP[223]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10947.785 1046.435 10948.065 1047.435 ;
    END
  END Data_COMP[223]
  PIN Data_COMP[224]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10946.665 1046.435 10946.945 1047.435 ;
    END
  END Data_COMP[224]
  PIN nTOK_COMP[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10941.345 1046.435 10941.625 1047.435 ;
    END
  END nTOK_COMP[10]
  PIN BcidMtx[735]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10939.105 1046.435 10939.385 1047.435 ;
    END
  END BcidMtx[735]
  PIN BcidMtx[734]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10911.945 1046.435 10912.225 1047.435 ;
    END
  END BcidMtx[734]
  PIN Data_HV[1063]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18613.065 1046.435 18613.345 1047.435 ;
    END
  END Data_HV[1063]
  PIN Data_COMP[212]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10908.025 1046.435 10908.305 1047.435 ;
    END
  END Data_COMP[212]
  PIN Data_COMP[225]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10906.905 1046.435 10907.185 1047.435 ;
    END
  END Data_COMP[225]
  PIN Data_COMP[221]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10904.665 1046.435 10904.945 1047.435 ;
    END
  END Data_COMP[221]
  PIN Data_COMP[227]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10902.985 1046.435 10903.265 1047.435 ;
    END
  END Data_COMP[227]
  PIN MASKH[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10901.865 1046.435 10902.145 1047.435 ;
    END
  END MASKH[122]
  PIN DIG_MON_SEL[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10885.625 1046.435 10885.905 1047.435 ;
    END
  END DIG_MON_SEL[244]
  PIN DIG_MON_COMP[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10882.825 1046.435 10883.105 1047.435 ;
    END
  END DIG_MON_COMP[19]
  PIN MASKV[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10881.145 1046.435 10881.425 1047.435 ;
    END
  END MASKV[243]
  PIN Data_COMP[208]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10878.905 1046.435 10879.185 1047.435 ;
    END
  END Data_COMP[208]
  PIN Data_COMP[209]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10877.225 1046.435 10877.505 1047.435 ;
    END
  END Data_COMP[209]
  PIN Data_COMP[196]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10876.105 1046.435 10876.385 1047.435 ;
    END
  END Data_COMP[196]
  PIN BcidMtx[731]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10832.985 1046.435 10833.265 1047.435 ;
    END
  END BcidMtx[731]
  PIN FREEZE_COMP[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10831.305 1046.435 10831.585 1047.435 ;
    END
  END FREEZE_COMP[9]
  PIN BcidMtx[728]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10830.185 1046.435 10830.465 1047.435 ;
    END
  END BcidMtx[728]
  PIN Data_HV[1099]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18786.105 1046.435 18786.385 1047.435 ;
    END
  END Data_HV[1099]
  PIN Data_COMP[198]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10825.705 1046.435 10825.985 1047.435 ;
    END
  END Data_COMP[198]
  PIN Data_COMP[204]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10825.145 1046.435 10825.425 1047.435 ;
    END
  END Data_COMP[204]
  PIN Data_COMP[200]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10822.905 1046.435 10823.185 1047.435 ;
    END
  END Data_COMP[200]
  PIN Data_COMP[206]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10821.225 1046.435 10821.505 1047.435 ;
    END
  END Data_COMP[206]
  PIN MASKH[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10811.705 1046.435 10811.985 1047.435 ;
    END
  END MASKH[121]
  PIN DIG_MON_SEL[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10808.345 1046.435 10808.625 1047.435 ;
    END
  END DIG_MON_SEL[242]
  PIN DIG_MON_COMP[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10805.545 1046.435 10805.825 1047.435 ;
    END
  END DIG_MON_COMP[17]
  PIN MASKV[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10801.905 1046.435 10802.185 1047.435 ;
    END
  END MASKV[241]
  PIN Data_COMP[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10799.665 1046.435 10799.945 1047.435 ;
    END
  END Data_COMP[187]
  PIN Data_COMP[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10772.505 1046.435 10772.785 1047.435 ;
    END
  END Data_COMP[188]
  PIN Data_COMP[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10771.385 1046.435 10771.665 1047.435 ;
    END
  END Data_COMP[175]
  PIN BcidMtx[725]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10767.465 1046.435 10767.745 1047.435 ;
    END
  END BcidMtx[725]
  PIN FREEZE_COMP[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10765.785 1046.435 10766.065 1047.435 ;
    END
  END FREEZE_COMP[8]
  PIN BcidMtx[722]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10764.665 1046.435 10764.945 1047.435 ;
    END
  END BcidMtx[722]
  PIN Data_HV[1098]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18785.545 1046.435 18785.825 1047.435 ;
    END
  END Data_HV[1098]
  PIN Data_COMP[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10760.185 1046.435 10760.465 1047.435 ;
    END
  END Data_COMP[177]
  PIN Data_COMP[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10746.185 1046.435 10746.465 1047.435 ;
    END
  END Data_COMP[178]
  PIN Data_HV[1054]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18585.625 1046.435 18585.905 1047.435 ;
    END
  END Data_HV[1054]
  PIN Data_COMP[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10743.385 1046.435 10743.665 1047.435 ;
    END
  END Data_COMP[168]
  PIN MASKV[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10742.265 1046.435 10742.545 1047.435 ;
    END
  END MASKV[240]
  PIN MASKD[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10736.665 1046.435 10736.945 1047.435 ;
    END
  END MASKD[239]
  PIN INJ_ROW[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10734.425 1046.435 10734.705 1047.435 ;
    END
  END INJ_ROW[119]
  PIN Data_COMP[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10692.425 1046.435 10692.705 1047.435 ;
    END
  END Data_COMP[159]
  PIN Data_COMP[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10690.745 1046.435 10691.025 1047.435 ;
    END
  END Data_COMP[160]
  PIN Data_COMP[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10689.625 1046.435 10689.905 1047.435 ;
    END
  END Data_COMP[161]
  PIN nTOK_COMP[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10686.265 1046.435 10686.545 1047.435 ;
    END
  END nTOK_COMP[7]
  PIN BcidMtx[717]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10684.025 1046.435 10684.305 1047.435 ;
    END
  END BcidMtx[717]
  PIN Read_COMP[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10682.905 1046.435 10683.185 1047.435 ;
    END
  END Read_COMP[7]
  PIN INJ_IN[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10671.705 1046.435 10671.985 1047.435 ;
    END
  END INJ_IN[238]
  PIN Data_COMP[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10669.465 1046.435 10669.745 1047.435 ;
    END
  END Data_COMP[156]
  PIN Data_COMP[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10668.345 1046.435 10668.625 1047.435 ;
    END
  END Data_COMP[157]
  PIN Data_PMOS[1046]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9544.985 1046.435 9545.265 1047.435 ;
    END
  END Data_PMOS[1046]
  PIN Data_HV[1100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18790.025 1046.435 18790.305 1047.435 ;
    END
  END Data_HV[1100]
  PIN FREEZE_PMOS[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9793.065 1046.435 9793.345 1047.435 ;
    END
  END FREEZE_PMOS[52]
  PIN DIG_MON_SEL[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10631.945 1046.435 10632.225 1047.435 ;
    END
  END DIG_MON_SEL[237]
  PIN Data_COMP[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10627.465 1046.435 10627.745 1047.435 ;
    END
  END Data_COMP[144]
  PIN Data_COMP[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10625.785 1046.435 10626.065 1047.435 ;
    END
  END Data_COMP[145]
  PIN Data_COMP[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10624.665 1046.435 10624.945 1047.435 ;
    END
  END Data_COMP[139]
  PIN INJ_IN[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10621.305 1046.435 10621.585 1047.435 ;
    END
  END INJ_IN[237]
  PIN BcidMtx[713]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10605.625 1046.435 10605.905 1047.435 ;
    END
  END BcidMtx[713]
  PIN BcidMtx[711]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10604.505 1046.435 10604.785 1047.435 ;
    END
  END BcidMtx[711]
  PIN BcidMtx[708]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10601.705 1046.435 10601.985 1047.435 ;
    END
  END BcidMtx[708]
  PIN Data_COMP[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10599.465 1046.435 10599.745 1047.435 ;
    END
  END Data_COMP[129]
  PIN Data_COMP[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10598.345 1046.435 10598.625 1047.435 ;
    END
  END Data_COMP[135]
  PIN Data_COMP[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10595.545 1046.435 10595.825 1047.435 ;
    END
  END Data_COMP[137]
  PIN Data_COMP[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10594.425 1046.435 10594.705 1047.435 ;
    END
  END Data_COMP[126]
  PIN MASKV[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10554.665 1046.435 10554.945 1047.435 ;
    END
  END MASKV[236]
  PIN DIG_MON_SEL[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10550.745 1046.435 10551.025 1047.435 ;
    END
  END DIG_MON_SEL[236]
  PIN Data_HV[1104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18789.465 1046.435 18789.745 1047.435 ;
    END
  END Data_HV[1104]
  PIN DIG_MON_COMP[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10547.945 1046.435 10548.225 1047.435 ;
    END
  END DIG_MON_COMP[11]
  PIN Data_COMP[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10544.585 1046.435 10544.865 1047.435 ;
    END
  END Data_COMP[117]
  PIN Data_COMP[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10543.465 1046.435 10543.745 1047.435 ;
    END
  END Data_COMP[110]
  PIN Data_COMP[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10542.345 1046.435 10542.625 1047.435 ;
    END
  END Data_COMP[125]
  PIN nTOK_COMP[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10530.025 1046.435 10530.305 1047.435 ;
    END
  END nTOK_COMP[5]
  PIN BcidMtx[706]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10528.345 1046.435 10528.625 1047.435 ;
    END
  END BcidMtx[706]
  PIN FREEZE_COMP[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10527.225 1046.435 10527.505 1047.435 ;
    END
  END FREEZE_COMP[5]
  PIN INJ_IN[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10521.905 1046.435 10522.185 1047.435 ;
    END
  END INJ_IN[234]
  PIN Data_COMP[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10520.225 1046.435 10520.505 1047.435 ;
    END
  END Data_COMP[107]
  PIN Data_COMP[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10519.105 1046.435 10519.385 1047.435 ;
    END
  END Data_COMP[120]
  PIN Data_COMP[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10490.825 1046.435 10491.105 1047.435 ;
    END
  END Data_COMP[106]
  PIN Data_COMP[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10489.705 1046.435 10489.985 1047.435 ;
    END
  END Data_COMP[122]
  PIN MASKH[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10488.585 1046.435 10488.865 1047.435 ;
    END
  END MASKH[117]
  PIN DIG_MON_SEL[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10484.665 1046.435 10484.945 1047.435 ;
    END
  END DIG_MON_SEL[233]
  PIN INJ_ROW[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10481.305 1046.435 10481.585 1047.435 ;
    END
  END INJ_ROW[116]
  PIN Data_COMP[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10480.185 1046.435 10480.465 1047.435 ;
    END
  END Data_COMP[102]
  PIN Data_COMP[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10465.065 1046.435 10465.345 1047.435 ;
    END
  END Data_COMP[89]
  PIN Data_COMP[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10463.385 1046.435 10463.665 1047.435 ;
    END
  END Data_COMP[98]
  PIN Data_COMP[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10462.265 1046.435 10462.545 1047.435 ;
    END
  END Data_COMP[90]
  PIN BcidMtx[699]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10457.785 1046.435 10458.065 1047.435 ;
    END
  END BcidMtx[699]
  PIN Read_COMP[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10456.665 1046.435 10456.945 1047.435 ;
    END
  END Read_COMP[4]
  PIN BcidMtx[697]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10455.545 1046.435 10455.825 1047.435 ;
    END
  END BcidMtx[697]
  PIN Data_COMP[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10412.985 1046.435 10413.265 1047.435 ;
    END
  END Data_COMP[93]
  PIN Data_COMP[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10411.865 1046.435 10412.145 1047.435 ;
    END
  END Data_COMP[94]
  PIN Data_COMP[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10410.745 1046.435 10411.025 1047.435 ;
    END
  END Data_COMP[100]
  PIN MASKV[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10407.945 1046.435 10408.225 1047.435 ;
    END
  END MASKV[232]
  PIN MASKD[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10406.825 1046.435 10407.105 1047.435 ;
    END
  END MASKD[232]
  PIN INJ_ROW[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10391.705 1046.435 10391.985 1047.435 ;
    END
  END INJ_ROW[115]
  PIN Data_COMP[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10390.585 1046.435 10390.865 1047.435 ;
    END
  END Data_COMP[81]
  PIN Data_COMP[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10389.465 1046.435 10389.745 1047.435 ;
    END
  END Data_COMP[75]
  PIN Data_COMP[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10386.665 1046.435 10386.945 1047.435 ;
    END
  END Data_COMP[77]
  PIN Data_COMP[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10385.545 1046.435 10385.825 1047.435 ;
    END
  END Data_COMP[69]
  PIN nTOK_COMP[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10381.345 1046.435 10381.625 1047.435 ;
    END
  END nTOK_COMP[3]
  PIN BcidMtx[692]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10351.945 1046.435 10352.225 1047.435 ;
    END
  END BcidMtx[692]
  PIN BcidMtx[690]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10350.825 1046.435 10351.105 1047.435 ;
    END
  END BcidMtx[690]
  PIN Data_COMP[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10348.585 1046.435 10348.865 1047.435 ;
    END
  END Data_COMP[66]
  PIN INJ_ROW[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18791.705 1046.435 18791.985 1047.435 ;
    END
  END INJ_ROW[220]
  PIN Data_COMP[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10345.225 1046.435 10345.505 1047.435 ;
    END
  END Data_COMP[79]
  PIN Data_COMP[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10344.105 1046.435 10344.385 1047.435 ;
    END
  END Data_COMP[64]
  PIN MASKD[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10341.305 1046.435 10341.585 1047.435 ;
    END
  END MASKD[230]
  PIN DIG_MON_SEL[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10325.065 1046.435 10325.345 1047.435 ;
    END
  END DIG_MON_SEL[229]
  PIN Data_COMP[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10320.585 1046.435 10320.865 1047.435 ;
    END
  END Data_COMP[60]
  PIN Data_COMP[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10319.465 1046.435 10319.745 1047.435 ;
    END
  END Data_COMP[54]
  PIN Data_COMP[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10318.345 1046.435 10318.625 1047.435 ;
    END
  END Data_COMP[47]
  PIN Data_COMP[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10315.545 1046.435 10315.825 1047.435 ;
    END
  END Data_COMP[48]
  PIN nTOK_COMP[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10274.105 1046.435 10274.385 1047.435 ;
    END
  END nTOK_COMP[2]
  PIN BcidMtx[688]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10272.425 1046.435 10272.705 1047.435 ;
    END
  END BcidMtx[688]
  PIN BcidMtx[685]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10269.625 1046.435 10269.905 1047.435 ;
    END
  END BcidMtx[685]
  PIN Data_COMP[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10266.825 1046.435 10267.105 1047.435 ;
    END
  END Data_COMP[45]
  PIN Data_COMP[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10265.145 1046.435 10265.425 1047.435 ;
    END
  END Data_COMP[57]
  PIN Data_COMP[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10263.465 1046.435 10263.745 1047.435 ;
    END
  END Data_COMP[58]
  PIN Data_COMP[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10262.345 1046.435 10262.625 1047.435 ;
    END
  END Data_COMP[43]
  PIN Data_HV[1105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18787.785 1046.435 18788.065 1047.435 ;
    END
  END Data_HV[1105]
  PIN MASKD[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10251.145 1046.435 10251.425 1047.435 ;
    END
  END MASKD[228]
  PIN DIG_MON_SEL[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10248.345 1046.435 10248.625 1047.435 ;
    END
  END DIG_MON_SEL[228]
  PIN DIG_MON_COMP[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10245.545 1046.435 10245.825 1047.435 ;
    END
  END DIG_MON_COMP[3]
  PIN Data_COMP[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10241.345 1046.435 10241.625 1047.435 ;
    END
  END Data_COMP[39]
  PIN Data_COMP[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10239.665 1046.435 10239.945 1047.435 ;
    END
  END Data_COMP[40]
  PIN Data_COMP[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10212.505 1046.435 10212.785 1047.435 ;
    END
  END Data_COMP[41]
  PIN Data_COMP[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10210.825 1046.435 10211.105 1047.435 ;
    END
  END Data_COMP[27]
  PIN BcidMtx[681]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10206.345 1046.435 10206.625 1047.435 ;
    END
  END BcidMtx[681]
  PIN BcidMtx[680]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10204.665 1046.435 10204.945 1047.435 ;
    END
  END BcidMtx[680]
  PIN BcidMtx[678]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10203.545 1046.435 10203.825 1047.435 ;
    END
  END BcidMtx[678]
  PIN Data_COMP[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10200.185 1046.435 10200.465 1047.435 ;
    END
  END Data_COMP[30]
  PIN Data_COMP[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10185.625 1046.435 10185.905 1047.435 ;
    END
  END Data_COMP[25]
  PIN Data_HV[1097]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18788.345 1046.435 18788.625 1047.435 ;
    END
  END Data_HV[1097]
  PIN Data_COMP[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10182.825 1046.435 10183.105 1047.435 ;
    END
  END Data_COMP[38]
  PIN MASKD[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10181.145 1046.435 10181.425 1047.435 ;
    END
  END MASKD[226]
  PIN DIG_MON_COMP[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10180.025 1046.435 10180.305 1047.435 ;
    END
  END DIG_MON_COMP[2]
  PIN MASKD[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10176.665 1046.435 10176.945 1047.435 ;
    END
  END MASKD[225]
  PIN MASKV[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10173.865 1046.435 10174.145 1047.435 ;
    END
  END MASKV[225]
  PIN Data_COMP[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10132.985 1046.435 10133.265 1047.435 ;
    END
  END Data_COMP[8]
  PIN Data_COMP[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10130.745 1046.435 10131.025 1047.435 ;
    END
  END Data_COMP[13]
  PIN Data_COMP[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10129.065 1046.435 10129.345 1047.435 ;
    END
  END Data_COMP[7]
  PIN INJ_IN[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10127.385 1046.435 10127.665 1047.435 ;
    END
  END INJ_IN[225]
  PIN BcidMtx[677]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10125.145 1046.435 10125.425 1047.435 ;
    END
  END BcidMtx[677]
  PIN FREEZE_COMP[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10123.465 1046.435 10123.745 1047.435 ;
    END
  END FREEZE_COMP[0]
  PIN BcidMtx[673]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10121.785 1046.435 10122.065 1047.435 ;
    END
  END BcidMtx[673]
  PIN Data_COMP[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10110.585 1046.435 10110.865 1047.435 ;
    END
  END Data_COMP[3]
  PIN Data_COMP[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10108.905 1046.435 10109.185 1047.435 ;
    END
  END Data_COMP[15]
  PIN Data_COMP[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10107.225 1046.435 10107.505 1047.435 ;
    END
  END Data_COMP[16]
  PIN Data_COMP[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10105.545 1046.435 10105.825 1047.435 ;
    END
  END Data_COMP[0]
  PIN BcidMtx[1220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17402.345 1046.435 17402.625 1047.435 ;
    END
  END BcidMtx[1220]
  PIN INJ_IN[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17391.705 1046.435 17391.985 1047.435 ;
    END
  END INJ_IN[406]
  PIN Data_HV[737]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17390.025 1046.435 17390.305 1047.435 ;
    END
  END Data_HV[737]
  PIN Data_HV[739]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17387.785 1046.435 17388.065 1047.435 ;
    END
  END Data_HV[739]
  PIN Data_HV[736]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17386.105 1046.435 17386.385 1047.435 ;
    END
  END Data_HV[736]
  PIN Data_HV[752]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17384.985 1046.435 17385.265 1047.435 ;
    END
  END Data_HV[752]
  PIN DIG_MON_HV[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17380.225 1046.435 17380.505 1047.435 ;
    END
  END DIG_MON_HV[70]
  PIN FREEZE_HV[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17633.065 1046.435 17633.345 1047.435 ;
    END
  END FREEZE_HV[38]
  PIN MASKD[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18470.825 1046.435 18471.105 1047.435 ;
    END
  END MASKD[433]
  PIN Data_HV[1026]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18467.465 1046.435 18467.745 1047.435 ;
    END
  END Data_HV[1026]
  PIN Data_HV[1027]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18465.785 1046.435 18466.065 1047.435 ;
    END
  END Data_HV[1027]
  PIN Data_HV[1028]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18464.105 1046.435 18464.385 1047.435 ;
    END
  END Data_HV[1028]
  PIN Data_HV[1014]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18462.425 1046.435 18462.705 1047.435 ;
    END
  END Data_HV[1014]
  PIN BcidMtx[1301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18445.625 1046.435 18445.905 1047.435 ;
    END
  END BcidMtx[1301]
  PIN FREEZE_HV[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18443.945 1046.435 18444.225 1047.435 ;
    END
  END FREEZE_HV[48]
  PIN BcidMtx[1297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18442.265 1046.435 18442.545 1047.435 ;
    END
  END BcidMtx[1297]
  PIN Data_HV[1011]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18439.465 1046.435 18439.745 1047.435 ;
    END
  END Data_HV[1011]
  PIN Data_HV[1023]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18437.785 1046.435 18438.065 1047.435 ;
    END
  END Data_HV[1023]
  PIN Data_HV[1024]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18436.105 1046.435 18436.385 1047.435 ;
    END
  END Data_HV[1024]
  PIN Data_HV[1008]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18434.425 1046.435 18434.705 1047.435 ;
    END
  END Data_HV[1008]
  PIN MASKH[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18394.105 1046.435 18394.385 1047.435 ;
    END
  END MASKH[216]
  PIN MASKD[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18389.065 1046.435 18389.345 1047.435 ;
    END
  END MASKD[431]
  PIN MASKV[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18386.265 1046.435 18386.545 1047.435 ;
    END
  END MASKV[431]
  PIN Data_HV[999]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18384.585 1046.435 18384.865 1047.435 ;
    END
  END Data_HV[999]
  PIN Data_HV[1000]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18382.905 1046.435 18383.185 1047.435 ;
    END
  END Data_HV[1000]
  PIN Data_HV[994]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18381.225 1046.435 18381.505 1047.435 ;
    END
  END Data_HV[994]
  PIN nTOK_HV[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18370.025 1046.435 18370.305 1047.435 ;
    END
  END nTOK_HV[47]
  PIN BcidMtx[1293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18367.785 1046.435 18368.065 1047.435 ;
    END
  END BcidMtx[1293]
  PIN BcidMtx[1292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18366.105 1046.435 18366.385 1047.435 ;
    END
  END BcidMtx[1292]
  PIN INJ_IN[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18361.905 1046.435 18362.185 1047.435 ;
    END
  END INJ_IN[430]
  PIN Data_HV[996]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18359.665 1046.435 18359.945 1047.435 ;
    END
  END Data_HV[996]
  PIN Data_HV[991]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18332.505 1046.435 18332.785 1047.435 ;
    END
  END Data_HV[991]
  PIN Data_HV[988]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18330.825 1046.435 18331.105 1047.435 ;
    END
  END Data_HV[988]
  PIN MASKV[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18329.145 1046.435 18329.425 1047.435 ;
    END
  END MASKV[430]
  PIN DIG_MON_HV[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18326.905 1046.435 18327.185 1047.435 ;
    END
  END DIG_MON_HV[94]
  PIN DIG_MON_SEL[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18324.665 1046.435 18324.945 1047.435 ;
    END
  END DIG_MON_SEL[429]
  PIN INJ_ROW[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18321.305 1046.435 18321.585 1047.435 ;
    END
  END INJ_ROW[214]
  PIN Data_HV[974]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18319.625 1046.435 18319.905 1047.435 ;
    END
  END Data_HV[974]
  PIN Data_HV[971]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18305.065 1046.435 18305.345 1047.435 ;
    END
  END Data_HV[971]
  PIN Data_HV[980]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18303.385 1046.435 18303.665 1047.435 ;
    END
  END Data_HV[980]
  PIN INJ_IN[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18301.145 1046.435 18301.425 1047.435 ;
    END
  END INJ_IN[429]
  PIN BcidMtx[1287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18297.785 1046.435 18298.065 1047.435 ;
    END
  END BcidMtx[1287]
  PIN BcidMtx[1286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18296.105 1046.435 18296.385 1047.435 ;
    END
  END BcidMtx[1286]
  PIN BcidMtx[1284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18294.985 1046.435 18295.265 1047.435 ;
    END
  END BcidMtx[1284]
  PIN Data_HV[975]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18252.985 1046.435 18253.265 1047.435 ;
    END
  END Data_HV[975]
  PIN Data_HV[970]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18251.305 1046.435 18251.585 1047.435 ;
    END
  END Data_HV[970]
  PIN Data_HV[977]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18250.185 1046.435 18250.465 1047.435 ;
    END
  END Data_HV[977]
  PIN MASKV[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18247.945 1046.435 18248.225 1047.435 ;
    END
  END MASKV[428]
  PIN MASKD[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18246.825 1046.435 18247.105 1047.435 ;
    END
  END MASKD[428]
  PIN DIG_MON_HV[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18245.705 1046.435 18245.985 1047.435 ;
    END
  END DIG_MON_HV[92]
  PIN MASKD[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18242.345 1046.435 18242.625 1047.435 ;
    END
  END MASKD[427]
  PIN MASKV[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18231.145 1046.435 18231.425 1047.435 ;
    END
  END MASKV[427]
  PIN Data_HV[953]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18230.025 1046.435 18230.305 1047.435 ;
    END
  END Data_HV[953]
  PIN Data_HV[958]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18227.785 1046.435 18228.065 1047.435 ;
    END
  END Data_HV[958]
  PIN Data_HV[952]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18226.105 1046.435 18226.385 1047.435 ;
    END
  END Data_HV[952]
  PIN INJ_IN[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18222.465 1046.435 18222.745 1047.435 ;
    END
  END INJ_IN[427]
  PIN BcidMtx[1281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18219.105 1046.435 18219.385 1047.435 ;
    END
  END BcidMtx[1281]
  PIN BcidMtx[1279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18191.385 1046.435 18191.665 1047.435 ;
    END
  END BcidMtx[1279]
  PIN INJ_IN[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18189.705 1046.435 18189.985 1047.435 ;
    END
  END INJ_IN[426]
  PIN Data_HV[955]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18186.345 1046.435 18186.625 1047.435 ;
    END
  END Data_HV[955]
  PIN Data_HV[956]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18184.665 1046.435 18184.945 1047.435 ;
    END
  END Data_HV[956]
  PIN Data_HV[945]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18183.545 1046.435 18183.825 1047.435 ;
    END
  END Data_HV[945]
  PIN DIG_MON_HV[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18180.185 1046.435 18180.465 1047.435 ;
    END
  END DIG_MON_HV[90]
  PIN Data_HV[1073]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18666.265 1046.435 18666.545 1047.435 ;
    END
  END Data_HV[1073]
  PIN DIG_MON_SEL[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18165.065 1046.435 18165.345 1047.435 ;
    END
  END DIG_MON_SEL[425]
  PIN MASKV[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18161.145 1046.435 18161.425 1047.435 ;
    END
  END MASKV[425]
  PIN Data_HV[936]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18159.465 1046.435 18159.745 1047.435 ;
    END
  END Data_HV[936]
  PIN Data_HV[943]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18158.905 1046.435 18159.185 1047.435 ;
    END
  END Data_HV[943]
  PIN Data_HV[931]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18156.105 1046.435 18156.385 1047.435 ;
    END
  END Data_HV[931]
  PIN nTOK_HV[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18114.105 1046.435 18114.385 1047.435 ;
    END
  END nTOK_HV[44]
  PIN BcidMtx[1277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18112.985 1046.435 18113.265 1047.435 ;
    END
  END BcidMtx[1277]
  PIN BcidMtx[1274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18110.185 1046.435 18110.465 1047.435 ;
    END
  END BcidMtx[1274]
  PIN INJ_IN[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18107.945 1046.435 18108.225 1047.435 ;
    END
  END INJ_IN[424]
  PIN Data_HV[927]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18106.825 1046.435 18107.105 1047.435 ;
    END
  END Data_HV[927]
  PIN Data_HV[928]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18104.025 1046.435 18104.305 1047.435 ;
    END
  END Data_HV[928]
  PIN Data_HV[925]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18102.345 1046.435 18102.625 1047.435 ;
    END
  END Data_HV[925]
  PIN Data_HV[924]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18101.785 1046.435 18102.065 1047.435 ;
    END
  END Data_HV[924]
  PIN Data_HV[1080]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18665.705 1046.435 18665.985 1047.435 ;
    END
  END Data_HV[1080]
  PIN DIG_MON_SEL[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18088.345 1046.435 18088.625 1047.435 ;
    END
  END DIG_MON_SEL[424]
  PIN DIG_MON_SEL[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18087.785 1046.435 18088.065 1047.435 ;
    END
  END DIG_MON_SEL[423]
  PIN MASKV[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18081.905 1046.435 18082.185 1047.435 ;
    END
  END MASKV[423]
  PIN Data_HV[915]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18080.225 1046.435 18080.505 1047.435 ;
    END
  END Data_HV[915]
  PIN Data_HV[908]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18079.105 1046.435 18079.385 1047.435 ;
    END
  END Data_HV[908]
  PIN Data_HV[909]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18050.825 1046.435 18051.105 1047.435 ;
    END
  END Data_HV[909]
  PIN nTOK_HV[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18048.585 1046.435 18048.865 1047.435 ;
    END
  END nTOK_HV[43]
  PIN BcidMtx[1270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18046.905 1046.435 18047.185 1047.435 ;
    END
  END BcidMtx[1270]
  PIN BcidMtx[1267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18044.105 1046.435 18044.385 1047.435 ;
    END
  END BcidMtx[1267]
  PIN Data_HV[906]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18041.305 1046.435 18041.585 1047.435 ;
    END
  END Data_HV[906]
  PIN Data_HV[912]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18040.185 1046.435 18040.465 1047.435 ;
    END
  END Data_HV[912]
  PIN Data_HV[919]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18025.065 1046.435 18025.345 1047.435 ;
    END
  END Data_HV[919]
  PIN Data_HV[903]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18023.385 1046.435 18023.665 1047.435 ;
    END
  END Data_HV[903]
  PIN MASKV[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18022.265 1046.435 18022.545 1047.435 ;
    END
  END MASKV[422]
  PIN DIG_MON_SEL[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18017.785 1046.435 18018.065 1047.435 ;
    END
  END DIG_MON_SEL[421]
  PIN DIG_MON_HV[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18015.545 1046.435 18015.825 1047.435 ;
    END
  END DIG_MON_HV[85]
  PIN Data_HV[890]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17972.985 1046.435 17973.265 1047.435 ;
    END
  END Data_HV[890]
  PIN Data_HV[887]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17971.305 1046.435 17971.585 1047.435 ;
    END
  END Data_HV[887]
  PIN Data_HV[902]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17970.185 1046.435 17970.465 1047.435 ;
    END
  END Data_HV[902]
  PIN INJ_IN[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17967.385 1046.435 17967.665 1047.435 ;
    END
  END INJ_IN[421]
  PIN BcidMtx[1264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17964.585 1046.435 17964.865 1047.435 ;
    END
  END BcidMtx[1264]
  PIN FREEZE_HV[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17963.465 1046.435 17963.745 1047.435 ;
    END
  END FREEZE_HV[42]
  PIN BcidMtx[1176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16841.225 1046.435 16841.505 1047.435 ;
    END
  END BcidMtx[1176]
  PIN Data_HV[590]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16830.025 1046.435 16830.305 1047.435 ;
    END
  END Data_HV[590]
  PIN Data_HV[603]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16828.905 1046.435 16829.185 1047.435 ;
    END
  END Data_HV[603]
  PIN Data_HV[599]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16826.665 1046.435 16826.945 1047.435 ;
    END
  END Data_HV[599]
  PIN Data_HV[605]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16824.985 1046.435 16825.265 1047.435 ;
    END
  END Data_HV[605]
  PIN MASKH[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16821.905 1046.435 16822.185 1047.435 ;
    END
  END MASKH[196]
  PIN DIG_MON_SEL[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16818.545 1046.435 16818.825 1047.435 ;
    END
  END DIG_MON_SEL[392]
  PIN MASKD[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17910.825 1046.435 17911.105 1047.435 ;
    END
  END MASKD[419]
  PIN INJ_ROW[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17908.585 1046.435 17908.865 1047.435 ;
    END
  END INJ_ROW[209]
  PIN Data_HV[873]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17906.345 1046.435 17906.625 1047.435 ;
    END
  END Data_HV[873]
  PIN Data_HV[874]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17904.665 1046.435 17904.945 1047.435 ;
    END
  END Data_HV[874]
  PIN Data_HV[875]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17903.545 1046.435 17903.825 1047.435 ;
    END
  END Data_HV[875]
  PIN INJ_IN[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17901.305 1046.435 17901.585 1047.435 ;
    END
  END INJ_IN[419]
  PIN BcidMtx[1258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17885.065 1046.435 17885.345 1047.435 ;
    END
  END BcidMtx[1258]
  PIN FREEZE_HV[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17883.945 1046.435 17884.225 1047.435 ;
    END
  END FREEZE_HV[41]
  PIN BcidMtx[1254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17881.705 1046.435 17881.985 1047.435 ;
    END
  END BcidMtx[1254]
  PIN Data_HV[863]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17878.905 1046.435 17879.185 1047.435 ;
    END
  END Data_HV[863]
  PIN Data_HV[876]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17877.785 1046.435 17878.065 1047.435 ;
    END
  END Data_HV[876]
  PIN Data_HV[872]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17875.545 1046.435 17875.825 1047.435 ;
    END
  END Data_HV[872]
  PIN Data_HV[878]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17873.865 1046.435 17874.145 1047.435 ;
    END
  END Data_HV[878]
  PIN MASKH[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17834.105 1046.435 17834.385 1047.435 ;
    END
  END MASKH[209]
  PIN DIG_MON_SEL[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17830.745 1046.435 17831.025 1047.435 ;
    END
  END DIG_MON_SEL[418]
  PIN DIG_MON_HV[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17827.945 1046.435 17828.225 1047.435 ;
    END
  END DIG_MON_HV[81]
  PIN MASKV[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17826.265 1046.435 17826.545 1047.435 ;
    END
  END MASKV[417]
  PIN Data_HV[859]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17824.025 1046.435 17824.305 1047.435 ;
    END
  END Data_HV[859]
  PIN Data_HV[860]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17822.345 1046.435 17822.625 1047.435 ;
    END
  END Data_HV[860]
  PIN Data_HV[847]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17821.225 1046.435 17821.505 1047.435 ;
    END
  END Data_HV[847]
  PIN BcidMtx[1253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17808.905 1046.435 17809.185 1047.435 ;
    END
  END BcidMtx[1253]
  PIN FREEZE_HV[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17807.225 1046.435 17807.505 1047.435 ;
    END
  END FREEZE_HV[40]
  PIN BcidMtx[1250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17806.105 1046.435 17806.385 1047.435 ;
    END
  END BcidMtx[1250]
  PIN Data_HV[843]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17800.785 1046.435 17801.065 1047.435 ;
    END
  END Data_HV[843]
  PIN Data_HV[855]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17799.105 1046.435 17799.385 1047.435 ;
    END
  END Data_HV[855]
  PIN Data_HV[844]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17772.505 1046.435 17772.785 1047.435 ;
    END
  END Data_HV[844]
  PIN Data_HV[840]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17770.265 1046.435 17770.545 1047.435 ;
    END
  END Data_HV[840]
  PIN MASKH[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17768.585 1046.435 17768.865 1047.435 ;
    END
  END MASKH[208]
  PIN DIG_MON_HV[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17766.905 1046.435 17767.185 1047.435 ;
    END
  END DIG_MON_HV[80]
  PIN DIG_MON_SEL[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17764.665 1046.435 17764.945 1047.435 ;
    END
  END DIG_MON_SEL[415]
  PIN INJ_ROW[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17761.305 1046.435 17761.585 1047.435 ;
    END
  END INJ_ROW[207]
  PIN Data_HV[837]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17760.185 1046.435 17760.465 1047.435 ;
    END
  END Data_HV[837]
  PIN Data_HV[824]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17745.065 1046.435 17745.345 1047.435 ;
    END
  END Data_HV[824]
  PIN Data_HV[833]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17743.385 1046.435 17743.665 1047.435 ;
    END
  END Data_HV[833]
  PIN Data_HV[825]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17742.265 1046.435 17742.545 1047.435 ;
    END
  END Data_HV[825]
  PIN BcidMtx[1246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17738.345 1046.435 17738.625 1047.435 ;
    END
  END BcidMtx[1246]
  PIN Read_HV[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17736.665 1046.435 17736.945 1047.435 ;
    END
  END Read_HV[39]
  PIN BcidMtx[1243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17735.545 1046.435 17735.825 1047.435 ;
    END
  END BcidMtx[1243]
  PIN Data_HV[821]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17693.545 1046.435 17693.825 1047.435 ;
    END
  END Data_HV[821]
  PIN Data_HV[829]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17691.865 1046.435 17692.145 1047.435 ;
    END
  END Data_HV[829]
  PIN Data_HV[835]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17690.745 1046.435 17691.025 1047.435 ;
    END
  END Data_HV[835]
  PIN Data_HV[836]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17688.505 1046.435 17688.785 1047.435 ;
    END
  END Data_HV[836]
  PIN MASKD[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17686.825 1046.435 17687.105 1047.435 ;
    END
  END MASKD[414]
  PIN BcidMtx[1315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18669.625 1046.435 18669.905 1047.435 ;
    END
  END BcidMtx[1315]
  PIN INJ_ROW[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17671.705 1046.435 17671.985 1047.435 ;
    END
  END INJ_ROW[206]
  PIN Data_HV[816]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17670.585 1046.435 17670.865 1047.435 ;
    END
  END Data_HV[816]
  PIN Data_HV[803]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17668.345 1046.435 17668.625 1047.435 ;
    END
  END Data_HV[803]
  PIN Data_HV[812]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17666.665 1046.435 17666.945 1047.435 ;
    END
  END Data_HV[812]
  PIN Data_HV[804]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17665.545 1046.435 17665.825 1047.435 ;
    END
  END Data_HV[804]
  PIN BcidMtx[1240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17659.665 1046.435 17659.945 1047.435 ;
    END
  END BcidMtx[1240]
  PIN BcidMtx[1238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17631.945 1046.435 17632.225 1047.435 ;
    END
  END BcidMtx[1238]
  PIN BcidMtx[1236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17630.825 1046.435 17631.105 1047.435 ;
    END
  END BcidMtx[1236]
  PIN Data_HV[807]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17627.465 1046.435 17627.745 1047.435 ;
    END
  END Data_HV[807]
  PIN Data_HV[802]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17625.785 1046.435 17626.065 1047.435 ;
    END
  END Data_HV[802]
  PIN Data_HV[809]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17624.665 1046.435 17624.945 1047.435 ;
    END
  END Data_HV[809]
  PIN MASKV[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17622.425 1046.435 17622.705 1047.435 ;
    END
  END MASKV[412]
  PIN DIG_MON_HV[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17620.185 1046.435 17620.465 1047.435 ;
    END
  END DIG_MON_HV[76]
  PIN DIG_MON_SEL[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17605.625 1046.435 17605.905 1047.435 ;
    END
  END DIG_MON_SEL[412]
  PIN DIG_MON_HV[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17602.825 1046.435 17603.105 1047.435 ;
    END
  END DIG_MON_HV[75]
  PIN INJ_ROW[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17601.705 1046.435 17601.985 1047.435 ;
    END
  END INJ_ROW[205]
  PIN Data_HV[795]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17600.585 1046.435 17600.865 1047.435 ;
    END
  END Data_HV[795]
  PIN Data_HV[782]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17598.345 1046.435 17598.625 1047.435 ;
    END
  END Data_HV[782]
  PIN Data_HV[791]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17596.665 1046.435 17596.945 1047.435 ;
    END
  END Data_HV[791]
  PIN INJ_IN[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17594.425 1046.435 17594.705 1047.435 ;
    END
  END INJ_IN[411]
  PIN BcidMtx[1234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17552.425 1046.435 17552.705 1047.435 ;
    END
  END BcidMtx[1234]
  PIN Read_HV[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17550.745 1046.435 17551.025 1047.435 ;
    END
  END Read_HV[37]
  PIN BcidMtx[1231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17549.625 1046.435 17549.905 1047.435 ;
    END
  END BcidMtx[1231]
  PIN Data_HV[779]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17546.265 1046.435 17546.545 1047.435 ;
    END
  END Data_HV[779]
  PIN Data_HV[787]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17544.585 1046.435 17544.865 1047.435 ;
    END
  END Data_HV[787]
  PIN Data_HV[793]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17543.465 1046.435 17543.745 1047.435 ;
    END
  END Data_HV[793]
  PIN Data_HV[794]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17541.225 1046.435 17541.505 1047.435 ;
    END
  END Data_HV[794]
  PIN MASKD[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17531.145 1046.435 17531.425 1047.435 ;
    END
  END MASKD[410]
  PIN DIG_MON_HV[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17525.545 1046.435 17525.825 1047.435 ;
    END
  END DIG_MON_HV[73]
  PIN Data_HV[774]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17521.345 1046.435 17521.625 1047.435 ;
    END
  END Data_HV[774]
  PIN Data_HV[768]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17520.225 1046.435 17520.505 1047.435 ;
    END
  END Data_HV[768]
  PIN Data_HV[776]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17492.505 1046.435 17492.785 1047.435 ;
    END
  END Data_HV[776]
  PIN Data_HV[762]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17490.825 1046.435 17491.105 1047.435 ;
    END
  END Data_HV[762]
  PIN nTOK_HV[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17488.585 1046.435 17488.865 1047.435 ;
    END
  END nTOK_HV[36]
  PIN FREEZE_HV[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17485.785 1046.435 17486.065 1047.435 ;
    END
  END FREEZE_HV[36]
  PIN BcidMtx[1225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17484.105 1046.435 17484.385 1047.435 ;
    END
  END BcidMtx[1225]
  PIN INJ_IN[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17482.425 1046.435 17482.705 1047.435 ;
    END
  END INJ_IN[408]
  PIN Data_HV[771]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17466.745 1046.435 17467.025 1047.435 ;
    END
  END Data_HV[771]
  PIN Data_HV[772]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17465.065 1046.435 17465.345 1047.435 ;
    END
  END Data_HV[772]
  PIN Data_HV[757]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17463.945 1046.435 17464.225 1047.435 ;
    END
  END Data_HV[757]
  PIN MASKH[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17461.705 1046.435 17461.985 1047.435 ;
    END
  END MASKH[204]
  PIN DIG_MON_SEL[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17457.785 1046.435 17458.065 1047.435 ;
    END
  END DIG_MON_SEL[407]
  PIN MASKV[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17453.865 1046.435 17454.145 1047.435 ;
    END
  END MASKV[407]
  PIN Data_HV[747]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17412.425 1046.435 17412.705 1047.435 ;
    END
  END Data_HV[747]
  PIN Data_HV[740]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17411.305 1046.435 17411.585 1047.435 ;
    END
  END Data_HV[740]
  PIN Data_HV[742]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17409.065 1046.435 17409.345 1047.435 ;
    END
  END Data_HV[742]
  PIN nTOK_HV[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17406.265 1046.435 17406.545 1047.435 ;
    END
  END nTOK_HV[35]
  PIN BcidMtx[1222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17404.585 1046.435 17404.865 1047.435 ;
    END
  END BcidMtx[1222]
  PIN Data_COMP[1030]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14026.105 1046.435 14026.385 1047.435 ;
    END
  END Data_COMP[1030]
  PIN MASKD[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14021.345 1046.435 14021.625 1047.435 ;
    END
  END MASKD[322]
  PIN DIG_MON_COMP[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14020.225 1046.435 14020.505 1047.435 ;
    END
  END DIG_MON_COMP[98]
  PIN DIG_MON_SEL[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14018.545 1046.435 14018.825 1047.435 ;
    END
  END DIG_MON_SEL[322]
  PIN MASKD[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15110.825 1046.435 15111.105 1047.435 ;
    END
  END MASKD[349]
  PIN MASKV[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15108.025 1046.435 15108.305 1047.435 ;
    END
  END MASKV[349]
  PIN Data_HV[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15106.345 1046.435 15106.625 1047.435 ;
    END
  END Data_HV[138]
  PIN Data_HV[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15104.665 1046.435 15104.945 1047.435 ;
    END
  END Data_HV[139]
  PIN Data_HV[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15102.985 1046.435 15103.265 1047.435 ;
    END
  END Data_HV[133]
  PIN BcidMtx[1049]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15085.625 1046.435 15085.905 1047.435 ;
    END
  END BcidMtx[1049]
  PIN BcidMtx[1047]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15084.505 1046.435 15084.785 1047.435 ;
    END
  END BcidMtx[1047]
  PIN BcidMtx[1046]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15082.825 1046.435 15083.105 1047.435 ;
    END
  END BcidMtx[1046]
  PIN Data_HV[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15079.465 1046.435 15079.745 1047.435 ;
    END
  END Data_HV[129]
  PIN Data_HV[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15077.785 1046.435 15078.065 1047.435 ;
    END
  END Data_HV[141]
  PIN Data_HV[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15076.665 1046.435 15076.945 1047.435 ;
    END
  END Data_HV[130]
  PIN Data_HV[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15074.425 1046.435 15074.705 1047.435 ;
    END
  END Data_HV[126]
  PIN MASKH[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15034.105 1046.435 15034.385 1047.435 ;
    END
  END MASKH[174]
  PIN DIG_MON_HV[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15032.425 1046.435 15032.705 1047.435 ;
    END
  END DIG_MON_HV[12]
  PIN MASKD[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15029.065 1046.435 15029.345 1047.435 ;
    END
  END MASKD[347]
  PIN MASKV[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15026.265 1046.435 15026.545 1047.435 ;
    END
  END MASKV[347]
  PIN Data_HV[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15024.585 1046.435 15024.865 1047.435 ;
    END
  END Data_HV[117]
  PIN Data_HV[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15022.905 1046.435 15023.185 1047.435 ;
    END
  END Data_HV[118]
  PIN Data_HV[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15021.225 1046.435 15021.505 1047.435 ;
    END
  END Data_HV[112]
  PIN nTOK_HV[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15010.025 1046.435 15010.305 1047.435 ;
    END
  END nTOK_HV[5]
  PIN FREEZE_HV[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15007.225 1046.435 15007.505 1047.435 ;
    END
  END FREEZE_HV[5]
  PIN BcidMtx[1040]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15006.105 1046.435 15006.385 1047.435 ;
    END
  END BcidMtx[1040]
  PIN INJ_IN[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15001.905 1046.435 15002.185 1047.435 ;
    END
  END INJ_IN[346]
  PIN Data_HV[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14999.665 1046.435 14999.945 1047.435 ;
    END
  END Data_HV[114]
  PIN Data_HV[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14972.505 1046.435 14972.785 1047.435 ;
    END
  END Data_HV[109]
  PIN Data_HV[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14970.825 1046.435 14971.105 1047.435 ;
    END
  END Data_HV[106]
  PIN MASKH[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14968.585 1046.435 14968.865 1047.435 ;
    END
  END MASKH[173]
  PIN DIG_MON_HV[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14966.905 1046.435 14967.185 1047.435 ;
    END
  END DIG_MON_HV[10]
  PIN DIG_MON_SEL[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14964.665 1046.435 14964.945 1047.435 ;
    END
  END DIG_MON_SEL[345]
  PIN MASKV[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14960.745 1046.435 14961.025 1047.435 ;
    END
  END MASKV[345]
  PIN Data_HV[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14959.625 1046.435 14959.905 1047.435 ;
    END
  END Data_HV[92]
  PIN Data_HV[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14945.065 1046.435 14945.345 1047.435 ;
    END
  END Data_HV[89]
  PIN Data_HV[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14943.385 1046.435 14943.665 1047.435 ;
    END
  END Data_HV[98]
  PIN INJ_IN[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14941.145 1046.435 14941.425 1047.435 ;
    END
  END INJ_IN[345]
  PIN BcidMtx[1036]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14938.345 1046.435 14938.625 1047.435 ;
    END
  END BcidMtx[1036]
  PIN Read_HV[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14936.665 1046.435 14936.945 1047.435 ;
    END
  END Read_HV[4]
  PIN BcidMtx[1032]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14934.985 1046.435 14935.265 1047.435 ;
    END
  END BcidMtx[1032]
  PIN Data_HV[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14893.545 1046.435 14893.825 1047.435 ;
    END
  END Data_HV[86]
  PIN Data_HV[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14891.865 1046.435 14892.145 1047.435 ;
    END
  END Data_HV[94]
  PIN Data_HV[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14890.745 1046.435 14891.025 1047.435 ;
    END
  END Data_HV[100]
  PIN Data_HV[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14889.065 1046.435 14889.345 1047.435 ;
    END
  END Data_HV[84]
  PIN MASKH[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14887.385 1046.435 14887.665 1047.435 ;
    END
  END MASKH[172]
  PIN MASKD[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14882.345 1046.435 14882.625 1047.435 ;
    END
  END MASKD[343]
  PIN MASKV[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14871.145 1046.435 14871.425 1047.435 ;
    END
  END MASKV[343]
  PIN Data_HV[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14869.465 1046.435 14869.745 1047.435 ;
    END
  END Data_HV[75]
  PIN Data_HV[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14867.785 1046.435 14868.065 1047.435 ;
    END
  END Data_HV[76]
  PIN Data_HV[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14866.105 1046.435 14866.385 1047.435 ;
    END
  END Data_HV[70]
  PIN nTOK_HV[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14861.345 1046.435 14861.625 1047.435 ;
    END
  END nTOK_HV[3]
  PIN BcidMtx[1029]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14859.105 1046.435 14859.385 1047.435 ;
    END
  END BcidMtx[1029]
  PIN BcidMtx[1026]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14830.825 1046.435 14831.105 1047.435 ;
    END
  END BcidMtx[1026]
  PIN Data_HV[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14828.585 1046.435 14828.865 1047.435 ;
    END
  END Data_HV[66]
  PIN Data_HV[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14826.905 1046.435 14827.185 1047.435 ;
    END
  END Data_HV[78]
  PIN Data_HV[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14824.665 1046.435 14824.945 1047.435 ;
    END
  END Data_HV[74]
  PIN Data_HV[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14823.545 1046.435 14823.825 1047.435 ;
    END
  END Data_HV[63]
  PIN MASKH[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14821.865 1046.435 14822.145 1047.435 ;
    END
  END MASKH[171]
  PIN MASKD[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14803.945 1046.435 14804.225 1047.435 ;
    END
  END MASKD[341]
  PIN MASKV[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14801.145 1046.435 14801.425 1047.435 ;
    END
  END MASKV[341]
  PIN Data_HV[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14799.465 1046.435 14799.745 1047.435 ;
    END
  END Data_HV[54]
  PIN Data_HV[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14797.785 1046.435 14798.065 1047.435 ;
    END
  END Data_HV[55]
  PIN Data_HV[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14796.105 1046.435 14796.385 1047.435 ;
    END
  END Data_HV[49]
  PIN nTOK_HV[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14754.105 1046.435 14754.385 1047.435 ;
    END
  END nTOK_HV[2]
  PIN BcidMtx[1023]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14751.865 1046.435 14752.145 1047.435 ;
    END
  END BcidMtx[1023]
  PIN BcidMtx[1022]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14750.185 1046.435 14750.465 1047.435 ;
    END
  END BcidMtx[1022]
  PIN INJ_IN[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14747.945 1046.435 14748.225 1047.435 ;
    END
  END INJ_IN[340]
  PIN Data_HV[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14746.265 1046.435 14746.545 1047.435 ;
    END
  END Data_HV[44]
  PIN Data_HV[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14744.585 1046.435 14744.865 1047.435 ;
    END
  END Data_HV[52]
  PIN Data_HV[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14743.465 1046.435 14743.745 1047.435 ;
    END
  END Data_HV[58]
  PIN Data_HV[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14742.345 1046.435 14742.625 1047.435 ;
    END
  END Data_HV[43]
  PIN MASKV[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14732.265 1046.435 14732.545 1047.435 ;
    END
  END MASKV[340]
  PIN DIG_MON_SEL[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14727.785 1046.435 14728.065 1047.435 ;
    END
  END DIG_MON_SEL[339]
  PIN DIG_MON_HV[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14725.545 1046.435 14725.825 1047.435 ;
    END
  END DIG_MON_HV[3]
  PIN Data_HV[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14721.345 1046.435 14721.625 1047.435 ;
    END
  END Data_HV[39]
  PIN Data_HV[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14719.105 1046.435 14719.385 1047.435 ;
    END
  END Data_HV[26]
  PIN Data_HV[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14692.505 1046.435 14692.785 1047.435 ;
    END
  END Data_HV[41]
  PIN Data_HV[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14690.825 1046.435 14691.105 1047.435 ;
    END
  END Data_HV[27]
  PIN nTOK_HV[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14688.585 1046.435 14688.865 1047.435 ;
    END
  END nTOK_HV[1]
  PIN BcidMtx[1017]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14686.345 1046.435 14686.625 1047.435 ;
    END
  END BcidMtx[1017]
  PIN Read_HV[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14685.225 1046.435 14685.505 1047.435 ;
    END
  END Read_HV[1]
  PIN INJ_IN[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14682.425 1046.435 14682.705 1047.435 ;
    END
  END INJ_IN[338]
  PIN Data_HV[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14680.745 1046.435 14681.025 1047.435 ;
    END
  END Data_HV[23]
  PIN Data_HV[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14666.185 1046.435 14666.465 1047.435 ;
    END
  END Data_HV[31]
  PIN Data_HV[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14665.065 1046.435 14665.345 1047.435 ;
    END
  END Data_HV[37]
  PIN Data_HV[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14663.385 1046.435 14663.665 1047.435 ;
    END
  END Data_HV[21]
  PIN MASKH[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14661.705 1046.435 14661.985 1047.435 ;
    END
  END MASKH[169]
  PIN DIG_MON_SEL[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14657.785 1046.435 14658.065 1047.435 ;
    END
  END DIG_MON_SEL[337]
  PIN MASKV[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14653.865 1046.435 14654.145 1047.435 ;
    END
  END MASKV[337]
  PIN Data_HV[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14612.425 1046.435 14612.705 1047.435 ;
    END
  END Data_HV[12]
  PIN Data_HV[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14611.305 1046.435 14611.585 1047.435 ;
    END
  END Data_HV[5]
  PIN Data_HV[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14610.185 1046.435 14610.465 1047.435 ;
    END
  END Data_HV[20]
  PIN nTOK_HV[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14606.265 1046.435 14606.545 1047.435 ;
    END
  END nTOK_HV[0]
  PIN BcidMtx[1012]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14604.585 1046.435 14604.865 1047.435 ;
    END
  END BcidMtx[1012]
  PIN FREEZE_HV[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14603.465 1046.435 14603.745 1047.435 ;
    END
  END FREEZE_HV[0]
  PIN BcidMtx[1009]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14601.785 1046.435 14602.065 1047.435 ;
    END
  END BcidMtx[1009]
  PIN Data_HV[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14590.025 1046.435 14590.305 1047.435 ;
    END
  END Data_HV[2]
  PIN Data_HV[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14588.345 1046.435 14588.625 1047.435 ;
    END
  END Data_HV[10]
  PIN Data_COMP[735]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12905.545 1046.435 12905.825 1047.435 ;
    END
  END Data_COMP[735]
  PIN MASKH[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12901.905 1046.435 12902.185 1047.435 ;
    END
  END MASKH[147]
  PIN DIG_MON_SEL[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13991.945 1046.435 13992.225 1047.435 ;
    END
  END DIG_MON_SEL[321]
  PIN INJ_ROW[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13988.585 1046.435 13988.865 1047.435 ;
    END
  END INJ_ROW[160]
  PIN Data_COMP[1016]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13986.905 1046.435 13987.185 1047.435 ;
    END
  END Data_COMP[1016]
  PIN Data_COMP[1027]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13985.785 1046.435 13986.065 1047.435 ;
    END
  END Data_COMP[1027]
  PIN Data_COMP[1028]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13984.105 1046.435 13984.385 1047.435 ;
    END
  END Data_COMP[1028]
  PIN Data_COMP[1014]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13982.425 1046.435 13982.705 1047.435 ;
    END
  END Data_COMP[1014]
  PIN BcidMtx[965]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13965.625 1046.435 13965.905 1047.435 ;
    END
  END BcidMtx[965]
  PIN FREEZE_COMP[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13963.945 1046.435 13964.225 1047.435 ;
    END
  END FREEZE_COMP[48]
  PIN BcidMtx[961]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13962.265 1046.435 13962.545 1047.435 ;
    END
  END BcidMtx[961]
  PIN Data_COMP[1011]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13959.465 1046.435 13959.745 1047.435 ;
    END
  END Data_COMP[1011]
  PIN Data_COMP[1023]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13957.785 1046.435 13958.065 1047.435 ;
    END
  END Data_COMP[1023]
  PIN Data_COMP[1024]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13956.105 1046.435 13956.385 1047.435 ;
    END
  END Data_COMP[1024]
  PIN Data_COMP[1008]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13954.425 1046.435 13954.705 1047.435 ;
    END
  END Data_COMP[1008]
  PIN MASKH[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13914.105 1046.435 13914.385 1047.435 ;
    END
  END MASKH[160]
  PIN MASKD[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13909.065 1046.435 13909.345 1047.435 ;
    END
  END MASKD[319]
  PIN MASKV[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13906.265 1046.435 13906.545 1047.435 ;
    END
  END MASKV[319]
  PIN Data_COMP[999]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13904.585 1046.435 13904.865 1047.435 ;
    END
  END Data_COMP[999]
  PIN Data_COMP[1000]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13902.905 1046.435 13903.185 1047.435 ;
    END
  END Data_COMP[1000]
  PIN Data_COMP[994]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13901.225 1046.435 13901.505 1047.435 ;
    END
  END Data_COMP[994]
  PIN nTOK_COMP[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13890.025 1046.435 13890.305 1047.435 ;
    END
  END nTOK_COMP[47]
  PIN BcidMtx[957]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13887.785 1046.435 13888.065 1047.435 ;
    END
  END BcidMtx[957]
  PIN BcidMtx[956]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13886.105 1046.435 13886.385 1047.435 ;
    END
  END BcidMtx[956]
  PIN INJ_IN[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13881.905 1046.435 13882.185 1047.435 ;
    END
  END INJ_IN[318]
  PIN Data_COMP[996]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13879.665 1046.435 13879.945 1047.435 ;
    END
  END Data_COMP[996]
  PIN Data_COMP[991]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13852.505 1046.435 13852.785 1047.435 ;
    END
  END Data_COMP[991]
  PIN Data_COMP[988]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13850.825 1046.435 13851.105 1047.435 ;
    END
  END Data_COMP[988]
  PIN MASKV[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13849.145 1046.435 13849.425 1047.435 ;
    END
  END MASKV[318]
  PIN DIG_MON_COMP[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13846.905 1046.435 13847.185 1047.435 ;
    END
  END DIG_MON_COMP[94]
  PIN DIG_MON_SEL[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13844.665 1046.435 13844.945 1047.435 ;
    END
  END DIG_MON_SEL[317]
  PIN INJ_ROW[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13841.305 1046.435 13841.585 1047.435 ;
    END
  END INJ_ROW[158]
  PIN Data_COMP[974]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13839.625 1046.435 13839.905 1047.435 ;
    END
  END Data_COMP[974]
  PIN Data_COMP[971]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13825.065 1046.435 13825.345 1047.435 ;
    END
  END Data_COMP[971]
  PIN Data_COMP[980]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13823.385 1046.435 13823.665 1047.435 ;
    END
  END Data_COMP[980]
  PIN INJ_IN[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13821.145 1046.435 13821.425 1047.435 ;
    END
  END INJ_IN[317]
  PIN BcidMtx[952]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13818.345 1046.435 13818.625 1047.435 ;
    END
  END BcidMtx[952]
  PIN Read_COMP[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13816.665 1046.435 13816.945 1047.435 ;
    END
  END Read_COMP[46]
  PIN BcidMtx[948]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13814.985 1046.435 13815.265 1047.435 ;
    END
  END BcidMtx[948]
  PIN Data_COMP[968]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13773.545 1046.435 13773.825 1047.435 ;
    END
  END Data_COMP[968]
  PIN Data_COMP[976]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13771.865 1046.435 13772.145 1047.435 ;
    END
  END Data_COMP[976]
  PIN Data_COMP[977]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13770.185 1046.435 13770.465 1047.435 ;
    END
  END Data_COMP[977]
  PIN Data_COMP[983]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13768.505 1046.435 13768.785 1047.435 ;
    END
  END Data_COMP[983]
  PIN MASKD[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13766.825 1046.435 13767.105 1047.435 ;
    END
  END MASKD[316]
  PIN DIG_MON_SEL[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13764.025 1046.435 13764.305 1047.435 ;
    END
  END DIG_MON_SEL[316]
  PIN DIG_MON_COMP[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13761.225 1046.435 13761.505 1047.435 ;
    END
  END DIG_MON_COMP[91]
  PIN Data_COMP[963]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13750.585 1046.435 13750.865 1047.435 ;
    END
  END Data_COMP[963]
  PIN Data_COMP[964]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13748.905 1046.435 13749.185 1047.435 ;
    END
  END Data_COMP[964]
  PIN Data_COMP[965]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13747.225 1046.435 13747.505 1047.435 ;
    END
  END Data_COMP[965]
  PIN Data_COMP[951]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13745.545 1046.435 13745.825 1047.435 ;
    END
  END Data_COMP[951]
  PIN BcidMtx[947]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13740.225 1046.435 13740.505 1047.435 ;
    END
  END BcidMtx[947]
  PIN Read_COMP[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13712.505 1046.435 13712.785 1047.435 ;
    END
  END Read_COMP[45]
  PIN BcidMtx[942]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13710.825 1046.435 13711.105 1047.435 ;
    END
  END BcidMtx[942]
  PIN Data_COMP[947]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13708.025 1046.435 13708.305 1047.435 ;
    END
  END Data_COMP[947]
  PIN Data_COMP[955]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13706.345 1046.435 13706.625 1047.435 ;
    END
  END Data_COMP[955]
  PIN Data_COMP[956]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13704.665 1046.435 13704.945 1047.435 ;
    END
  END Data_COMP[956]
  PIN Data_COMP[962]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13702.985 1046.435 13703.265 1047.435 ;
    END
  END Data_COMP[962]
  PIN MASKD[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13701.305 1046.435 13701.585 1047.435 ;
    END
  END MASKD[314]
  PIN MASKV[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18742.425 1046.435 18742.705 1047.435 ;
    END
  END MASKV[440]
  PIN INJ_ROW[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13681.705 1046.435 13681.985 1047.435 ;
    END
  END INJ_ROW[156]
  PIN Data_COMP[932]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13680.025 1046.435 13680.305 1047.435 ;
    END
  END Data_COMP[932]
  PIN Data_COMP[929]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13678.345 1046.435 13678.625 1047.435 ;
    END
  END Data_COMP[929]
  PIN Data_COMP[938]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13676.665 1046.435 13676.945 1047.435 ;
    END
  END Data_COMP[938]
  PIN INJ_IN[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13674.425 1046.435 13674.705 1047.435 ;
    END
  END INJ_IN[313]
  PIN BcidMtx[940]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13632.425 1046.435 13632.705 1047.435 ;
    END
  END BcidMtx[940]
  PIN Read_COMP[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13630.745 1046.435 13631.025 1047.435 ;
    END
  END Read_COMP[44]
  PIN BcidMtx[936]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13629.065 1046.435 13629.345 1047.435 ;
    END
  END BcidMtx[936]
  PIN Data_COMP[926]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13626.265 1046.435 13626.545 1047.435 ;
    END
  END Data_COMP[926]
  PIN Data_COMP[934]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13624.585 1046.435 13624.865 1047.435 ;
    END
  END Data_COMP[934]
  PIN Data_COMP[935]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13622.905 1046.435 13623.185 1047.435 ;
    END
  END Data_COMP[935]
  PIN Data_COMP[941]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13621.225 1046.435 13621.505 1047.435 ;
    END
  END Data_COMP[941]
  PIN MASKD[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13611.145 1046.435 13611.425 1047.435 ;
    END
  END MASKD[312]
  PIN MASKD[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13606.665 1046.435 13606.945 1047.435 ;
    END
  END MASKD[311]
  PIN INJ_ROW[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13602.465 1046.435 13602.745 1047.435 ;
    END
  END INJ_ROW[155]
  PIN Data_COMP[911]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13600.785 1046.435 13601.065 1047.435 ;
    END
  END Data_COMP[911]
  PIN Data_COMP[908]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13599.105 1046.435 13599.385 1047.435 ;
    END
  END Data_COMP[908]
  PIN Data_COMP[917]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13571.945 1046.435 13572.225 1047.435 ;
    END
  END Data_COMP[917]
  PIN INJ_IN[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13569.705 1046.435 13569.985 1047.435 ;
    END
  END INJ_IN[311]
  PIN BcidMtx[934]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13566.905 1046.435 13567.185 1047.435 ;
    END
  END BcidMtx[934]
  PIN Read_COMP[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13565.225 1046.435 13565.505 1047.435 ;
    END
  END Read_COMP[43]
  PIN BcidMtx[930]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13563.545 1046.435 13563.825 1047.435 ;
    END
  END BcidMtx[930]
  PIN Data_COMP[905]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13560.745 1046.435 13561.025 1047.435 ;
    END
  END Data_COMP[905]
  PIN Data_COMP[913]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13546.185 1046.435 13546.465 1047.435 ;
    END
  END Data_COMP[913]
  PIN Data_COMP[914]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13544.505 1046.435 13544.785 1047.435 ;
    END
  END Data_COMP[914]
  PIN Data_COMP[920]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13542.825 1046.435 13543.105 1047.435 ;
    END
  END Data_COMP[920]
  PIN MASKD[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13541.145 1046.435 13541.425 1047.435 ;
    END
  END MASKD[310]
  PIN DIG_MON_SEL[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13538.345 1046.435 13538.625 1047.435 ;
    END
  END DIG_MON_SEL[310]
  PIN MASKD[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13536.665 1046.435 13536.945 1047.435 ;
    END
  END MASKD[309]
  PIN MASKV[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13533.865 1046.435 13534.145 1047.435 ;
    END
  END MASKV[309]
  PIN Data_COMP[894]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13492.425 1046.435 13492.705 1047.435 ;
    END
  END Data_COMP[894]
  PIN Data_COMP[895]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13490.745 1046.435 13491.025 1047.435 ;
    END
  END Data_COMP[895]
  PIN Data_COMP[889]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13489.065 1046.435 13489.345 1047.435 ;
    END
  END Data_COMP[889]
  PIN nTOK_COMP[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13486.265 1046.435 13486.545 1047.435 ;
    END
  END nTOK_COMP[42]
  PIN BcidMtx[927]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13484.025 1046.435 13484.305 1047.435 ;
    END
  END BcidMtx[927]
  PIN Read_COMP[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13482.905 1046.435 13483.185 1047.435 ;
    END
  END Read_COMP[42]
  PIN INJ_IN[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13471.705 1046.435 13471.985 1047.435 ;
    END
  END INJ_IN[308]
  PIN Data_COMP[884]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13470.025 1046.435 13470.305 1047.435 ;
    END
  END Data_COMP[884]
  PIN Data_COMP[897]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13468.905 1046.435 13469.185 1047.435 ;
    END
  END Data_COMP[897]
  PIN Data_COMP[893]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13466.665 1046.435 13466.945 1047.435 ;
    END
  END Data_COMP[893]
  PIN Data_COMP[899]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13464.985 1046.435 13465.265 1047.435 ;
    END
  END Data_COMP[899]
  PIN MASKH[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13461.905 1046.435 13462.185 1047.435 ;
    END
  END MASKH[154]
  PIN DIG_MON_SEL[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13458.545 1046.435 13458.825 1047.435 ;
    END
  END DIG_MON_SEL[308]
  PIN MASKD[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14550.825 1046.435 14551.105 1047.435 ;
    END
  END MASKD[335]
  PIN DIG_MON_COMP[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14549.705 1046.435 14549.985 1047.435 ;
    END
  END DIG_MON_COMP[111]
  PIN Data_COMP[1163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14546.905 1046.435 14547.185 1047.435 ;
    END
  END Data_COMP[1163]
  PIN Data_COMP[1160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14545.225 1046.435 14545.505 1047.435 ;
    END
  END Data_COMP[1160]
  PIN Data_COMP[1175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14544.105 1046.435 14544.385 1047.435 ;
    END
  END Data_COMP[1175]
  PIN Data_COMP[1161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14542.425 1046.435 14542.705 1047.435 ;
    END
  END Data_COMP[1161]
  PIN BcidMtx[1007]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14525.625 1046.435 14525.905 1047.435 ;
    END
  END BcidMtx[1007]
  PIN FREEZE_COMP[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14523.945 1046.435 14524.225 1047.435 ;
    END
  END FREEZE_COMP[55]
  PIN BcidMtx[1003]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14522.265 1046.435 14522.545 1047.435 ;
    END
  END BcidMtx[1003]
  PIN Data_COMP[1158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14519.465 1046.435 14519.745 1047.435 ;
    END
  END Data_COMP[1158]
  PIN Data_COMP[1170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14517.785 1046.435 14518.065 1047.435 ;
    END
  END Data_COMP[1170]
  PIN Data_COMP[1171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14516.105 1046.435 14516.385 1047.435 ;
    END
  END Data_COMP[1171]
  PIN Data_COMP[1155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14514.425 1046.435 14514.705 1047.435 ;
    END
  END Data_COMP[1155]
  PIN MASKH[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14474.105 1046.435 14474.385 1047.435 ;
    END
  END MASKH[167]
  PIN MASKD[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14469.065 1046.435 14469.345 1047.435 ;
    END
  END MASKD[333]
  PIN MASKV[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14466.265 1046.435 14466.545 1047.435 ;
    END
  END MASKV[333]
  PIN Data_COMP[1146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14464.585 1046.435 14464.865 1047.435 ;
    END
  END Data_COMP[1146]
  PIN Data_COMP[1147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14462.905 1046.435 14463.185 1047.435 ;
    END
  END Data_COMP[1147]
  PIN Data_COMP[1141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14461.225 1046.435 14461.505 1047.435 ;
    END
  END Data_COMP[1141]
  PIN BcidMtx[1000]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14448.345 1046.435 14448.625 1047.435 ;
    END
  END BcidMtx[1000]
  PIN Read_COMP[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14446.665 1046.435 14446.945 1047.435 ;
    END
  END Read_COMP[54]
  PIN BcidMtx[998]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14446.105 1046.435 14446.385 1047.435 ;
    END
  END BcidMtx[998]
  PIN Data_COMP[1136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14440.225 1046.435 14440.505 1047.435 ;
    END
  END Data_COMP[1136]
  PIN Data_COMP[1144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14438.545 1046.435 14438.825 1047.435 ;
    END
  END Data_COMP[1144]
  PIN Data_COMP[1138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14412.505 1046.435 14412.785 1047.435 ;
    END
  END Data_COMP[1138]
  PIN Data_COMP[1151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14409.705 1046.435 14409.985 1047.435 ;
    END
  END Data_COMP[1151]
  PIN MASKD[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14408.025 1046.435 14408.305 1047.435 ;
    END
  END MASKD[332]
  PIN DIG_MON_COMP[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14406.905 1046.435 14407.185 1047.435 ;
    END
  END DIG_MON_COMP[108]
  PIN DIG_MON_COMP[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14402.425 1046.435 14402.705 1047.435 ;
    END
  END DIG_MON_COMP[107]
  PIN Data_COMP[1131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14400.185 1046.435 14400.465 1047.435 ;
    END
  END Data_COMP[1131]
  PIN Data_COMP[1121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14399.625 1046.435 14399.905 1047.435 ;
    END
  END Data_COMP[1121]
  PIN Data_COMP[1133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14383.945 1046.435 14384.225 1047.435 ;
    END
  END Data_COMP[1133]
  PIN Data_COMP[1119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14382.265 1046.435 14382.545 1047.435 ;
    END
  END Data_COMP[1119]
  PIN INJ_IN[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14381.145 1046.435 14381.425 1047.435 ;
    END
  END INJ_IN[331]
  PIN FREEZE_COMP[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14377.225 1046.435 14377.505 1047.435 ;
    END
  END FREEZE_COMP[53]
  PIN BcidMtx[991]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14375.545 1046.435 14375.825 1047.435 ;
    END
  END BcidMtx[991]
  PIN BcidMtx[990]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14374.985 1046.435 14375.265 1047.435 ;
    END
  END BcidMtx[990]
  PIN Data_COMP[1128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14332.425 1046.435 14332.705 1047.435 ;
    END
  END Data_COMP[1128]
  PIN Data_COMP[1129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14330.745 1046.435 14331.025 1047.435 ;
    END
  END Data_COMP[1129]
  PIN Data_COMP[1124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14330.185 1046.435 14330.465 1047.435 ;
    END
  END Data_COMP[1124]
  PIN MASKH[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14327.385 1046.435 14327.665 1047.435 ;
    END
  END MASKH[165]
  PIN DIG_MON_SEL[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14324.025 1046.435 14324.305 1047.435 ;
    END
  END DIG_MON_SEL[330]
  PIN MASKV[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14311.145 1046.435 14311.425 1047.435 ;
    END
  END MASKV[329]
  PIN Data_COMP[1104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14309.465 1046.435 14309.745 1047.435 ;
    END
  END Data_COMP[1104]
  PIN Data_COMP[1111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14308.905 1046.435 14309.185 1047.435 ;
    END
  END Data_COMP[1111]
  PIN Data_COMP[1099]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14306.105 1046.435 14306.385 1047.435 ;
    END
  END Data_COMP[1099]
  PIN nTOK_COMP[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14301.345 1046.435 14301.625 1047.435 ;
    END
  END nTOK_COMP[52]
  PIN BcidMtx[989]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14300.225 1046.435 14300.505 1047.435 ;
    END
  END BcidMtx[989]
  PIN BcidMtx[985]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14271.385 1046.435 14271.665 1047.435 ;
    END
  END BcidMtx[985]
  PIN INJ_IN[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14269.705 1046.435 14269.985 1047.435 ;
    END
  END INJ_IN[328]
  PIN Data_COMP[1094]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14268.025 1046.435 14268.305 1047.435 ;
    END
  END Data_COMP[1094]
  PIN Data_COMP[1108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14265.225 1046.435 14265.505 1047.435 ;
    END
  END Data_COMP[1108]
  PIN Data_COMP[1092]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14263.545 1046.435 14263.825 1047.435 ;
    END
  END Data_COMP[1092]
  PIN Data_COMP[1109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14262.985 1046.435 14263.265 1047.435 ;
    END
  END Data_COMP[1109]
  PIN DIG_MON_COMP[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14260.185 1046.435 14260.465 1047.435 ;
    END
  END DIG_MON_COMP[104]
  PIN DIG_MON_SEL[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14245.065 1046.435 14245.345 1047.435 ;
    END
  END DIG_MON_SEL[327]
  PIN MASKD[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14243.945 1046.435 14244.225 1047.435 ;
    END
  END MASKD[327]
  PIN Data_COMP[1079]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14240.025 1046.435 14240.305 1047.435 ;
    END
  END Data_COMP[1079]
  PIN Data_COMP[1076]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14238.345 1046.435 14238.625 1047.435 ;
    END
  END Data_COMP[1076]
  PIN Data_COMP[1084]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14237.785 1046.435 14238.065 1047.435 ;
    END
  END Data_COMP[1084]
  PIN INJ_IN[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14234.425 1046.435 14234.705 1047.435 ;
    END
  END INJ_IN[327]
  PIN BcidMtx[982]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14192.425 1046.435 14192.705 1047.435 ;
    END
  END BcidMtx[982]
  PIN BcidMtx[981]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14191.865 1046.435 14192.145 1047.435 ;
    END
  END BcidMtx[981]
  PIN BcidMtx[978]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14189.065 1046.435 14189.345 1047.435 ;
    END
  END BcidMtx[978]
  PIN Data_COMP[1073]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14186.265 1046.435 14186.545 1047.435 ;
    END
  END Data_COMP[1073]
  PIN Data_COMP[1080]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14185.705 1046.435 14185.985 1047.435 ;
    END
  END Data_COMP[1080]
  PIN Data_COMP[1082]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14182.905 1046.435 14183.185 1047.435 ;
    END
  END Data_COMP[1082]
  PIN Data_COMP[1088]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14181.225 1046.435 14181.505 1047.435 ;
    END
  END Data_COMP[1088]
  PIN MASKV[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14172.265 1046.435 14172.545 1047.435 ;
    END
  END MASKV[326]
  PIN MASKD[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14166.665 1046.435 14166.945 1047.435 ;
    END
  END MASKD[325]
  PIN DIG_MON_COMP[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14165.545 1046.435 14165.825 1047.435 ;
    END
  END DIG_MON_COMP[101]
  PIN Data_COMP[1062]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14160.225 1046.435 14160.505 1047.435 ;
    END
  END Data_COMP[1062]
  PIN Data_COMP[1063]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14133.065 1046.435 14133.345 1047.435 ;
    END
  END Data_COMP[1063]
  PIN Data_COMP[1070]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14132.505 1046.435 14132.785 1047.435 ;
    END
  END Data_COMP[1070]
  PIN nTOK_COMP[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14128.585 1046.435 14128.865 1047.435 ;
    END
  END nTOK_COMP[50]
  PIN BcidMtx[975]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14126.345 1046.435 14126.625 1047.435 ;
    END
  END BcidMtx[975]
  PIN FREEZE_COMP[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14125.785 1046.435 14126.065 1047.435 ;
    END
  END FREEZE_COMP[50]
  PIN INJ_IN[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14122.425 1046.435 14122.705 1047.435 ;
    END
  END INJ_IN[324]
  PIN Data_COMP[1059]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14120.185 1046.435 14120.465 1047.435 ;
    END
  END Data_COMP[1059]
  PIN Data_COMP[1065]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14106.745 1046.435 14107.025 1047.435 ;
    END
  END Data_COMP[1065]
  PIN Data_COMP[1051]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14103.945 1046.435 14104.225 1047.435 ;
    END
  END Data_COMP[1051]
  PIN MASKV[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14102.265 1046.435 14102.545 1047.435 ;
    END
  END MASKV[324]
  PIN MASKH[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14101.705 1046.435 14101.985 1047.435 ;
    END
  END MASKH[162]
  PIN DIG_MON_SEL[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14098.345 1046.435 14098.625 1047.435 ;
    END
  END DIG_MON_SEL[324]
  PIN DIG_MON_COMP[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14095.545 1046.435 14095.825 1047.435 ;
    END
  END DIG_MON_COMP[99]
  PIN INJ_ROW[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14094.425 1046.435 14094.705 1047.435 ;
    END
  END INJ_ROW[161]
  PIN Data_COMP[1048]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14051.865 1046.435 14052.145 1047.435 ;
    END
  END Data_COMP[1048]
  PIN Data_COMP[1049]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14050.185 1046.435 14050.465 1047.435 ;
    END
  END Data_COMP[1049]
  PIN Data_COMP[1043]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14049.625 1046.435 14049.905 1047.435 ;
    END
  END Data_COMP[1043]
  PIN BcidMtx[971]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14045.145 1046.435 14045.425 1047.435 ;
    END
  END BcidMtx[971]
  PIN FREEZE_COMP[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14043.465 1046.435 14043.745 1047.435 ;
    END
  END FREEZE_COMP[49]
  PIN BcidMtx[968]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14042.345 1046.435 14042.625 1047.435 ;
    END
  END BcidMtx[968]
  PIN Data_COMP[1031]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14030.025 1046.435 14030.305 1047.435 ;
    END
  END Data_COMP[1031]
  PIN Data_COMP[1044]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14028.905 1046.435 14029.185 1047.435 ;
    END
  END Data_COMP[1044]
  PIN Data_COMP[1033]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14027.785 1046.435 14028.065 1047.435 ;
    END
  END Data_COMP[1033]
  PIN BcidMtx[1134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16281.225 1046.435 16281.505 1047.435 ;
    END
  END BcidMtx[1134]
  PIN Data_HV[443]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16270.025 1046.435 16270.305 1047.435 ;
    END
  END Data_HV[443]
  PIN Data_HV[451]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16268.345 1046.435 16268.625 1047.435 ;
    END
  END Data_HV[451]
  PIN Data_HV[452]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16266.665 1046.435 16266.945 1047.435 ;
    END
  END Data_HV[452]
  PIN Data_HV[458]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16264.985 1046.435 16265.265 1047.435 ;
    END
  END Data_HV[458]
  PIN DIG_MON_SEL[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17351.945 1046.435 17352.225 1047.435 ;
    END
  END DIG_MON_SEL[405]
  PIN DIG_MON_HV[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17349.705 1046.435 17349.985 1047.435 ;
    END
  END DIG_MON_HV[69]
  PIN Data_HV[722]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17346.905 1046.435 17347.185 1047.435 ;
    END
  END Data_HV[722]
  PIN Data_HV[719]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17345.225 1046.435 17345.505 1047.435 ;
    END
  END Data_HV[719]
  PIN Data_HV[734]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17344.105 1046.435 17344.385 1047.435 ;
    END
  END Data_HV[734]
  PIN INJ_IN[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17341.305 1046.435 17341.585 1047.435 ;
    END
  END INJ_IN[405]
  PIN BcidMtx[1216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17325.065 1046.435 17325.345 1047.435 ;
    END
  END BcidMtx[1216]
  PIN FREEZE_HV[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17323.945 1046.435 17324.225 1047.435 ;
    END
  END FREEZE_HV[34]
  PIN BcidMtx[1212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17321.705 1046.435 17321.985 1047.435 ;
    END
  END BcidMtx[1212]
  PIN Data_HV[716]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17318.905 1046.435 17319.185 1047.435 ;
    END
  END Data_HV[716]
  PIN Data_HV[729]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17317.785 1046.435 17318.065 1047.435 ;
    END
  END Data_HV[729]
  PIN Data_HV[725]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17315.545 1046.435 17315.825 1047.435 ;
    END
  END Data_HV[725]
  PIN Data_HV[731]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17313.865 1046.435 17314.145 1047.435 ;
    END
  END Data_HV[731]
  PIN MASKH[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17274.105 1046.435 17274.385 1047.435 ;
    END
  END MASKH[202]
  PIN DIG_MON_HV[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17272.425 1046.435 17272.705 1047.435 ;
    END
  END DIG_MON_HV[68]
  PIN DIG_MON_SEL[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17270.185 1046.435 17270.465 1047.435 ;
    END
  END DIG_MON_SEL[403]
  PIN INJ_ROW[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17266.825 1046.435 17267.105 1047.435 ;
    END
  END INJ_ROW[201]
  PIN Data_HV[701]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17265.145 1046.435 17265.425 1047.435 ;
    END
  END Data_HV[701]
  PIN Data_HV[698]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17263.465 1046.435 17263.745 1047.435 ;
    END
  END Data_HV[698]
  PIN Data_HV[707]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17261.785 1046.435 17262.065 1047.435 ;
    END
  END Data_HV[707]
  PIN Data_HV[699]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17252.265 1046.435 17252.545 1047.435 ;
    END
  END Data_HV[699]
  PIN BcidMtx[1210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17248.345 1046.435 17248.625 1047.435 ;
    END
  END BcidMtx[1210]
  PIN Read_HV[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17246.665 1046.435 17246.945 1047.435 ;
    END
  END Read_HV[33]
  PIN BcidMtx[1207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17245.545 1046.435 17245.825 1047.435 ;
    END
  END BcidMtx[1207]
  PIN Data_HV[695]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17240.225 1046.435 17240.505 1047.435 ;
    END
  END Data_HV[695]
  PIN Data_HV[703]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17238.545 1046.435 17238.825 1047.435 ;
    END
  END Data_HV[703]
  PIN Data_HV[709]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17211.945 1046.435 17212.225 1047.435 ;
    END
  END Data_HV[709]
  PIN Data_HV[710]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17209.705 1046.435 17209.985 1047.435 ;
    END
  END Data_HV[710]
  PIN MASKD[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17208.025 1046.435 17208.305 1047.435 ;
    END
  END MASKD[402]
  PIN DIG_MON_HV[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17202.425 1046.435 17202.705 1047.435 ;
    END
  END DIG_MON_HV[65]
  PIN MASKV[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17200.745 1046.435 17201.025 1047.435 ;
    END
  END MASKV[401]
  PIN Data_HV[680]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17199.625 1046.435 17199.905 1047.435 ;
    END
  END Data_HV[680]
  PIN Data_HV[685]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17184.505 1046.435 17184.785 1047.435 ;
    END
  END Data_HV[685]
  PIN Data_HV[679]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17182.825 1046.435 17183.105 1047.435 ;
    END
  END Data_HV[679]
  PIN INJ_IN[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17181.145 1046.435 17181.425 1047.435 ;
    END
  END INJ_IN[401]
  PIN BcidMtx[1203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17177.785 1046.435 17178.065 1047.435 ;
    END
  END BcidMtx[1203]
  PIN BcidMtx[1202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17176.105 1046.435 17176.385 1047.435 ;
    END
  END BcidMtx[1202]
  PIN BcidMtx[1200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17174.985 1046.435 17175.265 1047.435 ;
    END
  END BcidMtx[1200]
  PIN Data_HV[681]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17132.985 1046.435 17133.265 1047.435 ;
    END
  END Data_HV[681]
  PIN Data_HV[676]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17131.305 1046.435 17131.585 1047.435 ;
    END
  END Data_HV[676]
  PIN Data_HV[683]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17130.185 1046.435 17130.465 1047.435 ;
    END
  END Data_HV[683]
  PIN MASKV[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17127.945 1046.435 17128.225 1047.435 ;
    END
  END MASKV[400]
  PIN DIG_MON_HV[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17125.705 1046.435 17125.985 1047.435 ;
    END
  END DIG_MON_HV[64]
  PIN DIG_MON_SEL[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17124.025 1046.435 17124.305 1047.435 ;
    END
  END DIG_MON_SEL[400]
  PIN INJ_ROW[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17111.705 1046.435 17111.985 1047.435 ;
    END
  END INJ_ROW[199]
  PIN Data_HV[659]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17110.025 1046.435 17110.305 1047.435 ;
    END
  END Data_HV[659]
  PIN Data_HV[670]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17108.905 1046.435 17109.185 1047.435 ;
    END
  END Data_HV[670]
  PIN Data_HV[665]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17106.665 1046.435 17106.945 1047.435 ;
    END
  END Data_HV[665]
  PIN INJ_IN[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17102.465 1046.435 17102.745 1047.435 ;
    END
  END INJ_IN[399]
  PIN BcidMtx[1199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17100.225 1046.435 17100.505 1047.435 ;
    END
  END BcidMtx[1199]
  PIN BcidMtx[1196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17071.945 1046.435 17072.225 1047.435 ;
    END
  END BcidMtx[1196]
  PIN INJ_IN[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17069.705 1046.435 17069.985 1047.435 ;
    END
  END INJ_IN[398]
  PIN Data_HV[653]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17068.025 1046.435 17068.305 1047.435 ;
    END
  END Data_HV[653]
  PIN Data_HV[655]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17065.785 1046.435 17066.065 1047.435 ;
    END
  END Data_HV[655]
  PIN Data_HV[652]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17064.105 1046.435 17064.385 1047.435 ;
    END
  END Data_HV[652]
  PIN Data_HV[668]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17062.985 1046.435 17063.265 1047.435 ;
    END
  END Data_HV[668]
  PIN DIG_MON_HV[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17060.185 1046.435 17060.465 1047.435 ;
    END
  END DIG_MON_HV[62]
  PIN DIG_MON_SEL[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17045.065 1046.435 17045.345 1047.435 ;
    END
  END DIG_MON_SEL[397]
  PIN DIG_MON_HV[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17042.825 1046.435 17043.105 1047.435 ;
    END
  END DIG_MON_HV[61]
  PIN Data_HV[648]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17040.585 1046.435 17040.865 1047.435 ;
    END
  END Data_HV[648]
  PIN Data_HV[649]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17038.905 1046.435 17039.185 1047.435 ;
    END
  END Data_HV[649]
  PIN Data_HV[643]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17037.785 1046.435 17038.065 1047.435 ;
    END
  END Data_HV[643]
  PIN Data_HV[637]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17036.105 1046.435 17036.385 1047.435 ;
    END
  END Data_HV[637]
  PIN nTOK_HV[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16994.105 1046.435 16994.385 1047.435 ;
    END
  END nTOK_HV[30]
  PIN BcidMtx[1192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16992.425 1046.435 16992.705 1047.435 ;
    END
  END BcidMtx[1192]
  PIN BcidMtx[1190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16990.185 1046.435 16990.465 1047.435 ;
    END
  END BcidMtx[1190]
  PIN INJ_IN[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16987.945 1046.435 16988.225 1047.435 ;
    END
  END INJ_IN[396]
  PIN Data_HV[632]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16986.265 1046.435 16986.545 1047.435 ;
    END
  END Data_HV[632]
  PIN Data_HV[634]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16984.025 1046.435 16984.305 1047.435 ;
    END
  END Data_HV[634]
  PIN Data_HV[631]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16982.345 1046.435 16982.625 1047.435 ;
    END
  END Data_HV[631]
  PIN Data_HV[647]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16981.225 1046.435 16981.505 1047.435 ;
    END
  END Data_HV[647]
  PIN DIG_MON_HV[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16970.025 1046.435 16970.305 1047.435 ;
    END
  END DIG_MON_HV[60]
  PIN DIG_MON_SEL[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16967.785 1046.435 16968.065 1047.435 ;
    END
  END DIG_MON_SEL[395]
  PIN DIG_MON_HV[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16965.545 1046.435 16965.825 1047.435 ;
    END
  END DIG_MON_HV[59]
  PIN Data_HV[617]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16960.785 1046.435 16961.065 1047.435 ;
    END
  END Data_HV[617]
  PIN Data_HV[628]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16959.665 1046.435 16959.945 1047.435 ;
    END
  END Data_HV[628]
  PIN Data_HV[622]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16933.065 1046.435 16933.345 1047.435 ;
    END
  END Data_HV[622]
  PIN Data_HV[615]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16930.825 1046.435 16931.105 1047.435 ;
    END
  END Data_HV[615]
  PIN BcidMtx[1187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16927.465 1046.435 16927.745 1047.435 ;
    END
  END BcidMtx[1187]
  PIN BcidMtx[1185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16926.345 1046.435 16926.625 1047.435 ;
    END
  END BcidMtx[1185]
  PIN BcidMtx[1183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16924.105 1046.435 16924.385 1047.435 ;
    END
  END BcidMtx[1183]
  PIN Data_HV[612]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16921.305 1046.435 16921.585 1047.435 ;
    END
  END Data_HV[612]
  PIN Data_HV[618]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16920.185 1046.435 16920.465 1047.435 ;
    END
  END Data_HV[618]
  PIN Data_HV[625]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16905.065 1046.435 16905.345 1047.435 ;
    END
  END Data_HV[625]
  PIN Data_HV[609]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16903.385 1046.435 16903.665 1047.435 ;
    END
  END Data_HV[609]
  PIN MASKV[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16902.265 1046.435 16902.545 1047.435 ;
    END
  END MASKV[394]
  PIN MASKD[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16896.665 1046.435 16896.945 1047.435 ;
    END
  END MASKD[393]
  PIN INJ_ROW[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16894.425 1046.435 16894.705 1047.435 ;
    END
  END INJ_ROW[196]
  PIN Data_HV[600]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16852.425 1046.435 16852.705 1047.435 ;
    END
  END Data_HV[600]
  PIN Data_HV[601]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16850.745 1046.435 16851.025 1047.435 ;
    END
  END Data_HV[601]
  PIN Data_HV[608]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16850.185 1046.435 16850.465 1047.435 ;
    END
  END Data_HV[608]
  PIN INJ_IN[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16847.385 1046.435 16847.665 1047.435 ;
    END
  END INJ_IN[393]
  PIN BcidMtx[1180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16844.585 1046.435 16844.865 1047.435 ;
    END
  END BcidMtx[1180]
  PIN FREEZE_HV[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16843.465 1046.435 16843.745 1047.435 ;
    END
  END FREEZE_HV[28]
  PIN Data_HV[303]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15709.465 1046.435 15709.745 1047.435 ;
    END
  END Data_HV[303]
  PIN Data_HV[304]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15708.345 1046.435 15708.625 1047.435 ;
    END
  END Data_HV[304]
  PIN Data_HV[310]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15707.225 1046.435 15707.505 1047.435 ;
    END
  END Data_HV[310]
  PIN MASKV[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15702.465 1046.435 15702.745 1047.435 ;
    END
  END MASKV[364]
  PIN MASKD[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15701.345 1046.435 15701.625 1047.435 ;
    END
  END MASKD[364]
  PIN DIG_MON_HV[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16789.705 1046.435 16789.985 1047.435 ;
    END
  END DIG_MON_HV[55]
  PIN MASKV[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16788.025 1046.435 16788.305 1047.435 ;
    END
  END MASKV[391]
  PIN Data_HV[575]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16786.905 1046.435 16787.185 1047.435 ;
    END
  END Data_HV[575]
  PIN Data_HV[587]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16784.105 1046.435 16784.385 1047.435 ;
    END
  END Data_HV[587]
  PIN Data_HV[574]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16782.985 1046.435 16783.265 1047.435 ;
    END
  END Data_HV[574]
  PIN INJ_IN[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16781.305 1046.435 16781.585 1047.435 ;
    END
  END INJ_IN[391]
  PIN FREEZE_HV[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16763.945 1046.435 16764.225 1047.435 ;
    END
  END FREEZE_HV[27]
  PIN BcidMtx[1172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16762.825 1046.435 16763.105 1047.435 ;
    END
  END BcidMtx[1172]
  PIN BcidMtx[1171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16762.265 1046.435 16762.545 1047.435 ;
    END
  END BcidMtx[1171]
  PIN Data_HV[576]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16758.345 1046.435 16758.625 1047.435 ;
    END
  END Data_HV[576]
  PIN Data_HV[571]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16756.665 1046.435 16756.945 1047.435 ;
    END
  END Data_HV[571]
  PIN Data_HV[583]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16756.105 1046.435 16756.385 1047.435 ;
    END
  END Data_HV[583]
  PIN MASKV[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16714.665 1046.435 16714.945 1047.435 ;
    END
  END MASKV[390]
  PIN DIG_MON_HV[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16712.425 1046.435 16712.705 1047.435 ;
    END
  END DIG_MON_HV[54]
  PIN INJ_ROW[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16706.825 1046.435 16707.105 1047.435 ;
    END
  END INJ_ROW[194]
  PIN Data_HV[554]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16705.145 1046.435 16705.425 1047.435 ;
    END
  END Data_HV[554]
  PIN Data_HV[558]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16704.585 1046.435 16704.865 1047.435 ;
    END
  END Data_HV[558]
  PIN Data_HV[560]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16701.785 1046.435 16702.065 1047.435 ;
    END
  END Data_HV[560]
  PIN INJ_IN[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16691.145 1046.435 16691.425 1047.435 ;
    END
  END INJ_IN[389]
  PIN nTOK_HV[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16690.025 1046.435 16690.305 1047.435 ;
    END
  END nTOK_HV[26]
  PIN Read_HV[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16686.665 1046.435 16686.945 1047.435 ;
    END
  END Read_HV[26]
  PIN BcidMtx[1164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16684.985 1046.435 16685.265 1047.435 ;
    END
  END BcidMtx[1164]
  PIN Data_HV[549]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16680.785 1046.435 16681.065 1047.435 ;
    END
  END Data_HV[549]
  PIN Data_HV[550]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16652.505 1046.435 16652.785 1047.435 ;
    END
  END Data_HV[550]
  PIN Data_HV[557]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16651.385 1046.435 16651.665 1047.435 ;
    END
  END Data_HV[557]
  PIN Data_HV[547]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16650.825 1046.435 16651.105 1047.435 ;
    END
  END Data_HV[547]
  PIN MASKD[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16648.025 1046.435 16648.305 1047.435 ;
    END
  END MASKD[388]
  PIN DIG_MON_SEL[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16645.225 1046.435 16645.505 1047.435 ;
    END
  END DIG_MON_SEL[388]
  PIN DIG_MON_SEL[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16644.665 1046.435 16644.945 1047.435 ;
    END
  END DIG_MON_SEL[387]
  PIN MASKV[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16640.745 1046.435 16641.025 1047.435 ;
    END
  END MASKV[387]
  PIN Data_HV[533]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16639.625 1046.435 16639.905 1047.435 ;
    END
  END Data_HV[533]
  PIN Data_HV[544]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16625.625 1046.435 16625.905 1047.435 ;
    END
  END Data_HV[544]
  PIN Data_HV[539]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16623.385 1046.435 16623.665 1047.435 ;
    END
  END Data_HV[539]
  PIN Data_HV[531]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16622.265 1046.435 16622.545 1047.435 ;
    END
  END Data_HV[531]
  PIN nTOK_HV[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16620.025 1046.435 16620.305 1047.435 ;
    END
  END nTOK_HV[25]
  PIN Read_HV[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16616.665 1046.435 16616.945 1047.435 ;
    END
  END Read_HV[25]
  PIN BcidMtx[1159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16615.545 1046.435 16615.825 1047.435 ;
    END
  END BcidMtx[1159]
  PIN INJ_IN[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16613.865 1046.435 16614.145 1047.435 ;
    END
  END INJ_IN[386]
  PIN Data_HV[535]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16571.865 1046.435 16572.145 1047.435 ;
    END
  END Data_HV[535]
  PIN Data_HV[541]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16570.745 1046.435 16571.025 1047.435 ;
    END
  END Data_HV[541]
  PIN Data_HV[526]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16569.625 1046.435 16569.905 1047.435 ;
    END
  END Data_HV[526]
  PIN MASKD[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16566.825 1046.435 16567.105 1047.435 ;
    END
  END MASKD[386]
  PIN DIG_MON_SEL[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16563.465 1046.435 16563.745 1047.435 ;
    END
  END DIG_MON_SEL[385]
  PIN Data_HV[522]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16550.585 1046.435 16550.865 1047.435 ;
    END
  END Data_HV[522]
  PIN Data_HV[516]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16549.465 1046.435 16549.745 1047.435 ;
    END
  END Data_HV[516]
  PIN Data_HV[509]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16548.345 1046.435 16548.625 1047.435 ;
    END
  END Data_HV[509]
  PIN Data_HV[511]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16546.105 1046.435 16546.385 1047.435 ;
    END
  END Data_HV[511]
  PIN Data_HV[510]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16545.545 1046.435 16545.825 1047.435 ;
    END
  END Data_HV[510]
  PIN nTOK_HV[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16541.345 1046.435 16541.625 1047.435 ;
    END
  END nTOK_HV[24]
  PIN BcidMtx[1154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16511.945 1046.435 16512.225 1047.435 ;
    END
  END BcidMtx[1154]
  PIN BcidMtx[1152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16510.825 1046.435 16511.105 1047.435 ;
    END
  END BcidMtx[1152]
  PIN Data_HV[507]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16508.585 1046.435 16508.865 1047.435 ;
    END
  END Data_HV[507]
  PIN Data_HV[508]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16505.785 1046.435 16506.065 1047.435 ;
    END
  END Data_HV[508]
  PIN Data_HV[515]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16504.665 1046.435 16504.945 1047.435 ;
    END
  END Data_HV[515]
  PIN Data_HV[504]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16503.545 1046.435 16503.825 1047.435 ;
    END
  END Data_HV[504]
  PIN DIG_MON_HV[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16500.185 1046.435 16500.465 1047.435 ;
    END
  END DIG_MON_HV[48]
  PIN DIG_MON_SEL[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16485.625 1046.435 16485.905 1047.435 ;
    END
  END DIG_MON_SEL[384]
  PIN MASKD[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16483.945 1046.435 16484.225 1047.435 ;
    END
  END MASKD[383]
  PIN Data_HV[491]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16480.025 1046.435 16480.305 1047.435 ;
    END
  END Data_HV[491]
  PIN Data_HV[502]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16478.905 1046.435 16479.185 1047.435 ;
    END
  END Data_HV[502]
  PIN Data_HV[496]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16477.785 1046.435 16478.065 1047.435 ;
    END
  END Data_HV[496]
  PIN INJ_IN[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16474.425 1046.435 16474.705 1047.435 ;
    END
  END INJ_IN[383]
  PIN nTOK_HV[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16434.105 1046.435 16434.385 1047.435 ;
    END
  END nTOK_HV[23]
  PIN BcidMtx[1150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16432.425 1046.435 16432.705 1047.435 ;
    END
  END BcidMtx[1150]
  PIN BcidMtx[1147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16429.625 1046.435 16429.905 1047.435 ;
    END
  END BcidMtx[1147]
  PIN INJ_IN[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16427.945 1046.435 16428.225 1047.435 ;
    END
  END INJ_IN[382]
  PIN Data_HV[485]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16426.265 1046.435 16426.545 1047.435 ;
    END
  END Data_HV[485]
  PIN Data_HV[499]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16423.465 1046.435 16423.745 1047.435 ;
    END
  END Data_HV[499]
  PIN Data_HV[484]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16422.345 1046.435 16422.625 1047.435 ;
    END
  END Data_HV[484]
  PIN Data_HV[500]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16421.225 1046.435 16421.505 1047.435 ;
    END
  END Data_HV[500]
  PIN DIG_MON_SEL[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16407.785 1046.435 16408.065 1047.435 ;
    END
  END DIG_MON_SEL[381]
  PIN DIG_MON_HV[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16405.545 1046.435 16405.825 1047.435 ;
    END
  END DIG_MON_HV[45]
  PIN Data_HV[474]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16400.225 1046.435 16400.505 1047.435 ;
    END
  END Data_HV[474]
  PIN Data_HV[467]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16399.105 1046.435 16399.385 1047.435 ;
    END
  END Data_HV[467]
  PIN Data_HV[482]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16372.505 1046.435 16372.785 1047.435 ;
    END
  END Data_HV[482]
  PIN nTOK_HV[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16368.585 1046.435 16368.865 1047.435 ;
    END
  END nTOK_HV[22]
  PIN BcidMtx[1144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16366.905 1046.435 16367.185 1047.435 ;
    END
  END BcidMtx[1144]
  PIN FREEZE_HV[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16365.785 1046.435 16366.065 1047.435 ;
    END
  END FREEZE_HV[22]
  PIN INJ_IN[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16362.425 1046.435 16362.705 1047.435 ;
    END
  END INJ_IN[380]
  PIN Data_HV[464]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16360.745 1046.435 16361.025 1047.435 ;
    END
  END Data_HV[464]
  PIN Data_HV[477]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16346.745 1046.435 16347.025 1047.435 ;
    END
  END Data_HV[477]
  PIN Data_HV[463]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16343.945 1046.435 16344.225 1047.435 ;
    END
  END Data_HV[463]
  PIN MASKV[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16342.265 1046.435 16342.545 1047.435 ;
    END
  END MASKV[380]
  PIN DIG_MON_HV[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16340.025 1046.435 16340.305 1047.435 ;
    END
  END DIG_MON_HV[44]
  PIN DIG_MON_SEL[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16337.785 1046.435 16338.065 1047.435 ;
    END
  END DIG_MON_SEL[379]
  PIN INJ_ROW[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16334.425 1046.435 16334.705 1047.435 ;
    END
  END INJ_ROW[189]
  PIN Data_HV[449]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16292.985 1046.435 16293.265 1047.435 ;
    END
  END Data_HV[449]
  PIN Data_HV[446]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16291.305 1046.435 16291.585 1047.435 ;
    END
  END Data_HV[446]
  PIN Data_HV[461]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16290.185 1046.435 16290.465 1047.435 ;
    END
  END Data_HV[461]
  PIN Data_HV[448]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16289.065 1046.435 16289.345 1047.435 ;
    END
  END Data_HV[448]
  PIN BcidMtx[1139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16285.145 1046.435 16285.425 1047.435 ;
    END
  END BcidMtx[1139]
  PIN BcidMtx[1137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16284.025 1046.435 16284.305 1047.435 ;
    END
  END BcidMtx[1137]
  PIN Read_HV[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16282.905 1046.435 16283.185 1047.435 ;
    END
  END Read_HV[21]
  PIN DIG_MON_SEL[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8391.945 1046.435 8392.225 1047.435 ;
    END
  END DIG_MON_SEL[181]
  PIN MASKD[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8390.825 1046.435 8391.105 1047.435 ;
    END
  END MASKD[181]
  PIN Data_PMOS[722]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8386.905 1046.435 8387.185 1047.435 ;
    END
  END Data_PMOS[722]
  PIN Data_PMOS[719]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8385.225 1046.435 8385.505 1047.435 ;
    END
  END Data_PMOS[719]
  PIN Data_PMOS[727]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8384.665 1046.435 8384.945 1047.435 ;
    END
  END Data_PMOS[727]
  PIN INJ_IN[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8381.305 1046.435 8381.585 1047.435 ;
    END
  END INJ_IN[181]
  PIN BcidMtx[544]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8365.065 1046.435 8365.345 1047.435 ;
    END
  END BcidMtx[544]
  PIN BcidMtx[543]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8364.505 1046.435 8364.785 1047.435 ;
    END
  END BcidMtx[543]
  PIN BcidMtx[540]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8361.705 1046.435 8361.985 1047.435 ;
    END
  END BcidMtx[540]
  PIN Data_PMOS[716]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8358.905 1046.435 8359.185 1047.435 ;
    END
  END Data_PMOS[716]
  PIN Data_PMOS[723]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8358.345 1046.435 8358.625 1047.435 ;
    END
  END Data_PMOS[723]
  PIN Data_PMOS[725]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8355.545 1046.435 8355.825 1047.435 ;
    END
  END Data_PMOS[725]
  PIN Data_PMOS[731]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8353.865 1046.435 8354.145 1047.435 ;
    END
  END Data_PMOS[731]
  PIN MASKV[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8314.665 1046.435 8314.945 1047.435 ;
    END
  END MASKV[180]
  PIN DIG_MON_SEL[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8310.745 1046.435 8311.025 1047.435 ;
    END
  END DIG_MON_SEL[180]
  PIN DIG_MON_PMOS[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8307.945 1046.435 8308.225 1047.435 ;
    END
  END DIG_MON_PMOS[67]
  PIN INJ_ROW[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8306.825 1046.435 8307.105 1047.435 ;
    END
  END INJ_ROW[89]
  PIN Data_PMOS[712]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8304.025 1046.435 8304.305 1047.435 ;
    END
  END Data_PMOS[712]
  PIN Data_PMOS[713]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8302.345 1046.435 8302.625 1047.435 ;
    END
  END Data_PMOS[713]
  PIN Data_PMOS[707]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8301.785 1046.435 8302.065 1047.435 ;
    END
  END Data_PMOS[707]
  PIN BcidMtx[539]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8288.905 1046.435 8289.185 1047.435 ;
    END
  END BcidMtx[539]
  PIN FREEZE_PMOS[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8287.225 1046.435 8287.505 1047.435 ;
    END
  END FREEZE_PMOS[33]
  PIN Read_PMOS[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8286.665 1046.435 8286.945 1047.435 ;
    END
  END Read_PMOS[33]
  PIN INJ_IN[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8281.905 1046.435 8282.185 1047.435 ;
    END
  END INJ_IN[178]
  PIN Data_PMOS[702]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8279.665 1046.435 8279.945 1047.435 ;
    END
  END Data_PMOS[702]
  PIN Data_PMOS[708]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8279.105 1046.435 8279.385 1047.435 ;
    END
  END Data_PMOS[708]
  PIN Data_PMOS[694]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8250.825 1046.435 8251.105 1047.435 ;
    END
  END Data_PMOS[694]
  PIN MASKV[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8249.145 1046.435 8249.425 1047.435 ;
    END
  END MASKV[178]
  PIN MASKH[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8248.585 1046.435 8248.865 1047.435 ;
    END
  END MASKH[89]
  PIN DIG_MON_SEL[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8244.665 1046.435 8244.945 1047.435 ;
    END
  END DIG_MON_SEL[177]
  PIN INJ_ROW[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8241.305 1046.435 8241.585 1047.435 ;
    END
  END INJ_ROW[88]
  PIN MASKV[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8240.745 1046.435 8241.025 1047.435 ;
    END
  END MASKV[177]
  PIN Data_PMOS[677]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8225.065 1046.435 8225.345 1047.435 ;
    END
  END Data_PMOS[677]
  PIN Data_PMOS[686]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8223.385 1046.435 8223.665 1047.435 ;
    END
  END Data_PMOS[686]
  PIN Data_PMOS[679]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8222.825 1046.435 8223.105 1047.435 ;
    END
  END Data_PMOS[679]
  PIN BcidMtx[532]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8218.345 1046.435 8218.625 1047.435 ;
    END
  END BcidMtx[532]
  PIN Read_PMOS[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8216.665 1046.435 8216.945 1047.435 ;
    END
  END Read_PMOS[32]
  PIN BcidMtx[529]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8215.545 1046.435 8215.825 1047.435 ;
    END
  END BcidMtx[529]
  PIN Data_PMOS[681]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8172.985 1046.435 8173.265 1047.435 ;
    END
  END Data_PMOS[681]
  PIN Data_PMOS[676]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8171.305 1046.435 8171.585 1047.435 ;
    END
  END Data_PMOS[676]
  PIN Data_PMOS[688]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8170.745 1046.435 8171.025 1047.435 ;
    END
  END Data_PMOS[688]
  PIN MASKV[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8167.945 1046.435 8168.225 1047.435 ;
    END
  END MASKV[176]
  PIN DIG_MON_PMOS[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8165.705 1046.435 8165.985 1047.435 ;
    END
  END DIG_MON_PMOS[64]
  PIN INJ_ROW[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8151.705 1046.435 8151.985 1047.435 ;
    END
  END INJ_ROW[87]
  PIN Data_PMOS[659]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8150.025 1046.435 8150.305 1047.435 ;
    END
  END Data_PMOS[659]
  PIN Data_PMOS[663]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8149.465 1046.435 8149.745 1047.435 ;
    END
  END Data_PMOS[663]
  PIN Data_PMOS[665]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8146.665 1046.435 8146.945 1047.435 ;
    END
  END Data_PMOS[665]
  PIN INJ_IN[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8142.465 1046.435 8142.745 1047.435 ;
    END
  END INJ_IN[175]
  PIN nTOK_PMOS[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8141.345 1046.435 8141.625 1047.435 ;
    END
  END nTOK_PMOS[31]
  PIN BcidMtx[524]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8111.945 1046.435 8112.225 1047.435 ;
    END
  END BcidMtx[524]
  PIN BcidMtx[522]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8110.825 1046.435 8111.105 1047.435 ;
    END
  END BcidMtx[522]
  PIN Data_PMOS[654]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8108.585 1046.435 8108.865 1047.435 ;
    END
  END Data_PMOS[654]
  PIN Data_PMOS[655]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8105.785 1046.435 8106.065 1047.435 ;
    END
  END Data_PMOS[655]
  PIN Data_PMOS[652]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8104.105 1046.435 8104.385 1047.435 ;
    END
  END Data_PMOS[652]
  PIN Data_PMOS[651]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8103.545 1046.435 8103.825 1047.435 ;
    END
  END Data_PMOS[651]
  PIN DIG_MON_PMOS[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8100.185 1046.435 8100.465 1047.435 ;
    END
  END DIG_MON_PMOS[62]
  PIN DIG_MON_SEL[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8085.065 1046.435 8085.345 1047.435 ;
    END
  END DIG_MON_SEL[173]
  PIN MASKD[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8083.945 1046.435 8084.225 1047.435 ;
    END
  END MASKD[173]
  PIN Data_PMOS[638]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8080.025 1046.435 8080.305 1047.435 ;
    END
  END Data_PMOS[638]
  PIN Data_PMOS[635]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8078.345 1046.435 8078.625 1047.435 ;
    END
  END Data_PMOS[635]
  PIN Data_PMOS[643]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8077.785 1046.435 8078.065 1047.435 ;
    END
  END Data_PMOS[643]
  PIN INJ_IN[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8074.425 1046.435 8074.705 1047.435 ;
    END
  END INJ_IN[173]
  PIN BcidMtx[520]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8032.425 1046.435 8032.705 1047.435 ;
    END
  END BcidMtx[520]
  PIN BcidMtx[519]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8031.865 1046.435 8032.145 1047.435 ;
    END
  END BcidMtx[519]
  PIN BcidMtx[516]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8029.065 1046.435 8029.345 1047.435 ;
    END
  END BcidMtx[516]
  PIN Data_PMOS[632]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8026.265 1046.435 8026.545 1047.435 ;
    END
  END Data_PMOS[632]
  PIN Data_PMOS[639]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8025.705 1046.435 8025.985 1047.435 ;
    END
  END Data_PMOS[639]
  PIN Data_PMOS[641]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8022.905 1046.435 8023.185 1047.435 ;
    END
  END Data_PMOS[641]
  PIN Data_PMOS[647]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8021.225 1046.435 8021.505 1047.435 ;
    END
  END Data_PMOS[647]
  PIN MASKV[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8012.265 1046.435 8012.545 1047.435 ;
    END
  END MASKV[172]
  PIN DIG_MON_SEL[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8008.345 1046.435 8008.625 1047.435 ;
    END
  END DIG_MON_SEL[172]
  PIN DIG_MON_PMOS[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8005.545 1046.435 8005.825 1047.435 ;
    END
  END DIG_MON_PMOS[59]
  PIN MASKV[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8001.905 1046.435 8002.185 1047.435 ;
    END
  END MASKV[171]
  PIN Data_PMOS[614]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7999.105 1046.435 7999.385 1047.435 ;
    END
  END Data_PMOS[614]
  PIN Data_PMOS[629]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7972.505 1046.435 7972.785 1047.435 ;
    END
  END Data_PMOS[629]
  PIN Data_PMOS[616]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7971.385 1046.435 7971.665 1047.435 ;
    END
  END Data_PMOS[616]
  PIN MASKH[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18807.385 1046.435 18807.665 1047.435 ;
    END
  END MASKH[221]
  PIN FREEZE_PMOS[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7965.785 1046.435 7966.065 1047.435 ;
    END
  END FREEZE_PMOS[29]
  PIN Read_PMOS[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7965.225 1046.435 7965.505 1047.435 ;
    END
  END Read_PMOS[29]
  PIN BcidMtx[510]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7963.545 1046.435 7963.825 1047.435 ;
    END
  END BcidMtx[510]
  PIN Data_PMOS[611]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7960.745 1046.435 7961.025 1047.435 ;
    END
  END Data_PMOS[611]
  PIN Data_PMOS[619]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7946.185 1046.435 7946.465 1047.435 ;
    END
  END Data_PMOS[619]
  PIN Data_PMOS[620]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7944.505 1046.435 7944.785 1047.435 ;
    END
  END Data_PMOS[620]
  PIN Data_PMOS[626]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7942.825 1046.435 7943.105 1047.435 ;
    END
  END Data_PMOS[626]
  PIN MASKD[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7941.145 1046.435 7941.425 1047.435 ;
    END
  END MASKD[170]
  PIN DIG_MON_SEL[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7937.785 1046.435 7938.065 1047.435 ;
    END
  END DIG_MON_SEL[169]
  PIN DIG_MON_PMOS[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7935.545 1046.435 7935.825 1047.435 ;
    END
  END DIG_MON_PMOS[57]
  PIN Data_PMOS[606]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7893.545 1046.435 7893.825 1047.435 ;
    END
  END Data_PMOS[606]
  PIN Data_PMOS[593]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7891.305 1046.435 7891.585 1047.435 ;
    END
  END Data_PMOS[593]
  PIN Data_PMOS[602]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7889.625 1046.435 7889.905 1047.435 ;
    END
  END Data_PMOS[602]
  PIN Data_PMOS[594]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7888.505 1046.435 7888.785 1047.435 ;
    END
  END Data_PMOS[594]
  PIN MASKD[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18806.825 1046.435 18807.105 1047.435 ;
    END
  END MASKD[442]
  PIN FREEZE_PMOS[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7883.465 1046.435 7883.745 1047.435 ;
    END
  END FREEZE_PMOS[28]
  PIN BcidMtx[506]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7882.345 1046.435 7882.625 1047.435 ;
    END
  END BcidMtx[506]
  PIN Data_PMOS[591]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7870.585 1046.435 7870.865 1047.435 ;
    END
  END Data_PMOS[591]
  PIN Data_PMOS[603]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7868.905 1046.435 7869.185 1047.435 ;
    END
  END Data_PMOS[603]
  PIN Data_PMOS[604]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7867.225 1046.435 7867.505 1047.435 ;
    END
  END Data_PMOS[604]
  PIN Data_PMOS[588]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7865.545 1046.435 7865.825 1047.435 ;
    END
  END Data_PMOS[588]
  PIN MASKH[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7861.905 1046.435 7862.185 1047.435 ;
    END
  END MASKH[84]
  PIN MASKD[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8950.825 1046.435 8951.105 1047.435 ;
    END
  END MASKD[195]
  PIN DIG_MON_PMOS[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8980.225 1046.435 8980.505 1047.435 ;
    END
  END DIG_MON_PMOS[84]
  PIN FREEZE_PMOS[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9233.065 1046.435 9233.345 1047.435 ;
    END
  END FREEZE_PMOS[45]
  PIN DIG_MON_HV[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18801.225 1046.435 18801.505 1047.435 ;
    END
  END DIG_MON_HV[105]
  PIN MASKV[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10068.025 1046.435 10068.305 1047.435 ;
    END
  END MASKV[223]
  PIN Data_PMOS[1167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10066.345 1046.435 10066.625 1047.435 ;
    END
  END Data_PMOS[1167]
  PIN Data_PMOS[1168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10064.665 1046.435 10064.945 1047.435 ;
    END
  END Data_PMOS[1168]
  PIN Data_PMOS[1162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10062.985 1046.435 10063.265 1047.435 ;
    END
  END Data_PMOS[1162]
  PIN nTOK_PMOS[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10060.185 1046.435 10060.465 1047.435 ;
    END
  END nTOK_PMOS[55]
  PIN BcidMtx[669]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10044.505 1046.435 10044.785 1047.435 ;
    END
  END BcidMtx[669]
  PIN BcidMtx[668]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10042.825 1046.435 10043.105 1047.435 ;
    END
  END BcidMtx[668]
  PIN INJ_IN[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10040.585 1046.435 10040.865 1047.435 ;
    END
  END INJ_IN[222]
  PIN Data_PMOS[1164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10038.345 1046.435 10038.625 1047.435 ;
    END
  END Data_PMOS[1164]
  PIN Data_PMOS[1159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10036.665 1046.435 10036.945 1047.435 ;
    END
  END Data_PMOS[1159]
  PIN Data_PMOS[1156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10034.985 1046.435 10035.265 1047.435 ;
    END
  END Data_PMOS[1156]
  PIN MASKV[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9994.665 1046.435 9994.945 1047.435 ;
    END
  END MASKV[222]
  PIN DIG_MON_PMOS[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9992.425 1046.435 9992.705 1047.435 ;
    END
  END DIG_MON_PMOS[110]
  PIN DIG_MON_SEL[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9990.185 1046.435 9990.465 1047.435 ;
    END
  END DIG_MON_SEL[221]
  PIN INJ_ROW[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9986.825 1046.435 9987.105 1047.435 ;
    END
  END INJ_ROW[110]
  PIN Data_PMOS[1152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9985.705 1046.435 9985.985 1047.435 ;
    END
  END Data_PMOS[1152]
  PIN Data_PMOS[1153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9984.025 1046.435 9984.305 1047.435 ;
    END
  END Data_PMOS[1153]
  PIN Data_PMOS[1154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9982.345 1046.435 9982.625 1047.435 ;
    END
  END Data_PMOS[1154]
  PIN Data_PMOS[1140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9972.265 1046.435 9972.545 1047.435 ;
    END
  END Data_PMOS[1140]
  PIN BcidMtx[665]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9968.905 1046.435 9969.185 1047.435 ;
    END
  END BcidMtx[665]
  PIN FREEZE_PMOS[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9967.225 1046.435 9967.505 1047.435 ;
    END
  END FREEZE_PMOS[54]
  PIN BcidMtx[661]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9965.545 1046.435 9965.825 1047.435 ;
    END
  END BcidMtx[661]
  PIN Data_PMOS[1137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9960.785 1046.435 9961.065 1047.435 ;
    END
  END Data_PMOS[1137]
  PIN Data_PMOS[1149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9959.105 1046.435 9959.385 1047.435 ;
    END
  END Data_PMOS[1149]
  PIN Data_PMOS[1150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9931.945 1046.435 9932.225 1047.435 ;
    END
  END Data_PMOS[1150]
  PIN Data_PMOS[1134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9930.265 1046.435 9930.545 1047.435 ;
    END
  END Data_PMOS[1134]
  PIN MASKH[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9928.585 1046.435 9928.865 1047.435 ;
    END
  END MASKH[110]
  PIN DIG_MON_SEL[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9925.225 1046.435 9925.505 1047.435 ;
    END
  END DIG_MON_SEL[220]
  PIN MASKD[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9923.545 1046.435 9923.825 1047.435 ;
    END
  END MASKD[219]
  PIN MASKV[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9920.745 1046.435 9921.025 1047.435 ;
    END
  END MASKV[219]
  PIN Data_PMOS[1125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9906.185 1046.435 9906.465 1047.435 ;
    END
  END Data_PMOS[1125]
  PIN Data_PMOS[1118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9905.065 1046.435 9905.345 1047.435 ;
    END
  END Data_PMOS[1118]
  PIN Data_PMOS[1120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9902.825 1046.435 9903.105 1047.435 ;
    END
  END Data_PMOS[1120]
  PIN nTOK_PMOS[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9900.025 1046.435 9900.305 1047.435 ;
    END
  END nTOK_PMOS[53]
  PIN FREEZE_PMOS[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9897.225 1046.435 9897.505 1047.435 ;
    END
  END FREEZE_PMOS[53]
  PIN BcidMtx[656]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9896.105 1046.435 9896.385 1047.435 ;
    END
  END BcidMtx[656]
  PIN INJ_IN[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9893.865 1046.435 9894.145 1047.435 ;
    END
  END INJ_IN[218]
  PIN Data_PMOS[1122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9852.985 1046.435 9853.265 1047.435 ;
    END
  END Data_PMOS[1122]
  PIN Data_PMOS[1117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9851.305 1046.435 9851.585 1047.435 ;
    END
  END Data_PMOS[1117]
  PIN Data_PMOS[1114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9849.625 1046.435 9849.905 1047.435 ;
    END
  END Data_PMOS[1114]
  PIN MASKV[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9847.945 1046.435 9848.225 1047.435 ;
    END
  END MASKV[218]
  PIN DIG_MON_PMOS[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9845.705 1046.435 9845.985 1047.435 ;
    END
  END DIG_MON_PMOS[106]
  PIN DIG_MON_SEL[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9844.025 1046.435 9844.305 1047.435 ;
    END
  END DIG_MON_SEL[218]
  PIN INJ_ROW[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9831.705 1046.435 9831.985 1047.435 ;
    END
  END INJ_ROW[108]
  PIN Data_PMOS[1100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9830.025 1046.435 9830.305 1047.435 ;
    END
  END Data_PMOS[1100]
  PIN Data_PMOS[1111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9828.905 1046.435 9829.185 1047.435 ;
    END
  END Data_PMOS[1111]
  PIN Data_PMOS[1105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9827.785 1046.435 9828.065 1047.435 ;
    END
  END Data_PMOS[1105]
  PIN INJ_IN[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9822.465 1046.435 9822.745 1047.435 ;
    END
  END INJ_IN[217]
  PIN BcidMtx[653]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9820.225 1046.435 9820.505 1047.435 ;
    END
  END BcidMtx[653]
  PIN BcidMtx[650]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9791.945 1046.435 9792.225 1047.435 ;
    END
  END BcidMtx[650]
  PIN INJ_IN[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9789.705 1046.435 9789.985 1047.435 ;
    END
  END INJ_IN[216]
  PIN Data_PMOS[1094]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9788.025 1046.435 9788.305 1047.435 ;
    END
  END Data_PMOS[1094]
  PIN Data_PMOS[1096]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9785.785 1046.435 9786.065 1047.435 ;
    END
  END Data_PMOS[1096]
  PIN Data_PMOS[1093]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9784.105 1046.435 9784.385 1047.435 ;
    END
  END Data_PMOS[1093]
  PIN Data_PMOS[1109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9782.985 1046.435 9783.265 1047.435 ;
    END
  END Data_PMOS[1109]
  PIN Data_HV[1062]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18640.225 1046.435 18640.505 1047.435 ;
    END
  END Data_HV[1062]
  PIN DIG_MON_SEL[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9765.065 1046.435 9765.345 1047.435 ;
    END
  END DIG_MON_SEL[215]
  PIN MASKV[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9761.145 1046.435 9761.425 1047.435 ;
    END
  END MASKV[215]
  PIN Data_PMOS[1083]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9759.465 1046.435 9759.745 1047.435 ;
    END
  END Data_PMOS[1083]
  PIN Data_PMOS[1076]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9758.345 1046.435 9758.625 1047.435 ;
    END
  END Data_PMOS[1076]
  PIN Data_PMOS[1078]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9756.105 1046.435 9756.385 1047.435 ;
    END
  END Data_PMOS[1078]
  PIN nTOK_PMOS[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9714.105 1046.435 9714.385 1047.435 ;
    END
  END nTOK_PMOS[51]
  PIN BcidMtx[646]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9712.425 1046.435 9712.705 1047.435 ;
    END
  END BcidMtx[646]
  PIN BcidMtx[644]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9710.185 1046.435 9710.465 1047.435 ;
    END
  END BcidMtx[644]
  PIN INJ_IN[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9707.945 1046.435 9708.225 1047.435 ;
    END
  END INJ_IN[214]
  PIN Data_PMOS[1073]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9706.265 1046.435 9706.545 1047.435 ;
    END
  END Data_PMOS[1073]
  PIN Data_PMOS[1075]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9704.025 1046.435 9704.305 1047.435 ;
    END
  END Data_PMOS[1075]
  PIN Data_PMOS[1072]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9702.345 1046.435 9702.625 1047.435 ;
    END
  END Data_PMOS[1072]
  PIN Data_PMOS[1088]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9701.225 1046.435 9701.505 1047.435 ;
    END
  END Data_PMOS[1088]
  PIN DIG_MON_PMOS[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9690.025 1046.435 9690.305 1047.435 ;
    END
  END DIG_MON_PMOS[102]
  PIN DIG_MON_SEL[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9688.345 1046.435 9688.625 1047.435 ;
    END
  END DIG_MON_SEL[214]
  PIN DIG_MON_PMOS[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9685.545 1046.435 9685.825 1047.435 ;
    END
  END DIG_MON_PMOS[101]
  PIN Data_PMOS[1058]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9680.785 1046.435 9681.065 1047.435 ;
    END
  END Data_PMOS[1058]
  PIN Data_PMOS[1055]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9679.105 1046.435 9679.385 1047.435 ;
    END
  END Data_PMOS[1055]
  PIN Data_PMOS[1070]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9652.505 1046.435 9652.785 1047.435 ;
    END
  END Data_PMOS[1070]
  PIN INJ_IN[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9649.705 1046.435 9649.985 1047.435 ;
    END
  END INJ_IN[213]
  PIN BcidMtx[641]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9647.465 1046.435 9647.745 1047.435 ;
    END
  END BcidMtx[641]
  PIN BcidMtx[639]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9646.345 1046.435 9646.625 1047.435 ;
    END
  END BcidMtx[639]
  PIN BcidMtx[636]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9643.545 1046.435 9643.825 1047.435 ;
    END
  END BcidMtx[636]
  PIN Data_PMOS[1053]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9641.305 1046.435 9641.585 1047.435 ;
    END
  END Data_PMOS[1053]
  PIN Data_PMOS[1059]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9640.185 1046.435 9640.465 1047.435 ;
    END
  END Data_PMOS[1059]
  PIN Data_PMOS[1061]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9624.505 1046.435 9624.785 1047.435 ;
    END
  END Data_PMOS[1061]
  PIN Data_PMOS[1050]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9623.385 1046.435 9623.665 1047.435 ;
    END
  END Data_PMOS[1050]
  PIN MASKV[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9622.265 1046.435 9622.545 1047.435 ;
    END
  END MASKV[212]
  PIN DIG_MON_SEL[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9617.785 1046.435 9618.065 1047.435 ;
    END
  END DIG_MON_SEL[211]
  PIN Data_HV[1110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18790.585 1046.435 18790.865 1047.435 ;
    END
  END Data_HV[1110]
  PIN Data_PMOS[1037]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9572.985 1046.435 9573.265 1047.435 ;
    END
  END Data_PMOS[1037]
  PIN Data_PMOS[1048]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9571.865 1046.435 9572.145 1047.435 ;
    END
  END Data_PMOS[1048]
  PIN Data_PMOS[1034]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9571.305 1046.435 9571.585 1047.435 ;
    END
  END Data_PMOS[1034]
  PIN Data_PMOS[1035]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9568.505 1046.435 9568.785 1047.435 ;
    END
  END Data_PMOS[1035]
  PIN BcidMtx[635]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9565.145 1046.435 9565.425 1047.435 ;
    END
  END BcidMtx[635]
  PIN BcidMtx[634]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9564.585 1046.435 9564.865 1047.435 ;
    END
  END BcidMtx[634]
  PIN BcidMtx[631]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9561.785 1046.435 9562.065 1047.435 ;
    END
  END BcidMtx[631]
  PIN Data_PMOS[1032]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9550.585 1046.435 9550.865 1047.435 ;
    END
  END Data_PMOS[1032]
  PIN Data_PMOS[1031]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9550.025 1046.435 9550.305 1047.435 ;
    END
  END Data_PMOS[1031]
  PIN Data_PMOS[1045]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9547.225 1046.435 9547.505 1047.435 ;
    END
  END Data_PMOS[1045]
  PIN Data_PMOS[1029]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9545.545 1046.435 9545.825 1047.435 ;
    END
  END Data_PMOS[1029]
  PIN MASKD[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8421.345 1046.435 8421.625 1047.435 ;
    END
  END MASKD[182]
  PIN DIG_MON_SEL[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8418.545 1046.435 8418.825 1047.435 ;
    END
  END DIG_MON_SEL[182]
  PIN MASKD[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9510.825 1046.435 9511.105 1047.435 ;
    END
  END MASKD[209]
  PIN INJ_ROW[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9508.585 1046.435 9508.865 1047.435 ;
    END
  END INJ_ROW[104]
  PIN Data_PMOS[1027]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9505.785 1046.435 9506.065 1047.435 ;
    END
  END Data_PMOS[1027]
  PIN Data_PMOS[1021]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9504.665 1046.435 9504.945 1047.435 ;
    END
  END Data_PMOS[1021]
  PIN Data_PMOS[1014]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9502.425 1046.435 9502.705 1047.435 ;
    END
  END Data_PMOS[1014]
  PIN BcidMtx[629]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9485.625 1046.435 9485.905 1047.435 ;
    END
  END BcidMtx[629]
  PIN BcidMtx[627]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9484.505 1046.435 9484.785 1047.435 ;
    END
  END BcidMtx[627]
  PIN BcidMtx[625]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9482.265 1046.435 9482.545 1047.435 ;
    END
  END BcidMtx[625]
  PIN Data_PMOS[1011]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9479.465 1046.435 9479.745 1047.435 ;
    END
  END Data_PMOS[1011]
  PIN Data_PMOS[1017]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9478.345 1046.435 9478.625 1047.435 ;
    END
  END Data_PMOS[1017]
  PIN Data_PMOS[1024]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9476.105 1046.435 9476.385 1047.435 ;
    END
  END Data_PMOS[1024]
  PIN Data_PMOS[1008]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9474.425 1046.435 9474.705 1047.435 ;
    END
  END Data_PMOS[1008]
  PIN MASKV[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9434.665 1046.435 9434.945 1047.435 ;
    END
  END MASKV[208]
  PIN MASKD[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9433.545 1046.435 9433.825 1047.435 ;
    END
  END MASKD[208]
  PIN MASKD[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9429.065 1046.435 9429.345 1047.435 ;
    END
  END MASKD[207]
  PIN INJ_ROW[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9426.825 1046.435 9427.105 1047.435 ;
    END
  END INJ_ROW[103]
  PIN Data_PMOS[995]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9425.145 1046.435 9425.425 1047.435 ;
    END
  END Data_PMOS[995]
  PIN Data_PMOS[1000]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9422.905 1046.435 9423.185 1047.435 ;
    END
  END Data_PMOS[1000]
  PIN DIG_MON_SEL[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18804.025 1046.435 18804.305 1047.435 ;
    END
  END DIG_MON_SEL[442]
  PIN INJ_IN[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9411.145 1046.435 9411.425 1047.435 ;
    END
  END INJ_IN[207]
  PIN BcidMtx[622]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9408.345 1046.435 9408.625 1047.435 ;
    END
  END BcidMtx[622]
  PIN Read_PMOS[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9406.665 1046.435 9406.945 1047.435 ;
    END
  END Read_PMOS[47]
  PIN BcidMtx[618]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9404.985 1046.435 9405.265 1047.435 ;
    END
  END BcidMtx[618]
  PIN Data_PMOS[989]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9400.225 1046.435 9400.505 1047.435 ;
    END
  END Data_PMOS[989]
  PIN Data_PMOS[1002]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9399.105 1046.435 9399.385 1047.435 ;
    END
  END Data_PMOS[1002]
  PIN Data_PMOS[1003]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9371.945 1046.435 9372.225 1047.435 ;
    END
  END Data_PMOS[1003]
  PIN Data_PMOS[987]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9370.265 1046.435 9370.545 1047.435 ;
    END
  END Data_PMOS[987]
  PIN MASKH[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9368.585 1046.435 9368.865 1047.435 ;
    END
  END MASKH[103]
  PIN MASKD[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9363.545 1046.435 9363.825 1047.435 ;
    END
  END MASKD[205]
  PIN MASKV[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9360.745 1046.435 9361.025 1047.435 ;
    END
  END MASKV[205]
  PIN Data_PMOS[978]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9346.185 1046.435 9346.465 1047.435 ;
    END
  END Data_PMOS[978]
  PIN Data_PMOS[979]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9344.505 1046.435 9344.785 1047.435 ;
    END
  END Data_PMOS[979]
  PIN Data_PMOS[973]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9342.825 1046.435 9343.105 1047.435 ;
    END
  END Data_PMOS[973]
  PIN INJ_IN[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9341.145 1046.435 9341.425 1047.435 ;
    END
  END INJ_IN[205]
  PIN BcidMtx[615]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9337.785 1046.435 9338.065 1047.435 ;
    END
  END BcidMtx[615]
  PIN BcidMtx[614]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9336.105 1046.435 9336.385 1047.435 ;
    END
  END BcidMtx[614]
  PIN BcidMtx[612]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9334.985 1046.435 9335.265 1047.435 ;
    END
  END BcidMtx[612]
  PIN Data_PMOS[975]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9292.985 1046.435 9293.265 1047.435 ;
    END
  END Data_PMOS[975]
  PIN Data_PMOS[970]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9291.305 1046.435 9291.585 1047.435 ;
    END
  END Data_PMOS[970]
  PIN Data_PMOS[977]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9290.185 1046.435 9290.465 1047.435 ;
    END
  END Data_PMOS[977]
  PIN MASKV[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9287.945 1046.435 9288.225 1047.435 ;
    END
  END MASKV[204]
  PIN DIG_MON_PMOS[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9285.705 1046.435 9285.985 1047.435 ;
    END
  END DIG_MON_PMOS[92]
  PIN DIG_MON_SEL[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9283.465 1046.435 9283.745 1047.435 ;
    END
  END DIG_MON_SEL[203]
  PIN INJ_ROW[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9271.705 1046.435 9271.985 1047.435 ;
    END
  END INJ_ROW[101]
  PIN Data_PMOS[953]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9270.025 1046.435 9270.305 1047.435 ;
    END
  END Data_PMOS[953]
  PIN Data_PMOS[950]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9268.345 1046.435 9268.625 1047.435 ;
    END
  END Data_PMOS[950]
  PIN Data_PMOS[959]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9266.665 1046.435 9266.945 1047.435 ;
    END
  END Data_PMOS[959]
  PIN INJ_IN[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9262.465 1046.435 9262.745 1047.435 ;
    END
  END INJ_IN[203]
  PIN BcidMtx[611]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9260.225 1046.435 9260.505 1047.435 ;
    END
  END BcidMtx[611]
  PIN BcidMtx[608]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9231.945 1046.435 9232.225 1047.435 ;
    END
  END BcidMtx[608]
  PIN INJ_IN[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9229.705 1046.435 9229.985 1047.435 ;
    END
  END INJ_IN[202]
  PIN Data_PMOS[954]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9227.465 1046.435 9227.745 1047.435 ;
    END
  END Data_PMOS[954]
  PIN Data_PMOS[949]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9225.785 1046.435 9226.065 1047.435 ;
    END
  END Data_PMOS[949]
  PIN Data_PMOS[946]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9224.105 1046.435 9224.385 1047.435 ;
    END
  END Data_PMOS[946]
  PIN MASKV[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9222.425 1046.435 9222.705 1047.435 ;
    END
  END MASKV[202]
  PIN DIG_MON_PMOS[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9220.185 1046.435 9220.465 1047.435 ;
    END
  END DIG_MON_PMOS[90]
  PIN DIG_MON_SEL[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9205.065 1046.435 9205.345 1047.435 ;
    END
  END DIG_MON_SEL[201]
  PIN MASKD[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9203.945 1046.435 9204.225 1047.435 ;
    END
  END MASKD[201]
  PIN Data_PMOS[942]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9200.585 1046.435 9200.865 1047.435 ;
    END
  END Data_PMOS[942]
  PIN Data_PMOS[943]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9198.905 1046.435 9199.185 1047.435 ;
    END
  END Data_PMOS[943]
  PIN Data_PMOS[937]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9197.785 1046.435 9198.065 1047.435 ;
    END
  END Data_PMOS[937]
  PIN Data_PMOS[930]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9195.545 1046.435 9195.825 1047.435 ;
    END
  END Data_PMOS[930]
  PIN BcidMtx[605]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9152.985 1046.435 9153.265 1047.435 ;
    END
  END BcidMtx[605]
  PIN FREEZE_PMOS[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9151.305 1046.435 9151.585 1047.435 ;
    END
  END FREEZE_PMOS[44]
  PIN BcidMtx[601]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9149.625 1046.435 9149.905 1047.435 ;
    END
  END BcidMtx[601]
  PIN Data_PMOS[927]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9146.825 1046.435 9147.105 1047.435 ;
    END
  END Data_PMOS[927]
  PIN Data_PMOS[939]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9145.145 1046.435 9145.425 1047.435 ;
    END
  END Data_PMOS[939]
  PIN Data_PMOS[940]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9143.465 1046.435 9143.745 1047.435 ;
    END
  END Data_PMOS[940]
  PIN Data_PMOS[924]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9141.785 1046.435 9142.065 1047.435 ;
    END
  END Data_PMOS[924]
  PIN MASKV[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9132.265 1046.435 9132.545 1047.435 ;
    END
  END MASKV[200]
  PIN MASKD[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9126.665 1046.435 9126.945 1047.435 ;
    END
  END MASKD[199]
  PIN DIG_MON_PMOS[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9125.545 1046.435 9125.825 1047.435 ;
    END
  END DIG_MON_PMOS[87]
  PIN Data_PMOS[921]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9121.345 1046.435 9121.625 1047.435 ;
    END
  END Data_PMOS[921]
  PIN Data_PMOS[922]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9119.665 1046.435 9119.945 1047.435 ;
    END
  END Data_PMOS[922]
  PIN Data_PMOS[916]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9093.065 1046.435 9093.345 1047.435 ;
    END
  END Data_PMOS[916]
  PIN Data_PMOS[909]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9090.825 1046.435 9091.105 1047.435 ;
    END
  END Data_PMOS[909]
  PIN BcidMtx[599]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9087.465 1046.435 9087.745 1047.435 ;
    END
  END BcidMtx[599]
  PIN BcidMtx[597]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9086.345 1046.435 9086.625 1047.435 ;
    END
  END BcidMtx[597]
  PIN BcidMtx[595]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9084.105 1046.435 9084.385 1047.435 ;
    END
  END BcidMtx[595]
  PIN Data_PMOS[906]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9081.305 1046.435 9081.585 1047.435 ;
    END
  END Data_PMOS[906]
  PIN Data_PMOS[912]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9080.185 1046.435 9080.465 1047.435 ;
    END
  END Data_PMOS[912]
  PIN Data_PMOS[919]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9065.065 1046.435 9065.345 1047.435 ;
    END
  END Data_PMOS[919]
  PIN Data_PMOS[903]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9063.385 1046.435 9063.665 1047.435 ;
    END
  END Data_PMOS[903]
  PIN MASKH[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9061.705 1046.435 9061.985 1047.435 ;
    END
  END MASKH[99]
  PIN MASKD[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9056.665 1046.435 9056.945 1047.435 ;
    END
  END MASKD[197]
  PIN MASKV[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9053.865 1046.435 9054.145 1047.435 ;
    END
  END MASKV[197]
  PIN Data_PMOS[894]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9012.425 1046.435 9012.705 1047.435 ;
    END
  END Data_PMOS[894]
  PIN Data_PMOS[895]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9010.745 1046.435 9011.025 1047.435 ;
    END
  END Data_PMOS[895]
  PIN Data_PMOS[889]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9009.065 1046.435 9009.345 1047.435 ;
    END
  END Data_PMOS[889]
  PIN nTOK_PMOS[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9006.265 1046.435 9006.545 1047.435 ;
    END
  END nTOK_PMOS[42]
  PIN BcidMtx[591]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9004.025 1046.435 9004.305 1047.435 ;
    END
  END BcidMtx[591]
  PIN BcidMtx[590]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9002.345 1046.435 9002.625 1047.435 ;
    END
  END BcidMtx[590]
  PIN INJ_IN[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8991.705 1046.435 8991.985 1047.435 ;
    END
  END INJ_IN[196]
  PIN Data_PMOS[891]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8989.465 1046.435 8989.745 1047.435 ;
    END
  END Data_PMOS[891]
  PIN Data_PMOS[898]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8987.225 1046.435 8987.505 1047.435 ;
    END
  END Data_PMOS[898]
  PIN Data_PMOS[883]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8986.105 1046.435 8986.385 1047.435 ;
    END
  END Data_PMOS[883]
  PIN MASKV[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8982.465 1046.435 8982.745 1047.435 ;
    END
  END MASKV[196]
  PIN Data_HV[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15150.025 1046.435 15150.305 1047.435 ;
    END
  END Data_HV[149]
  PIN Data_HV[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15148.345 1046.435 15148.625 1047.435 ;
    END
  END Data_HV[157]
  PIN Data_HV[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15146.665 1046.435 15146.945 1047.435 ;
    END
  END Data_HV[158]
  PIN Data_HV[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15145.545 1046.435 15145.825 1047.435 ;
    END
  END Data_HV[147]
  PIN MASKD[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15141.345 1046.435 15141.625 1047.435 ;
    END
  END MASKD[350]
  PIN DIG_MON_SEL[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15138.545 1046.435 15138.825 1047.435 ;
    END
  END DIG_MON_SEL[350]
  PIN DIG_MON_SEL[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16231.945 1046.435 16232.225 1047.435 ;
    END
  END DIG_MON_SEL[377]
  PIN MASKV[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16228.025 1046.435 16228.305 1047.435 ;
    END
  END MASKV[377]
  PIN Data_HV[432]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16226.345 1046.435 16226.625 1047.435 ;
    END
  END Data_HV[432]
  PIN Data_HV[433]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16224.665 1046.435 16224.945 1047.435 ;
    END
  END Data_HV[433]
  PIN Data_HV[427]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16222.985 1046.435 16223.265 1047.435 ;
    END
  END Data_HV[427]
  PIN nTOK_HV[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16220.185 1046.435 16220.465 1047.435 ;
    END
  END nTOK_HV[20]
  PIN BcidMtx[1131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16204.505 1046.435 16204.785 1047.435 ;
    END
  END BcidMtx[1131]
  PIN BcidMtx[1130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16202.825 1046.435 16203.105 1047.435 ;
    END
  END BcidMtx[1130]
  PIN INJ_IN[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16200.585 1046.435 16200.865 1047.435 ;
    END
  END INJ_IN[376]
  PIN Data_HV[429]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16198.345 1046.435 16198.625 1047.435 ;
    END
  END Data_HV[429]
  PIN Data_HV[424]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16196.665 1046.435 16196.945 1047.435 ;
    END
  END Data_HV[424]
  PIN Data_HV[421]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16194.985 1046.435 16195.265 1047.435 ;
    END
  END Data_HV[421]
  PIN MASKV[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16154.665 1046.435 16154.945 1047.435 ;
    END
  END MASKV[376]
  PIN DIG_MON_HV[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16152.425 1046.435 16152.705 1047.435 ;
    END
  END DIG_MON_HV[40]
  PIN DIG_MON_SEL[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16150.185 1046.435 16150.465 1047.435 ;
    END
  END DIG_MON_SEL[375]
  PIN MASKV[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16146.265 1046.435 16146.545 1047.435 ;
    END
  END MASKV[375]
  PIN Data_HV[407]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16145.145 1046.435 16145.425 1047.435 ;
    END
  END Data_HV[407]
  PIN Data_HV[404]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16143.465 1046.435 16143.745 1047.435 ;
    END
  END Data_HV[404]
  PIN Data_HV[413]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16141.785 1046.435 16142.065 1047.435 ;
    END
  END Data_HV[413]
  PIN INJ_IN[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16131.145 1046.435 16131.425 1047.435 ;
    END
  END INJ_IN[375]
  PIN BcidMtx[1126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16128.345 1046.435 16128.625 1047.435 ;
    END
  END BcidMtx[1126]
  PIN Read_HV[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16126.665 1046.435 16126.945 1047.435 ;
    END
  END Read_HV[19]
  PIN BcidMtx[1122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16124.985 1046.435 16125.265 1047.435 ;
    END
  END BcidMtx[1122]
  PIN Data_HV[401]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16120.225 1046.435 16120.505 1047.435 ;
    END
  END Data_HV[401]
  PIN Data_HV[409]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16118.545 1046.435 16118.825 1047.435 ;
    END
  END Data_HV[409]
  PIN Data_HV[410]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16091.385 1046.435 16091.665 1047.435 ;
    END
  END Data_HV[410]
  PIN Data_HV[416]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16089.705 1046.435 16089.985 1047.435 ;
    END
  END Data_HV[416]
  PIN MASKD[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16088.025 1046.435 16088.305 1047.435 ;
    END
  END MASKD[374]
  PIN DIG_MON_SEL[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16085.225 1046.435 16085.505 1047.435 ;
    END
  END DIG_MON_SEL[374]
  PIN DIG_MON_HV[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16082.425 1046.435 16082.705 1047.435 ;
    END
  END DIG_MON_HV[37]
  PIN Data_HV[396]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16080.185 1046.435 16080.465 1047.435 ;
    END
  END Data_HV[396]
  PIN Data_HV[386]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16079.625 1046.435 16079.905 1047.435 ;
    END
  END Data_HV[386]
  PIN Data_HV[398]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16063.945 1046.435 16064.225 1047.435 ;
    END
  END Data_HV[398]
  PIN Data_HV[384]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16062.265 1046.435 16062.545 1047.435 ;
    END
  END Data_HV[384]
  PIN BcidMtx[1121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16058.905 1046.435 16059.185 1047.435 ;
    END
  END BcidMtx[1121]
  PIN FREEZE_HV[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16057.225 1046.435 16057.505 1047.435 ;
    END
  END FREEZE_HV[18]
  PIN BcidMtx[1117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16055.545 1046.435 16055.825 1047.435 ;
    END
  END BcidMtx[1117]
  PIN Data_HV[381]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16014.105 1046.435 16014.385 1047.435 ;
    END
  END Data_HV[381]
  PIN Data_HV[393]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16012.425 1046.435 16012.705 1047.435 ;
    END
  END Data_HV[393]
  PIN Data_HV[394]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16010.745 1046.435 16011.025 1047.435 ;
    END
  END Data_HV[394]
  PIN Data_HV[378]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16009.065 1046.435 16009.345 1047.435 ;
    END
  END Data_HV[378]
  PIN MASKH[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16007.385 1046.435 16007.665 1047.435 ;
    END
  END MASKH[186]
  PIN MASKD[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16002.345 1046.435 16002.625 1047.435 ;
    END
  END MASKD[371]
  PIN MASKV[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15991.145 1046.435 15991.425 1047.435 ;
    END
  END MASKV[371]
  PIN Data_HV[376]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15988.905 1046.435 15989.185 1047.435 ;
    END
  END Data_HV[376]
  PIN Data_HV[371]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15986.665 1046.435 15986.945 1047.435 ;
    END
  END Data_HV[371]
  PIN INJ_IN[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15982.465 1046.435 15982.745 1047.435 ;
    END
  END INJ_IN[371]
  PIN BcidMtx[1115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15980.225 1046.435 15980.505 1047.435 ;
    END
  END BcidMtx[1115]
  PIN BcidMtx[1113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15979.105 1046.435 15979.385 1047.435 ;
    END
  END BcidMtx[1113]
  PIN BcidMtx[1111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15951.385 1046.435 15951.665 1047.435 ;
    END
  END BcidMtx[1111]
  PIN Data_HV[360]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15948.585 1046.435 15948.865 1047.435 ;
    END
  END Data_HV[360]
  PIN Data_HV[372]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15946.905 1046.435 15947.185 1047.435 ;
    END
  END Data_HV[372]
  PIN Data_HV[368]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15944.665 1046.435 15944.945 1047.435 ;
    END
  END Data_HV[368]
  PIN Data_HV[374]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15942.985 1046.435 15943.265 1047.435 ;
    END
  END Data_HV[374]
  PIN MASKH[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15941.865 1046.435 15942.145 1047.435 ;
    END
  END MASKH[185]
  PIN MASKD[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15923.945 1046.435 15924.225 1047.435 ;
    END
  END MASKD[369]
  PIN MASKV[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15921.145 1046.435 15921.425 1047.435 ;
    END
  END MASKV[369]
  PIN Data_HV[344]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15920.025 1046.435 15920.305 1047.435 ;
    END
  END Data_HV[344]
  PIN Data_HV[349]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15917.785 1046.435 15918.065 1047.435 ;
    END
  END Data_HV[349]
  PIN Data_HV[343]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15916.105 1046.435 15916.385 1047.435 ;
    END
  END Data_HV[343]
  PIN Data_HV[1076]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18718.345 1046.435 18718.625 1047.435 ;
    END
  END Data_HV[1076]
  PIN BcidMtx[1108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15872.425 1046.435 15872.705 1047.435 ;
    END
  END BcidMtx[1108]
  PIN Read_HV[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15870.745 1046.435 15871.025 1047.435 ;
    END
  END Read_HV[16]
  PIN BcidMtx[1106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15870.185 1046.435 15870.465 1047.435 ;
    END
  END BcidMtx[1106]
  PIN Data_HV[339]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15866.825 1046.435 15867.105 1047.435 ;
    END
  END Data_HV[339]
  PIN Data_HV[351]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15865.145 1046.435 15865.425 1047.435 ;
    END
  END Data_HV[351]
  PIN Data_HV[340]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15864.025 1046.435 15864.305 1047.435 ;
    END
  END Data_HV[340]
  PIN Data_HV[336]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15861.785 1046.435 15862.065 1047.435 ;
    END
  END Data_HV[336]
  PIN MASKV[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15852.265 1046.435 15852.545 1047.435 ;
    END
  END MASKV[368]
  PIN DIG_MON_HV[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15850.025 1046.435 15850.305 1047.435 ;
    END
  END DIG_MON_HV[32]
  PIN MASKD[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15846.665 1046.435 15846.945 1047.435 ;
    END
  END MASKD[367]
  PIN MASKV[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15841.905 1046.435 15842.185 1047.435 ;
    END
  END MASKV[367]
  PIN Data_HV[323]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15840.785 1046.435 15841.065 1047.435 ;
    END
  END Data_HV[323]
  PIN Data_HV[328]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15813.065 1046.435 15813.345 1047.435 ;
    END
  END Data_HV[328]
  PIN Data_HV[322]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15811.385 1046.435 15811.665 1047.435 ;
    END
  END Data_HV[322]
  PIN INJ_IN[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15809.705 1046.435 15809.985 1047.435 ;
    END
  END INJ_IN[367]
  PIN Data_HV[1085]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18716.665 1046.435 18716.945 1047.435 ;
    END
  END Data_HV[1085]
  PIN Read_HV[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15805.225 1046.435 15805.505 1047.435 ;
    END
  END Read_HV[15]
  PIN BcidMtx[1099]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15804.105 1046.435 15804.385 1047.435 ;
    END
  END BcidMtx[1099]
  PIN Data_HV[317]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15800.745 1046.435 15801.025 1047.435 ;
    END
  END Data_HV[317]
  PIN Data_HV[325]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15786.185 1046.435 15786.465 1047.435 ;
    END
  END Data_HV[325]
  PIN Data_HV[331]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15785.065 1046.435 15785.345 1047.435 ;
    END
  END Data_HV[331]
  PIN Data_HV[332]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15782.825 1046.435 15783.105 1047.435 ;
    END
  END Data_HV[332]
  PIN MASKD[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15781.145 1046.435 15781.425 1047.435 ;
    END
  END MASKD[366]
  PIN DIG_MON_HV[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15775.545 1046.435 15775.825 1047.435 ;
    END
  END DIG_MON_HV[29]
  PIN Data_HV[312]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15733.545 1046.435 15733.825 1047.435 ;
    END
  END Data_HV[312]
  PIN Data_HV[306]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15732.425 1046.435 15732.705 1047.435 ;
    END
  END Data_HV[306]
  PIN Data_HV[314]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15730.185 1046.435 15730.465 1047.435 ;
    END
  END Data_HV[314]
  PIN Data_HV[300]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15728.505 1046.435 15728.785 1047.435 ;
    END
  END Data_HV[300]
  PIN nTOK_HV[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15726.265 1046.435 15726.545 1047.435 ;
    END
  END nTOK_HV[14]
  PIN FREEZE_HV[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15723.465 1046.435 15723.745 1047.435 ;
    END
  END FREEZE_HV[14]
  PIN BcidMtx[1309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18604.105 1046.435 18604.385 1047.435 ;
    END
  END BcidMtx[1309]
  PIN BcidMtx[1092]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15721.225 1046.435 15721.505 1047.435 ;
    END
  END BcidMtx[1092]
  PIN Data_HV[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14587.225 1046.435 14587.505 1047.435 ;
    END
  END Data_HV[16]
  PIN Data_HV[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14584.985 1046.435 14585.265 1047.435 ;
    END
  END Data_HV[17]
  PIN MASKH[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14581.905 1046.435 14582.185 1047.435 ;
    END
  END MASKH[168]
  PIN DIG_MON_HV[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14580.225 1046.435 14580.505 1047.435 ;
    END
  END DIG_MON_HV[0]
  PIN FREEZE_HV[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14833.065 1046.435 14833.345 1047.435 ;
    END
  END FREEZE_HV[3]
  PIN DIG_MON_HV[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15669.705 1046.435 15669.985 1047.435 ;
    END
  END DIG_MON_HV[27]
  PIN Data_HV[291]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15667.465 1046.435 15667.745 1047.435 ;
    END
  END Data_HV[291]
  PIN Data_HV[292]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15665.785 1046.435 15666.065 1047.435 ;
    END
  END Data_HV[292]
  PIN Data_HV[286]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15664.665 1046.435 15664.945 1047.435 ;
    END
  END Data_HV[286]
  PIN Data_HV[287]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15663.545 1046.435 15663.825 1047.435 ;
    END
  END Data_HV[287]
  PIN BcidMtx[1091]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15645.625 1046.435 15645.905 1047.435 ;
    END
  END BcidMtx[1091]
  PIN BcidMtx[1089]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15644.505 1046.435 15644.785 1047.435 ;
    END
  END BcidMtx[1089]
  PIN BcidMtx[1087]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15642.265 1046.435 15642.545 1047.435 ;
    END
  END BcidMtx[1087]
  PIN Data_HV[276]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15639.465 1046.435 15639.745 1047.435 ;
    END
  END Data_HV[276]
  PIN Data_HV[282]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15638.345 1046.435 15638.625 1047.435 ;
    END
  END Data_HV[282]
  PIN Data_HV[277]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15636.665 1046.435 15636.945 1047.435 ;
    END
  END Data_HV[277]
  PIN Data_HV[273]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15634.425 1046.435 15634.705 1047.435 ;
    END
  END Data_HV[273]
  PIN MASKV[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15594.665 1046.435 15594.945 1047.435 ;
    END
  END MASKV[362]
  PIN DIG_MON_HV[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15592.425 1046.435 15592.705 1047.435 ;
    END
  END DIG_MON_HV[26]
  PIN MASKD[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15589.065 1046.435 15589.345 1047.435 ;
    END
  END MASKD[361]
  PIN INJ_ROW[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15586.825 1046.435 15587.105 1047.435 ;
    END
  END INJ_ROW[180]
  PIN Data_HV[264]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15584.585 1046.435 15584.865 1047.435 ;
    END
  END Data_HV[264]
  PIN Data_HV[265]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15582.905 1046.435 15583.185 1047.435 ;
    END
  END Data_HV[265]
  PIN Data_HV[266]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15581.785 1046.435 15582.065 1047.435 ;
    END
  END Data_HV[266]
  PIN nTOK_HV[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15570.025 1046.435 15570.305 1047.435 ;
    END
  END nTOK_HV[12]
  PIN BcidMtx[1083]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15567.785 1046.435 15568.065 1047.435 ;
    END
  END BcidMtx[1083]
  PIN BcidMtx[1082]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15566.105 1046.435 15566.385 1047.435 ;
    END
  END BcidMtx[1082]
  PIN BcidMtx[1080]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15564.985 1046.435 15565.265 1047.435 ;
    END
  END BcidMtx[1080]
  PIN Data_HV[261]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15559.665 1046.435 15559.945 1047.435 ;
    END
  END Data_HV[261]
  PIN Data_HV[256]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15532.505 1046.435 15532.785 1047.435 ;
    END
  END Data_HV[256]
  PIN Data_HV[253]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15530.825 1046.435 15531.105 1047.435 ;
    END
  END Data_HV[253]
  PIN MASKV[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15529.145 1046.435 15529.425 1047.435 ;
    END
  END MASKV[360]
  PIN DIG_MON_HV[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15526.905 1046.435 15527.185 1047.435 ;
    END
  END DIG_MON_HV[24]
  PIN DIG_MON_SEL[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15524.665 1046.435 15524.945 1047.435 ;
    END
  END DIG_MON_SEL[359]
  PIN INJ_ROW[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15521.305 1046.435 15521.585 1047.435 ;
    END
  END INJ_ROW[179]
  PIN Data_HV[239]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15519.625 1046.435 15519.905 1047.435 ;
    END
  END Data_HV[239]
  PIN Data_HV[236]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15505.065 1046.435 15505.345 1047.435 ;
    END
  END Data_HV[236]
  PIN Data_HV[245]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15503.385 1046.435 15503.665 1047.435 ;
    END
  END Data_HV[245]
  PIN INJ_IN[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15501.145 1046.435 15501.425 1047.435 ;
    END
  END INJ_IN[359]
  PIN nTOK_HV[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15500.025 1046.435 15500.305 1047.435 ;
    END
  END nTOK_HV[11]
  PIN Read_HV[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15496.665 1046.435 15496.945 1047.435 ;
    END
  END Read_HV[11]
  PIN BcidMtx[1311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18606.345 1046.435 18606.625 1047.435 ;
    END
  END BcidMtx[1311]
  PIN BcidMtx[1074]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15494.985 1046.435 15495.265 1047.435 ;
    END
  END BcidMtx[1074]
  PIN Data_HV[240]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15452.985 1046.435 15453.265 1047.435 ;
    END
  END Data_HV[240]
  PIN Data_HV[235]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15451.305 1046.435 15451.585 1047.435 ;
    END
  END Data_HV[235]
  PIN Data_HV[232]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15449.625 1046.435 15449.905 1047.435 ;
    END
  END Data_HV[232]
  PIN MASKV[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15447.945 1046.435 15448.225 1047.435 ;
    END
  END MASKV[358]
  PIN DIG_MON_HV[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15445.705 1046.435 15445.985 1047.435 ;
    END
  END DIG_MON_HV[22]
  PIN DIG_MON_SEL[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15443.465 1046.435 15443.745 1047.435 ;
    END
  END DIG_MON_SEL[357]
  PIN INJ_ROW[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15431.705 1046.435 15431.985 1047.435 ;
    END
  END INJ_ROW[178]
  PIN Data_HV[218]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15430.025 1046.435 15430.305 1047.435 ;
    END
  END Data_HV[218]
  PIN Data_HV[215]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15428.345 1046.435 15428.625 1047.435 ;
    END
  END Data_HV[215]
  PIN Data_HV[224]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15426.665 1046.435 15426.945 1047.435 ;
    END
  END Data_HV[224]
  PIN INJ_IN[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15422.465 1046.435 15422.745 1047.435 ;
    END
  END INJ_IN[357]
  PIN BcidMtx[1072]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15419.665 1046.435 15419.945 1047.435 ;
    END
  END BcidMtx[1072]
  PIN BcidMtx[1070]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15391.945 1046.435 15392.225 1047.435 ;
    END
  END BcidMtx[1070]
  PIN BcidMtx[1068]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15390.825 1046.435 15391.105 1047.435 ;
    END
  END BcidMtx[1068]
  PIN INJ_IN[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15389.705 1046.435 15389.985 1047.435 ;
    END
  END INJ_IN[356]
  PIN Data_HV[219]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15387.465 1046.435 15387.745 1047.435 ;
    END
  END Data_HV[219]
  PIN Data_HV[214]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15385.785 1046.435 15386.065 1047.435 ;
    END
  END Data_HV[214]
  PIN Data_HV[221]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15384.665 1046.435 15384.945 1047.435 ;
    END
  END Data_HV[221]
  PIN MASKV[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15382.425 1046.435 15382.705 1047.435 ;
    END
  END MASKV[356]
  PIN DIG_MON_HV[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15380.185 1046.435 15380.465 1047.435 ;
    END
  END DIG_MON_HV[20]
  PIN DIG_MON_SEL[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15365.625 1046.435 15365.905 1047.435 ;
    END
  END DIG_MON_SEL[356]
  PIN INJ_ROW[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15361.705 1046.435 15361.985 1047.435 ;
    END
  END INJ_ROW[177]
  PIN Data_HV[197]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15360.025 1046.435 15360.305 1047.435 ;
    END
  END Data_HV[197]
  PIN Data_HV[208]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15358.905 1046.435 15359.185 1047.435 ;
    END
  END Data_HV[208]
  PIN Data_HV[203]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15356.665 1046.435 15356.945 1047.435 ;
    END
  END Data_HV[203]
  PIN INJ_IN[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15354.425 1046.435 15354.705 1047.435 ;
    END
  END INJ_IN[355]
  PIN BcidMtx[1066]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15312.425 1046.435 15312.705 1047.435 ;
    END
  END BcidMtx[1066]
  PIN Read_HV[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15310.745 1046.435 15311.025 1047.435 ;
    END
  END Read_HV[9]
  PIN BcidMtx[1063]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15309.625 1046.435 15309.905 1047.435 ;
    END
  END BcidMtx[1063]
  PIN Data_HV[192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15306.825 1046.435 15307.105 1047.435 ;
    END
  END Data_HV[192]
  PIN Data_HV[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15306.265 1046.435 15306.545 1047.435 ;
    END
  END Data_HV[191]
  PIN Data_HV[199]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15304.585 1046.435 15304.865 1047.435 ;
    END
  END Data_HV[199]
  PIN Data_HV[205]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15303.465 1046.435 15303.745 1047.435 ;
    END
  END Data_HV[205]
  PIN Data_HV[206]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15301.225 1046.435 15301.505 1047.435 ;
    END
  END Data_HV[206]
  PIN MASKD[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15291.145 1046.435 15291.425 1047.435 ;
    END
  END MASKD[354]
  PIN DIG_MON_SEL[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15288.345 1046.435 15288.625 1047.435 ;
    END
  END DIG_MON_SEL[354]
  PIN DIG_MON_HV[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15285.545 1046.435 15285.825 1047.435 ;
    END
  END DIG_MON_HV[17]
  PIN Data_HV[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15281.345 1046.435 15281.625 1047.435 ;
    END
  END Data_HV[186]
  PIN Data_HV[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15279.665 1046.435 15279.945 1047.435 ;
    END
  END Data_HV[187]
  PIN Data_HV[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15252.505 1046.435 15252.785 1047.435 ;
    END
  END Data_HV[188]
  PIN Data_HV[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15250.825 1046.435 15251.105 1047.435 ;
    END
  END Data_HV[174]
  PIN nTOK_HV[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15248.585 1046.435 15248.865 1047.435 ;
    END
  END nTOK_HV[8]
  PIN FREEZE_HV[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15245.785 1046.435 15246.065 1047.435 ;
    END
  END FREEZE_HV[8]
  PIN BcidMtx[1057]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15244.105 1046.435 15244.385 1047.435 ;
    END
  END BcidMtx[1057]
  PIN INJ_IN[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15242.425 1046.435 15242.705 1047.435 ;
    END
  END INJ_IN[352]
  PIN Data_HV[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15226.745 1046.435 15227.025 1047.435 ;
    END
  END Data_HV[183]
  PIN Data_HV[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15225.065 1046.435 15225.345 1047.435 ;
    END
  END Data_HV[184]
  PIN Data_HV[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15223.385 1046.435 15223.665 1047.435 ;
    END
  END Data_HV[168]
  PIN MASKH[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15221.705 1046.435 15221.985 1047.435 ;
    END
  END MASKH[176]
  PIN MASKD[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15216.665 1046.435 15216.945 1047.435 ;
    END
  END MASKD[351]
  PIN MASKV[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15213.865 1046.435 15214.145 1047.435 ;
    END
  END MASKV[351]
  PIN Data_HV[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15172.425 1046.435 15172.705 1047.435 ;
    END
  END Data_HV[159]
  PIN Data_HV[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15171.305 1046.435 15171.585 1047.435 ;
    END
  END Data_HV[152]
  PIN Data_HV[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15169.065 1046.435 15169.345 1047.435 ;
    END
  END Data_HV[154]
  PIN nTOK_HV[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15166.265 1046.435 15166.545 1047.435 ;
    END
  END nTOK_HV[7]
  PIN BcidMtx[1054]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15164.585 1046.435 15164.865 1047.435 ;
    END
  END BcidMtx[1054]
  PIN BcidMtx[1052]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15162.345 1046.435 15162.625 1047.435 ;
    END
  END BcidMtx[1052]
  PIN INJ_IN[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15151.705 1046.435 15151.985 1047.435 ;
    END
  END INJ_IN[350]
  PIN Data_PMOS_NOSF[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1667.465 1046.435 1667.745 1047.435 ;
    END
  END Data_PMOS_NOSF[144]
  PIN Data_PMOS_NOSF[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1665.785 1046.435 1666.065 1047.435 ;
    END
  END Data_PMOS_NOSF[145]
  PIN Data_PMOS_NOSF[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1664.105 1046.435 1664.385 1047.435 ;
    END
  END Data_PMOS_NOSF[146]
  PIN Data_PMOS_NOSF[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1662.425 1046.435 1662.705 1047.435 ;
    END
  END Data_PMOS_NOSF[132]
  PIN BcidMtx[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1645.625 1046.435 1645.905 1047.435 ;
    END
  END BcidMtx[41]
  PIN FREEZE_PMOS_NOSF[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1643.945 1046.435 1644.225 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[6]
  PIN BcidMtx[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1642.265 1046.435 1642.545 1047.435 ;
    END
  END BcidMtx[37]
  PIN Data_PMOS_NOSF[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1639.465 1046.435 1639.745 1047.435 ;
    END
  END Data_PMOS_NOSF[129]
  PIN Data_PMOS_NOSF[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1637.785 1046.435 1638.065 1047.435 ;
    END
  END Data_PMOS_NOSF[141]
  PIN Data_PMOS_NOSF[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1636.105 1046.435 1636.385 1047.435 ;
    END
  END Data_PMOS_NOSF[142]
  PIN Data_PMOS_NOSF[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1634.425 1046.435 1634.705 1047.435 ;
    END
  END Data_PMOS_NOSF[126]
  PIN MASKH[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1594.105 1046.435 1594.385 1047.435 ;
    END
  END MASKH[6]
  PIN MASKV[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18889.145 1046.435 18889.425 1047.435 ;
    END
  END MASKV[444]
  PIN DIG_MON_SEL[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1590.185 1046.435 1590.465 1047.435 ;
    END
  END DIG_MON_SEL[11]
  PIN INJ_ROW[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1586.825 1046.435 1587.105 1047.435 ;
    END
  END INJ_ROW[5]
  PIN Data_PMOS_NOSF[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1585.145 1046.435 1585.425 1047.435 ;
    END
  END Data_PMOS_NOSF[113]
  PIN Data_PMOS_NOSF[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1583.465 1046.435 1583.745 1047.435 ;
    END
  END Data_PMOS_NOSF[110]
  PIN Data_PMOS_NOSF[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1581.785 1046.435 1582.065 1047.435 ;
    END
  END Data_PMOS_NOSF[119]
  PIN INJ_IN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1571.145 1046.435 1571.425 1047.435 ;
    END
  END INJ_IN[11]
  PIN BcidMtx[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1568.345 1046.435 1568.625 1047.435 ;
    END
  END BcidMtx[34]
  PIN Read_PMOS_NOSF[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1566.665 1046.435 1566.945 1047.435 ;
    END
  END Read_PMOS_NOSF[5]
  PIN BcidMtx[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1564.985 1046.435 1565.265 1047.435 ;
    END
  END BcidMtx[30]
  PIN Data_PMOS_NOSF[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1560.225 1046.435 1560.505 1047.435 ;
    END
  END Data_PMOS_NOSF[107]
  PIN Data_PMOS_NOSF[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1558.545 1046.435 1558.825 1047.435 ;
    END
  END Data_PMOS_NOSF[115]
  PIN Data_PMOS_NOSF[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1531.385 1046.435 1531.665 1047.435 ;
    END
  END Data_PMOS_NOSF[116]
  PIN Data_PMOS_NOSF[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1529.705 1046.435 1529.985 1047.435 ;
    END
  END Data_PMOS_NOSF[122]
  PIN MASKD[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1528.025 1046.435 1528.305 1047.435 ;
    END
  END MASKD[10]
  PIN MASKD[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1523.545 1046.435 1523.825 1047.435 ;
    END
  END MASKD[9]
  PIN MASKV[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1520.745 1046.435 1521.025 1047.435 ;
    END
  END MASKV[9]
  PIN Data_PMOS_NOSF[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1506.185 1046.435 1506.465 1047.435 ;
    END
  END Data_PMOS_NOSF[96]
  PIN Data_PMOS_NOSF[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1504.505 1046.435 1504.785 1047.435 ;
    END
  END Data_PMOS_NOSF[97]
  PIN Data_PMOS_NOSF[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1502.825 1046.435 1503.105 1047.435 ;
    END
  END Data_PMOS_NOSF[91]
  PIN nTOK_PMOS_NOSF[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1500.025 1046.435 1500.305 1047.435 ;
    END
  END nTOK_PMOS_NOSF[4]
  PIN BcidMtx[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1497.785 1046.435 1498.065 1047.435 ;
    END
  END BcidMtx[27]
  PIN BcidMtx[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1496.105 1046.435 1496.385 1047.435 ;
    END
  END BcidMtx[26]
  PIN INJ_IN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1493.865 1046.435 1494.145 1047.435 ;
    END
  END INJ_IN[8]
  PIN Data_PMOS_NOSF[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1452.985 1046.435 1453.265 1047.435 ;
    END
  END Data_PMOS_NOSF[93]
  PIN Data_PMOS_NOSF[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1451.305 1046.435 1451.585 1047.435 ;
    END
  END Data_PMOS_NOSF[88]
  PIN Data_PMOS_NOSF[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1449.625 1046.435 1449.905 1047.435 ;
    END
  END Data_PMOS_NOSF[85]
  PIN MASKV[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1447.945 1046.435 1448.225 1047.435 ;
    END
  END MASKV[8]
  PIN Data_HV[1134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18890.265 1046.435 18890.545 1047.435 ;
    END
  END Data_HV[1134]
  PIN DIG_MON_SEL[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1444.025 1046.435 1444.305 1047.435 ;
    END
  END DIG_MON_SEL[8]
  PIN DIG_MON_PMOS_NOSF[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1441.225 1046.435 1441.505 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[7]
  PIN Data_PMOS_NOSF[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1430.585 1046.435 1430.865 1047.435 ;
    END
  END Data_PMOS_NOSF[81]
  PIN Data_PMOS_NOSF[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1428.905 1046.435 1429.185 1047.435 ;
    END
  END Data_PMOS_NOSF[82]
  PIN Data_PMOS_NOSF[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1427.225 1046.435 1427.505 1047.435 ;
    END
  END Data_PMOS_NOSF[83]
  PIN Data_PMOS_NOSF[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1425.545 1046.435 1425.825 1047.435 ;
    END
  END Data_PMOS_NOSF[69]
  PIN nTOK_PMOS_NOSF[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1421.345 1046.435 1421.625 1047.435 ;
    END
  END nTOK_PMOS_NOSF[3]
  PIN BcidMtx[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1419.105 1046.435 1419.385 1047.435 ;
    END
  END BcidMtx[21]
  PIN BcidMtx[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1391.385 1046.435 1391.665 1047.435 ;
    END
  END BcidMtx[19]
  PIN Data_PMOS_NOSF[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1388.585 1046.435 1388.865 1047.435 ;
    END
  END Data_PMOS_NOSF[66]
  PIN Data_PMOS_NOSF[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1387.465 1046.435 1387.745 1047.435 ;
    END
  END Data_PMOS_NOSF[72]
  PIN Data_PMOS_NOSF[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1385.225 1046.435 1385.505 1047.435 ;
    END
  END Data_PMOS_NOSF[79]
  PIN Data_PMOS_NOSF[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1383.545 1046.435 1383.825 1047.435 ;
    END
  END Data_PMOS_NOSF[63]
  PIN MASKV[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1382.425 1046.435 1382.705 1047.435 ;
    END
  END MASKV[6]
  PIN DIG_MON_PMOS_NOSF[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1380.185 1046.435 1380.465 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[6]
  PIN DIG_MON_SEL[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1365.065 1046.435 1365.345 1047.435 ;
    END
  END DIG_MON_SEL[5]
  PIN DIG_MON_PMOS_NOSF[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1362.825 1046.435 1363.105 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[5]
  PIN Data_PMOS_NOSF[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1360.025 1046.435 1360.305 1047.435 ;
    END
  END Data_PMOS_NOSF[50]
  PIN Data_PMOS_NOSF[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1358.345 1046.435 1358.625 1047.435 ;
    END
  END Data_PMOS_NOSF[47]
  PIN Data_PMOS_NOSF[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1357.225 1046.435 1357.505 1047.435 ;
    END
  END Data_PMOS_NOSF[62]
  PIN INJ_IN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1354.425 1046.435 1354.705 1047.435 ;
    END
  END INJ_IN[5]
  PIN BcidMtx[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1312.425 1046.435 1312.705 1047.435 ;
    END
  END BcidMtx[16]
  PIN FREEZE_PMOS_NOSF[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1311.305 1046.435 1311.585 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[2]
  PIN BcidMtx[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1309.065 1046.435 1309.345 1047.435 ;
    END
  END BcidMtx[12]
  PIN Data_PMOS_NOSF[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1306.265 1046.435 1306.545 1047.435 ;
    END
  END Data_PMOS_NOSF[44]
  PIN Data_PMOS_NOSF[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1304.585 1046.435 1304.865 1047.435 ;
    END
  END Data_PMOS_NOSF[52]
  PIN Data_PMOS_NOSF[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1302.905 1046.435 1303.185 1047.435 ;
    END
  END Data_PMOS_NOSF[53]
  PIN Data_PMOS_NOSF[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1301.225 1046.435 1301.505 1047.435 ;
    END
  END Data_PMOS_NOSF[59]
  PIN MASKD[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1291.145 1046.435 1291.425 1047.435 ;
    END
  END MASKD[4]
  PIN MASKD[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1286.665 1046.435 1286.945 1047.435 ;
    END
  END MASKD[3]
  PIN MASKV[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1281.905 1046.435 1282.185 1047.435 ;
    END
  END MASKV[3]
  PIN Data_PMOS_NOSF[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1280.225 1046.435 1280.505 1047.435 ;
    END
  END Data_PMOS_NOSF[33]
  PIN Data_PMOS_NOSF[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1253.065 1046.435 1253.345 1047.435 ;
    END
  END Data_PMOS_NOSF[34]
  PIN Data_PMOS_NOSF[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1251.385 1046.435 1251.665 1047.435 ;
    END
  END Data_PMOS_NOSF[28]
  PIN BcidMtx[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1247.465 1046.435 1247.745 1047.435 ;
    END
  END BcidMtx[11]
  PIN FREEZE_PMOS_NOSF[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1245.785 1046.435 1246.065 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[1]
  PIN BcidMtx[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1244.665 1046.435 1244.945 1047.435 ;
    END
  END BcidMtx[8]
  PIN Data_PMOS_NOSF[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1240.745 1046.435 1241.025 1047.435 ;
    END
  END Data_PMOS_NOSF[23]
  PIN Data_PMOS_NOSF[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1226.185 1046.435 1226.465 1047.435 ;
    END
  END Data_PMOS_NOSF[31]
  PIN Data_PMOS_NOSF[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1225.625 1046.435 1225.905 1047.435 ;
    END
  END Data_PMOS_NOSF[25]
  PIN Data_PMOS_NOSF[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1222.825 1046.435 1223.105 1047.435 ;
    END
  END Data_PMOS_NOSF[38]
  PIN Data_HV[1150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18891.945 1046.435 18892.225 1047.435 ;
    END
  END Data_HV[1150]
  PIN MASKD[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1221.145 1046.435 1221.425 1047.435 ;
    END
  END MASKD[2]
  PIN MASKD[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1216.665 1046.435 1216.945 1047.435 ;
    END
  END MASKD[1]
  PIN MASKV[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1213.865 1046.435 1214.145 1047.435 ;
    END
  END MASKV[1]
  PIN Data_PMOS_NOSF[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1173.545 1046.435 1173.825 1047.435 ;
    END
  END Data_PMOS_NOSF[18]
  PIN Data_PMOS_NOSF[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1170.745 1046.435 1171.025 1047.435 ;
    END
  END Data_PMOS_NOSF[13]
  PIN Data_PMOS_NOSF[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1169.065 1046.435 1169.345 1047.435 ;
    END
  END Data_PMOS_NOSF[7]
  PIN Data_PMOS_NOSF[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1168.505 1046.435 1168.785 1047.435 ;
    END
  END Data_PMOS_NOSF[6]
  PIN BcidMtx[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1164.025 1046.435 1164.305 1047.435 ;
    END
  END BcidMtx[3]
  PIN BcidMtx[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1162.345 1046.435 1162.625 1047.435 ;
    END
  END BcidMtx[2]
  PIN BcidMtx[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1161.785 1046.435 1162.065 1047.435 ;
    END
  END BcidMtx[1]
  PIN Data_PMOS_NOSF[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1149.465 1046.435 1149.745 1047.435 ;
    END
  END Data_PMOS_NOSF[9]
  PIN Data_PMOS_NOSF[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1147.785 1046.435 1148.065 1047.435 ;
    END
  END Data_PMOS_NOSF[4]
  PIN Data_PMOS_NOSF[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1147.225 1046.435 1147.505 1047.435 ;
    END
  END Data_PMOS_NOSF[16]
  PIN Data_HV[1138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18892.505 1046.435 18892.785 1047.435 ;
    END
  END Data_HV[1138]
  PIN MASKH[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1141.905 1046.435 1142.185 1047.435 ;
    END
  END MASKH[0]
  PIN DIG_MON_PMOS_NOSF[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1140.225 1046.435 1140.505 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[0]
  PIN MASKH[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18581.705 1046.435 18581.985 1047.435 ;
    END
  END MASKH[218]
  PIN Data_COMP[942]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13680.585 1046.435 13680.865 1047.435 ;
    END
  END Data_COMP[942]
  PIN Data_COMP[936]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13679.465 1046.435 13679.745 1047.435 ;
    END
  END Data_COMP[936]
  PIN Data_COMP[937]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13677.785 1046.435 13678.065 1047.435 ;
    END
  END Data_COMP[937]
  PIN Data_COMP[930]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13675.545 1046.435 13675.825 1047.435 ;
    END
  END Data_COMP[930]
  PIN nTOK_COMP[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13634.105 1046.435 13634.385 1047.435 ;
    END
  END nTOK_COMP[44]
  PIN BcidMtx[939]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13631.865 1046.435 13632.145 1047.435 ;
    END
  END BcidMtx[939]
  PIN BcidMtx[937]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13629.625 1046.435 13629.905 1047.435 ;
    END
  END BcidMtx[937]
  PIN INJ_IN[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13627.945 1046.435 13628.225 1047.435 ;
    END
  END INJ_IN[312]
  PIN Data_COMP[933]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13625.705 1046.435 13625.985 1047.435 ;
    END
  END Data_COMP[933]
  PIN Data_COMP[940]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13623.465 1046.435 13623.745 1047.435 ;
    END
  END Data_COMP[940]
  PIN Data_COMP[925]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13622.345 1046.435 13622.625 1047.435 ;
    END
  END Data_COMP[925]
  PIN MASKV[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13612.265 1046.435 13612.545 1047.435 ;
    END
  END MASKV[312]
  PIN Data_HV[1109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18742.985 1046.435 18743.265 1047.435 ;
    END
  END Data_HV[1109]
  PIN DIG_MON_SEL[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13608.345 1046.435 13608.625 1047.435 ;
    END
  END DIG_MON_SEL[312]
  PIN MASKH[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18741.865 1046.435 18742.145 1047.435 ;
    END
  END MASKH[220]
  PIN Data_COMP[921]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13601.345 1046.435 13601.625 1047.435 ;
    END
  END Data_COMP[921]
  PIN Data_COMP[915]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13600.225 1046.435 13600.505 1047.435 ;
    END
  END Data_COMP[915]
  PIN Data_COMP[916]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13573.065 1046.435 13573.345 1047.435 ;
    END
  END Data_COMP[916]
  PIN Data_COMP[909]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13570.825 1046.435 13571.105 1047.435 ;
    END
  END Data_COMP[909]
  PIN nTOK_COMP[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13568.585 1046.435 13568.865 1047.435 ;
    END
  END nTOK_COMP[43]
  PIN BcidMtx[933]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13566.345 1046.435 13566.625 1047.435 ;
    END
  END BcidMtx[933]
  PIN BcidMtx[931]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13564.105 1046.435 13564.385 1047.435 ;
    END
  END BcidMtx[931]
  PIN INJ_IN[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13562.425 1046.435 13562.705 1047.435 ;
    END
  END INJ_IN[310]
  PIN Data_COMP[912]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13560.185 1046.435 13560.465 1047.435 ;
    END
  END Data_COMP[912]
  PIN Data_COMP[919]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13545.065 1046.435 13545.345 1047.435 ;
    END
  END Data_COMP[919]
  PIN Data_COMP[904]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13543.945 1046.435 13544.225 1047.435 ;
    END
  END Data_COMP[904]
  PIN MASKV[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13542.265 1046.435 13542.545 1047.435 ;
    END
  END MASKV[310]
  PIN DIG_MON_SEL[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13537.785 1046.435 13538.065 1047.435 ;
    END
  END DIG_MON_SEL[309]
  PIN DIG_MON_COMP[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13535.545 1046.435 13535.825 1047.435 ;
    END
  END DIG_MON_COMP[85]
  PIN Data_COMP[890]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13492.985 1046.435 13493.265 1047.435 ;
    END
  END Data_COMP[890]
  PIN Data_COMP[901]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13491.865 1046.435 13492.145 1047.435 ;
    END
  END Data_COMP[901]
  PIN Data_COMP[902]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13490.185 1046.435 13490.465 1047.435 ;
    END
  END Data_COMP[902]
  PIN INJ_IN[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13487.385 1046.435 13487.665 1047.435 ;
    END
  END INJ_IN[309]
  PIN BcidMtx[929]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13485.145 1046.435 13485.425 1047.435 ;
    END
  END BcidMtx[929]
  PIN FREEZE_COMP[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13483.465 1046.435 13483.745 1047.435 ;
    END
  END FREEZE_COMP[42]
  PIN BcidMtx[925]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13481.785 1046.435 13482.065 1047.435 ;
    END
  END BcidMtx[925]
  PIN Data_COMP[891]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13469.465 1046.435 13469.745 1047.435 ;
    END
  END Data_COMP[891]
  PIN Data_COMP[892]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13468.345 1046.435 13468.625 1047.435 ;
    END
  END Data_COMP[892]
  PIN Data_COMP[883]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13466.105 1046.435 13466.385 1047.435 ;
    END
  END Data_COMP[883]
  PIN MASKV[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13462.465 1046.435 13462.745 1047.435 ;
    END
  END MASKV[308]
  PIN DIG_MON_COMP[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13460.225 1046.435 13460.505 1047.435 ;
    END
  END DIG_MON_COMP[84]
  PIN FREEZE_COMP[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13713.065 1046.435 13713.345 1047.435 ;
    END
  END FREEZE_COMP[45]
  PIN BcidMtx[1313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18607.465 1046.435 18607.745 1047.435 ;
    END
  END BcidMtx[1313]
  PIN MASKV[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14548.025 1046.435 14548.305 1047.435 ;
    END
  END MASKV[335]
  PIN Data_COMP[1167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14546.345 1046.435 14546.625 1047.435 ;
    END
  END Data_COMP[1167]
  PIN Data_COMP[1168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14544.665 1046.435 14544.945 1047.435 ;
    END
  END Data_COMP[1168]
  PIN Data_COMP[1169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14543.545 1046.435 14543.825 1047.435 ;
    END
  END Data_COMP[1169]
  PIN INJ_IN[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14541.305 1046.435 14541.585 1047.435 ;
    END
  END INJ_IN[335]
  PIN BcidMtx[1006]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14525.065 1046.435 14525.345 1047.435 ;
    END
  END BcidMtx[1006]
  PIN Read_COMP[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14523.385 1046.435 14523.665 1047.435 ;
    END
  END Read_COMP[55]
  PIN BcidMtx[1002]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14521.705 1046.435 14521.985 1047.435 ;
    END
  END BcidMtx[1002]
  PIN Data_COMP[1157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14518.905 1046.435 14519.185 1047.435 ;
    END
  END Data_COMP[1157]
  PIN Data_COMP[1165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14517.225 1046.435 14517.505 1047.435 ;
    END
  END Data_COMP[1165]
  PIN Data_COMP[1166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14515.545 1046.435 14515.825 1047.435 ;
    END
  END Data_COMP[1166]
  PIN Data_COMP[1172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14513.865 1046.435 14514.145 1047.435 ;
    END
  END Data_COMP[1172]
  PIN MASKD[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14473.545 1046.435 14473.825 1047.435 ;
    END
  END MASKD[334]
  PIN DIG_MON_SEL[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14470.745 1046.435 14471.025 1047.435 ;
    END
  END DIG_MON_SEL[334]
  PIN DIG_MON_COMP[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14467.945 1046.435 14468.225 1047.435 ;
    END
  END DIG_MON_COMP[109]
  PIN Data_COMP[1152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14465.705 1046.435 14465.985 1047.435 ;
    END
  END Data_COMP[1152]
  PIN Data_COMP[1153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14464.025 1046.435 14464.305 1047.435 ;
    END
  END Data_COMP[1153]
  PIN Data_COMP[1154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14462.345 1046.435 14462.625 1047.435 ;
    END
  END Data_COMP[1154]
  PIN Data_COMP[1140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14452.265 1046.435 14452.545 1047.435 ;
    END
  END Data_COMP[1140]
  PIN nTOK_COMP[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14450.025 1046.435 14450.305 1047.435 ;
    END
  END nTOK_COMP[54]
  PIN BcidMtx[999]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14447.785 1046.435 14448.065 1047.435 ;
    END
  END BcidMtx[999]
  PIN BcidMtx[997]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14445.545 1046.435 14445.825 1047.435 ;
    END
  END BcidMtx[997]
  PIN INJ_IN[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14441.905 1046.435 14442.185 1047.435 ;
    END
  END INJ_IN[332]
  PIN Data_COMP[1143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14439.665 1046.435 14439.945 1047.435 ;
    END
  END Data_COMP[1143]
  PIN Data_COMP[1150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14411.945 1046.435 14412.225 1047.435 ;
    END
  END Data_COMP[1150]
  PIN Data_COMP[1135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14410.825 1046.435 14411.105 1047.435 ;
    END
  END Data_COMP[1135]
  PIN MASKV[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14409.145 1046.435 14409.425 1047.435 ;
    END
  END MASKV[332]
  PIN DIG_MON_SEL[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14404.665 1046.435 14404.945 1047.435 ;
    END
  END DIG_MON_SEL[331]
  PIN INJ_ROW[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14401.305 1046.435 14401.585 1047.435 ;
    END
  END INJ_ROW[165]
  PIN Data_COMP[1125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14386.185 1046.435 14386.465 1047.435 ;
    END
  END Data_COMP[1125]
  PIN Data_COMP[1118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14385.065 1046.435 14385.345 1047.435 ;
    END
  END Data_COMP[1118]
  PIN Data_COMP[1127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14383.385 1046.435 14383.665 1047.435 ;
    END
  END Data_COMP[1127]
  PIN nTOK_COMP[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14380.025 1046.435 14380.305 1047.435 ;
    END
  END nTOK_COMP[53]
  PIN BcidMtx[994]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14378.345 1046.435 14378.625 1047.435 ;
    END
  END BcidMtx[994]
  PIN Read_COMP[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14376.665 1046.435 14376.945 1047.435 ;
    END
  END Read_COMP[53]
  PIN INJ_IN[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14373.865 1046.435 14374.145 1047.435 ;
    END
  END INJ_IN[330]
  PIN Data_COMP[1115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14333.545 1046.435 14333.825 1047.435 ;
    END
  END Data_COMP[1115]
  PIN Data_COMP[1123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14331.865 1046.435 14332.145 1047.435 ;
    END
  END Data_COMP[1123]
  PIN Data_COMP[1114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14329.625 1046.435 14329.905 1047.435 ;
    END
  END Data_COMP[1114]
  PIN Data_COMP[1130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14328.505 1046.435 14328.785 1047.435 ;
    END
  END Data_COMP[1130]
  PIN MASKD[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14326.825 1046.435 14327.105 1047.435 ;
    END
  END MASKD[330]
  PIN DIG_MON_SEL[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14323.465 1046.435 14323.745 1047.435 ;
    END
  END DIG_MON_SEL[329]
  PIN DIG_MON_COMP[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14321.225 1046.435 14321.505 1047.435 ;
    END
  END DIG_MON_COMP[105]
  PIN Data_COMP[1110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14310.585 1046.435 14310.865 1047.435 ;
    END
  END Data_COMP[1110]
  PIN Data_COMP[1097]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14308.345 1046.435 14308.625 1047.435 ;
    END
  END Data_COMP[1097]
  PIN Data_COMP[1112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14307.225 1046.435 14307.505 1047.435 ;
    END
  END Data_COMP[1112]
  PIN Data_COMP[1098]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14305.545 1046.435 14305.825 1047.435 ;
    END
  END Data_COMP[1098]
  PIN BcidMtx[988]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14299.665 1046.435 14299.945 1047.435 ;
    END
  END BcidMtx[988]
  PIN Read_COMP[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14272.505 1046.435 14272.785 1047.435 ;
    END
  END Read_COMP[52]
  PIN BcidMtx[984]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14270.825 1046.435 14271.105 1047.435 ;
    END
  END BcidMtx[984]
  PIN Data_COMP[1101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14267.465 1046.435 14267.745 1047.435 ;
    END
  END Data_COMP[1101]
  PIN Data_COMP[1102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14266.345 1046.435 14266.625 1047.435 ;
    END
  END Data_COMP[1102]
  PIN Data_COMP[1103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14264.665 1046.435 14264.945 1047.435 ;
    END
  END Data_COMP[1103]
  PIN MASKV[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14262.425 1046.435 14262.705 1047.435 ;
    END
  END MASKV[328]
  PIN BcidMtx[1312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18606.905 1046.435 18607.185 1047.435 ;
    END
  END BcidMtx[1312]
  PIN DIG_MON_COMP[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14242.825 1046.435 14243.105 1047.435 ;
    END
  END DIG_MON_COMP[103]
  PIN DIG_MON_HV[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14802.825 1046.435 14803.105 1047.435 ;
    END
  END DIG_MON_HV[5]
  PIN Data_HV[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14800.585 1046.435 14800.865 1047.435 ;
    END
  END Data_HV[60]
  PIN Data_HV[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14798.905 1046.435 14799.185 1047.435 ;
    END
  END Data_HV[61]
  PIN Data_HV[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14797.225 1046.435 14797.505 1047.435 ;
    END
  END Data_HV[62]
  PIN Data_HV[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14795.545 1046.435 14795.825 1047.435 ;
    END
  END Data_HV[48]
  PIN BcidMtx[1025]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14752.985 1046.435 14753.265 1047.435 ;
    END
  END BcidMtx[1025]
  PIN FREEZE_HV[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14751.305 1046.435 14751.585 1047.435 ;
    END
  END FREEZE_HV[2]
  PIN BcidMtx[1021]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14749.625 1046.435 14749.905 1047.435 ;
    END
  END BcidMtx[1021]
  PIN Data_HV[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14746.825 1046.435 14747.105 1047.435 ;
    END
  END Data_HV[45]
  PIN Data_HV[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14745.705 1046.435 14745.985 1047.435 ;
    END
  END Data_HV[51]
  PIN Data_HV[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14744.025 1046.435 14744.305 1047.435 ;
    END
  END Data_HV[46]
  PIN Data_HV[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14741.785 1046.435 14742.065 1047.435 ;
    END
  END Data_HV[42]
  PIN MASKH[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14731.705 1046.435 14731.985 1047.435 ;
    END
  END MASKH[170]
  PIN DIG_MON_HV[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14730.025 1046.435 14730.305 1047.435 ;
    END
  END DIG_MON_HV[4]
  PIN INJ_ROW[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14722.465 1046.435 14722.745 1047.435 ;
    END
  END INJ_ROW[169]
  PIN Data_HV[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14720.785 1046.435 14721.065 1047.435 ;
    END
  END Data_HV[29]
  PIN Data_HV[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14720.225 1046.435 14720.505 1047.435 ;
    END
  END Data_HV[33]
  PIN Data_HV[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14691.945 1046.435 14692.225 1047.435 ;
    END
  END Data_HV[35]
  PIN INJ_IN[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14689.705 1046.435 14689.985 1047.435 ;
    END
  END INJ_IN[339]
  PIN BcidMtx[1019]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14687.465 1046.435 14687.745 1047.435 ;
    END
  END BcidMtx[1019]
  PIN BcidMtx[1016]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14684.665 1046.435 14684.945 1047.435 ;
    END
  END BcidMtx[1016]
  PIN BcidMtx[1014]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14683.545 1046.435 14683.825 1047.435 ;
    END
  END BcidMtx[1014]
  PIN Data_HV[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14680.185 1046.435 14680.465 1047.435 ;
    END
  END Data_HV[30]
  PIN DIG_MON_HV[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18722.825 1046.435 18723.105 1047.435 ;
    END
  END DIG_MON_HV[103]
  PIN Data_HV[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14664.505 1046.435 14664.785 1047.435 ;
    END
  END Data_HV[32]
  PIN Data_HV[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14662.825 1046.435 14663.105 1047.435 ;
    END
  END Data_HV[38]
  PIN MASKD[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14661.145 1046.435 14661.425 1047.435 ;
    END
  END MASKD[338]
  PIN DIG_MON_SEL[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14658.345 1046.435 14658.625 1047.435 ;
    END
  END DIG_MON_SEL[338]
  PIN MASKD[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14656.665 1046.435 14656.945 1047.435 ;
    END
  END MASKD[337]
  PIN Data_HV[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14613.545 1046.435 14613.825 1047.435 ;
    END
  END Data_HV[18]
  PIN Data_HV[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14611.865 1046.435 14612.145 1047.435 ;
    END
  END Data_HV[19]
  PIN Data_HV[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14609.625 1046.435 14609.905 1047.435 ;
    END
  END Data_HV[14]
  PIN Data_HV[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14608.505 1046.435 14608.785 1047.435 ;
    END
  END Data_HV[6]
  PIN BcidMtx[1013]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14605.145 1046.435 14605.425 1047.435 ;
    END
  END BcidMtx[1013]
  PIN Read_HV[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14602.905 1046.435 14603.185 1047.435 ;
    END
  END Read_HV[0]
  PIN BcidMtx[1008]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14601.225 1046.435 14601.505 1047.435 ;
    END
  END BcidMtx[1008]
  PIN Data_HV[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14590.585 1046.435 14590.865 1047.435 ;
    END
  END Data_HV[3]
  PIN Data_HV[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14589.465 1046.435 14589.745 1047.435 ;
    END
  END Data_HV[9]
  PIN Data_HV[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14586.665 1046.435 14586.945 1047.435 ;
    END
  END Data_HV[11]
  PIN FREEZE_HV[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18605.785 1046.435 18606.065 1047.435 ;
    END
  END FREEZE_HV[50]
  PIN MASKV[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14582.465 1046.435 14582.745 1047.435 ;
    END
  END MASKV[336]
  PIN DIG_MON_SEL[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15671.945 1046.435 15672.225 1047.435 ;
    END
  END DIG_MON_SEL[363]
  PIN INJ_ROW[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15668.585 1046.435 15668.865 1047.435 ;
    END
  END INJ_ROW[181]
  PIN Data_HV[281]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15666.905 1046.435 15667.185 1047.435 ;
    END
  END Data_HV[281]
  PIN Data_HV[278]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15665.225 1046.435 15665.505 1047.435 ;
    END
  END Data_HV[278]
  PIN Data_HV[280]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15662.985 1046.435 15663.265 1047.435 ;
    END
  END Data_HV[280]
  PIN INJ_IN[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15661.305 1046.435 15661.585 1047.435 ;
    END
  END INJ_IN[363]
  PIN BcidMtx[1090]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15645.065 1046.435 15645.345 1047.435 ;
    END
  END BcidMtx[1090]
  PIN FREEZE_HV[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15643.945 1046.435 15644.225 1047.435 ;
    END
  END FREEZE_HV[13]
  PIN BcidMtx[1086]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15641.705 1046.435 15641.985 1047.435 ;
    END
  END BcidMtx[1086]
  PIN Data_HV[275]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15638.905 1046.435 15639.185 1047.435 ;
    END
  END Data_HV[275]
  PIN Data_HV[288]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15637.785 1046.435 15638.065 1047.435 ;
    END
  END Data_HV[288]
  PIN Data_HV[284]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15635.545 1046.435 15635.825 1047.435 ;
    END
  END Data_HV[284]
  PIN Data_HV[290]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15633.865 1046.435 15634.145 1047.435 ;
    END
  END Data_HV[290]
  PIN MASKH[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15594.105 1046.435 15594.385 1047.435 ;
    END
  END MASKH[181]
  PIN DIG_MON_SEL[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15590.745 1046.435 15591.025 1047.435 ;
    END
  END DIG_MON_SEL[362]
  PIN DIG_MON_HV[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15587.945 1046.435 15588.225 1047.435 ;
    END
  END DIG_MON_HV[25]
  PIN MASKV[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15586.265 1046.435 15586.545 1047.435 ;
    END
  END MASKV[361]
  PIN Data_HV[271]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15584.025 1046.435 15584.305 1047.435 ;
    END
  END Data_HV[271]
  PIN Data_HV[272]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15582.345 1046.435 15582.625 1047.435 ;
    END
  END Data_HV[272]
  PIN Data_HV[259]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15581.225 1046.435 15581.505 1047.435 ;
    END
  END Data_HV[259]
  PIN BcidMtx[1085]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15568.905 1046.435 15569.185 1047.435 ;
    END
  END BcidMtx[1085]
  PIN FREEZE_HV[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15567.225 1046.435 15567.505 1047.435 ;
    END
  END FREEZE_HV[12]
  PIN INJ_IN[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15561.905 1046.435 15562.185 1047.435 ;
    END
  END INJ_IN[360]
  PIN Data_HV[255]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15560.785 1046.435 15561.065 1047.435 ;
    END
  END Data_HV[255]
  PIN Data_HV[267]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15559.105 1046.435 15559.385 1047.435 ;
    END
  END Data_HV[267]
  PIN Data_HV[268]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15531.945 1046.435 15532.225 1047.435 ;
    END
  END Data_HV[268]
  PIN Data_HV[252]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15530.265 1046.435 15530.545 1047.435 ;
    END
  END Data_HV[252]
  PIN MASKH[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15528.585 1046.435 15528.865 1047.435 ;
    END
  END MASKH[180]
  PIN MASKD[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15523.545 1046.435 15523.825 1047.435 ;
    END
  END MASKD[359]
  PIN MASKV[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15520.745 1046.435 15521.025 1047.435 ;
    END
  END MASKV[359]
  PIN Data_HV[243]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15506.185 1046.435 15506.465 1047.435 ;
    END
  END Data_HV[243]
  PIN Data_HV[244]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15504.505 1046.435 15504.785 1047.435 ;
    END
  END Data_HV[244]
  PIN Data_HV[238]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15502.825 1046.435 15503.105 1047.435 ;
    END
  END Data_HV[238]
  PIN BcidMtx[1079]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15498.905 1046.435 15499.185 1047.435 ;
    END
  END BcidMtx[1079]
  PIN BcidMtx[1077]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15497.785 1046.435 15498.065 1047.435 ;
    END
  END BcidMtx[1077]
  PIN BcidMtx[1076]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15496.105 1046.435 15496.385 1047.435 ;
    END
  END BcidMtx[1076]
  PIN BcidMtx[1075]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15495.545 1046.435 15495.825 1047.435 ;
    END
  END BcidMtx[1075]
  PIN Data_HV[234]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15454.105 1046.435 15454.385 1047.435 ;
    END
  END Data_HV[234]
  PIN Data_HV[246]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15452.425 1046.435 15452.705 1047.435 ;
    END
  END Data_HV[246]
  PIN Data_HV[247]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15450.745 1046.435 15451.025 1047.435 ;
    END
  END Data_HV[247]
  PIN Data_HV[231]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15449.065 1046.435 15449.345 1047.435 ;
    END
  END Data_HV[231]
  PIN MASKH[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15447.385 1046.435 15447.665 1047.435 ;
    END
  END MASKH[179]
  PIN MASKD[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15442.345 1046.435 15442.625 1047.435 ;
    END
  END MASKD[357]
  PIN MASKV[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15431.145 1046.435 15431.425 1047.435 ;
    END
  END MASKV[357]
  PIN Data_HV[222]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15429.465 1046.435 15429.745 1047.435 ;
    END
  END Data_HV[222]
  PIN Data_HV[223]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15427.785 1046.435 15428.065 1047.435 ;
    END
  END Data_HV[223]
  PIN Data_HV[217]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15426.105 1046.435 15426.385 1047.435 ;
    END
  END Data_HV[217]
  PIN nTOK_HV[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15421.345 1046.435 15421.625 1047.435 ;
    END
  END nTOK_HV[10]
  PIN BcidMtx[1071]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15419.105 1046.435 15419.385 1047.435 ;
    END
  END BcidMtx[1071]
  PIN INJ_ROW[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18721.705 1046.435 18721.985 1047.435 ;
    END
  END INJ_ROW[219]
  PIN Data_HV[1089]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18720.585 1046.435 18720.865 1047.435 ;
    END
  END Data_HV[1089]
  PIN Data_HV[213]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15388.585 1046.435 15388.865 1047.435 ;
    END
  END Data_HV[213]
  PIN Data_HV[225]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15386.905 1046.435 15387.185 1047.435 ;
    END
  END Data_HV[225]
  PIN Data_HV[226]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15385.225 1046.435 15385.505 1047.435 ;
    END
  END Data_HV[226]
  PIN Data_HV[210]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15383.545 1046.435 15383.825 1047.435 ;
    END
  END Data_HV[210]
  PIN MASKH[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15381.865 1046.435 15382.145 1047.435 ;
    END
  END MASKH[178]
  PIN Data_COMP[795]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13120.585 1046.435 13120.865 1047.435 ;
    END
  END Data_COMP[795]
  PIN Data_COMP[796]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13118.905 1046.435 13119.185 1047.435 ;
    END
  END Data_COMP[796]
  PIN Data_COMP[797]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13117.225 1046.435 13117.505 1047.435 ;
    END
  END Data_COMP[797]
  PIN INJ_IN[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13114.425 1046.435 13114.705 1047.435 ;
    END
  END INJ_IN[299]
  PIN BcidMtx[899]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13072.985 1046.435 13073.265 1047.435 ;
    END
  END BcidMtx[899]
  PIN FREEZE_COMP[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13071.305 1046.435 13071.585 1047.435 ;
    END
  END FREEZE_COMP[37]
  PIN BcidMtx[894]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13069.065 1046.435 13069.345 1047.435 ;
    END
  END BcidMtx[894]
  PIN Data_COMP[780]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13066.825 1046.435 13067.105 1047.435 ;
    END
  END Data_COMP[780]
  PIN Data_COMP[792]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13065.145 1046.435 13065.425 1047.435 ;
    END
  END Data_COMP[792]
  PIN Data_COMP[793]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13063.465 1046.435 13063.745 1047.435 ;
    END
  END Data_COMP[793]
  PIN Data_COMP[777]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13061.785 1046.435 13062.065 1047.435 ;
    END
  END Data_COMP[777]
  PIN MASKH[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13051.705 1046.435 13051.985 1047.435 ;
    END
  END MASKH[149]
  PIN DIG_MON_SEL[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13048.345 1046.435 13048.625 1047.435 ;
    END
  END DIG_MON_SEL[298]
  PIN DIG_MON_COMP[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13045.545 1046.435 13045.825 1047.435 ;
    END
  END DIG_MON_COMP[73]
  PIN INJ_ROW[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13042.465 1046.435 13042.745 1047.435 ;
    END
  END INJ_ROW[148]
  PIN Data_COMP[764]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13040.785 1046.435 13041.065 1047.435 ;
    END
  END Data_COMP[764]
  PIN Data_HV[1103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18744.665 1046.435 18744.945 1047.435 ;
    END
  END Data_HV[1103]
  PIN Data_COMP[769]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13013.065 1046.435 13013.345 1047.435 ;
    END
  END Data_COMP[769]
  PIN Data_COMP[762]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13010.825 1046.435 13011.105 1047.435 ;
    END
  END Data_COMP[762]
  PIN nTOK_COMP[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13008.585 1046.435 13008.865 1047.435 ;
    END
  END nTOK_COMP[36]
  PIN BcidMtx[891]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13006.345 1046.435 13006.625 1047.435 ;
    END
  END BcidMtx[891]
  PIN BcidMtx[889]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13004.105 1046.435 13004.385 1047.435 ;
    END
  END BcidMtx[889]
  PIN INJ_IN[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13002.425 1046.435 13002.705 1047.435 ;
    END
  END INJ_IN[296]
  PIN Data_COMP[765]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13000.185 1046.435 13000.465 1047.435 ;
    END
  END Data_COMP[765]
  PIN Data_COMP[772]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12985.065 1046.435 12985.345 1047.435 ;
    END
  END Data_COMP[772]
  PIN Data_COMP[757]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12983.945 1046.435 12984.225 1047.435 ;
    END
  END Data_COMP[757]
  PIN MASKV[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12982.265 1046.435 12982.545 1047.435 ;
    END
  END MASKV[296]
  PIN DIG_MON_SEL[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12977.785 1046.435 12978.065 1047.435 ;
    END
  END DIG_MON_SEL[295]
  PIN INJ_ROW[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12974.425 1046.435 12974.705 1047.435 ;
    END
  END INJ_ROW[147]
  PIN Data_COMP[747]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12932.425 1046.435 12932.705 1047.435 ;
    END
  END Data_COMP[747]
  PIN Data_COMP[740]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12931.305 1046.435 12931.585 1047.435 ;
    END
  END Data_COMP[740]
  PIN Data_COMP[749]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12929.625 1046.435 12929.905 1047.435 ;
    END
  END Data_COMP[749]
  PIN nTOK_COMP[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12926.265 1046.435 12926.545 1047.435 ;
    END
  END nTOK_COMP[35]
  PIN BcidMtx[886]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12924.585 1046.435 12924.865 1047.435 ;
    END
  END BcidMtx[886]
  PIN Read_COMP[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12922.905 1046.435 12923.185 1047.435 ;
    END
  END Read_COMP[35]
  PIN INJ_IN[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12911.705 1046.435 12911.985 1047.435 ;
    END
  END INJ_IN[294]
  PIN Data_COMP[737]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12910.025 1046.435 12910.305 1047.435 ;
    END
  END Data_COMP[737]
  PIN Data_COMP[745]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12908.345 1046.435 12908.625 1047.435 ;
    END
  END Data_COMP[745]
  PIN Data_COMP[736]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12906.105 1046.435 12906.385 1047.435 ;
    END
  END Data_COMP[736]
  PIN Data_COMP[752]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12904.985 1046.435 12905.265 1047.435 ;
    END
  END Data_COMP[752]
  PIN MASKD[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12901.345 1046.435 12901.625 1047.435 ;
    END
  END MASKD[294]
  PIN FREEZE_COMP[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13153.065 1046.435 13153.345 1047.435 ;
    END
  END FREEZE_COMP[38]
  PIN MASKD[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13990.825 1046.435 13991.105 1047.435 ;
    END
  END MASKD[321]
  PIN MASKV[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13988.025 1046.435 13988.305 1047.435 ;
    END
  END MASKV[321]
  PIN Data_COMP[1020]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13986.345 1046.435 13986.625 1047.435 ;
    END
  END Data_COMP[1020]
  PIN Data_COMP[1013]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13985.225 1046.435 13985.505 1047.435 ;
    END
  END Data_COMP[1013]
  PIN Data_COMP[1022]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13983.545 1046.435 13983.825 1047.435 ;
    END
  END Data_COMP[1022]
  PIN nTOK_COMP[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13980.185 1046.435 13980.465 1047.435 ;
    END
  END nTOK_COMP[48]
  PIN BcidMtx[964]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13965.065 1046.435 13965.345 1047.435 ;
    END
  END BcidMtx[964]
  PIN Read_COMP[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13963.385 1046.435 13963.665 1047.435 ;
    END
  END Read_COMP[48]
  PIN INJ_IN[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13960.585 1046.435 13960.865 1047.435 ;
    END
  END INJ_IN[320]
  PIN Data_COMP[1010]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13958.905 1046.435 13959.185 1047.435 ;
    END
  END Data_COMP[1010]
  PIN Data_COMP[1018]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13957.225 1046.435 13957.505 1047.435 ;
    END
  END Data_COMP[1018]
  PIN Data_COMP[1009]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13954.985 1046.435 13955.265 1047.435 ;
    END
  END Data_COMP[1009]
  PIN Data_COMP[1025]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13953.865 1046.435 13954.145 1047.435 ;
    END
  END Data_COMP[1025]
  PIN MASKD[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13913.545 1046.435 13913.825 1047.435 ;
    END
  END MASKD[320]
  PIN DIG_MON_SEL[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13910.185 1046.435 13910.465 1047.435 ;
    END
  END DIG_MON_SEL[319]
  PIN DIG_MON_COMP[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13907.945 1046.435 13908.225 1047.435 ;
    END
  END DIG_MON_COMP[95]
  PIN Data_COMP[1005]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13905.705 1046.435 13905.985 1047.435 ;
    END
  END Data_COMP[1005]
  PIN Data_COMP[992]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13903.465 1046.435 13903.745 1047.435 ;
    END
  END Data_COMP[992]
  PIN Data_COMP[1007]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13902.345 1046.435 13902.625 1047.435 ;
    END
  END Data_COMP[1007]
  PIN Data_COMP[993]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13892.265 1046.435 13892.545 1047.435 ;
    END
  END Data_COMP[993]
  PIN BcidMtx[958]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13888.345 1046.435 13888.625 1047.435 ;
    END
  END BcidMtx[958]
  PIN FREEZE_COMP[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13887.225 1046.435 13887.505 1047.435 ;
    END
  END FREEZE_COMP[47]
  PIN BcidMtx[955]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13885.545 1046.435 13885.825 1047.435 ;
    END
  END BcidMtx[955]
  PIN Data_COMP[989]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13880.225 1046.435 13880.505 1047.435 ;
    END
  END Data_COMP[989]
  PIN Data_COMP[1002]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13879.105 1046.435 13879.385 1047.435 ;
    END
  END Data_COMP[1002]
  PIN Data_COMP[1003]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13851.945 1046.435 13852.225 1047.435 ;
    END
  END Data_COMP[1003]
  PIN Data_COMP[1004]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13849.705 1046.435 13849.985 1047.435 ;
    END
  END Data_COMP[1004]
  PIN MASKH[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13848.585 1046.435 13848.865 1047.435 ;
    END
  END MASKH[159]
  PIN DIG_MON_COMP[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13842.425 1046.435 13842.705 1047.435 ;
    END
  END DIG_MON_COMP[93]
  PIN MASKV[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13840.745 1046.435 13841.025 1047.435 ;
    END
  END MASKV[317]
  PIN Data_COMP[978]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13826.185 1046.435 13826.465 1047.435 ;
    END
  END Data_COMP[978]
  PIN Data_COMP[986]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13823.945 1046.435 13824.225 1047.435 ;
    END
  END Data_COMP[986]
  PIN Data_COMP[973]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13822.825 1046.435 13823.105 1047.435 ;
    END
  END Data_COMP[973]
  PIN nTOK_COMP[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13820.025 1046.435 13820.305 1047.435 ;
    END
  END nTOK_COMP[46]
  PIN FREEZE_COMP[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13817.225 1046.435 13817.505 1047.435 ;
    END
  END FREEZE_COMP[46]
  PIN BcidMtx[950]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13816.105 1046.435 13816.385 1047.435 ;
    END
  END BcidMtx[950]
  PIN INJ_IN[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13813.865 1046.435 13814.145 1047.435 ;
    END
  END INJ_IN[316]
  PIN Data_COMP[981]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13772.425 1046.435 13772.705 1047.435 ;
    END
  END Data_COMP[981]
  PIN Data_COMP[970]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13771.305 1046.435 13771.585 1047.435 ;
    END
  END Data_COMP[970]
  PIN Data_COMP[967]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13769.625 1046.435 13769.905 1047.435 ;
    END
  END Data_COMP[967]
  PIN MASKH[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13767.385 1046.435 13767.665 1047.435 ;
    END
  END MASKH[158]
  PIN DIG_MON_COMP[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13765.705 1046.435 13765.985 1047.435 ;
    END
  END DIG_MON_COMP[92]
  PIN DIG_MON_SEL[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13763.465 1046.435 13763.745 1047.435 ;
    END
  END DIG_MON_SEL[315]
  PIN MASKV[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13751.145 1046.435 13751.425 1047.435 ;
    END
  END MASKV[315]
  PIN Data_COMP[953]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13750.025 1046.435 13750.305 1047.435 ;
    END
  END Data_COMP[953]
  PIN Data_COMP[950]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13748.345 1046.435 13748.625 1047.435 ;
    END
  END Data_COMP[950]
  PIN Data_COMP[952]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13746.105 1046.435 13746.385 1047.435 ;
    END
  END Data_COMP[952]
  PIN INJ_IN[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13742.465 1046.435 13742.745 1047.435 ;
    END
  END INJ_IN[315]
  PIN BcidMtx[946]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13739.665 1046.435 13739.945 1047.435 ;
    END
  END BcidMtx[946]
  PIN BcidMtx[943]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13711.385 1046.435 13711.665 1047.435 ;
    END
  END BcidMtx[943]
  PIN INJ_IN[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13709.705 1046.435 13709.985 1047.435 ;
    END
  END INJ_IN[314]
  PIN Data_COMP[954]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13707.465 1046.435 13707.745 1047.435 ;
    END
  END Data_COMP[954]
  PIN Data_COMP[961]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13705.225 1046.435 13705.505 1047.435 ;
    END
  END Data_COMP[961]
  PIN Data_COMP[946]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13704.105 1046.435 13704.385 1047.435 ;
    END
  END Data_COMP[946]
  PIN MASKV[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13702.425 1046.435 13702.705 1047.435 ;
    END
  END MASKV[314]
  PIN Data_HV[1092]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18743.545 1046.435 18743.825 1047.435 ;
    END
  END Data_HV[1092]
  PIN DIG_MON_SEL[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13685.625 1046.435 13685.905 1047.435 ;
    END
  END DIG_MON_SEL[314]
  PIN MASKD[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13683.945 1046.435 13684.225 1047.435 ;
    END
  END MASKD[313]
  PIN Data_COMP[635]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12558.345 1046.435 12558.625 1047.435 ;
    END
  END Data_COMP[635]
  PIN Data_COMP[644]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12556.665 1046.435 12556.945 1047.435 ;
    END
  END Data_COMP[644]
  PIN Data_COMP[636]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12555.545 1046.435 12555.825 1047.435 ;
    END
  END Data_COMP[636]
  PIN BcidMtx[857]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12512.985 1046.435 12513.265 1047.435 ;
    END
  END BcidMtx[857]
  PIN FREEZE_COMP[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12511.305 1046.435 12511.585 1047.435 ;
    END
  END FREEZE_COMP[30]
  PIN BcidMtx[853]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12509.625 1046.435 12509.905 1047.435 ;
    END
  END BcidMtx[853]
  PIN Data_COMP[632]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12506.265 1046.435 12506.545 1047.435 ;
    END
  END Data_COMP[632]
  PIN Data_COMP[645]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12505.145 1046.435 12505.425 1047.435 ;
    END
  END Data_COMP[645]
  PIN Data_COMP[646]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12503.465 1046.435 12503.745 1047.435 ;
    END
  END Data_COMP[646]
  PIN Data_COMP[647]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12501.225 1046.435 12501.505 1047.435 ;
    END
  END Data_COMP[647]
  PIN MASKH[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12491.705 1046.435 12491.985 1047.435 ;
    END
  END MASKH[142]
  PIN DIG_MON_COMP[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12485.545 1046.435 12485.825 1047.435 ;
    END
  END DIG_MON_COMP[59]
  PIN MASKV[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12481.905 1046.435 12482.185 1047.435 ;
    END
  END MASKV[283]
  PIN Data_COMP[621]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12480.225 1046.435 12480.505 1047.435 ;
    END
  END Data_COMP[621]
  PIN Data_COMP[614]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12479.105 1046.435 12479.385 1047.435 ;
    END
  END Data_COMP[614]
  PIN Data_COMP[623]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12451.945 1046.435 12452.225 1047.435 ;
    END
  END Data_COMP[623]
  PIN INJ_IN[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12449.705 1046.435 12449.985 1047.435 ;
    END
  END INJ_IN[283]
  PIN BcidMtx[850]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12446.905 1046.435 12447.185 1047.435 ;
    END
  END BcidMtx[850]
  PIN Read_COMP[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12445.225 1046.435 12445.505 1047.435 ;
    END
  END Read_COMP[29]
  PIN BcidMtx[846]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12443.545 1046.435 12443.825 1047.435 ;
    END
  END BcidMtx[846]
  PIN Data_COMP[618]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12440.185 1046.435 12440.465 1047.435 ;
    END
  END Data_COMP[618]
  PIN Data_COMP[619]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12426.185 1046.435 12426.465 1047.435 ;
    END
  END Data_COMP[619]
  PIN Data_COMP[620]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12424.505 1046.435 12424.785 1047.435 ;
    END
  END Data_COMP[620]
  PIN Data_COMP[626]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12422.825 1046.435 12423.105 1047.435 ;
    END
  END Data_COMP[626]
  PIN MASKD[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12421.145 1046.435 12421.425 1047.435 ;
    END
  END MASKD[282]
  PIN DIG_MON_SEL[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12418.345 1046.435 12418.625 1047.435 ;
    END
  END DIG_MON_SEL[282]
  PIN DIG_MON_COMP[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12415.545 1046.435 12415.825 1047.435 ;
    END
  END DIG_MON_COMP[57]
  PIN Data_COMP[606]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12373.545 1046.435 12373.825 1047.435 ;
    END
  END Data_COMP[606]
  PIN Data_COMP[607]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12371.865 1046.435 12372.145 1047.435 ;
    END
  END Data_COMP[607]
  PIN Data_HV[1101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18747.465 1046.435 18747.745 1047.435 ;
    END
  END Data_HV[1101]
  PIN Data_COMP[595]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12369.065 1046.435 12369.345 1047.435 ;
    END
  END Data_COMP[595]
  PIN nTOK_COMP[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12366.265 1046.435 12366.545 1047.435 ;
    END
  END nTOK_COMP[28]
  PIN FREEZE_COMP[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12363.465 1046.435 12363.745 1047.435 ;
    END
  END FREEZE_COMP[28]
  PIN BcidMtx[842]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12362.345 1046.435 12362.625 1047.435 ;
    END
  END BcidMtx[842]
  PIN INJ_IN[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12351.705 1046.435 12351.985 1047.435 ;
    END
  END INJ_IN[280]
  PIN Data_COMP[597]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12349.465 1046.435 12349.745 1047.435 ;
    END
  END Data_COMP[597]
  PIN Data_COMP[592]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12347.785 1046.435 12348.065 1047.435 ;
    END
  END Data_COMP[592]
  PIN Data_COMP[589]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12346.105 1046.435 12346.385 1047.435 ;
    END
  END Data_COMP[589]
  PIN MASKV[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12342.465 1046.435 12342.745 1047.435 ;
    END
  END MASKV[280]
  PIN DIG_MON_COMP[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12340.225 1046.435 12340.505 1047.435 ;
    END
  END DIG_MON_COMP[56]
  PIN FREEZE_COMP[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12593.065 1046.435 12593.345 1047.435 ;
    END
  END FREEZE_COMP[31]
  PIN INJ_ROW[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13428.585 1046.435 13428.865 1047.435 ;
    END
  END INJ_ROW[153]
  PIN Data_COMP[879]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13427.465 1046.435 13427.745 1047.435 ;
    END
  END Data_COMP[879]
  PIN Data_COMP[880]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13425.785 1046.435 13426.065 1047.435 ;
    END
  END Data_COMP[880]
  PIN Data_COMP[875]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13423.545 1046.435 13423.825 1047.435 ;
    END
  END Data_COMP[875]
  PIN Data_HV[1107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18746.905 1046.435 18747.185 1047.435 ;
    END
  END Data_HV[1107]
  PIN nTOK_COMP[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13420.185 1046.435 13420.465 1047.435 ;
    END
  END nTOK_COMP[41]
  PIN FREEZE_COMP[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13403.945 1046.435 13404.225 1047.435 ;
    END
  END FREEZE_COMP[41]
  PIN BcidMtx[920]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13402.825 1046.435 13403.105 1047.435 ;
    END
  END BcidMtx[920]
  PIN INJ_IN[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13400.585 1046.435 13400.865 1047.435 ;
    END
  END INJ_IN[306]
  PIN Data_COMP[876]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13397.785 1046.435 13398.065 1047.435 ;
    END
  END Data_COMP[876]
  PIN Data_COMP[865]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13396.665 1046.435 13396.945 1047.435 ;
    END
  END Data_COMP[865]
  PIN Data_COMP[862]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13394.985 1046.435 13395.265 1047.435 ;
    END
  END Data_COMP[862]
  PIN MASKH[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13354.105 1046.435 13354.385 1047.435 ;
    END
  END MASKH[153]
  PIN DIG_MON_COMP[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13352.425 1046.435 13352.705 1047.435 ;
    END
  END DIG_MON_COMP[82]
  PIN DIG_MON_SEL[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13350.185 1046.435 13350.465 1047.435 ;
    END
  END DIG_MON_SEL[305]
  PIN INJ_ROW[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13346.825 1046.435 13347.105 1047.435 ;
    END
  END INJ_ROW[152]
  PIN Data_COMP[848]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13345.145 1046.435 13345.425 1047.435 ;
    END
  END Data_COMP[848]
  PIN Data_COMP[845]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13343.465 1046.435 13343.745 1047.435 ;
    END
  END Data_COMP[845]
  PIN Data_COMP[854]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13341.785 1046.435 13342.065 1047.435 ;
    END
  END Data_COMP[854]
  PIN INJ_IN[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13331.145 1046.435 13331.425 1047.435 ;
    END
  END INJ_IN[305]
  PIN BcidMtx[916]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13328.345 1046.435 13328.625 1047.435 ;
    END
  END BcidMtx[916]
  PIN BcidMtx[914]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13326.105 1046.435 13326.385 1047.435 ;
    END
  END BcidMtx[914]
  PIN BcidMtx[912]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13324.985 1046.435 13325.265 1047.435 ;
    END
  END BcidMtx[912]
  PIN Data_COMP[842]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13320.225 1046.435 13320.505 1047.435 ;
    END
  END Data_COMP[842]
  PIN Data_COMP[844]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13292.505 1046.435 13292.785 1047.435 ;
    END
  END Data_COMP[844]
  PIN Data_COMP[851]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13291.385 1046.435 13291.665 1047.435 ;
    END
  END Data_COMP[851]
  PIN MASKH[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13288.585 1046.435 13288.865 1047.435 ;
    END
  END MASKH[152]
  PIN MASKD[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13288.025 1046.435 13288.305 1047.435 ;
    END
  END MASKD[304]
  PIN DIG_MON_SEL[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13285.225 1046.435 13285.505 1047.435 ;
    END
  END DIG_MON_SEL[304]
  PIN DIG_MON_COMP[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13282.425 1046.435 13282.705 1047.435 ;
    END
  END DIG_MON_COMP[79]
  PIN Data_COMP[827]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13279.625 1046.435 13279.905 1047.435 ;
    END
  END Data_COMP[827]
  PIN Data_COMP[838]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13265.625 1046.435 13265.905 1047.435 ;
    END
  END Data_COMP[838]
  PIN Data_COMP[839]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13263.945 1046.435 13264.225 1047.435 ;
    END
  END Data_COMP[839]
  PIN INJ_IN[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13261.145 1046.435 13261.425 1047.435 ;
    END
  END INJ_IN[303]
  PIN BcidMtx[911]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13258.905 1046.435 13259.185 1047.435 ;
    END
  END BcidMtx[911]
  PIN FREEZE_COMP[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13257.225 1046.435 13257.505 1047.435 ;
    END
  END FREEZE_COMP[39]
  PIN BcidMtx[907]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13255.545 1046.435 13255.825 1047.435 ;
    END
  END BcidMtx[907]
  PIN Data_COMP[822]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13214.105 1046.435 13214.385 1047.435 ;
    END
  END Data_COMP[822]
  PIN Data_COMP[834]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13212.425 1046.435 13212.705 1047.435 ;
    END
  END Data_COMP[834]
  PIN Data_COMP[830]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13210.185 1046.435 13210.465 1047.435 ;
    END
  END Data_COMP[830]
  PIN Data_COMP[819]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13209.065 1046.435 13209.345 1047.435 ;
    END
  END Data_COMP[819]
  PIN MASKH[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13207.385 1046.435 13207.665 1047.435 ;
    END
  END MASKH[151]
  PIN DIG_MON_SEL[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13204.025 1046.435 13204.305 1047.435 ;
    END
  END DIG_MON_SEL[302]
  PIN Data_HV[1072]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18662.345 1046.435 18662.625 1047.435 ;
    END
  END Data_HV[1072]
  PIN DIG_MON_COMP[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13201.225 1046.435 13201.505 1047.435 ;
    END
  END DIG_MON_COMP[77]
  PIN Data_COMP[806]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13190.025 1046.435 13190.305 1047.435 ;
    END
  END Data_COMP[806]
  PIN Data_COMP[817]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13188.905 1046.435 13189.185 1047.435 ;
    END
  END Data_COMP[817]
  PIN Data_COMP[818]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13187.225 1046.435 13187.505 1047.435 ;
    END
  END Data_COMP[818]
  PIN INJ_IN[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13182.465 1046.435 13182.745 1047.435 ;
    END
  END INJ_IN[301]
  PIN BcidMtx[905]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13180.225 1046.435 13180.505 1047.435 ;
    END
  END BcidMtx[905]
  PIN Read_COMP[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13152.505 1046.435 13152.785 1047.435 ;
    END
  END Read_COMP[38]
  PIN INJ_IN[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13149.705 1046.435 13149.985 1047.435 ;
    END
  END INJ_IN[300]
  PIN Data_COMP[800]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13148.025 1046.435 13148.305 1047.435 ;
    END
  END Data_COMP[800]
  PIN Data_COMP[808]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13146.345 1046.435 13146.625 1047.435 ;
    END
  END Data_COMP[808]
  PIN Data_COMP[799]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13144.105 1046.435 13144.385 1047.435 ;
    END
  END Data_COMP[799]
  PIN Data_COMP[815]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13142.985 1046.435 13143.265 1047.435 ;
    END
  END Data_COMP[815]
  PIN MASKD[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13141.305 1046.435 13141.585 1047.435 ;
    END
  END MASKD[300]
  PIN DIG_MON_SEL[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13125.065 1046.435 13125.345 1047.435 ;
    END
  END DIG_MON_SEL[299]
  PIN Data_HV[1102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18746.345 1046.435 18746.625 1047.435 ;
    END
  END Data_HV[1102]
  PIN MASKV[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13121.145 1046.435 13121.425 1047.435 ;
    END
  END MASKV[299]
  PIN MASKV[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14241.145 1046.435 14241.425 1047.435 ;
    END
  END MASKV[327]
  PIN Data_COMP[1083]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14239.465 1046.435 14239.745 1047.435 ;
    END
  END Data_COMP[1083]
  PIN Data_COMP[1091]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14237.225 1046.435 14237.505 1047.435 ;
    END
  END Data_COMP[1091]
  PIN Data_COMP[1078]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14236.105 1046.435 14236.385 1047.435 ;
    END
  END Data_COMP[1078]
  PIN nTOK_COMP[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14194.105 1046.435 14194.385 1047.435 ;
    END
  END nTOK_COMP[51]
  PIN FREEZE_COMP[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14191.305 1046.435 14191.585 1047.435 ;
    END
  END FREEZE_COMP[51]
  PIN BcidMtx[980]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14190.185 1046.435 14190.465 1047.435 ;
    END
  END BcidMtx[980]
  PIN INJ_IN[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14187.945 1046.435 14188.225 1047.435 ;
    END
  END INJ_IN[326]
  PIN Data_COMP[1086]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14185.145 1046.435 14185.425 1047.435 ;
    END
  END Data_COMP[1086]
  PIN Data_COMP[1075]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14184.025 1046.435 14184.305 1047.435 ;
    END
  END Data_COMP[1075]
  PIN Data_COMP[1072]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14182.345 1046.435 14182.625 1047.435 ;
    END
  END Data_COMP[1072]
  PIN MASKH[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14171.705 1046.435 14171.985 1047.435 ;
    END
  END MASKH[163]
  PIN DIG_MON_COMP[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14170.025 1046.435 14170.305 1047.435 ;
    END
  END DIG_MON_COMP[102]
  PIN DIG_MON_SEL[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14168.345 1046.435 14168.625 1047.435 ;
    END
  END DIG_MON_SEL[326]
  PIN INJ_ROW[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14162.465 1046.435 14162.745 1047.435 ;
    END
  END INJ_ROW[162]
  PIN Data_COMP[1068]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14161.345 1046.435 14161.625 1047.435 ;
    END
  END Data_COMP[1068]
  PIN Data_COMP[1069]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14159.665 1046.435 14159.945 1047.435 ;
    END
  END Data_COMP[1069]
  PIN Data_COMP[1064]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14131.945 1046.435 14132.225 1047.435 ;
    END
  END Data_COMP[1064]
  PIN Data_COMP[1056]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14130.825 1046.435 14131.105 1047.435 ;
    END
  END Data_COMP[1056]
  PIN BcidMtx[977]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14127.465 1046.435 14127.745 1047.435 ;
    END
  END BcidMtx[977]
  PIN Read_COMP[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14125.225 1046.435 14125.505 1047.435 ;
    END
  END Read_COMP[50]
  PIN BcidMtx[973]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14124.105 1046.435 14124.385 1047.435 ;
    END
  END BcidMtx[973]
  PIN Data_COMP[1053]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14121.305 1046.435 14121.585 1047.435 ;
    END
  END Data_COMP[1053]
  PIN Data_COMP[1060]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14106.185 1046.435 14106.465 1047.435 ;
    END
  END Data_COMP[1060]
  PIN Data_COMP[1066]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14105.065 1046.435 14105.345 1047.435 ;
    END
  END Data_COMP[1066]
  PIN Data_COMP[1050]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14103.385 1046.435 14103.665 1047.435 ;
    END
  END Data_COMP[1050]
  PIN DIG_MON_SEL[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18725.625 1046.435 18725.905 1047.435 ;
    END
  END DIG_MON_SEL[440]
  PIN DIG_MON_COMP[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14100.025 1046.435 14100.305 1047.435 ;
    END
  END DIG_MON_COMP[100]
  PIN DIG_MON_SEL[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14097.785 1046.435 14098.065 1047.435 ;
    END
  END DIG_MON_SEL[323]
  PIN MASKV[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14093.865 1046.435 14094.145 1047.435 ;
    END
  END MASKV[323]
  PIN Data_COMP[1037]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14052.985 1046.435 14053.265 1047.435 ;
    END
  END Data_COMP[1037]
  PIN Data_COMP[1034]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14051.305 1046.435 14051.585 1047.435 ;
    END
  END Data_COMP[1034]
  PIN Data_COMP[1036]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14049.065 1046.435 14049.345 1047.435 ;
    END
  END Data_COMP[1036]
  PIN INJ_IN[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14047.385 1046.435 14047.665 1047.435 ;
    END
  END INJ_IN[323]
  PIN BcidMtx[970]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14044.585 1046.435 14044.865 1047.435 ;
    END
  END BcidMtx[970]
  PIN Read_COMP[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14042.905 1046.435 14043.185 1047.435 ;
    END
  END Read_COMP[49]
  PIN BcidMtx[967]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14041.785 1046.435 14042.065 1047.435 ;
    END
  END BcidMtx[967]
  PIN INJ_IN[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14031.705 1046.435 14031.985 1047.435 ;
    END
  END INJ_IN[322]
  PIN Data_COMP[1039]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14028.345 1046.435 14028.625 1047.435 ;
    END
  END Data_COMP[1039]
  PIN Data_COMP[1045]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14027.225 1046.435 14027.505 1047.435 ;
    END
  END Data_COMP[1045]
  PIN Data_COMP[1029]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14025.545 1046.435 14025.825 1047.435 ;
    END
  END Data_COMP[1029]
  PIN MASKV[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14022.465 1046.435 14022.745 1047.435 ;
    END
  END MASKV[322]
  PIN DIG_MON_SEL[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18725.065 1046.435 18725.345 1047.435 ;
    END
  END DIG_MON_SEL[439]
  PIN FREEZE_COMP[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14273.065 1046.435 14273.345 1047.435 ;
    END
  END FREEZE_COMP[52]
  PIN DIG_MON_HV[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15109.705 1046.435 15109.985 1047.435 ;
    END
  END DIG_MON_HV[13]
  PIN Data_HV[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15107.465 1046.435 15107.745 1047.435 ;
    END
  END Data_HV[144]
  PIN Data_HV[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15105.785 1046.435 15106.065 1047.435 ;
    END
  END Data_HV[145]
  PIN Data_HV[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15104.105 1046.435 15104.385 1047.435 ;
    END
  END Data_HV[146]
  PIN Data_HV[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15102.425 1046.435 15102.705 1047.435 ;
    END
  END Data_HV[132]
  PIN INJ_IN[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15101.305 1046.435 15101.585 1047.435 ;
    END
  END INJ_IN[349]
  PIN FREEZE_HV[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15083.945 1046.435 15084.225 1047.435 ;
    END
  END FREEZE_HV[6]
  PIN BcidMtx[1045]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15082.265 1046.435 15082.545 1047.435 ;
    END
  END BcidMtx[1045]
  PIN BcidMtx[1044]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15081.705 1046.435 15081.985 1047.435 ;
    END
  END BcidMtx[1044]
  PIN Data_HV[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15078.905 1046.435 15079.185 1047.435 ;
    END
  END Data_HV[128]
  PIN Data_HV[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15076.105 1046.435 15076.385 1047.435 ;
    END
  END Data_HV[142]
  PIN Data_HV[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15075.545 1046.435 15075.825 1047.435 ;
    END
  END Data_HV[137]
  PIN Data_HV[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15073.865 1046.435 15074.145 1047.435 ;
    END
  END Data_HV[143]
  PIN DIG_MON_SEL[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15030.745 1046.435 15031.025 1047.435 ;
    END
  END DIG_MON_SEL[348]
  PIN DIG_MON_HV[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15027.945 1046.435 15028.225 1047.435 ;
    END
  END DIG_MON_HV[11]
  PIN Data_HV[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15025.705 1046.435 15025.985 1047.435 ;
    END
  END Data_HV[123]
  PIN Data_HV[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15024.025 1046.435 15024.305 1047.435 ;
    END
  END Data_HV[124]
  PIN Data_HV[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15022.345 1046.435 15022.625 1047.435 ;
    END
  END Data_HV[125]
  PIN Data_HV[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15012.265 1046.435 15012.545 1047.435 ;
    END
  END Data_HV[111]
  PIN BcidMtx[1043]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15008.905 1046.435 15009.185 1047.435 ;
    END
  END BcidMtx[1043]
  PIN BcidMtx[1042]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15008.345 1046.435 15008.625 1047.435 ;
    END
  END BcidMtx[1042]
  PIN BcidMtx[1039]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15005.545 1046.435 15005.825 1047.435 ;
    END
  END BcidMtx[1039]
  PIN Data_HV[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15000.785 1046.435 15001.065 1047.435 ;
    END
  END Data_HV[108]
  PIN Data_HV[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14999.105 1046.435 14999.385 1047.435 ;
    END
  END Data_HV[120]
  PIN Data_HV[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14971.945 1046.435 14972.225 1047.435 ;
    END
  END Data_HV[121]
  PIN Data_HV[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14970.265 1046.435 14970.545 1047.435 ;
    END
  END Data_HV[105]
  PIN Data_HV[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14969.705 1046.435 14969.985 1047.435 ;
    END
  END Data_HV[122]
  PIN MASKD[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14963.545 1046.435 14963.825 1047.435 ;
    END
  END MASKD[345]
  PIN DIG_MON_HV[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14962.425 1046.435 14962.705 1047.435 ;
    END
  END DIG_MON_HV[9]
  PIN Data_HV[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14946.185 1046.435 14946.465 1047.435 ;
    END
  END Data_HV[96]
  PIN Data_HV[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14944.505 1046.435 14944.785 1047.435 ;
    END
  END Data_HV[97]
  PIN Data_HV[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14942.825 1046.435 14943.105 1047.435 ;
    END
  END Data_HV[91]
  PIN nTOK_HV[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14940.025 1046.435 14940.305 1047.435 ;
    END
  END nTOK_HV[4]
  PIN BcidMtx[1035]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14937.785 1046.435 14938.065 1047.435 ;
    END
  END BcidMtx[1035]
  PIN BcidMtx[1034]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14936.105 1046.435 14936.385 1047.435 ;
    END
  END BcidMtx[1034]
  PIN INJ_IN[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14933.865 1046.435 14934.145 1047.435 ;
    END
  END INJ_IN[344]
  PIN DIG_MON_HV[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18740.185 1046.435 18740.465 1047.435 ;
    END
  END DIG_MON_HV[104]
  PIN Data_HV[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14892.985 1046.435 14893.265 1047.435 ;
    END
  END Data_HV[93]
  PIN Data_HV[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14890.185 1046.435 14890.465 1047.435 ;
    END
  END Data_HV[95]
  PIN Data_HV[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14888.505 1046.435 14888.785 1047.435 ;
    END
  END Data_HV[101]
  PIN MASKD[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14886.825 1046.435 14887.105 1047.435 ;
    END
  END MASKD[344]
  PIN DIG_MON_SEL[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14884.025 1046.435 14884.305 1047.435 ;
    END
  END DIG_MON_SEL[344]
  PIN DIG_MON_HV[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14881.225 1046.435 14881.505 1047.435 ;
    END
  END DIG_MON_HV[7]
  PIN Data_HV[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14870.585 1046.435 14870.865 1047.435 ;
    END
  END Data_HV[81]
  PIN Data_HV[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14868.905 1046.435 14869.185 1047.435 ;
    END
  END Data_HV[82]
  PIN Data_HV[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14867.225 1046.435 14867.505 1047.435 ;
    END
  END Data_HV[83]
  PIN Data_HV[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14865.545 1046.435 14865.825 1047.435 ;
    END
  END Data_HV[69]
  PIN BcidMtx[1031]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14860.225 1046.435 14860.505 1047.435 ;
    END
  END BcidMtx[1031]
  PIN Read_HV[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14832.505 1046.435 14832.785 1047.435 ;
    END
  END Read_HV[3]
  PIN BcidMtx[1028]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14831.945 1046.435 14832.225 1047.435 ;
    END
  END BcidMtx[1028]
  PIN Data_HV[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14828.025 1046.435 14828.305 1047.435 ;
    END
  END Data_HV[65]
  PIN Data_HV[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14826.345 1046.435 14826.625 1047.435 ;
    END
  END Data_HV[73]
  PIN Data_HV[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14825.785 1046.435 14826.065 1047.435 ;
    END
  END Data_HV[67]
  PIN Data_HV[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14822.985 1046.435 14823.265 1047.435 ;
    END
  END Data_HV[80]
  PIN MASKD[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14821.305 1046.435 14821.585 1047.435 ;
    END
  END MASKD[342]
  PIN DIG_MON_SEL[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14805.625 1046.435 14805.905 1047.435 ;
    END
  END DIG_MON_SEL[342]
  PIN MASKD[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15363.945 1046.435 15364.225 1047.435 ;
    END
  END MASKD[355]
  PIN MASKV[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15361.145 1046.435 15361.425 1047.435 ;
    END
  END MASKV[355]
  PIN Data_HV[201]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15359.465 1046.435 15359.745 1047.435 ;
    END
  END Data_HV[201]
  PIN Data_HV[202]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15357.785 1046.435 15358.065 1047.435 ;
    END
  END Data_HV[202]
  PIN Data_HV[196]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15356.105 1046.435 15356.385 1047.435 ;
    END
  END Data_HV[196]
  PIN nTOK_HV[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15314.105 1046.435 15314.385 1047.435 ;
    END
  END nTOK_HV[9]
  PIN BcidMtx[1065]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15311.865 1046.435 15312.145 1047.435 ;
    END
  END BcidMtx[1065]
  PIN MASKV[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18721.145 1046.435 18721.425 1047.435 ;
    END
  END MASKV[439]
  PIN BcidMtx[1062]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15309.065 1046.435 15309.345 1047.435 ;
    END
  END BcidMtx[1062]
  PIN Data_HV[1079]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18720.025 1046.435 18720.305 1047.435 ;
    END
  END Data_HV[1079]
  PIN Data_HV[198]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15305.705 1046.435 15305.985 1047.435 ;
    END
  END Data_HV[198]
  PIN Data_HV[193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15304.025 1046.435 15304.305 1047.435 ;
    END
  END Data_HV[193]
  PIN Data_HV[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15302.345 1046.435 15302.625 1047.435 ;
    END
  END Data_HV[190]
  PIN MASKV[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15292.265 1046.435 15292.545 1047.435 ;
    END
  END MASKV[354]
  PIN DIG_MON_HV[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15290.025 1046.435 15290.305 1047.435 ;
    END
  END DIG_MON_HV[18]
  PIN DIG_MON_SEL[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15287.785 1046.435 15288.065 1047.435 ;
    END
  END DIG_MON_SEL[353]
  PIN INJ_ROW[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15282.465 1046.435 15282.745 1047.435 ;
    END
  END INJ_ROW[176]
  PIN Data_HV[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15280.785 1046.435 15281.065 1047.435 ;
    END
  END Data_HV[176]
  PIN Data_HV[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15279.105 1046.435 15279.385 1047.435 ;
    END
  END Data_HV[173]
  PIN Data_HV[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15251.945 1046.435 15252.225 1047.435 ;
    END
  END Data_HV[182]
  PIN INJ_IN[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15249.705 1046.435 15249.985 1047.435 ;
    END
  END INJ_IN[353]
  PIN BcidMtx[1060]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15246.905 1046.435 15247.185 1047.435 ;
    END
  END BcidMtx[1060]
  PIN Read_HV[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15245.225 1046.435 15245.505 1047.435 ;
    END
  END Read_HV[8]
  PIN BcidMtx[1056]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15243.545 1046.435 15243.825 1047.435 ;
    END
  END BcidMtx[1056]
  PIN Data_HV[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15240.745 1046.435 15241.025 1047.435 ;
    END
  END Data_HV[170]
  PIN Data_HV[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15226.185 1046.435 15226.465 1047.435 ;
    END
  END Data_HV[178]
  PIN Data_HV[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15224.505 1046.435 15224.785 1047.435 ;
    END
  END Data_HV[179]
  PIN Data_HV[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15222.825 1046.435 15223.105 1047.435 ;
    END
  END Data_HV[185]
  PIN MASKD[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15221.145 1046.435 15221.425 1047.435 ;
    END
  END MASKD[352]
  PIN DIG_MON_SEL[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15218.345 1046.435 15218.625 1047.435 ;
    END
  END DIG_MON_SEL[352]
  PIN DIG_MON_HV[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15215.545 1046.435 15215.825 1047.435 ;
    END
  END DIG_MON_HV[15]
  PIN Data_HV[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15173.545 1046.435 15173.825 1047.435 ;
    END
  END Data_HV[165]
  PIN Data_HV[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15171.865 1046.435 15172.145 1047.435 ;
    END
  END Data_HV[166]
  PIN Data_HV[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15170.185 1046.435 15170.465 1047.435 ;
    END
  END Data_HV[167]
  PIN Data_HV[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15168.505 1046.435 15168.785 1047.435 ;
    END
  END Data_HV[153]
  PIN BcidMtx[1055]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15165.145 1046.435 15165.425 1047.435 ;
    END
  END BcidMtx[1055]
  PIN FREEZE_HV[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15163.465 1046.435 15163.745 1047.435 ;
    END
  END FREEZE_HV[7]
  PIN BcidMtx[1051]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15161.785 1046.435 15162.065 1047.435 ;
    END
  END BcidMtx[1051]
  PIN Data_HV[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15150.585 1046.435 15150.865 1047.435 ;
    END
  END Data_HV[150]
  PIN Data_HV[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15149.465 1046.435 15149.745 1047.435 ;
    END
  END Data_HV[156]
  PIN Data_HV[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15147.785 1046.435 15148.065 1047.435 ;
    END
  END Data_HV[151]
  PIN Data_HV[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15146.105 1046.435 15146.385 1047.435 ;
    END
  END Data_HV[148]
  PIN MASKV[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15142.465 1046.435 15142.745 1047.435 ;
    END
  END MASKV[350]
  PIN DIG_MON_HV[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15140.225 1046.435 15140.505 1047.435 ;
    END
  END DIG_MON_HV[14]
  PIN FREEZE_HV[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15393.065 1046.435 15393.345 1047.435 ;
    END
  END FREEZE_HV[10]
  PIN DIG_MON_HV[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16229.705 1046.435 16229.985 1047.435 ;
    END
  END DIG_MON_HV[41]
  PIN Data_HV[438]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16227.465 1046.435 16227.745 1047.435 ;
    END
  END Data_HV[438]
  PIN Data_HV[439]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16225.785 1046.435 16226.065 1047.435 ;
    END
  END Data_HV[439]
  PIN Data_HV[440]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16224.105 1046.435 16224.385 1047.435 ;
    END
  END Data_HV[440]
  PIN Data_HV[426]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16222.425 1046.435 16222.705 1047.435 ;
    END
  END Data_HV[426]
  PIN BcidMtx[1133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16205.625 1046.435 16205.905 1047.435 ;
    END
  END BcidMtx[1133]
  PIN FREEZE_HV[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16203.945 1046.435 16204.225 1047.435 ;
    END
  END FREEZE_HV[20]
  PIN BcidMtx[1129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16202.265 1046.435 16202.545 1047.435 ;
    END
  END BcidMtx[1129]
  PIN Data_HV[423]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16199.465 1046.435 16199.745 1047.435 ;
    END
  END Data_HV[423]
  PIN Data_HV[430]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16197.225 1046.435 16197.505 1047.435 ;
    END
  END Data_HV[430]
  PIN Data_HV[436]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16196.105 1046.435 16196.385 1047.435 ;
    END
  END Data_HV[436]
  PIN Data_HV[420]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16194.425 1046.435 16194.705 1047.435 ;
    END
  END Data_HV[420]
  PIN MASKD[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16153.545 1046.435 16153.825 1047.435 ;
    END
  END MASKD[376]
  PIN MASKD[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16149.065 1046.435 16149.345 1047.435 ;
    END
  END MASKD[375]
  PIN Data_HV[417]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16145.705 1046.435 16145.985 1047.435 ;
    END
  END Data_HV[417]
  PIN Data_HV[411]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16144.585 1046.435 16144.865 1047.435 ;
    END
  END Data_HV[411]
  PIN Data_HV[412]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16142.905 1046.435 16143.185 1047.435 ;
    END
  END Data_HV[412]
  PIN Data_HV[405]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16132.265 1046.435 16132.545 1047.435 ;
    END
  END Data_HV[405]
  PIN nTOK_HV[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16130.025 1046.435 16130.305 1047.435 ;
    END
  END nTOK_HV[19]
  PIN BcidMtx[1125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16127.785 1046.435 16128.065 1047.435 ;
    END
  END BcidMtx[1125]
  PIN BcidMtx[1123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16125.545 1046.435 16125.825 1047.435 ;
    END
  END BcidMtx[1123]
  PIN INJ_IN[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16121.905 1046.435 16122.185 1047.435 ;
    END
  END INJ_IN[374]
  PIN Data_HV[408]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16119.665 1046.435 16119.945 1047.435 ;
    END
  END Data_HV[408]
  PIN Data_HV[403]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16092.505 1046.435 16092.785 1047.435 ;
    END
  END Data_HV[403]
  PIN Data_HV[400]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16090.825 1046.435 16091.105 1047.435 ;
    END
  END Data_HV[400]
  PIN MASKV[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16089.145 1046.435 16089.425 1047.435 ;
    END
  END MASKV[374]
  PIN DIG_MON_SEL[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16084.665 1046.435 16084.945 1047.435 ;
    END
  END DIG_MON_SEL[373]
  PIN INJ_ROW[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16081.305 1046.435 16081.585 1047.435 ;
    END
  END INJ_ROW[186]
  PIN Data_HV[390]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16066.185 1046.435 16066.465 1047.435 ;
    END
  END Data_HV[390]
  PIN Data_HV[383]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16065.065 1046.435 16065.345 1047.435 ;
    END
  END Data_HV[383]
  PIN Data_HV[392]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16063.385 1046.435 16063.665 1047.435 ;
    END
  END Data_HV[392]
  PIN INJ_IN[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16061.145 1046.435 16061.425 1047.435 ;
    END
  END INJ_IN[373]
  PIN BcidMtx[1120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16058.345 1046.435 16058.625 1047.435 ;
    END
  END BcidMtx[1120]
  PIN Read_HV[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16056.665 1046.435 16056.945 1047.435 ;
    END
  END Read_HV[18]
  PIN BcidMtx[1116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16054.985 1046.435 16055.265 1047.435 ;
    END
  END BcidMtx[1116]
  PIN Data_HV[380]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16013.545 1046.435 16013.825 1047.435 ;
    END
  END Data_HV[380]
  PIN Data_HV[388]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16011.865 1046.435 16012.145 1047.435 ;
    END
  END Data_HV[388]
  PIN Data_HV[379]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16009.625 1046.435 16009.905 1047.435 ;
    END
  END Data_HV[379]
  PIN Data_HV[395]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16008.505 1046.435 16008.785 1047.435 ;
    END
  END Data_HV[395]
  PIN MASKD[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16006.825 1046.435 16007.105 1047.435 ;
    END
  END MASKD[372]
  PIN DIG_MON_SEL[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16003.465 1046.435 16003.745 1047.435 ;
    END
  END DIG_MON_SEL[371]
  PIN DIG_MON_HV[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16001.225 1046.435 16001.505 1047.435 ;
    END
  END DIG_MON_HV[35]
  PIN Data_HV[375]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15990.585 1046.435 15990.865 1047.435 ;
    END
  END Data_HV[375]
  PIN Data_HV[362]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15988.345 1046.435 15988.625 1047.435 ;
    END
  END Data_HV[362]
  PIN Data_HV[370]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15987.785 1046.435 15988.065 1047.435 ;
    END
  END Data_HV[370]
  PIN Data_HV[364]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15986.105 1046.435 15986.385 1047.435 ;
    END
  END Data_HV[364]
  PIN nTOK_HV[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15981.345 1046.435 15981.625 1047.435 ;
    END
  END nTOK_HV[17]
  PIN Data_HV[1084]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18717.785 1046.435 18718.065 1047.435 ;
    END
  END Data_HV[1084]
  PIN Read_HV[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15952.505 1046.435 15952.785 1047.435 ;
    END
  END Read_HV[17]
  PIN INJ_IN[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15949.705 1046.435 15949.985 1047.435 ;
    END
  END INJ_IN[370]
  PIN Data_HV[359]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15948.025 1046.435 15948.305 1047.435 ;
    END
  END Data_HV[359]
  PIN Data_HV[367]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15946.345 1046.435 15946.625 1047.435 ;
    END
  END Data_HV[367]
  PIN Data_HV[358]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15944.105 1046.435 15944.385 1047.435 ;
    END
  END Data_HV[358]
  PIN MASKV[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15942.425 1046.435 15942.705 1047.435 ;
    END
  END MASKV[370]
  PIN MASKD[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15941.305 1046.435 15941.585 1047.435 ;
    END
  END MASKD[370]
  PIN INJ_IN[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2061.145 1046.435 2061.425 1047.435 ;
    END
  END INJ_IN[23]
  PIN BcidMtx[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2058.905 1046.435 2059.185 1047.435 ;
    END
  END BcidMtx[71]
  PIN FREEZE_PMOS_NOSF[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2057.225 1046.435 2057.505 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[11]
  PIN BcidMtx[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2056.105 1046.435 2056.385 1047.435 ;
    END
  END BcidMtx[68]
  PIN INJ_IN[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2053.865 1046.435 2054.145 1047.435 ;
    END
  END INJ_IN[22]
  PIN Data_PMOS_NOSF[233]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2013.545 1046.435 2013.825 1047.435 ;
    END
  END Data_PMOS_NOSF[233]
  PIN Data_PMOS_NOSF[241]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2011.865 1046.435 2012.145 1047.435 ;
    END
  END Data_PMOS_NOSF[241]
  PIN Data_PMOS_NOSF[232]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2009.625 1046.435 2009.905 1047.435 ;
    END
  END Data_PMOS_NOSF[232]
  PIN Data_PMOS_NOSF[248]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2008.505 1046.435 2008.785 1047.435 ;
    END
  END Data_PMOS_NOSF[248]
  PIN MASKD[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2006.825 1046.435 2007.105 1047.435 ;
    END
  END MASKD[22]
  PIN DIG_MON_SEL[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2004.025 1046.435 2004.305 1047.435 ;
    END
  END DIG_MON_SEL[22]
  PIN MASKD[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2002.345 1046.435 2002.625 1047.435 ;
    END
  END MASKD[21]
  PIN MASKV[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1991.145 1046.435 1991.425 1047.435 ;
    END
  END MASKV[21]
  PIN Data_PMOS_NOSF[229]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1988.905 1046.435 1989.185 1047.435 ;
    END
  END Data_PMOS_NOSF[229]
  PIN Data_PMOS_NOSF[223]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1987.785 1046.435 1988.065 1047.435 ;
    END
  END Data_PMOS_NOSF[223]
  PIN Data_PMOS_NOSF[217]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1986.105 1046.435 1986.385 1047.435 ;
    END
  END Data_PMOS_NOSF[217]
  PIN BcidMtx[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1980.225 1046.435 1980.505 1047.435 ;
    END
  END BcidMtx[65]
  PIN BcidMtx[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1979.105 1046.435 1979.385 1047.435 ;
    END
  END BcidMtx[63]
  PIN BcidMtx[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1951.385 1046.435 1951.665 1047.435 ;
    END
  END BcidMtx[61]
  PIN INJ_IN[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1949.705 1046.435 1949.985 1047.435 ;
    END
  END INJ_IN[20]
  PIN Data_PMOS_NOSF[225]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1946.905 1046.435 1947.185 1047.435 ;
    END
  END Data_PMOS_NOSF[225]
  PIN Data_PMOS_NOSF[214]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1945.785 1046.435 1946.065 1047.435 ;
    END
  END Data_PMOS_NOSF[214]
  PIN Data_PMOS_NOSF[227]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1942.985 1046.435 1943.265 1047.435 ;
    END
  END Data_PMOS_NOSF[227]
  PIN DIG_MON_PMOS_NOSF[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1940.185 1046.435 1940.465 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[20]
  PIN DIG_MON_SEL[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1925.625 1046.435 1925.905 1047.435 ;
    END
  END DIG_MON_SEL[20]
  PIN INJ_ROW[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1921.705 1046.435 1921.985 1047.435 ;
    END
  END INJ_ROW[9]
  PIN Data_PMOS_NOSF[197]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1920.025 1046.435 1920.305 1047.435 ;
    END
  END Data_PMOS_NOSF[197]
  PIN Data_PMOS_NOSF[194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1918.345 1046.435 1918.625 1047.435 ;
    END
  END Data_PMOS_NOSF[194]
  PIN Data_PMOS_NOSF[203]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1916.665 1046.435 1916.945 1047.435 ;
    END
  END Data_PMOS_NOSF[203]
  PIN INJ_IN[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1914.425 1046.435 1914.705 1047.435 ;
    END
  END INJ_IN[19]
  PIN BcidMtx[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1872.425 1046.435 1872.705 1047.435 ;
    END
  END BcidMtx[58]
  PIN BcidMtx[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1870.185 1046.435 1870.465 1047.435 ;
    END
  END BcidMtx[56]
  PIN BcidMtx[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1869.065 1046.435 1869.345 1047.435 ;
    END
  END BcidMtx[54]
  PIN Data_PMOS_NOSF[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1866.265 1046.435 1866.545 1047.435 ;
    END
  END Data_PMOS_NOSF[191]
  PIN Data_PMOS_NOSF[193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1864.025 1046.435 1864.305 1047.435 ;
    END
  END Data_PMOS_NOSF[193]
  PIN Data_PMOS_NOSF[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1862.345 1046.435 1862.625 1047.435 ;
    END
  END Data_PMOS_NOSF[190]
  PIN Data_PMOS_NOSF[206]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1861.225 1046.435 1861.505 1047.435 ;
    END
  END Data_PMOS_NOSF[206]
  PIN DIG_MON_PMOS_NOSF[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1850.025 1046.435 1850.305 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[18]
  PIN DIG_MON_SEL[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1847.785 1046.435 1848.065 1047.435 ;
    END
  END DIG_MON_SEL[17]
  PIN DIG_MON_PMOS_NOSF[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1845.545 1046.435 1845.825 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[17]
  PIN Data_PMOS_NOSF[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1840.785 1046.435 1841.065 1047.435 ;
    END
  END Data_PMOS_NOSF[176]
  PIN Data_PMOS_NOSF[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1839.105 1046.435 1839.385 1047.435 ;
    END
  END Data_PMOS_NOSF[173]
  PIN Data_PMOS_NOSF[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1811.945 1046.435 1812.225 1047.435 ;
    END
  END Data_PMOS_NOSF[182]
  PIN INJ_IN[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1809.705 1046.435 1809.985 1047.435 ;
    END
  END INJ_IN[17]
  PIN BcidMtx[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1806.905 1046.435 1807.185 1047.435 ;
    END
  END BcidMtx[52]
  PIN Read_PMOS_NOSF[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1805.225 1046.435 1805.505 1047.435 ;
    END
  END Read_PMOS_NOSF[8]
  PIN INJ_IN[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1802.425 1046.435 1802.705 1047.435 ;
    END
  END INJ_IN[16]
  PIN Data_PMOS_NOSF[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1800.745 1046.435 1801.025 1047.435 ;
    END
  END Data_PMOS_NOSF[170]
  PIN Data_PMOS_NOSF[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1786.185 1046.435 1786.465 1047.435 ;
    END
  END Data_PMOS_NOSF[178]
  PIN Data_HV[1067]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18582.825 1046.435 18583.105 1047.435 ;
    END
  END Data_HV[1067]
  PIN Data_PMOS_NOSF[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1783.385 1046.435 1783.665 1047.435 ;
    END
  END Data_PMOS_NOSF[168]
  PIN MASKH[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1781.705 1046.435 1781.985 1047.435 ;
    END
  END MASKH[8]
  PIN DIG_MON_SEL[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1778.345 1046.435 1778.625 1047.435 ;
    END
  END DIG_MON_SEL[16]
  PIN DIG_MON_PMOS_NOSF[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1775.545 1046.435 1775.825 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[15]
  PIN Data_PMOS_NOSF[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1733.545 1046.435 1733.825 1047.435 ;
    END
  END Data_PMOS_NOSF[165]
  PIN Data_PMOS_NOSF[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1731.305 1046.435 1731.585 1047.435 ;
    END
  END Data_PMOS_NOSF[152]
  PIN Data_PMOS_NOSF[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1730.185 1046.435 1730.465 1047.435 ;
    END
  END Data_PMOS_NOSF[167]
  PIN Data_PMOS_NOSF[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1728.505 1046.435 1728.785 1047.435 ;
    END
  END Data_PMOS_NOSF[153]
  PIN BcidMtx[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1725.145 1046.435 1725.425 1047.435 ;
    END
  END BcidMtx[47]
  PIN FREEZE_PMOS_NOSF[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1723.465 1046.435 1723.745 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[7]
  PIN BcidMtx[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1721.785 1046.435 1722.065 1047.435 ;
    END
  END BcidMtx[43]
  PIN Data_PMOS_NOSF[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1710.585 1046.435 1710.865 1047.435 ;
    END
  END Data_PMOS_NOSF[150]
  PIN Data_PMOS_NOSF[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1708.905 1046.435 1709.185 1047.435 ;
    END
  END Data_PMOS_NOSF[162]
  PIN Data_PMOS_NOSF[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1707.225 1046.435 1707.505 1047.435 ;
    END
  END Data_PMOS_NOSF[163]
  PIN Data_PMOS_NOSF[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.985 1046.435 1705.265 1047.435 ;
    END
  END Data_PMOS_NOSF[164]
  PIN MASKH[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1701.905 1046.435 1702.185 1047.435 ;
    END
  END MASKH[7]
  PIN DIG_MON_PMOS_NOSF[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1700.225 1046.435 1700.505 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[14]
  PIN FREEZE_PMOS_NOSF[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1953.065 1046.435 1953.345 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[10]
  PIN DIG_MON_PMOS_NOSF[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2789.705 1046.435 2789.985 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[41]
  PIN Data_PMOS_NOSF[438]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2787.465 1046.435 2787.745 1047.435 ;
    END
  END Data_PMOS_NOSF[438]
  PIN Data_PMOS_NOSF[439]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2785.785 1046.435 2786.065 1047.435 ;
    END
  END Data_PMOS_NOSF[439]
  PIN Data_PMOS_NOSF[440]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2784.105 1046.435 2784.385 1047.435 ;
    END
  END Data_PMOS_NOSF[440]
  PIN Data_PMOS_NOSF[426]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2782.425 1046.435 2782.705 1047.435 ;
    END
  END Data_PMOS_NOSF[426]
  PIN BcidMtx[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2765.625 1046.435 2765.905 1047.435 ;
    END
  END BcidMtx[125]
  PIN FREEZE_PMOS_NOSF[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2763.945 1046.435 2764.225 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[20]
  PIN BcidMtx[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2762.265 1046.435 2762.545 1047.435 ;
    END
  END BcidMtx[121]
  PIN Data_PMOS_NOSF[422]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2758.905 1046.435 2759.185 1047.435 ;
    END
  END Data_PMOS_NOSF[422]
  PIN Data_PMOS_NOSF[435]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2757.785 1046.435 2758.065 1047.435 ;
    END
  END Data_PMOS_NOSF[435]
  PIN Data_PMOS_NOSF[436]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2756.105 1046.435 2756.385 1047.435 ;
    END
  END Data_PMOS_NOSF[436]
  PIN Data_PMOS_NOSF[437]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2753.865 1046.435 2754.145 1047.435 ;
    END
  END Data_PMOS_NOSF[437]
  PIN MASKV[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2714.665 1046.435 2714.945 1047.435 ;
    END
  END MASKV[40]
  PIN DIG_MON_PMOS_NOSF[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2712.425 1046.435 2712.705 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[40]
  PIN DIG_MON_SEL[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2710.185 1046.435 2710.465 1047.435 ;
    END
  END DIG_MON_SEL[39]
  PIN INJ_ROW[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2706.825 1046.435 2707.105 1047.435 ;
    END
  END INJ_ROW[19]
  PIN Data_PMOS_NOSF[411]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2704.585 1046.435 2704.865 1047.435 ;
    END
  END Data_PMOS_NOSF[411]
  PIN Data_PMOS_NOSF[418]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2704.025 1046.435 2704.305 1047.435 ;
    END
  END Data_PMOS_NOSF[418]
  PIN Data_PMOS_NOSF[406]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2701.225 1046.435 2701.505 1047.435 ;
    END
  END Data_PMOS_NOSF[406]
  PIN INJ_IN[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2691.145 1046.435 2691.425 1047.435 ;
    END
  END INJ_IN[39]
  PIN BcidMtx[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2688.345 1046.435 2688.625 1047.435 ;
    END
  END BcidMtx[118]
  PIN Read_PMOS_NOSF[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2686.665 1046.435 2686.945 1047.435 ;
    END
  END Read_PMOS_NOSF[19]
  PIN BcidMtx[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2684.985 1046.435 2685.265 1047.435 ;
    END
  END BcidMtx[114]
  PIN Data_PMOS_NOSF[355]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2478.905 1046.435 2479.185 1047.435 ;
    END
  END Data_PMOS_NOSF[355]
  PIN Data_PMOS_NOSF[414]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2679.105 1046.435 2679.385 1047.435 ;
    END
  END Data_PMOS_NOSF[414]
  PIN Data_PMOS_NOSF[415]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2651.945 1046.435 2652.225 1047.435 ;
    END
  END Data_PMOS_NOSF[415]
  PIN Data_PMOS_NOSF[399]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2650.265 1046.435 2650.545 1047.435 ;
    END
  END Data_PMOS_NOSF[399]
  PIN MASKV[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2649.145 1046.435 2649.425 1047.435 ;
    END
  END MASKV[38]
  PIN DIG_MON_PMOS_NOSF[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2646.905 1046.435 2647.185 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[38]
  PIN MASKD[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2643.545 1046.435 2643.825 1047.435 ;
    END
  END MASKD[37]
  PIN INJ_ROW[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2641.305 1046.435 2641.585 1047.435 ;
    END
  END INJ_ROW[18]
  PIN Data_PMOS_NOSF[386]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2639.625 1046.435 2639.905 1047.435 ;
    END
  END Data_PMOS_NOSF[386]
  PIN Data_PMOS_NOSF[398]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2623.945 1046.435 2624.225 1047.435 ;
    END
  END Data_PMOS_NOSF[398]
  PIN Data_PMOS_NOSF[385]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2622.825 1046.435 2623.105 1047.435 ;
    END
  END Data_PMOS_NOSF[385]
  PIN INJ_IN[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3181.145 1046.435 3181.425 1047.435 ;
    END
  END INJ_IN[51]
  PIN BcidMtx[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3178.345 1046.435 3178.625 1047.435 ;
    END
  END BcidMtx[154]
  PIN Read_PMOS_NOSF[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3176.665 1046.435 3176.945 1047.435 ;
    END
  END Read_PMOS_NOSF[25]
  PIN INJ_IN[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3173.865 1046.435 3174.145 1047.435 ;
    END
  END INJ_IN[50]
  PIN Data_PMOS_NOSF[527]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3133.545 1046.435 3133.825 1047.435 ;
    END
  END Data_PMOS_NOSF[527]
  PIN Data_PMOS_NOSF[535]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3131.865 1046.435 3132.145 1047.435 ;
    END
  END Data_PMOS_NOSF[535]
  PIN Data_PMOS_NOSF[525]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3129.065 1046.435 3129.345 1047.435 ;
    END
  END Data_PMOS_NOSF[525]
  PIN MASKH[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3127.385 1046.435 3127.665 1047.435 ;
    END
  END MASKH[25]
  PIN MASKD[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3122.345 1046.435 3122.625 1047.435 ;
    END
  END MASKD[49]
  PIN MASKV[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3111.145 1046.435 3111.425 1047.435 ;
    END
  END MASKV[49]
  PIN Data_PMOS_NOSF[516]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3109.465 1046.435 3109.745 1047.435 ;
    END
  END Data_PMOS_NOSF[516]
  PIN Data_PMOS_NOSF[517]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3107.785 1046.435 3108.065 1047.435 ;
    END
  END Data_PMOS_NOSF[517]
  PIN Data_PMOS_NOSF[511]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3106.105 1046.435 3106.385 1047.435 ;
    END
  END Data_PMOS_NOSF[511]
  PIN BcidMtx[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3100.225 1046.435 3100.505 1047.435 ;
    END
  END BcidMtx[149]
  PIN BcidMtx[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3099.105 1046.435 3099.385 1047.435 ;
    END
  END BcidMtx[147]
  PIN BcidMtx[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3071.385 1046.435 3071.665 1047.435 ;
    END
  END BcidMtx[145]
  PIN Data_PMOS_NOSF[506]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3068.025 1046.435 3068.305 1047.435 ;
    END
  END Data_PMOS_NOSF[506]
  PIN Data_PMOS_NOSF[519]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3066.905 1046.435 3067.185 1047.435 ;
    END
  END Data_PMOS_NOSF[519]
  PIN Data_PMOS_NOSF[520]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3065.225 1046.435 3065.505 1047.435 ;
    END
  END Data_PMOS_NOSF[520]
  PIN Data_PMOS_NOSF[521]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3062.985 1046.435 3063.265 1047.435 ;
    END
  END Data_PMOS_NOSF[521]
  PIN MASKH[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3061.865 1046.435 3062.145 1047.435 ;
    END
  END MASKH[24]
  PIN DIG_MON_PMOS_NOSF[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3042.825 1046.435 3043.105 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[47]
  PIN MASKV[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3041.145 1046.435 3041.425 1047.435 ;
    END
  END MASKV[47]
  PIN Data_PMOS_NOSF[495]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3039.465 1046.435 3039.745 1047.435 ;
    END
  END Data_PMOS_NOSF[495]
  PIN Data_PMOS_NOSF[503]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3037.225 1046.435 3037.505 1047.435 ;
    END
  END Data_PMOS_NOSF[503]
  PIN Data_PMOS_NOSF[490]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3036.105 1046.435 3036.385 1047.435 ;
    END
  END Data_PMOS_NOSF[490]
  PIN nTOK_PMOS_NOSF[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2994.105 1046.435 2994.385 1047.435 ;
    END
  END nTOK_PMOS_NOSF[23]
  PIN BcidMtx[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2991.865 1046.435 2992.145 1047.435 ;
    END
  END BcidMtx[141]
  PIN BcidMtx[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2990.185 1046.435 2990.465 1047.435 ;
    END
  END BcidMtx[140]
  PIN INJ_IN[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2987.945 1046.435 2988.225 1047.435 ;
    END
  END INJ_IN[46]
  PIN Data_PMOS_NOSF[492]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2985.705 1046.435 2985.985 1047.435 ;
    END
  END Data_PMOS_NOSF[492]
  PIN Data_PMOS_NOSF[487]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2984.025 1046.435 2984.305 1047.435 ;
    END
  END Data_PMOS_NOSF[487]
  PIN Data_PMOS_NOSF[484]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2982.345 1046.435 2982.625 1047.435 ;
    END
  END Data_PMOS_NOSF[484]
  PIN MASKV[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2972.265 1046.435 2972.545 1047.435 ;
    END
  END MASKV[46]
  PIN MASKD[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2971.145 1046.435 2971.425 1047.435 ;
    END
  END MASKD[46]
  PIN DIG_MON_SEL[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2967.785 1046.435 2968.065 1047.435 ;
    END
  END DIG_MON_SEL[45]
  PIN INJ_ROW[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2962.465 1046.435 2962.745 1047.435 ;
    END
  END INJ_ROW[22]
  PIN Data_PMOS_NOSF[480]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2961.345 1046.435 2961.625 1047.435 ;
    END
  END Data_PMOS_NOSF[480]
  PIN Data_PMOS_NOSF[467]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2959.105 1046.435 2959.385 1047.435 ;
    END
  END Data_PMOS_NOSF[467]
  PIN Data_PMOS_NOSF[476]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2931.945 1046.435 2932.225 1047.435 ;
    END
  END Data_PMOS_NOSF[476]
  PIN Data_PMOS_NOSF[469]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2931.385 1046.435 2931.665 1047.435 ;
    END
  END Data_PMOS_NOSF[469]
  PIN BcidMtx[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2926.905 1046.435 2927.185 1047.435 ;
    END
  END BcidMtx[136]
  PIN Read_PMOS_NOSF[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2925.225 1046.435 2925.505 1047.435 ;
    END
  END Read_PMOS_NOSF[22]
  PIN Data_HV[1086]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18665.145 1046.435 18665.425 1047.435 ;
    END
  END Data_HV[1086]
  PIN INJ_IN[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2922.425 1046.435 2922.705 1047.435 ;
    END
  END INJ_IN[44]
  PIN Data_PMOS_NOSF[471]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2920.185 1046.435 2920.465 1047.435 ;
    END
  END Data_PMOS_NOSF[471]
  PIN Data_PMOS_NOSF[472]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2906.185 1046.435 2906.465 1047.435 ;
    END
  END Data_PMOS_NOSF[472]
  PIN Data_PMOS_NOSF[463]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2903.945 1046.435 2904.225 1047.435 ;
    END
  END Data_PMOS_NOSF[463]
  PIN MASKV[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2902.265 1046.435 2902.545 1047.435 ;
    END
  END MASKV[44]
  PIN DIG_MON_PMOS_NOSF[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2900.025 1046.435 2900.305 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[44]
  PIN DIG_MON_SEL[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2897.785 1046.435 2898.065 1047.435 ;
    END
  END DIG_MON_SEL[43]
  PIN INJ_ROW[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2894.425 1046.435 2894.705 1047.435 ;
    END
  END INJ_ROW[21]
  PIN Data_PMOS_NOSF[459]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2853.545 1046.435 2853.825 1047.435 ;
    END
  END Data_PMOS_NOSF[459]
  PIN Data_PMOS_NOSF[446]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2851.305 1046.435 2851.585 1047.435 ;
    END
  END Data_PMOS_NOSF[446]
  PIN Data_PMOS_NOSF[455]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2849.625 1046.435 2849.905 1047.435 ;
    END
  END Data_PMOS_NOSF[455]
  PIN INJ_IN[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2847.385 1046.435 2847.665 1047.435 ;
    END
  END INJ_IN[43]
  PIN BcidMtx[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2844.585 1046.435 2844.865 1047.435 ;
    END
  END BcidMtx[130]
  PIN Read_PMOS_NOSF[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2842.905 1046.435 2843.185 1047.435 ;
    END
  END Read_PMOS_NOSF[21]
  PIN BcidMtx[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2841.785 1046.435 2842.065 1047.435 ;
    END
  END BcidMtx[127]
  PIN Data_PMOS_NOSF[444]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2830.585 1046.435 2830.865 1047.435 ;
    END
  END Data_PMOS_NOSF[444]
  PIN Data_PMOS_NOSF[456]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2828.905 1046.435 2829.185 1047.435 ;
    END
  END Data_PMOS_NOSF[456]
  PIN Data_PMOS_NOSF[457]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2827.225 1046.435 2827.505 1047.435 ;
    END
  END Data_PMOS_NOSF[457]
  PIN Data_PMOS_NOSF[441]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2825.545 1046.435 2825.825 1047.435 ;
    END
  END Data_PMOS_NOSF[441]
  PIN MASKH[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2821.905 1046.435 2822.185 1047.435 ;
    END
  END MASKH[21]
  PIN DIG_MON_PMOS_NOSF[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2820.225 1046.435 2820.505 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[42]
  PIN DIG_MON_SEL[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3911.945 1046.435 3912.225 1047.435 ;
    END
  END DIG_MON_SEL[69]
  PIN INJ_ROW[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3908.585 1046.435 3908.865 1047.435 ;
    END
  END INJ_ROW[34]
  PIN Data_PMOS_NOSF[732]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3907.465 1046.435 3907.745 1047.435 ;
    END
  END Data_PMOS_NOSF[732]
  PIN Data_PMOS_NOSF[719]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3905.225 1046.435 3905.505 1047.435 ;
    END
  END Data_PMOS_NOSF[719]
  PIN Data_PMOS_NOSF[728]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3903.545 1046.435 3903.825 1047.435 ;
    END
  END Data_PMOS_NOSF[728]
  PIN Data_PMOS_NOSF[720]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3902.425 1046.435 3902.705 1047.435 ;
    END
  END Data_PMOS_NOSF[720]
  PIN BcidMtx[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3885.065 1046.435 3885.345 1047.435 ;
    END
  END BcidMtx[208]
  PIN DIG_MON_SEL[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18884.665 1046.435 18884.945 1047.435 ;
    END
  END DIG_MON_SEL[443]
  PIN Read_PMOS_NOSF[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3883.385 1046.435 3883.665 1047.435 ;
    END
  END Read_PMOS_NOSF[34]
  PIN Data_PMOS_NOSF[717]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3879.465 1046.435 3879.745 1047.435 ;
    END
  END Data_PMOS_NOSF[717]
  PIN Data_PMOS_NOSF[729]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3877.785 1046.435 3878.065 1047.435 ;
    END
  END Data_PMOS_NOSF[729]
  PIN Data_PMOS_NOSF[718]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3876.665 1046.435 3876.945 1047.435 ;
    END
  END Data_PMOS_NOSF[718]
  PIN Data_PMOS_NOSF[714]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3874.425 1046.435 3874.705 1047.435 ;
    END
  END Data_PMOS_NOSF[714]
  PIN MASKH[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3834.105 1046.435 3834.385 1047.435 ;
    END
  END MASKH[34]
  PIN DIG_MON_PMOS_NOSF[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3832.425 1046.435 3832.705 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[68]
  PIN DIG_MON_SEL[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3830.745 1046.435 3831.025 1047.435 ;
    END
  END DIG_MON_SEL[68]
  PIN MASKV[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3826.265 1046.435 3826.545 1047.435 ;
    END
  END MASKV[67]
  PIN Data_PMOS_NOSF[705]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3824.585 1046.435 3824.865 1047.435 ;
    END
  END Data_PMOS_NOSF[705]
  PIN Data_PMOS_NOSF[706]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3822.905 1046.435 3823.185 1047.435 ;
    END
  END Data_PMOS_NOSF[706]
  PIN Data_PMOS_NOSF[699]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3812.265 1046.435 3812.545 1047.435 ;
    END
  END Data_PMOS_NOSF[699]
  PIN nTOK_PMOS_NOSF[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3810.025 1046.435 3810.305 1047.435 ;
    END
  END nTOK_PMOS_NOSF[33]
  PIN BcidMtx[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3807.785 1046.435 3808.065 1047.435 ;
    END
  END BcidMtx[201]
  PIN BcidMtx[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3805.545 1046.435 3805.825 1047.435 ;
    END
  END BcidMtx[199]
  PIN MASKD[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18883.545 1046.435 18883.825 1047.435 ;
    END
  END MASKD[443]
  PIN Data_PMOS_NOSF[696]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3800.785 1046.435 3801.065 1047.435 ;
    END
  END Data_PMOS_NOSF[696]
  PIN Data_PMOS_NOSF[703]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3798.545 1046.435 3798.825 1047.435 ;
    END
  END Data_PMOS_NOSF[703]
  PIN Data_PMOS_NOSF[709]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3771.945 1046.435 3772.225 1047.435 ;
    END
  END Data_PMOS_NOSF[709]
  PIN Data_PMOS_NOSF[693]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3770.265 1046.435 3770.545 1047.435 ;
    END
  END Data_PMOS_NOSF[693]
  PIN MASKD[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3768.025 1046.435 3768.305 1047.435 ;
    END
  END MASKD[66]
  PIN MASKD[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3763.545 1046.435 3763.825 1047.435 ;
    END
  END MASKD[65]
  PIN Data_PMOS_NOSF[690]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3760.185 1046.435 3760.465 1047.435 ;
    END
  END Data_PMOS_NOSF[690]
  PIN Data_PMOS_NOSF[691]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3745.625 1046.435 3745.905 1047.435 ;
    END
  END Data_PMOS_NOSF[691]
  PIN Data_PMOS_NOSF[692]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3743.945 1046.435 3744.225 1047.435 ;
    END
  END Data_PMOS_NOSF[692]
  PIN BcidMtx[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1498.345 1046.435 1498.625 1047.435 ;
    END
  END BcidMtx[28]
  PIN FREEZE_PMOS_NOSF[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1497.225 1046.435 1497.505 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[4]
  PIN BcidMtx[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1494.985 1046.435 1495.265 1047.435 ;
    END
  END BcidMtx[24]
  PIN Data_PMOS_NOSF[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1453.545 1046.435 1453.825 1047.435 ;
    END
  END Data_PMOS_NOSF[86]
  PIN Data_PMOS_NOSF[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1452.425 1046.435 1452.705 1047.435 ;
    END
  END Data_PMOS_NOSF[99]
  PIN Data_PMOS_NOSF[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1450.185 1046.435 1450.465 1047.435 ;
    END
  END Data_PMOS_NOSF[95]
  PIN Data_PMOS_NOSF[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1449.065 1046.435 1449.345 1047.435 ;
    END
  END Data_PMOS_NOSF[84]
  PIN MASKH[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1447.385 1046.435 1447.665 1047.435 ;
    END
  END MASKH[4]
  PIN MASKD[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1442.345 1046.435 1442.625 1047.435 ;
    END
  END MASKD[7]
  PIN INJ_ROW[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1431.705 1046.435 1431.985 1047.435 ;
    END
  END INJ_ROW[3]
  PIN Data_PMOS_NOSF[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1429.465 1046.435 1429.745 1047.435 ;
    END
  END Data_PMOS_NOSF[75]
  PIN Data_PMOS_NOSF[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1427.785 1046.435 1428.065 1047.435 ;
    END
  END Data_PMOS_NOSF[76]
  PIN Data_PMOS_NOSF[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1426.665 1046.435 1426.945 1047.435 ;
    END
  END Data_PMOS_NOSF[77]
  PIN BcidMtx[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1310.185 1046.435 1310.465 1047.435 ;
    END
  END BcidMtx[14]
  PIN BcidMtx[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1419.665 1046.435 1419.945 1047.435 ;
    END
  END BcidMtx[22]
  PIN Read_PMOS_NOSF[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1392.505 1046.435 1392.785 1047.435 ;
    END
  END Read_PMOS_NOSF[3]
  PIN INJ_IN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1389.705 1046.435 1389.985 1047.435 ;
    END
  END INJ_IN[6]
  PIN Data_PMOS_NOSF[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1386.905 1046.435 1387.185 1047.435 ;
    END
  END Data_PMOS_NOSF[78]
  PIN Data_PMOS_NOSF[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1385.785 1046.435 1386.065 1047.435 ;
    END
  END Data_PMOS_NOSF[67]
  PIN Data_PMOS_NOSF[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1384.105 1046.435 1384.385 1047.435 ;
    END
  END Data_PMOS_NOSF[64]
  PIN MASKH[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1381.865 1046.435 1382.145 1047.435 ;
    END
  END MASKH[3]
  PIN Data_HV[1135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18890.825 1046.435 18891.105 1047.435 ;
    END
  END Data_HV[1135]
  PIN DIG_MON_SEL[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1365.625 1046.435 1365.905 1047.435 ;
    END
  END DIG_MON_SEL[6]
  PIN INJ_ROW[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1361.705 1046.435 1361.985 1047.435 ;
    END
  END INJ_ROW[2]
  PIN Data_PMOS_NOSF[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1360.585 1046.435 1360.865 1047.435 ;
    END
  END Data_PMOS_NOSF[60]
  PIN Data_PMOS_NOSF[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1358.905 1046.435 1359.185 1047.435 ;
    END
  END Data_PMOS_NOSF[61]
  PIN Data_PMOS_NOSF[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1356.665 1046.435 1356.945 1047.435 ;
    END
  END Data_PMOS_NOSF[56]
  PIN Data_PMOS_NOSF[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1355.545 1046.435 1355.825 1047.435 ;
    END
  END Data_PMOS_NOSF[48]
  PIN BcidMtx[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1312.985 1046.435 1313.265 1047.435 ;
    END
  END BcidMtx[17]
  PIN BcidMtx[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1309.625 1046.435 1309.905 1047.435 ;
    END
  END BcidMtx[13]
  PIN Data_PMOS_NOSF[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1306.825 1046.435 1307.105 1047.435 ;
    END
  END Data_PMOS_NOSF[45]
  PIN Data_PMOS_NOSF[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1305.145 1046.435 1305.425 1047.435 ;
    END
  END Data_PMOS_NOSF[57]
  PIN Data_PMOS_NOSF[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1303.465 1046.435 1303.745 1047.435 ;
    END
  END Data_PMOS_NOSF[58]
  PIN Data_PMOS_NOSF[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1301.785 1046.435 1302.065 1047.435 ;
    END
  END Data_PMOS_NOSF[42]
  PIN MASKH[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1291.705 1046.435 1291.985 1047.435 ;
    END
  END MASKH[2]
  PIN DIG_MON_PMOS_NOSF[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1290.025 1046.435 1290.305 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[4]
  PIN DIG_MON_SEL[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1287.785 1046.435 1288.065 1047.435 ;
    END
  END DIG_MON_SEL[3]
  PIN INJ_ROW[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1282.465 1046.435 1282.745 1047.435 ;
    END
  END INJ_ROW[1]
  PIN Data_PMOS_NOSF[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1280.785 1046.435 1281.065 1047.435 ;
    END
  END Data_PMOS_NOSF[29]
  PIN Data_PMOS_NOSF[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1279.105 1046.435 1279.385 1047.435 ;
    END
  END Data_PMOS_NOSF[26]
  PIN Data_PMOS_NOSF[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1251.945 1046.435 1252.225 1047.435 ;
    END
  END Data_PMOS_NOSF[35]
  PIN nTOK_PMOS_NOSF[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1248.585 1046.435 1248.865 1047.435 ;
    END
  END nTOK_PMOS_NOSF[1]
  PIN BcidMtx[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1246.345 1046.435 1246.625 1047.435 ;
    END
  END BcidMtx[9]
  PIN Read_PMOS_NOSF[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1245.225 1046.435 1245.505 1047.435 ;
    END
  END Read_PMOS_NOSF[1]
  PIN BcidMtx[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1243.545 1046.435 1243.825 1047.435 ;
    END
  END BcidMtx[6]
  PIN Data_PMOS_NOSF[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1241.305 1046.435 1241.585 1047.435 ;
    END
  END Data_PMOS_NOSF[24]
  PIN Data_PMOS_NOSF[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1226.745 1046.435 1227.025 1047.435 ;
    END
  END Data_PMOS_NOSF[36]
  PIN Data_PMOS_NOSF[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1224.505 1046.435 1224.785 1047.435 ;
    END
  END Data_PMOS_NOSF[32]
  PIN Data_PMOS_NOSF[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1223.385 1046.435 1223.665 1047.435 ;
    END
  END Data_PMOS_NOSF[21]
  PIN MASKH[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1221.705 1046.435 1221.985 1047.435 ;
    END
  END MASKH[1]
  PIN DIG_MON_SEL[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1217.785 1046.435 1218.065 1047.435 ;
    END
  END DIG_MON_SEL[1]
  PIN INJ_ROW[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1214.425 1046.435 1214.705 1047.435 ;
    END
  END INJ_ROW[0]
  PIN Data_PMOS_NOSF[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1172.425 1046.435 1172.705 1047.435 ;
    END
  END Data_PMOS_NOSF[12]
  PIN Data_PMOS_NOSF[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1171.305 1046.435 1171.585 1047.435 ;
    END
  END Data_PMOS_NOSF[5]
  PIN Data_PMOS_NOSF[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1169.625 1046.435 1169.905 1047.435 ;
    END
  END Data_PMOS_NOSF[14]
  PIN nTOK_PMOS_NOSF[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1166.265 1046.435 1166.545 1047.435 ;
    END
  END nTOK_PMOS_NOSF[0]
  PIN BcidMtx[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1164.585 1046.435 1164.865 1047.435 ;
    END
  END BcidMtx[4]
  PIN Read_PMOS_NOSF[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1162.905 1046.435 1163.185 1047.435 ;
    END
  END Read_PMOS_NOSF[0]
  PIN INJ_IN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1151.705 1046.435 1151.985 1047.435 ;
    END
  END INJ_IN[0]
  PIN Data_PMOS_NOSF[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1150.025 1046.435 1150.305 1047.435 ;
    END
  END Data_PMOS_NOSF[2]
  PIN Data_PMOS_NOSF[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1148.345 1046.435 1148.625 1047.435 ;
    END
  END Data_PMOS_NOSF[10]
  PIN Data_PMOS_NOSF[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1146.105 1046.435 1146.385 1047.435 ;
    END
  END Data_PMOS_NOSF[1]
  PIN Data_PMOS_NOSF[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1144.985 1046.435 1145.265 1047.435 ;
    END
  END Data_PMOS_NOSF[17]
  PIN MASKV[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1142.465 1046.435 1142.745 1047.435 ;
    END
  END MASKV[0]
  PIN FREEZE_PMOS_NOSF[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1393.065 1046.435 1393.345 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[3]
  PIN MASKD[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2230.825 1046.435 2231.105 1047.435 ;
    END
  END MASKD[27]
  PIN Data_PMOS_NOSF[291]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2227.465 1046.435 2227.745 1047.435 ;
    END
  END Data_PMOS_NOSF[291]
  PIN Data_PMOS_NOSF[285]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2226.345 1046.435 2226.625 1047.435 ;
    END
  END Data_PMOS_NOSF[285]
  PIN Data_PMOS_NOSF[286]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2224.665 1046.435 2224.945 1047.435 ;
    END
  END Data_PMOS_NOSF[286]
  PIN Data_PMOS_NOSF[279]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2222.425 1046.435 2222.705 1047.435 ;
    END
  END Data_PMOS_NOSF[279]
  PIN nTOK_PMOS_NOSF[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2220.185 1046.435 2220.465 1047.435 ;
    END
  END nTOK_PMOS_NOSF[13]
  PIN BcidMtx[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2204.505 1046.435 2204.785 1047.435 ;
    END
  END BcidMtx[81]
  PIN BcidMtx[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2202.265 1046.435 2202.545 1047.435 ;
    END
  END BcidMtx[79]
  PIN INJ_IN[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2200.585 1046.435 2200.865 1047.435 ;
    END
  END INJ_IN[26]
  PIN Data_PMOS_NOSF[282]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2198.345 1046.435 2198.625 1047.435 ;
    END
  END Data_PMOS_NOSF[282]
  PIN Data_PMOS_NOSF[289]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2196.105 1046.435 2196.385 1047.435 ;
    END
  END Data_PMOS_NOSF[289]
  PIN Data_PMOS_NOSF[274]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2194.985 1046.435 2195.265 1047.435 ;
    END
  END Data_PMOS_NOSF[274]
  PIN MASKV[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2154.665 1046.435 2154.945 1047.435 ;
    END
  END MASKV[26]
  PIN DIG_MON_PMOS_NOSF[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2152.425 1046.435 2152.705 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[26]
  PIN DIG_MON_SEL[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2150.745 1046.435 2151.025 1047.435 ;
    END
  END DIG_MON_SEL[26]
  PIN MASKD[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2149.065 1046.435 2149.345 1047.435 ;
    END
  END MASKD[25]
  PIN MASKV[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2146.265 1046.435 2146.545 1047.435 ;
    END
  END MASKV[25]
  PIN Data_PMOS_NOSF[260]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2145.145 1046.435 2145.425 1047.435 ;
    END
  END Data_PMOS_NOSF[260]
  PIN Data_PMOS_NOSF[265]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2142.905 1046.435 2143.185 1047.435 ;
    END
  END Data_PMOS_NOSF[265]
  PIN Data_PMOS_NOSF[259]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2141.225 1046.435 2141.505 1047.435 ;
    END
  END Data_PMOS_NOSF[259]
  PIN nTOK_PMOS_NOSF[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2130.025 1046.435 2130.305 1047.435 ;
    END
  END nTOK_PMOS_NOSF[12]
  PIN BcidMtx[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2127.785 1046.435 2128.065 1047.435 ;
    END
  END BcidMtx[75]
  PIN BcidMtx[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2126.105 1046.435 2126.385 1047.435 ;
    END
  END BcidMtx[74]
  PIN INJ_IN[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2121.905 1046.435 2122.185 1047.435 ;
    END
  END INJ_IN[24]
  PIN Data_PMOS_NOSF[254]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2120.225 1046.435 2120.505 1047.435 ;
    END
  END Data_PMOS_NOSF[254]
  PIN Data_PMOS_NOSF[256]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2092.505 1046.435 2092.785 1047.435 ;
    END
  END Data_PMOS_NOSF[256]
  PIN Data_PMOS_NOSF[268]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2091.945 1046.435 2092.225 1047.435 ;
    END
  END Data_PMOS_NOSF[268]
  PIN Data_PMOS_NOSF[269]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2089.705 1046.435 2089.985 1047.435 ;
    END
  END Data_PMOS_NOSF[269]
  PIN DIG_MON_PMOS_NOSF[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2086.905 1046.435 2087.185 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[24]
  PIN DIG_MON_SEL[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2085.225 1046.435 2085.505 1047.435 ;
    END
  END DIG_MON_SEL[24]
  PIN DIG_MON_PMOS_NOSF[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2082.425 1046.435 2082.705 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[23]
  PIN Data_PMOS_NOSF[239]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2079.625 1046.435 2079.905 1047.435 ;
    END
  END Data_PMOS_NOSF[239]
  PIN Data_PMOS_NOSF[250]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2065.625 1046.435 2065.905 1047.435 ;
    END
  END Data_PMOS_NOSF[250]
  PIN Data_PMOS_NOSF[251]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2063.945 1046.435 2064.225 1047.435 ;
    END
  END Data_PMOS_NOSF[251]
  PIN DIG_MON_SEL[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17605.065 1046.435 17605.345 1047.435 ;
    END
  END DIG_MON_SEL[411]
  PIN BcidMtx[1314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18669.065 1046.435 18669.345 1047.435 ;
    END
  END BcidMtx[1314]
  PIN Data_HV[785]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17600.025 1046.435 17600.305 1047.435 ;
    END
  END Data_HV[785]
  PIN Data_HV[789]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17599.465 1046.435 17599.745 1047.435 ;
    END
  END Data_HV[789]
  PIN Data_HV[790]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17597.785 1046.435 17598.065 1047.435 ;
    END
  END Data_HV[790]
  PIN Data_HV[783]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17595.545 1046.435 17595.825 1047.435 ;
    END
  END Data_HV[783]
  PIN nTOK_HV[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17554.105 1046.435 17554.385 1047.435 ;
    END
  END nTOK_HV[37]
  PIN BcidMtx[1233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17551.865 1046.435 17552.145 1047.435 ;
    END
  END BcidMtx[1233]
  PIN BcidMtx[1230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17549.065 1046.435 17549.345 1047.435 ;
    END
  END BcidMtx[1230]
  PIN INJ_IN[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17547.945 1046.435 17548.225 1047.435 ;
    END
  END INJ_IN[410]
  PIN Data_HV[786]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17545.705 1046.435 17545.985 1047.435 ;
    END
  END Data_HV[786]
  PIN Data_HV[788]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17542.905 1046.435 17543.185 1047.435 ;
    END
  END Data_HV[788]
  PIN Data_HV[778]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17542.345 1046.435 17542.625 1047.435 ;
    END
  END Data_HV[778]
  PIN MASKV[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17532.265 1046.435 17532.545 1047.435 ;
    END
  END MASKV[410]
  PIN DIG_MON_SEL[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17528.345 1046.435 17528.625 1047.435 ;
    END
  END DIG_MON_SEL[410]
  PIN DIG_MON_SEL[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17527.785 1046.435 17528.065 1047.435 ;
    END
  END DIG_MON_SEL[409]
  PIN INJ_ROW[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17522.465 1046.435 17522.745 1047.435 ;
    END
  END INJ_ROW[204]
  PIN Data_HV[775]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17519.665 1046.435 17519.945 1047.435 ;
    END
  END Data_HV[775]
  PIN Data_HV[761]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17519.105 1046.435 17519.385 1047.435 ;
    END
  END Data_HV[761]
  PIN Data_HV[770]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17491.945 1046.435 17492.225 1047.435 ;
    END
  END Data_HV[770]
  PIN BcidMtx[1229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17487.465 1046.435 17487.745 1047.435 ;
    END
  END BcidMtx[1229]
  PIN BcidMtx[1228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17486.905 1046.435 17487.185 1047.435 ;
    END
  END BcidMtx[1228]
  PIN Read_HV[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17485.225 1046.435 17485.505 1047.435 ;
    END
  END Read_HV[36]
  PIN Data_HV[759]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17481.305 1046.435 17481.585 1047.435 ;
    END
  END Data_HV[759]
  PIN Data_HV[758]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17480.745 1046.435 17481.025 1047.435 ;
    END
  END Data_HV[758]
  PIN Data_HV[766]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17466.185 1046.435 17466.465 1047.435 ;
    END
  END Data_HV[766]
  PIN Data_HV[756]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17463.385 1046.435 17463.665 1047.435 ;
    END
  END Data_HV[756]
  PIN Data_HV[773]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17462.825 1046.435 17463.105 1047.435 ;
    END
  END Data_HV[773]
  PIN MASKD[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17461.145 1046.435 17461.425 1047.435 ;
    END
  END MASKD[408]
  PIN MASKD[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17456.665 1046.435 17456.945 1047.435 ;
    END
  END MASKD[407]
  PIN DIG_MON_HV[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17455.545 1046.435 17455.825 1047.435 ;
    END
  END DIG_MON_HV[71]
  PIN Data_HV[753]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17413.545 1046.435 17413.825 1047.435 ;
    END
  END Data_HV[753]
  PIN Data_HV[748]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17410.745 1046.435 17411.025 1047.435 ;
    END
  END Data_HV[748]
  PIN Data_HV[755]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17410.185 1046.435 17410.465 1047.435 ;
    END
  END Data_HV[755]
  PIN Data_HV[741]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17408.505 1046.435 17408.785 1047.435 ;
    END
  END Data_HV[741]
  PIN BcidMtx[1221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17404.025 1046.435 17404.305 1047.435 ;
    END
  END BcidMtx[1221]
  PIN FREEZE_HV[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17403.465 1046.435 17403.745 1047.435 ;
    END
  END FREEZE_HV[35]
  PIN BcidMtx[1219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17401.785 1046.435 17402.065 1047.435 ;
    END
  END BcidMtx[1219]
  PIN Data_HV[744]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17389.465 1046.435 17389.745 1047.435 ;
    END
  END Data_HV[744]
  PIN Data_HV[750]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17388.905 1046.435 17389.185 1047.435 ;
    END
  END Data_HV[750]
  PIN Data_HV[751]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17387.225 1046.435 17387.505 1047.435 ;
    END
  END Data_HV[751]
  PIN MASKV[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17382.465 1046.435 17382.745 1047.435 ;
    END
  END MASKV[406]
  PIN MASKH[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17381.905 1046.435 17382.185 1047.435 ;
    END
  END MASKH[203]
  PIN DIG_MON_HV[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18469.705 1046.435 18469.985 1047.435 ;
    END
  END DIG_MON_HV[97]
  PIN INJ_ROW[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18468.585 1046.435 18468.865 1047.435 ;
    END
  END INJ_ROW[216]
  PIN Data_HV[1016]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18466.905 1046.435 18467.185 1047.435 ;
    END
  END Data_HV[1016]
  PIN Data_HV[1013]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18465.225 1046.435 18465.505 1047.435 ;
    END
  END Data_HV[1013]
  PIN Data_HV[1022]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18463.545 1046.435 18463.825 1047.435 ;
    END
  END Data_HV[1022]
  PIN INJ_IN[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18461.305 1046.435 18461.585 1047.435 ;
    END
  END INJ_IN[433]
  PIN BcidMtx[1300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18445.065 1046.435 18445.345 1047.435 ;
    END
  END BcidMtx[1300]
  PIN Read_HV[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18443.385 1046.435 18443.665 1047.435 ;
    END
  END Read_HV[48]
  PIN BcidMtx[1296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18441.705 1046.435 18441.985 1047.435 ;
    END
  END BcidMtx[1296]
  PIN Data_HV[1010]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18438.905 1046.435 18439.185 1047.435 ;
    END
  END Data_HV[1010]
  PIN Data_HV[1018]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18437.225 1046.435 18437.505 1047.435 ;
    END
  END Data_HV[1018]
  PIN Data_HV[1019]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18435.545 1046.435 18435.825 1047.435 ;
    END
  END Data_HV[1019]
  PIN Data_HV[1025]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18433.865 1046.435 18434.145 1047.435 ;
    END
  END Data_HV[1025]
  PIN MASKD[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18393.545 1046.435 18393.825 1047.435 ;
    END
  END MASKD[432]
  PIN DIG_MON_SEL[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18390.745 1046.435 18391.025 1047.435 ;
    END
  END DIG_MON_SEL[432]
  PIN DIG_MON_HV[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18387.945 1046.435 18388.225 1047.435 ;
    END
  END DIG_MON_HV[95]
  PIN Data_HV[1005]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18385.705 1046.435 18385.985 1047.435 ;
    END
  END Data_HV[1005]
  PIN Data_HV[1006]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18384.025 1046.435 18384.305 1047.435 ;
    END
  END Data_HV[1006]
  PIN Data_HV[1007]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18382.345 1046.435 18382.625 1047.435 ;
    END
  END Data_HV[1007]
  PIN Data_HV[993]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18372.265 1046.435 18372.545 1047.435 ;
    END
  END Data_HV[993]
  PIN BcidMtx[1295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18368.905 1046.435 18369.185 1047.435 ;
    END
  END BcidMtx[1295]
  PIN FREEZE_HV[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18367.225 1046.435 18367.505 1047.435 ;
    END
  END FREEZE_HV[47]
  PIN BcidMtx[1291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18365.545 1046.435 18365.825 1047.435 ;
    END
  END BcidMtx[1291]
  PIN Data_HV[990]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18360.785 1046.435 18361.065 1047.435 ;
    END
  END Data_HV[990]
  PIN Data_HV[1002]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18359.105 1046.435 18359.385 1047.435 ;
    END
  END Data_HV[1002]
  PIN Data_HV[1003]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18331.945 1046.435 18332.225 1047.435 ;
    END
  END Data_HV[1003]
  PIN Data_HV[987]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18330.265 1046.435 18330.545 1047.435 ;
    END
  END Data_HV[987]
  PIN MASKH[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18328.585 1046.435 18328.865 1047.435 ;
    END
  END MASKH[215]
  PIN MASKD[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18323.545 1046.435 18323.825 1047.435 ;
    END
  END MASKD[429]
  PIN MASKV[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18320.745 1046.435 18321.025 1047.435 ;
    END
  END MASKV[429]
  PIN Data_HV[985]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18305.625 1046.435 18305.905 1047.435 ;
    END
  END Data_HV[985]
  PIN Data_HV[979]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18304.505 1046.435 18304.785 1047.435 ;
    END
  END Data_HV[979]
  PIN Data_HV[973]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18302.825 1046.435 18303.105 1047.435 ;
    END
  END Data_HV[973]
  PIN BcidMtx[1289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18298.905 1046.435 18299.185 1047.435 ;
    END
  END BcidMtx[1289]
  PIN FREEZE_HV[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18297.225 1046.435 18297.505 1047.435 ;
    END
  END FREEZE_HV[46]
  PIN BcidMtx[1285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18295.545 1046.435 18295.825 1047.435 ;
    END
  END BcidMtx[1285]
  PIN INJ_IN[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18293.865 1046.435 18294.145 1047.435 ;
    END
  END INJ_IN[428]
  PIN Data_HV[981]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18252.425 1046.435 18252.705 1047.435 ;
    END
  END Data_HV[981]
  PIN Data_HV[982]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18250.745 1046.435 18251.025 1047.435 ;
    END
  END Data_HV[982]
  PIN Data_HV[967]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18249.625 1046.435 18249.905 1047.435 ;
    END
  END Data_HV[967]
  PIN INJ_IN[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18667.945 1046.435 18668.225 1047.435 ;
    END
  END INJ_IN[438]
  PIN Data_HV[1074]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18666.825 1046.435 18667.105 1047.435 ;
    END
  END Data_HV[1074]
  PIN DIG_MON_HV[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18241.225 1046.435 18241.505 1047.435 ;
    END
  END DIG_MON_HV[91]
  PIN Data_HV[963]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18230.585 1046.435 18230.865 1047.435 ;
    END
  END Data_HV[963]
  PIN Data_HV[957]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18229.465 1046.435 18229.745 1047.435 ;
    END
  END Data_HV[957]
  PIN Data_HV[965]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18227.225 1046.435 18227.505 1047.435 ;
    END
  END Data_HV[965]
  PIN Data_HV[951]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18225.545 1046.435 18225.825 1047.435 ;
    END
  END Data_HV[951]
  PIN nTOK_HV[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18221.345 1046.435 18221.625 1047.435 ;
    END
  END nTOK_HV[45]
  PIN Read_HV[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18192.505 1046.435 18192.785 1047.435 ;
    END
  END Read_HV[45]
  PIN BcidMtx[1278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18190.825 1046.435 18191.105 1047.435 ;
    END
  END BcidMtx[1278]
  PIN Data_HV[948]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18188.585 1046.435 18188.865 1047.435 ;
    END
  END Data_HV[948]
  PIN Data_HV[954]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18187.465 1046.435 18187.745 1047.435 ;
    END
  END Data_HV[954]
  PIN Data_HV[949]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18185.785 1046.435 18186.065 1047.435 ;
    END
  END Data_HV[949]
  PIN Data_HV[946]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18184.105 1046.435 18184.385 1047.435 ;
    END
  END Data_HV[946]
  PIN Data_HV[962]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18182.985 1046.435 18183.265 1047.435 ;
    END
  END Data_HV[962]
  PIN MASKH[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18181.865 1046.435 18182.145 1047.435 ;
    END
  END MASKH[213]
  PIN DIG_MON_SEL[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18165.625 1046.435 18165.905 1047.435 ;
    END
  END DIG_MON_SEL[426]
  PIN DIG_MON_HV[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18162.825 1046.435 18163.105 1047.435 ;
    END
  END DIG_MON_HV[89]
  PIN Data_HV[942]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18160.585 1046.435 18160.865 1047.435 ;
    END
  END Data_HV[942]
  PIN Data_HV[929]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18158.345 1046.435 18158.625 1047.435 ;
    END
  END Data_HV[929]
  PIN Data_HV[944]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18157.225 1046.435 18157.505 1047.435 ;
    END
  END Data_HV[944]
  PIN Data_HV[930]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18155.545 1046.435 18155.825 1047.435 ;
    END
  END Data_HV[930]
  PIN BcidMtx[1276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18112.425 1046.435 18112.705 1047.435 ;
    END
  END BcidMtx[1276]
  PIN FREEZE_HV[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18111.305 1046.435 18111.585 1047.435 ;
    END
  END FREEZE_HV[44]
  PIN BcidMtx[1273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18109.625 1046.435 18109.905 1047.435 ;
    END
  END BcidMtx[1273]
  PIN Data_HV[926]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18106.265 1046.435 18106.545 1047.435 ;
    END
  END Data_HV[926]
  PIN Data_HV[939]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18105.145 1046.435 18105.425 1047.435 ;
    END
  END Data_HV[939]
  PIN Data_HV[940]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18103.465 1046.435 18103.745 1047.435 ;
    END
  END Data_HV[940]
  PIN Data_HV[941]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18101.225 1046.435 18101.505 1047.435 ;
    END
  END Data_HV[941]
  PIN MASKH[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18091.705 1046.435 18091.985 1047.435 ;
    END
  END MASKH[212]
  PIN DIG_MON_HV[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18090.025 1046.435 18090.305 1047.435 ;
    END
  END DIG_MON_HV[88]
  PIN MASKD[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18086.665 1046.435 18086.945 1047.435 ;
    END
  END MASKD[423]
  PIN Data_HV[921]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18081.345 1046.435 18081.625 1047.435 ;
    END
  END Data_HV[921]
  PIN Data_HV[922]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18079.665 1046.435 18079.945 1047.435 ;
    END
  END Data_HV[922]
  PIN Data_HV[916]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18053.065 1046.435 18053.345 1047.435 ;
    END
  END Data_HV[916]
  PIN Data_HV[917]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18051.945 1046.435 18052.225 1047.435 ;
    END
  END Data_HV[917]
  PIN BcidMtx[1271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18047.465 1046.435 18047.745 1047.435 ;
    END
  END BcidMtx[1271]
  PIN BcidMtx[1269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18046.345 1046.435 18046.625 1047.435 ;
    END
  END BcidMtx[1269]
  PIN Read_HV[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18045.225 1046.435 18045.505 1047.435 ;
    END
  END Read_HV[43]
  PIN BcidMtx[1266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18043.545 1046.435 18043.825 1047.435 ;
    END
  END BcidMtx[1266]
  PIN Data_HV[905]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18040.745 1046.435 18041.025 1047.435 ;
    END
  END Data_HV[905]
  PIN Data_HV[913]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18026.185 1046.435 18026.465 1047.435 ;
    END
  END Data_HV[913]
  PIN Data_HV[914]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18024.505 1046.435 18024.785 1047.435 ;
    END
  END Data_HV[914]
  PIN Data_HV[920]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18022.825 1046.435 18023.105 1047.435 ;
    END
  END Data_HV[920]
  PIN MASKD[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18021.145 1046.435 18021.425 1047.435 ;
    END
  END MASKD[422]
  PIN DIG_MON_SEL[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18018.345 1046.435 18018.625 1047.435 ;
    END
  END DIG_MON_SEL[422]
  PIN MASKD[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18016.665 1046.435 18016.945 1047.435 ;
    END
  END MASKD[421]
  PIN MASKV[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18013.865 1046.435 18014.145 1047.435 ;
    END
  END MASKV[421]
  PIN Data_HV[894]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17972.425 1046.435 17972.705 1047.435 ;
    END
  END Data_HV[894]
  PIN Data_HV[895]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17970.745 1046.435 17971.025 1047.435 ;
    END
  END Data_HV[895]
  PIN Data_HV[889]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17969.065 1046.435 17969.345 1047.435 ;
    END
  END Data_HV[889]
  PIN nTOK_HV[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17966.265 1046.435 17966.545 1047.435 ;
    END
  END nTOK_HV[42]
  PIN BcidMtx[1263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17964.025 1046.435 17964.305 1047.435 ;
    END
  END BcidMtx[1263]
  PIN BcidMtx[1261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17961.785 1046.435 17962.065 1047.435 ;
    END
  END BcidMtx[1261]
  PIN INJ_IN[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17951.705 1046.435 17951.985 1047.435 ;
    END
  END INJ_IN[420]
  PIN Data_HV[891]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17949.465 1046.435 17949.745 1047.435 ;
    END
  END Data_HV[891]
  PIN Data_HV[898]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17947.225 1046.435 17947.505 1047.435 ;
    END
  END Data_HV[898]
  PIN Data_HV[882]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17945.545 1046.435 17945.825 1047.435 ;
    END
  END Data_HV[882]
  PIN MASKV[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17942.465 1046.435 17942.745 1047.435 ;
    END
  END MASKV[420]
  PIN DIG_MON_SEL[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 19031.945 1046.435 19032.225 1047.435 ;
    END
  END DIG_MON_SEL[447]
  PIN DIG_MON_HV[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 19029.705 1046.435 19029.985 1047.435 ;
    END
  END DIG_MON_HV[111]
  PIN Data_HV[1163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 19026.905 1046.435 19027.185 1047.435 ;
    END
  END Data_HV[1163]
  PIN Data_HV[1160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 19025.225 1046.435 19025.505 1047.435 ;
    END
  END Data_HV[1160]
  PIN Data_HV[1175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 19024.105 1046.435 19024.385 1047.435 ;
    END
  END Data_HV[1175]
  PIN INJ_IN[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 19021.305 1046.435 19021.585 1047.435 ;
    END
  END INJ_IN[447]
  PIN BcidMtx[1342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 19005.065 1046.435 19005.345 1047.435 ;
    END
  END BcidMtx[1342]
  PIN FREEZE_HV[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 19003.945 1046.435 19004.225 1047.435 ;
    END
  END FREEZE_HV[55]
  PIN INJ_IN[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 19000.585 1046.435 19000.865 1047.435 ;
    END
  END INJ_IN[446]
  PIN Data_HV[1164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18998.345 1046.435 18998.625 1047.435 ;
    END
  END Data_HV[1164]
  PIN Data_HV[1170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18997.785 1046.435 18998.065 1047.435 ;
    END
  END Data_HV[1170]
  PIN Data_HV[1156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18994.985 1046.435 18995.265 1047.435 ;
    END
  END Data_HV[1156]
  PIN Data_HV[1172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18993.865 1046.435 18994.145 1047.435 ;
    END
  END Data_HV[1172]
  PIN MASKD[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18953.545 1046.435 18953.825 1047.435 ;
    END
  END MASKD[446]
  PIN DIG_MON_SEL[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18950.185 1046.435 18950.465 1047.435 ;
    END
  END DIG_MON_SEL[445]
  PIN INJ_ROW[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18946.825 1046.435 18947.105 1047.435 ;
    END
  END INJ_ROW[222]
  PIN Data_HV[1152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18945.705 1046.435 18945.985 1047.435 ;
    END
  END Data_HV[1152]
  PIN Data_HV[1139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18943.465 1046.435 18943.745 1047.435 ;
    END
  END Data_HV[1139]
  PIN Data_HV[1154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18942.345 1046.435 18942.625 1047.435 ;
    END
  END Data_HV[1154]
  PIN Data_HV[1140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18932.265 1046.435 18932.545 1047.435 ;
    END
  END Data_HV[1140]
  PIN BcidMtx[1335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18927.785 1046.435 18928.065 1047.435 ;
    END
  END BcidMtx[1335]
  PIN FREEZE_HV[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18927.225 1046.435 18927.505 1047.435 ;
    END
  END FREEZE_HV[54]
  PIN BcidMtx[1333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18925.545 1046.435 18925.825 1047.435 ;
    END
  END BcidMtx[1333]
  PIN DIG_MON_SEL[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1671.945 1046.435 1672.225 1047.435 ;
    END
  END DIG_MON_SEL[13]
  PIN MASKV[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1668.025 1046.435 1668.305 1047.435 ;
    END
  END MASKV[13]
  PIN Data_PMOS_NOSF[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1666.345 1046.435 1666.625 1047.435 ;
    END
  END Data_PMOS_NOSF[138]
  PIN Data_PMOS_NOSF[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1665.225 1046.435 1665.505 1047.435 ;
    END
  END Data_PMOS_NOSF[131]
  PIN Data_PMOS_NOSF[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1662.985 1046.435 1663.265 1047.435 ;
    END
  END Data_PMOS_NOSF[133]
  PIN nTOK_PMOS_NOSF[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1660.185 1046.435 1660.465 1047.435 ;
    END
  END nTOK_PMOS_NOSF[6]
  PIN BcidMtx[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1645.065 1046.435 1645.345 1047.435 ;
    END
  END BcidMtx[40]
  PIN BcidMtx[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1642.825 1046.435 1643.105 1047.435 ;
    END
  END BcidMtx[38]
  PIN INJ_IN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1640.585 1046.435 1640.865 1047.435 ;
    END
  END INJ_IN[12]
  PIN Data_PMOS_NOSF[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1638.905 1046.435 1639.185 1047.435 ;
    END
  END Data_PMOS_NOSF[128]
  PIN Data_PMOS_NOSF[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1636.665 1046.435 1636.945 1047.435 ;
    END
  END Data_PMOS_NOSF[130]
  PIN Data_PMOS_NOSF[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1634.985 1046.435 1635.265 1047.435 ;
    END
  END Data_PMOS_NOSF[127]
  PIN Data_PMOS_NOSF[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1633.865 1046.435 1634.145 1047.435 ;
    END
  END Data_PMOS_NOSF[143]
  PIN DIG_MON_PMOS_NOSF[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1592.425 1046.435 1592.705 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[12]
  PIN DIG_MON_SEL[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1590.745 1046.435 1591.025 1047.435 ;
    END
  END DIG_MON_SEL[12]
  PIN MASKD[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1589.065 1046.435 1589.345 1047.435 ;
    END
  END MASKD[11]
  PIN Data_PMOS_NOSF[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1585.705 1046.435 1585.985 1047.435 ;
    END
  END Data_PMOS_NOSF[123]
  PIN Data_PMOS_NOSF[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1584.025 1046.435 1584.305 1047.435 ;
    END
  END Data_PMOS_NOSF[124]
  PIN Data_PMOS_NOSF[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1582.905 1046.435 1583.185 1047.435 ;
    END
  END Data_PMOS_NOSF[118]
  PIN Data_PMOS_NOSF[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1572.265 1046.435 1572.545 1047.435 ;
    END
  END Data_PMOS_NOSF[111]
  PIN BcidMtx[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1568.905 1046.435 1569.185 1047.435 ;
    END
  END BcidMtx[35]
  PIN BcidMtx[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1567.785 1046.435 1568.065 1047.435 ;
    END
  END BcidMtx[33]
  PIN BcidMtx[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1565.545 1046.435 1565.825 1047.435 ;
    END
  END BcidMtx[31]
  PIN Data_PMOS_NOSF[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1560.785 1046.435 1561.065 1047.435 ;
    END
  END Data_PMOS_NOSF[108]
  PIN Data_PMOS_NOSF[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1559.665 1046.435 1559.945 1047.435 ;
    END
  END Data_PMOS_NOSF[114]
  PIN Data_PMOS_NOSF[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1531.945 1046.435 1532.225 1047.435 ;
    END
  END Data_PMOS_NOSF[121]
  PIN Data_PMOS_NOSF[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1530.265 1046.435 1530.545 1047.435 ;
    END
  END Data_PMOS_NOSF[105]
  PIN MASKV[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1529.145 1046.435 1529.425 1047.435 ;
    END
  END MASKV[10]
  PIN Data_HV[1151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18889.705 1046.435 18889.985 1047.435 ;
    END
  END Data_HV[1151]
  PIN DIG_MON_SEL[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1524.665 1046.435 1524.945 1047.435 ;
    END
  END DIG_MON_SEL[9]
  PIN DIG_MON_PMOS_NOSF[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1522.425 1046.435 1522.705 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[9]
  PIN Data_PMOS_NOSF[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1519.625 1046.435 1519.905 1047.435 ;
    END
  END Data_PMOS_NOSF[92]
  PIN Data_PMOS_NOSF[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1505.065 1046.435 1505.345 1047.435 ;
    END
  END Data_PMOS_NOSF[89]
  PIN Data_PMOS_NOSF[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1503.945 1046.435 1504.225 1047.435 ;
    END
  END Data_PMOS_NOSF[104]
  PIN INJ_IN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1501.145 1046.435 1501.425 1047.435 ;
    END
  END INJ_IN[9]
  PIN DIG_MON_SEL[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15925.625 1046.435 15925.905 1047.435 ;
    END
  END DIG_MON_SEL[370]
  PIN DIG_MON_HV[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15922.825 1046.435 15923.105 1047.435 ;
    END
  END DIG_MON_HV[33]
  PIN Data_HV[354]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15920.585 1046.435 15920.865 1047.435 ;
    END
  END Data_HV[354]
  PIN Data_HV[355]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15918.905 1046.435 15919.185 1047.435 ;
    END
  END Data_HV[355]
  PIN Data_HV[356]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15917.225 1046.435 15917.505 1047.435 ;
    END
  END Data_HV[356]
  PIN Data_HV[342]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15915.545 1046.435 15915.825 1047.435 ;
    END
  END Data_HV[342]
  PIN nTOK_HV[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15874.105 1046.435 15874.385 1047.435 ;
    END
  END nTOK_HV[16]
  PIN BcidMtx[1107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15871.865 1046.435 15872.145 1047.435 ;
    END
  END BcidMtx[1107]
  PIN Data_HV[1091]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18717.225 1046.435 18717.505 1047.435 ;
    END
  END Data_HV[1091]
  PIN BcidMtx[1104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15869.065 1046.435 15869.345 1047.435 ;
    END
  END BcidMtx[1104]
  PIN Data_HV[338]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15866.265 1046.435 15866.545 1047.435 ;
    END
  END Data_HV[338]
  PIN Data_HV[346]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15864.585 1046.435 15864.865 1047.435 ;
    END
  END Data_HV[346]
  PIN Data_HV[347]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15862.905 1046.435 15863.185 1047.435 ;
    END
  END Data_HV[347]
  PIN Data_HV[353]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15861.225 1046.435 15861.505 1047.435 ;
    END
  END Data_HV[353]
  PIN MASKH[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15851.705 1046.435 15851.985 1047.435 ;
    END
  END MASKH[184]
  PIN DIG_MON_SEL[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15848.345 1046.435 15848.625 1047.435 ;
    END
  END DIG_MON_SEL[368]
  PIN DIG_MON_HV[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15845.545 1046.435 15845.825 1047.435 ;
    END
  END DIG_MON_HV[31]
  PIN Data_HV[333]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15841.345 1046.435 15841.625 1047.435 ;
    END
  END Data_HV[333]
  PIN Data_HV[334]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15839.665 1046.435 15839.945 1047.435 ;
    END
  END Data_HV[334]
  PIN Data_HV[335]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15812.505 1046.435 15812.785 1047.435 ;
    END
  END Data_HV[335]
  PIN Data_HV[321]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15810.825 1046.435 15811.105 1047.435 ;
    END
  END Data_HV[321]
  PIN BcidMtx[1103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15807.465 1046.435 15807.745 1047.435 ;
    END
  END BcidMtx[1103]
  PIN BcidMtx[1101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15806.345 1046.435 15806.625 1047.435 ;
    END
  END BcidMtx[1101]
  PIN BcidMtx[1100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15804.665 1046.435 15804.945 1047.435 ;
    END
  END BcidMtx[1100]
  PIN INJ_IN[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15802.425 1046.435 15802.705 1047.435 ;
    END
  END INJ_IN[366]
  PIN Data_HV[324]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15800.185 1046.435 15800.465 1047.435 ;
    END
  END Data_HV[324]
  PIN Data_HV[319]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15785.625 1046.435 15785.905 1047.435 ;
    END
  END Data_HV[319]
  PIN Data_HV[316]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15783.945 1046.435 15784.225 1047.435 ;
    END
  END Data_HV[316]
  PIN MASKV[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15782.265 1046.435 15782.545 1047.435 ;
    END
  END MASKV[366]
  PIN DIG_MON_HV[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15780.025 1046.435 15780.305 1047.435 ;
    END
  END DIG_MON_HV[30]
  PIN DIG_MON_SEL[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15777.785 1046.435 15778.065 1047.435 ;
    END
  END DIG_MON_SEL[365]
  PIN INJ_ROW[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15774.425 1046.435 15774.705 1047.435 ;
    END
  END INJ_ROW[182]
  PIN Data_HV[302]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15732.985 1046.435 15733.265 1047.435 ;
    END
  END Data_HV[302]
  PIN Data_HV[299]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15731.305 1046.435 15731.585 1047.435 ;
    END
  END Data_HV[299]
  PIN Data_HV[308]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15729.625 1046.435 15729.905 1047.435 ;
    END
  END Data_HV[308]
  PIN INJ_IN[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15727.385 1046.435 15727.665 1047.435 ;
    END
  END INJ_IN[365]
  PIN BcidMtx[1096]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15724.585 1046.435 15724.865 1047.435 ;
    END
  END BcidMtx[1096]
  PIN Read_HV[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15722.905 1046.435 15723.185 1047.435 ;
    END
  END Read_HV[14]
  PIN BcidMtx[1093]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15721.785 1046.435 15722.065 1047.435 ;
    END
  END BcidMtx[1093]
  PIN Data_HV[297]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15710.585 1046.435 15710.865 1047.435 ;
    END
  END Data_HV[297]
  PIN Data_HV[298]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15707.785 1046.435 15708.065 1047.435 ;
    END
  END Data_HV[298]
  PIN Data_HV[305]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15706.665 1046.435 15706.945 1047.435 ;
    END
  END Data_HV[305]
  PIN Data_HV[294]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15705.545 1046.435 15705.825 1047.435 ;
    END
  END Data_HV[294]
  PIN DIG_MON_HV[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15700.225 1046.435 15700.505 1047.435 ;
    END
  END DIG_MON_HV[28]
  PIN DIG_MON_SEL[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15698.545 1046.435 15698.825 1047.435 ;
    END
  END DIG_MON_SEL[364]
  PIN DIG_MON_SEL[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16791.945 1046.435 16792.225 1047.435 ;
    END
  END DIG_MON_SEL[391]
  PIN Data_HV[585]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16787.465 1046.435 16787.745 1047.435 ;
    END
  END Data_HV[585]
  PIN Data_HV[579]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16786.345 1046.435 16786.625 1047.435 ;
    END
  END Data_HV[579]
  PIN Data_HV[572]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16785.225 1046.435 16785.505 1047.435 ;
    END
  END Data_HV[572]
  PIN Data_HV[573]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16782.425 1046.435 16782.705 1047.435 ;
    END
  END Data_HV[573]
  PIN nTOK_HV[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16780.185 1046.435 16780.465 1047.435 ;
    END
  END nTOK_HV[27]
  PIN BcidMtx[1174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16765.065 1046.435 16765.345 1047.435 ;
    END
  END BcidMtx[1174]
  PIN BcidMtx[1170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16761.705 1046.435 16761.985 1047.435 ;
    END
  END BcidMtx[1170]
  PIN Data_HV[570]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16759.465 1046.435 16759.745 1047.435 ;
    END
  END Data_HV[570]
  PIN Data_HV[582]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16757.785 1046.435 16758.065 1047.435 ;
    END
  END Data_HV[582]
  PIN Data_HV[578]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16755.545 1046.435 16755.825 1047.435 ;
    END
  END Data_HV[578]
  PIN Data_HV[567]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16754.425 1046.435 16754.705 1047.435 ;
    END
  END Data_HV[567]
  PIN MASKH[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16714.105 1046.435 16714.385 1047.435 ;
    END
  END MASKH[195]
  PIN DIG_MON_SEL[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16710.745 1046.435 16711.025 1047.435 ;
    END
  END DIG_MON_SEL[390]
  PIN MASKD[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16709.065 1046.435 16709.345 1047.435 ;
    END
  END MASKD[389]
  PIN MASKV[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16706.265 1046.435 16706.545 1047.435 ;
    END
  END MASKV[389]
  PIN Data_HV[565]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16704.025 1046.435 16704.305 1047.435 ;
    END
  END Data_HV[565]
  PIN Data_HV[559]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16702.905 1046.435 16703.185 1047.435 ;
    END
  END Data_HV[559]
  PIN Data_HV[553]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16701.225 1046.435 16701.505 1047.435 ;
    END
  END Data_HV[553]
  PIN BcidMtx[1169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16688.905 1046.435 16689.185 1047.435 ;
    END
  END BcidMtx[1169]
  PIN BcidMtx[1167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16687.785 1046.435 16688.065 1047.435 ;
    END
  END BcidMtx[1167]
  PIN BcidMtx[1166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16686.105 1046.435 16686.385 1047.435 ;
    END
  END BcidMtx[1166]
  PIN INJ_IN[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16681.905 1046.435 16682.185 1047.435 ;
    END
  END INJ_IN[388]
  PIN Data_HV[548]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16680.225 1046.435 16680.505 1047.435 ;
    END
  END Data_HV[548]
  PIN Data_HV[561]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16679.105 1046.435 16679.385 1047.435 ;
    END
  END Data_HV[561]
  PIN Data_HV[546]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16650.265 1046.435 16650.545 1047.435 ;
    END
  END Data_HV[546]
  PIN MASKV[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16649.145 1046.435 16649.425 1047.435 ;
    END
  END MASKV[388]
  PIN DIG_MON_HV[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16646.905 1046.435 16647.185 1047.435 ;
    END
  END DIG_MON_HV[52]
  PIN MASKD[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16643.545 1046.435 16643.825 1047.435 ;
    END
  END MASKD[387]
  PIN Data_HV[537]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16626.185 1046.435 16626.465 1047.435 ;
    END
  END Data_HV[537]
  PIN Data_HV[530]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16625.065 1046.435 16625.345 1047.435 ;
    END
  END Data_HV[530]
  PIN Data_HV[545]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16623.945 1046.435 16624.225 1047.435 ;
    END
  END Data_HV[545]
  PIN INJ_IN[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16621.145 1046.435 16621.425 1047.435 ;
    END
  END INJ_IN[387]
  PIN BcidMtx[1163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16618.905 1046.435 16619.185 1047.435 ;
    END
  END BcidMtx[1163]
  PIN BcidMtx[1161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16617.785 1046.435 16618.065 1047.435 ;
    END
  END BcidMtx[1161]
  PIN BcidMtx[1158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16614.985 1046.435 16615.265 1047.435 ;
    END
  END BcidMtx[1158]
  PIN Data_HV[528]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16574.105 1046.435 16574.385 1047.435 ;
    END
  END Data_HV[528]
  PIN Data_HV[534]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16572.985 1046.435 16573.265 1047.435 ;
    END
  END Data_HV[534]
  PIN Data_HV[536]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16570.185 1046.435 16570.465 1047.435 ;
    END
  END Data_HV[536]
  PIN Data_HV[525]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16569.065 1046.435 16569.345 1047.435 ;
    END
  END Data_HV[525]
  PIN MASKV[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16567.945 1046.435 16568.225 1047.435 ;
    END
  END MASKV[386]
  PIN DIG_MON_SEL[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16564.025 1046.435 16564.305 1047.435 ;
    END
  END DIG_MON_SEL[386]
  PIN MASKD[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16562.345 1046.435 16562.625 1047.435 ;
    END
  END MASKD[385]
  PIN INJ_ROW[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16551.705 1046.435 16551.985 1047.435 ;
    END
  END INJ_ROW[192]
  PIN Data_HV[523]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16548.905 1046.435 16549.185 1047.435 ;
    END
  END Data_HV[523]
  PIN Data_HV[1078]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18716.105 1046.435 18716.385 1047.435 ;
    END
  END Data_HV[1078]
  PIN Data_HV[524]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16547.225 1046.435 16547.505 1047.435 ;
    END
  END Data_HV[524]
  PIN INJ_IN[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16542.465 1046.435 16542.745 1047.435 ;
    END
  END INJ_IN[385]
  PIN BcidMtx[1157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16540.225 1046.435 16540.505 1047.435 ;
    END
  END BcidMtx[1157]
  PIN BcidMtx[1155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16539.105 1046.435 16539.385 1047.435 ;
    END
  END BcidMtx[1155]
  PIN INJ_IN[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16509.705 1046.435 16509.985 1047.435 ;
    END
  END INJ_IN[384]
  PIN Data_HV[506]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16508.025 1046.435 16508.305 1047.435 ;
    END
  END Data_HV[506]
  PIN Data_HV[519]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16506.905 1046.435 16507.185 1047.435 ;
    END
  END Data_HV[519]
  PIN Data_HV[505]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16504.105 1046.435 16504.385 1047.435 ;
    END
  END Data_HV[505]
  PIN Data_HV[521]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16502.985 1046.435 16503.265 1047.435 ;
    END
  END Data_HV[521]
  PIN MASKH[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16501.865 1046.435 16502.145 1047.435 ;
    END
  END MASKH[192]
  PIN DIG_MON_SEL[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16485.065 1046.435 16485.345 1047.435 ;
    END
  END DIG_MON_SEL[383]
  PIN INJ_ROW[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17041.705 1046.435 17041.985 1047.435 ;
    END
  END INJ_ROW[198]
  PIN Data_HV[638]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17040.025 1046.435 17040.305 1047.435 ;
    END
  END Data_HV[638]
  PIN BcidMtx[1318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18672.425 1046.435 18672.705 1047.435 ;
    END
  END BcidMtx[1318]
  PIN Data_HV[650]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17037.225 1046.435 17037.505 1047.435 ;
    END
  END Data_HV[650]
  PIN Data_HV[636]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17035.545 1046.435 17035.825 1047.435 ;
    END
  END Data_HV[636]
  PIN BcidMtx[1191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16991.865 1046.435 16992.145 1047.435 ;
    END
  END BcidMtx[1191]
  PIN FREEZE_HV[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16991.305 1046.435 16991.585 1047.435 ;
    END
  END FREEZE_HV[30]
  PIN BcidMtx[1189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16989.625 1046.435 16989.905 1047.435 ;
    END
  END BcidMtx[1189]
  PIN Data_HV[639]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16985.705 1046.435 16985.985 1047.435 ;
    END
  END Data_HV[639]
  PIN Data_HV[645]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16985.145 1046.435 16985.425 1047.435 ;
    END
  END Data_HV[645]
  PIN Data_HV[646]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16983.465 1046.435 16983.745 1047.435 ;
    END
  END Data_HV[646]
  PIN MASKV[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16972.265 1046.435 16972.545 1047.435 ;
    END
  END MASKV[396]
  PIN MASKH[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16971.705 1046.435 16971.985 1047.435 ;
    END
  END MASKH[198]
  PIN INJ_ROW[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16962.465 1046.435 16962.745 1047.435 ;
    END
  END INJ_ROW[197]
  PIN MASKV[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16961.905 1046.435 16962.185 1047.435 ;
    END
  END MASKV[395]
  PIN BcidMtx[1317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18671.865 1046.435 18672.145 1047.435 ;
    END
  END BcidMtx[1317]
  PIN Data_HV[629]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16932.505 1046.435 16932.785 1047.435 ;
    END
  END Data_HV[629]
  PIN Data_HV[623]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16931.945 1046.435 16932.225 1047.435 ;
    END
  END Data_HV[623]
  PIN INJ_IN[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16929.705 1046.435 16929.985 1047.435 ;
    END
  END INJ_IN[395]
  PIN FREEZE_HV[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16925.785 1046.435 16926.065 1047.435 ;
    END
  END FREEZE_HV[29]
  PIN Read_HV[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16925.225 1046.435 16925.505 1047.435 ;
    END
  END Read_HV[29]
  PIN BcidMtx[1182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16923.545 1046.435 16923.825 1047.435 ;
    END
  END BcidMtx[1182]
  PIN Data_HV[624]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16906.745 1046.435 16907.025 1047.435 ;
    END
  END Data_HV[624]
  PIN Data_HV[619]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16906.185 1046.435 16906.465 1047.435 ;
    END
  END Data_HV[619]
  PIN Data_HV[620]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16904.505 1046.435 16904.785 1047.435 ;
    END
  END Data_HV[620]
  PIN MASKH[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16901.705 1046.435 16901.985 1047.435 ;
    END
  END MASKH[197]
  PIN MASKD[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16901.145 1046.435 16901.425 1047.435 ;
    END
  END MASKD[394]
  PIN DIG_MON_SEL[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16898.345 1046.435 16898.625 1047.435 ;
    END
  END DIG_MON_SEL[394]
  PIN MASKV[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16893.865 1046.435 16894.145 1047.435 ;
    END
  END MASKV[393]
  PIN Data_HV[606]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16853.545 1046.435 16853.825 1047.435 ;
    END
  END Data_HV[606]
  PIN Data_HV[607]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16851.865 1046.435 16852.145 1047.435 ;
    END
  END Data_HV[607]
  PIN FREEZE_HV[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18671.305 1046.435 18671.585 1047.435 ;
    END
  END FREEZE_HV[51]
  PIN Data_HV[602]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16849.625 1046.435 16849.905 1047.435 ;
    END
  END Data_HV[602]
  PIN Data_HV[595]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16849.065 1046.435 16849.345 1047.435 ;
    END
  END Data_HV[595]
  PIN nTOK_HV[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16846.265 1046.435 16846.545 1047.435 ;
    END
  END nTOK_HV[28]
  PIN Read_HV[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16842.905 1046.435 16843.185 1047.435 ;
    END
  END Read_HV[28]
  PIN BcidMtx[1178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16842.345 1046.435 16842.625 1047.435 ;
    END
  END BcidMtx[1178]
  PIN INJ_IN[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16831.705 1046.435 16831.985 1047.435 ;
    END
  END INJ_IN[392]
  PIN Data_HV[598]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16828.345 1046.435 16828.625 1047.435 ;
    END
  END Data_HV[598]
  PIN Data_HV[592]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16827.785 1046.435 16828.065 1047.435 ;
    END
  END Data_HV[592]
  PIN Data_HV[589]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16826.105 1046.435 16826.385 1047.435 ;
    END
  END Data_HV[589]
  PIN MASKD[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16821.345 1046.435 16821.625 1047.435 ;
    END
  END MASKD[392]
  PIN DIG_MON_HV[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16820.225 1046.435 16820.505 1047.435 ;
    END
  END DIG_MON_HV[56]
  PIN FREEZE_HV[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17073.065 1046.435 17073.345 1047.435 ;
    END
  END FREEZE_HV[31]
  PIN MASKV[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17908.025 1046.435 17908.305 1047.435 ;
    END
  END MASKV[419]
  PIN Data_HV[879]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17907.465 1046.435 17907.745 1047.435 ;
    END
  END Data_HV[879]
  PIN Data_HV[880]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17905.785 1046.435 17906.065 1047.435 ;
    END
  END Data_HV[880]
  PIN Data_HV[868]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17902.985 1046.435 17903.265 1047.435 ;
    END
  END Data_HV[868]
  PIN nTOK_HV[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17900.185 1046.435 17900.465 1047.435 ;
    END
  END nTOK_HV[41]
  PIN Read_HV[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17883.385 1046.435 17883.665 1047.435 ;
    END
  END Read_HV[41]
  PIN BcidMtx[1256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17882.825 1046.435 17883.105 1047.435 ;
    END
  END BcidMtx[1256]
  PIN INJ_IN[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17880.585 1046.435 17880.865 1047.435 ;
    END
  END INJ_IN[418]
  PIN Data_HV[871]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17877.225 1046.435 17877.505 1047.435 ;
    END
  END Data_HV[871]
  PIN Data_HV[865]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17876.665 1046.435 17876.945 1047.435 ;
    END
  END Data_HV[865]
  PIN Data_HV[862]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17874.985 1046.435 17875.265 1047.435 ;
    END
  END Data_HV[862]
  PIN MASKD[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17833.545 1046.435 17833.825 1047.435 ;
    END
  END MASKD[418]
  PIN DIG_MON_HV[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17832.425 1046.435 17832.705 1047.435 ;
    END
  END DIG_MON_HV[82]
  PIN DIG_MON_SEL[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17830.185 1046.435 17830.465 1047.435 ;
    END
  END DIG_MON_SEL[417]
  PIN Data_HV[858]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17825.705 1046.435 17825.985 1047.435 ;
    END
  END Data_HV[858]
  PIN Data_HV[848]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17825.145 1046.435 17825.425 1047.435 ;
    END
  END Data_HV[848]
  PIN Data_HV[845]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17823.465 1046.435 17823.745 1047.435 ;
    END
  END Data_HV[845]
  PIN Data_HV[846]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17812.265 1046.435 17812.545 1047.435 ;
    END
  END Data_HV[846]
  PIN INJ_IN[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17811.145 1046.435 17811.425 1047.435 ;
    END
  END INJ_IN[417]
  PIN BcidMtx[1252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17808.345 1046.435 17808.625 1047.435 ;
    END
  END BcidMtx[1252]
  PIN BcidMtx[1249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17805.545 1046.435 17805.825 1047.435 ;
    END
  END BcidMtx[1249]
  PIN BcidMtx[1248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17804.985 1046.435 17805.265 1047.435 ;
    END
  END BcidMtx[1248]
  PIN Data_HV[842]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17800.225 1046.435 17800.505 1047.435 ;
    END
  END Data_HV[842]
  PIN Data_HV[856]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17771.945 1046.435 17772.225 1047.435 ;
    END
  END Data_HV[856]
  PIN Data_HV[851]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17771.385 1046.435 17771.665 1047.435 ;
    END
  END Data_HV[851]
  PIN Data_HV[857]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17769.705 1046.435 17769.985 1047.435 ;
    END
  END Data_HV[857]
  PIN DIG_MON_SEL[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17765.225 1046.435 17765.505 1047.435 ;
    END
  END DIG_MON_SEL[416]
  PIN MASKD[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17763.545 1046.435 17763.825 1047.435 ;
    END
  END MASKD[415]
  PIN Data_HV[827]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17759.625 1046.435 17759.905 1047.435 ;
    END
  END Data_HV[827]
  PIN Data_HV[831]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17746.185 1046.435 17746.465 1047.435 ;
    END
  END Data_HV[831]
  PIN Data_HV[832]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17744.505 1046.435 17744.785 1047.435 ;
    END
  END Data_HV[832]
  PIN INJ_IN[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17741.145 1046.435 17741.425 1047.435 ;
    END
  END INJ_IN[415]
  PIN nTOK_HV[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17740.025 1046.435 17740.305 1047.435 ;
    END
  END nTOK_HV[39]
  PIN BcidMtx[1245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17737.785 1046.435 17738.065 1047.435 ;
    END
  END BcidMtx[1245]
  PIN BcidMtx[1242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17734.985 1046.435 17735.265 1047.435 ;
    END
  END BcidMtx[1242]
  PIN INJ_IN[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17733.865 1046.435 17734.145 1047.435 ;
    END
  END INJ_IN[414]
  PIN Data_HV[828]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17692.985 1046.435 17693.265 1047.435 ;
    END
  END Data_HV[828]
  PIN Data_HV[830]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17690.185 1046.435 17690.465 1047.435 ;
    END
  END Data_HV[830]
  PIN Data_HV[820]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17689.625 1046.435 17689.905 1047.435 ;
    END
  END Data_HV[820]
  PIN MASKV[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17687.945 1046.435 17688.225 1047.435 ;
    END
  END MASKV[414]
  PIN Read_HV[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18670.745 1046.435 18671.025 1047.435 ;
    END
  END Read_HV[51]
  PIN DIG_MON_SEL[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17684.025 1046.435 17684.305 1047.435 ;
    END
  END DIG_MON_SEL[414]
  PIN MASKD[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17682.345 1046.435 17682.625 1047.435 ;
    END
  END MASKD[413]
  PIN Data_HV[806]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17670.025 1046.435 17670.305 1047.435 ;
    END
  END Data_HV[806]
  PIN Data_HV[810]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17669.465 1046.435 17669.745 1047.435 ;
    END
  END Data_HV[810]
  PIN Data_HV[811]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17667.785 1046.435 17668.065 1047.435 ;
    END
  END Data_HV[811]
  PIN INJ_IN[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17662.465 1046.435 17662.745 1047.435 ;
    END
  END INJ_IN[413]
  PIN nTOK_HV[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17661.345 1046.435 17661.625 1047.435 ;
    END
  END nTOK_HV[38]
  PIN BcidMtx[1239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17659.105 1046.435 17659.385 1047.435 ;
    END
  END BcidMtx[1239]
  PIN INJ_IN[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17629.705 1046.435 17629.985 1047.435 ;
    END
  END INJ_IN[412]
  PIN Data_HV[801]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17628.585 1046.435 17628.865 1047.435 ;
    END
  END Data_HV[801]
  PIN Data_HV[813]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17626.905 1046.435 17627.185 1047.435 ;
    END
  END Data_HV[813]
  PIN Data_HV[799]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17624.105 1046.435 17624.385 1047.435 ;
    END
  END Data_HV[799]
  PIN Data_HV[798]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17623.545 1046.435 17623.825 1047.435 ;
    END
  END Data_HV[798]
  PIN MASKH[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17621.865 1046.435 17622.145 1047.435 ;
    END
  END MASKH[206]
  PIN BcidMtx[1316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18670.185 1046.435 18670.465 1047.435 ;
    END
  END BcidMtx[1316]
  PIN DIG_MON_HV[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16482.825 1046.435 16483.105 1047.435 ;
    END
  END DIG_MON_HV[47]
  PIN MASKV[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16481.145 1046.435 16481.425 1047.435 ;
    END
  END MASKV[383]
  PIN Data_HV[488]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16478.345 1046.435 16478.625 1047.435 ;
    END
  END Data_HV[488]
  PIN Data_HV[503]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16477.225 1046.435 16477.505 1047.435 ;
    END
  END Data_HV[503]
  PIN Data_HV[490]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16476.105 1046.435 16476.385 1047.435 ;
    END
  END Data_HV[490]
  PIN BcidMtx[1151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16432.985 1046.435 16433.265 1047.435 ;
    END
  END BcidMtx[1151]
  PIN BcidMtx[1149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16431.865 1046.435 16432.145 1047.435 ;
    END
  END BcidMtx[1149]
  PIN Read_HV[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16430.745 1046.435 16431.025 1047.435 ;
    END
  END Read_HV[23]
  PIN Data_HV[486]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16426.825 1046.435 16427.105 1047.435 ;
    END
  END Data_HV[486]
  PIN Data_HV[492]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16425.705 1046.435 16425.985 1047.435 ;
    END
  END Data_HV[492]
  PIN Data_HV[493]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16424.585 1046.435 16424.865 1047.435 ;
    END
  END Data_HV[493]
  PIN Data_HV[483]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16421.785 1046.435 16422.065 1047.435 ;
    END
  END Data_HV[483]
  PIN MASKV[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16412.265 1046.435 16412.545 1047.435 ;
    END
  END MASKV[382]
  PIN MASKD[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16411.145 1046.435 16411.425 1047.435 ;
    END
  END MASKD[382]
  PIN MASKD[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16406.665 1046.435 16406.945 1047.435 ;
    END
  END MASKD[381]
  PIN INJ_ROW[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16402.465 1046.435 16402.745 1047.435 ;
    END
  END INJ_ROW[190]
  PIN Data_HV[480]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16401.345 1046.435 16401.625 1047.435 ;
    END
  END Data_HV[480]
  PIN Data_HV[475]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16373.065 1046.435 16373.345 1047.435 ;
    END
  END Data_HV[475]
  PIN Data_HV[476]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16371.945 1046.435 16372.225 1047.435 ;
    END
  END Data_HV[476]
  PIN Data_HV[468]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16370.825 1046.435 16371.105 1047.435 ;
    END
  END Data_HV[468]
  PIN BcidMtx[1143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16366.345 1046.435 16366.625 1047.435 ;
    END
  END BcidMtx[1143]
  PIN Read_HV[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16365.225 1046.435 16365.505 1047.435 ;
    END
  END Read_HV[22]
  PIN BcidMtx[1141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16364.105 1046.435 16364.385 1047.435 ;
    END
  END BcidMtx[1141]
  PIN Data_HV[471]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16360.185 1046.435 16360.465 1047.435 ;
    END
  END Data_HV[471]
  PIN Data_HV[472]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16346.185 1046.435 16346.465 1047.435 ;
    END
  END Data_HV[472]
  PIN Data_HV[478]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16345.065 1046.435 16345.345 1047.435 ;
    END
  END Data_HV[478]
  PIN Data_HV[479]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16342.825 1046.435 16343.105 1047.435 ;
    END
  END Data_HV[479]
  PIN MASKH[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16341.705 1046.435 16341.985 1047.435 ;
    END
  END MASKH[190]
  PIN DIG_MON_HV[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16335.545 1046.435 16335.825 1047.435 ;
    END
  END DIG_MON_HV[43]
  PIN MASKV[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16333.865 1046.435 16334.145 1047.435 ;
    END
  END MASKV[379]
  PIN Data_HV[453]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16292.425 1046.435 16292.705 1047.435 ;
    END
  END Data_HV[453]
  PIN Data_HV[455]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16289.625 1046.435 16289.905 1047.435 ;
    END
  END Data_HV[455]
  PIN Data_HV[447]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16288.505 1046.435 16288.785 1047.435 ;
    END
  END Data_HV[447]
  PIN nTOK_HV[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16286.265 1046.435 16286.545 1047.435 ;
    END
  END nTOK_HV[21]
  PIN FREEZE_HV[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16283.465 1046.435 16283.745 1047.435 ;
    END
  END FREEZE_HV[21]
  PIN BcidMtx[1136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16282.345 1046.435 16282.625 1047.435 ;
    END
  END BcidMtx[1136]
  PIN INJ_IN[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16271.705 1046.435 16271.985 1047.435 ;
    END
  END INJ_IN[378]
  PIN Data_HV[456]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16268.905 1046.435 16269.185 1047.435 ;
    END
  END Data_HV[456]
  PIN Data_HV[445]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16267.785 1046.435 16268.065 1047.435 ;
    END
  END Data_HV[445]
  PIN Data_HV[442]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16266.105 1046.435 16266.385 1047.435 ;
    END
  END Data_HV[442]
  PIN MASKH[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16261.905 1046.435 16262.185 1047.435 ;
    END
  END MASKH[189]
  PIN MASKD[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16261.345 1046.435 16261.625 1047.435 ;
    END
  END MASKD[378]
  PIN DIG_MON_SEL[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16258.545 1046.435 16258.825 1047.435 ;
    END
  END DIG_MON_SEL[378]
  PIN INJ_ROW[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17348.585 1046.435 17348.865 1047.435 ;
    END
  END INJ_ROW[202]
  PIN MASKV[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17348.025 1046.435 17348.305 1047.435 ;
    END
  END MASKV[405]
  PIN Data_HV[726]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17346.345 1046.435 17346.625 1047.435 ;
    END
  END Data_HV[726]
  PIN Data_HV[728]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17343.545 1046.435 17343.825 1047.435 ;
    END
  END Data_HV[728]
  PIN Data_HV[721]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17342.985 1046.435 17343.265 1047.435 ;
    END
  END Data_HV[721]
  PIN nTOK_HV[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17340.185 1046.435 17340.465 1047.435 ;
    END
  END nTOK_HV[34]
  PIN Read_HV[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17323.385 1046.435 17323.665 1047.435 ;
    END
  END Read_HV[34]
  PIN BcidMtx[1214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17322.825 1046.435 17323.105 1047.435 ;
    END
  END BcidMtx[1214]
  PIN INJ_IN[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17320.585 1046.435 17320.865 1047.435 ;
    END
  END INJ_IN[404]
  PIN Data_HV[724]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17317.225 1046.435 17317.505 1047.435 ;
    END
  END Data_HV[724]
  PIN Data_HV[718]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17316.665 1046.435 17316.945 1047.435 ;
    END
  END Data_HV[718]
  PIN Data_HV[715]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17314.985 1046.435 17315.265 1047.435 ;
    END
  END Data_HV[715]
  PIN MASKD[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17273.545 1046.435 17273.825 1047.435 ;
    END
  END MASKD[404]
  PIN MASKD[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17269.065 1046.435 17269.345 1047.435 ;
    END
  END MASKD[403]
  PIN Data_HV[711]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17265.705 1046.435 17265.985 1047.435 ;
    END
  END Data_HV[711]
  PIN Data_HV[705]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17264.585 1046.435 17264.865 1047.435 ;
    END
  END Data_HV[705]
  PIN Data_HV[706]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17262.905 1046.435 17263.185 1047.435 ;
    END
  END Data_HV[706]
  PIN INJ_IN[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17251.145 1046.435 17251.425 1047.435 ;
    END
  END INJ_IN[403]
  PIN nTOK_HV[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17250.025 1046.435 17250.305 1047.435 ;
    END
  END nTOK_HV[33]
  PIN BcidMtx[1209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17247.785 1046.435 17248.065 1047.435 ;
    END
  END BcidMtx[1209]
  PIN BcidMtx[1206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17244.985 1046.435 17245.265 1047.435 ;
    END
  END BcidMtx[1206]
  PIN INJ_IN[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17241.905 1046.435 17242.185 1047.435 ;
    END
  END INJ_IN[402]
  PIN Data_HV[702]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17239.665 1046.435 17239.945 1047.435 ;
    END
  END Data_HV[702]
  PIN Data_HV[704]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17211.385 1046.435 17211.665 1047.435 ;
    END
  END Data_HV[704]
  PIN Data_HV[694]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17210.825 1046.435 17211.105 1047.435 ;
    END
  END Data_HV[694]
  PIN MASKV[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17209.145 1046.435 17209.425 1047.435 ;
    END
  END MASKV[402]
  PIN DIG_MON_SEL[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17205.225 1046.435 17205.505 1047.435 ;
    END
  END DIG_MON_SEL[402]
  PIN DIG_MON_SEL[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17204.665 1046.435 17204.945 1047.435 ;
    END
  END DIG_MON_SEL[401]
  PIN INJ_ROW[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17201.305 1046.435 17201.585 1047.435 ;
    END
  END INJ_ROW[200]
  PIN Data_HV[684]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17186.185 1046.435 17186.465 1047.435 ;
    END
  END Data_HV[684]
  PIN Data_HV[691]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17185.625 1046.435 17185.905 1047.435 ;
    END
  END Data_HV[691]
  PIN Data_HV[692]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17183.945 1046.435 17184.225 1047.435 ;
    END
  END Data_HV[692]
  PIN nTOK_HV[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17180.025 1046.435 17180.305 1047.435 ;
    END
  END nTOK_HV[32]
  PIN BcidMtx[1205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17178.905 1046.435 17179.185 1047.435 ;
    END
  END BcidMtx[1205]
  PIN FREEZE_HV[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17177.225 1046.435 17177.505 1047.435 ;
    END
  END FREEZE_HV[32]
  PIN INJ_IN[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17173.865 1046.435 17174.145 1047.435 ;
    END
  END INJ_IN[400]
  PIN Data_HV[675]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17134.105 1046.435 17134.385 1047.435 ;
    END
  END Data_HV[675]
  PIN Data_HV[687]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17132.425 1046.435 17132.705 1047.435 ;
    END
  END Data_HV[687]
  PIN Data_HV[673]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17129.625 1046.435 17129.905 1047.435 ;
    END
  END Data_HV[673]
  PIN Data_HV[689]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17128.505 1046.435 17128.785 1047.435 ;
    END
  END Data_HV[689]
  PIN MASKH[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17127.385 1046.435 17127.665 1047.435 ;
    END
  END MASKH[200]
  PIN DIG_MON_SEL[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17123.465 1046.435 17123.745 1047.435 ;
    END
  END DIG_MON_SEL[399]
  PIN MASKD[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17122.345 1046.435 17122.625 1047.435 ;
    END
  END MASKD[399]
  PIN MASKV[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17111.145 1046.435 17111.425 1047.435 ;
    END
  END MASKV[399]
  PIN Data_HV[656]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17108.345 1046.435 17108.625 1047.435 ;
    END
  END Data_HV[656]
  PIN Data_HV[664]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17107.785 1046.435 17108.065 1047.435 ;
    END
  END Data_HV[664]
  PIN Data_HV[658]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17106.105 1046.435 17106.385 1047.435 ;
    END
  END Data_HV[658]
  PIN BcidMtx[1198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17099.665 1046.435 17099.945 1047.435 ;
    END
  END BcidMtx[1198]
  PIN BcidMtx[1197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17099.105 1046.435 17099.385 1047.435 ;
    END
  END BcidMtx[1197]
  PIN BcidMtx[1195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17071.385 1046.435 17071.665 1047.435 ;
    END
  END BcidMtx[1195]
  PIN Data_HV[660]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17067.465 1046.435 17067.745 1047.435 ;
    END
  END Data_HV[660]
  PIN Data_HV[666]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17066.905 1046.435 17067.185 1047.435 ;
    END
  END Data_HV[666]
  PIN Data_HV[667]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17065.225 1046.435 17065.505 1047.435 ;
    END
  END Data_HV[667]
  PIN MASKV[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17062.425 1046.435 17062.705 1047.435 ;
    END
  END MASKV[398]
  PIN MASKH[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17061.865 1046.435 17062.145 1047.435 ;
    END
  END MASKH[199]
  PIN BcidMtx[1319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18672.985 1046.435 18673.265 1047.435 ;
    END
  END BcidMtx[1319]
  PIN nTOK_PMOS_NOSF[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2620.025 1046.435 2620.305 1047.435 ;
    END
  END nTOK_PMOS_NOSF[18]
  PIN FREEZE_PMOS_NOSF[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2617.225 1046.435 2617.505 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[18]
  PIN BcidMtx[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2616.105 1046.435 2616.385 1047.435 ;
    END
  END BcidMtx[110]
  PIN INJ_IN[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2613.865 1046.435 2614.145 1047.435 ;
    END
  END INJ_IN[36]
  PIN Data_PMOS_NOSF[387]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2572.985 1046.435 2573.265 1047.435 ;
    END
  END Data_PMOS_NOSF[387]
  PIN Data_PMOS_NOSF[382]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2571.305 1046.435 2571.585 1047.435 ;
    END
  END Data_PMOS_NOSF[382]
  PIN Data_PMOS_NOSF[379]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2569.625 1046.435 2569.905 1047.435 ;
    END
  END Data_PMOS_NOSF[379]
  PIN MASKH[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2567.385 1046.435 2567.665 1047.435 ;
    END
  END MASKH[18]
  PIN DIG_MON_PMOS_NOSF[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2565.705 1046.435 2565.985 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[36]
  PIN DIG_MON_SEL[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2563.465 1046.435 2563.745 1047.435 ;
    END
  END DIG_MON_SEL[35]
  PIN Data_PMOS_NOSF[375]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2550.585 1046.435 2550.865 1047.435 ;
    END
  END Data_PMOS_NOSF[375]
  PIN Data_PMOS_NOSF[369]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2549.465 1046.435 2549.745 1047.435 ;
    END
  END Data_PMOS_NOSF[369]
  PIN Data_PMOS_NOSF[362]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2548.345 1046.435 2548.625 1047.435 ;
    END
  END Data_PMOS_NOSF[362]
  PIN Data_PMOS_NOSF[364]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2546.105 1046.435 2546.385 1047.435 ;
    END
  END Data_PMOS_NOSF[364]
  PIN nTOK_PMOS_NOSF[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2541.345 1046.435 2541.625 1047.435 ;
    END
  END nTOK_PMOS_NOSF[17]
  PIN BcidMtx[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2539.105 1046.435 2539.385 1047.435 ;
    END
  END BcidMtx[105]
  PIN BcidMtx[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2511.385 1046.435 2511.665 1047.435 ;
    END
  END BcidMtx[103]
  PIN Data_PMOS_NOSF[360]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2508.585 1046.435 2508.865 1047.435 ;
    END
  END Data_PMOS_NOSF[360]
  PIN Data_PMOS_NOSF[372]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2506.905 1046.435 2507.185 1047.435 ;
    END
  END Data_PMOS_NOSF[372]
  PIN Data_PMOS_NOSF[373]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2505.225 1046.435 2505.505 1047.435 ;
    END
  END Data_PMOS_NOSF[373]
  PIN Data_PMOS_NOSF[357]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2503.545 1046.435 2503.825 1047.435 ;
    END
  END Data_PMOS_NOSF[357]
  PIN MASKH[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2501.865 1046.435 2502.145 1047.435 ;
    END
  END MASKH[17]
  PIN DIG_MON_SEL[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2485.625 1046.435 2485.905 1047.435 ;
    END
  END DIG_MON_SEL[34]
  PIN MASKD[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2483.945 1046.435 2484.225 1047.435 ;
    END
  END MASKD[33]
  PIN MASKV[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2481.145 1046.435 2481.425 1047.435 ;
    END
  END MASKV[33]
  PIN Data_PMOS_NOSF[341]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2478.345 1046.435 2478.625 1047.435 ;
    END
  END Data_PMOS_NOSF[341]
  PIN Data_PMOS_NOSF[350]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2476.665 1046.435 2476.945 1047.435 ;
    END
  END Data_PMOS_NOSF[350]
  PIN Data_PMOS_NOSF[342]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2475.545 1046.435 2475.825 1047.435 ;
    END
  END Data_PMOS_NOSF[342]
  PIN BcidMtx[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2432.425 1046.435 2432.705 1047.435 ;
    END
  END BcidMtx[100]
  PIN FREEZE_PMOS_NOSF[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2431.305 1046.435 2431.585 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[16]
  PIN BcidMtx[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2429.625 1046.435 2429.905 1047.435 ;
    END
  END BcidMtx[97]
  PIN Data_PMOS_NOSF[345]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2425.705 1046.435 2425.985 1047.435 ;
    END
  END Data_PMOS_NOSF[345]
  PIN MASKV[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2333.865 1046.435 2334.145 1047.435 ;
    END
  END MASKV[29]
  PIN Data_PMOS_NOSF[340]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2424.025 1046.435 2424.305 1047.435 ;
    END
  END Data_PMOS_NOSF[340]
  PIN Data_PMOS_NOSF[353]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2421.225 1046.435 2421.505 1047.435 ;
    END
  END Data_PMOS_NOSF[353]
  PIN MASKV[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2412.265 1046.435 2412.545 1047.435 ;
    END
  END MASKV[32]
  PIN DIG_MON_PMOS_NOSF[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2410.025 1046.435 2410.305 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[32]
  PIN MASKD[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2406.665 1046.435 2406.945 1047.435 ;
    END
  END MASKD[31]
  PIN DIG_MON_PMOS_NOSF[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2405.545 1046.435 2405.825 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[31]
  PIN Data_PMOS_NOSF[333]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2401.345 1046.435 2401.625 1047.435 ;
    END
  END Data_PMOS_NOSF[333]
  PIN Data_PMOS_NOSF[334]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2399.665 1046.435 2399.945 1047.435 ;
    END
  END Data_PMOS_NOSF[334]
  PIN Data_PMOS_NOSF[335]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2372.505 1046.435 2372.785 1047.435 ;
    END
  END Data_PMOS_NOSF[335]
  PIN Data_PMOS_NOSF[329]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2371.945 1046.435 2372.225 1047.435 ;
    END
  END Data_PMOS_NOSF[329]
  PIN BcidMtx[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2366.905 1046.435 2367.185 1047.435 ;
    END
  END BcidMtx[94]
  PIN BcidMtx[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2366.345 1046.435 2366.625 1047.435 ;
    END
  END BcidMtx[93]
  PIN BcidMtx[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2364.665 1046.435 2364.945 1047.435 ;
    END
  END BcidMtx[92]
  PIN Data_PMOS_NOSF[324]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2360.185 1046.435 2360.465 1047.435 ;
    END
  END Data_PMOS_NOSF[324]
  PIN Data_PMOS_NOSF[325]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2346.185 1046.435 2346.465 1047.435 ;
    END
  END Data_PMOS_NOSF[325]
  PIN Data_PMOS_NOSF[316]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2343.945 1046.435 2344.225 1047.435 ;
    END
  END Data_PMOS_NOSF[316]
  PIN Data_PMOS_NOSF[332]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2342.825 1046.435 2343.105 1047.435 ;
    END
  END Data_PMOS_NOSF[332]
  PIN MASKD[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2341.145 1046.435 2341.425 1047.435 ;
    END
  END MASKD[30]
  PIN MASKD[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2336.665 1046.435 2336.945 1047.435 ;
    END
  END MASKD[29]
  PIN DIG_MON_PMOS_NOSF[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2335.545 1046.435 2335.825 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[29]
  PIN Data_PMOS_NOSF[302]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2292.985 1046.435 2293.265 1047.435 ;
    END
  END Data_PMOS_NOSF[302]
  PIN Data_PMOS_NOSF[314]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2290.185 1046.435 2290.465 1047.435 ;
    END
  END Data_PMOS_NOSF[314]
  PIN Data_PMOS_NOSF[308]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2289.625 1046.435 2289.905 1047.435 ;
    END
  END Data_PMOS_NOSF[308]
  PIN INJ_IN[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2287.385 1046.435 2287.665 1047.435 ;
    END
  END INJ_IN[29]
  PIN BcidMtx[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2284.025 1046.435 2284.305 1047.435 ;
    END
  END BcidMtx[87]
  PIN BcidMtx[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2282.345 1046.435 2282.625 1047.435 ;
    END
  END BcidMtx[86]
  PIN BcidMtx[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2281.225 1046.435 2281.505 1047.435 ;
    END
  END BcidMtx[84]
  PIN MASKH[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18888.585 1046.435 18888.865 1047.435 ;
    END
  END MASKH[222]
  PIN Data_PMOS_NOSF[304]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2268.345 1046.435 2268.625 1047.435 ;
    END
  END Data_PMOS_NOSF[304]
  PIN Data_PMOS_NOSF[310]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2267.225 1046.435 2267.505 1047.435 ;
    END
  END Data_PMOS_NOSF[310]
  PIN MASKV[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2262.465 1046.435 2262.745 1047.435 ;
    END
  END MASKV[28]
  PIN MASKH[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2261.905 1046.435 2262.185 1047.435 ;
    END
  END MASKH[14]
  PIN DIG_MON_SEL[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3351.945 1046.435 3352.225 1047.435 ;
    END
  END DIG_MON_SEL[55]
  PIN DIG_MON_PMOS_NOSF[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3349.705 1046.435 3349.985 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[55]
  PIN MASKV[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3348.025 1046.435 3348.305 1047.435 ;
    END
  END MASKV[55]
  PIN Data_PMOS_NOSF[572]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3345.225 1046.435 3345.505 1047.435 ;
    END
  END Data_PMOS_NOSF[572]
  PIN Data_PMOS_NOSF[581]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3343.545 1046.435 3343.825 1047.435 ;
    END
  END Data_PMOS_NOSF[581]
  PIN Data_PMOS_NOSF[574]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3342.985 1046.435 3343.265 1047.435 ;
    END
  END Data_PMOS_NOSF[574]
  PIN nTOK_PMOS_NOSF[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3340.185 1046.435 3340.465 1047.435 ;
    END
  END nTOK_PMOS_NOSF[27]
  PIN Read_PMOS_NOSF[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3323.385 1046.435 3323.665 1047.435 ;
    END
  END Read_PMOS_NOSF[27]
  PIN BcidMtx[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3322.825 1046.435 3323.105 1047.435 ;
    END
  END BcidMtx[164]
  PIN INJ_IN[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3320.585 1046.435 3320.865 1047.435 ;
    END
  END INJ_IN[54]
  PIN Data_PMOS_NOSF[582]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3317.785 1046.435 3318.065 1047.435 ;
    END
  END Data_PMOS_NOSF[582]
  PIN Data_PMOS_NOSF[577]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3317.225 1046.435 3317.505 1047.435 ;
    END
  END Data_PMOS_NOSF[577]
  PIN Data_PMOS_NOSF[578]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3315.545 1046.435 3315.825 1047.435 ;
    END
  END Data_PMOS_NOSF[578]
  PIN MASKV[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3274.665 1046.435 3274.945 1047.435 ;
    END
  END MASKV[54]
  PIN MASKD[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3273.545 1046.435 3273.825 1047.435 ;
    END
  END MASKD[54]
  PIN INJ_ROW[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3266.825 1046.435 3267.105 1047.435 ;
    END
  END INJ_ROW[26]
  PIN Data_PMOS_NOSF[564]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3265.705 1046.435 3265.985 1047.435 ;
    END
  END Data_PMOS_NOSF[564]
  PIN Data_PMOS_NOSF[558]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3264.585 1046.435 3264.865 1047.435 ;
    END
  END Data_PMOS_NOSF[558]
  PIN Data_PMOS_NOSF[560]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3261.785 1046.435 3262.065 1047.435 ;
    END
  END Data_PMOS_NOSF[560]
  PIN Data_PMOS_NOSF[552]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3252.265 1046.435 3252.545 1047.435 ;
    END
  END Data_PMOS_NOSF[552]
  PIN nTOK_PMOS_NOSF[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3250.025 1046.435 3250.305 1047.435 ;
    END
  END nTOK_PMOS_NOSF[26]
  PIN Read_PMOS_NOSF[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3246.665 1046.435 3246.945 1047.435 ;
    END
  END Read_PMOS_NOSF[26]
  PIN BcidMtx[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3244.985 1046.435 3245.265 1047.435 ;
    END
  END BcidMtx[156]
  PIN Data_PMOS_NOSF[548]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3240.225 1046.435 3240.505 1047.435 ;
    END
  END Data_PMOS_NOSF[548]
  PIN Data_PMOS_NOSF[561]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3239.105 1046.435 3239.385 1047.435 ;
    END
  END Data_PMOS_NOSF[561]
  PIN Data_PMOS_NOSF[550]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3212.505 1046.435 3212.785 1047.435 ;
    END
  END Data_PMOS_NOSF[550]
  PIN Data_PMOS_NOSF[547]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3210.825 1046.435 3211.105 1047.435 ;
    END
  END Data_PMOS_NOSF[547]
  PIN MASKD[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3208.025 1046.435 3208.305 1047.435 ;
    END
  END MASKD[52]
  PIN DIG_MON_SEL[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3204.665 1046.435 3204.945 1047.435 ;
    END
  END DIG_MON_SEL[51]
  PIN INJ_ROW[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3201.305 1046.435 3201.585 1047.435 ;
    END
  END INJ_ROW[25]
  PIN Data_PMOS_NOSF[533]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3199.625 1046.435 3199.905 1047.435 ;
    END
  END Data_PMOS_NOSF[533]
  PIN Data_PMOS_NOSF[530]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3185.065 1046.435 3185.345 1047.435 ;
    END
  END Data_PMOS_NOSF[530]
  PIN Data_PMOS_NOSF[539]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3183.385 1046.435 3183.665 1047.435 ;
    END
  END Data_PMOS_NOSF[539]
  PIN Data_PMOS_NOSF[678]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3742.265 1046.435 3742.545 1047.435 ;
    END
  END Data_PMOS_NOSF[678]
  PIN nTOK_PMOS_NOSF[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3740.025 1046.435 3740.305 1047.435 ;
    END
  END nTOK_PMOS_NOSF[32]
  PIN BcidMtx[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3737.785 1046.435 3738.065 1047.435 ;
    END
  END BcidMtx[195]
  PIN BcidMtx[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3735.545 1046.435 3735.825 1047.435 ;
    END
  END BcidMtx[193]
  PIN INJ_IN[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3733.865 1046.435 3734.145 1047.435 ;
    END
  END INJ_IN[64]
  PIN Data_PMOS_NOSF[681]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3692.985 1046.435 3693.265 1047.435 ;
    END
  END Data_PMOS_NOSF[681]
  PIN Data_PMOS_NOSF[688]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3690.745 1046.435 3691.025 1047.435 ;
    END
  END Data_PMOS_NOSF[688]
  PIN Data_PMOS_NOSF[673]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3689.625 1046.435 3689.905 1047.435 ;
    END
  END Data_PMOS_NOSF[673]
  PIN MASKV[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3687.945 1046.435 3688.225 1047.435 ;
    END
  END MASKV[64]
  PIN DIG_MON_SEL[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3683.465 1046.435 3683.745 1047.435 ;
    END
  END DIG_MON_SEL[63]
  PIN INJ_ROW[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3671.705 1046.435 3671.985 1047.435 ;
    END
  END INJ_ROW[31]
  PIN Data_PMOS_NOSF[663]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3669.465 1046.435 3669.745 1047.435 ;
    END
  END Data_PMOS_NOSF[663]
  PIN Data_PMOS_NOSF[656]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3668.345 1046.435 3668.625 1047.435 ;
    END
  END Data_PMOS_NOSF[656]
  PIN Data_PMOS_NOSF[671]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3667.225 1046.435 3667.505 1047.435 ;
    END
  END Data_PMOS_NOSF[671]
  PIN INJ_IN[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3662.465 1046.435 3662.745 1047.435 ;
    END
  END INJ_IN[63]
  PIN BcidMtx[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3660.225 1046.435 3660.505 1047.435 ;
    END
  END BcidMtx[191]
  PIN Read_PMOS_NOSF[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3632.505 1046.435 3632.785 1047.435 ;
    END
  END Read_PMOS_NOSF[31]
  PIN INJ_IN[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3629.705 1046.435 3629.985 1047.435 ;
    END
  END INJ_IN[62]
  PIN Data_PMOS_NOSF[653]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3628.025 1046.435 3628.305 1047.435 ;
    END
  END Data_PMOS_NOSF[653]
  PIN Data_PMOS_NOSF[661]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3626.345 1046.435 3626.625 1047.435 ;
    END
  END Data_PMOS_NOSF[661]
  PIN Data_PMOS_NOSF[652]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3624.105 1046.435 3624.385 1047.435 ;
    END
  END Data_PMOS_NOSF[652]
  PIN Data_PMOS_NOSF[668]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3622.985 1046.435 3623.265 1047.435 ;
    END
  END Data_PMOS_NOSF[668]
  PIN MASKH[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3621.865 1046.435 3622.145 1047.435 ;
    END
  END MASKH[31]
  PIN DIG_MON_SEL[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3605.065 1046.435 3605.345 1047.435 ;
    END
  END DIG_MON_SEL[61]
  PIN DIG_MON_PMOS_NOSF[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3602.825 1046.435 3603.105 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[61]
  PIN MASKV[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3601.145 1046.435 3601.425 1047.435 ;
    END
  END MASKV[61]
  PIN Data_PMOS_NOSF[635]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3598.345 1046.435 3598.625 1047.435 ;
    END
  END Data_PMOS_NOSF[635]
  PIN Data_PMOS_NOSF[650]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3597.225 1046.435 3597.505 1047.435 ;
    END
  END Data_PMOS_NOSF[650]
  PIN Data_PMOS_NOSF[637]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3596.105 1046.435 3596.385 1047.435 ;
    END
  END Data_PMOS_NOSF[637]
  PIN BcidMtx[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3552.425 1046.435 3552.705 1047.435 ;
    END
  END BcidMtx[184]
  PIN FREEZE_PMOS_NOSF[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3551.305 1046.435 3551.585 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[30]
  PIN BcidMtx[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3550.185 1046.435 3550.465 1047.435 ;
    END
  END BcidMtx[182]
  PIN Data_PMOS_NOSF[632]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3546.265 1046.435 3546.545 1047.435 ;
    END
  END Data_PMOS_NOSF[632]
  PIN Data_PMOS_NOSF[645]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3545.145 1046.435 3545.425 1047.435 ;
    END
  END Data_PMOS_NOSF[645]
  PIN Data_PMOS_NOSF[634]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3544.025 1046.435 3544.305 1047.435 ;
    END
  END Data_PMOS_NOSF[634]
  PIN Data_PMOS_NOSF[630]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3541.785 1046.435 3542.065 1047.435 ;
    END
  END Data_PMOS_NOSF[630]
  PIN MASKV[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3532.265 1046.435 3532.545 1047.435 ;
    END
  END MASKV[60]
  PIN DIG_MON_PMOS_NOSF[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3530.025 1046.435 3530.305 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[60]
  PIN DIG_MON_SEL[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3528.345 1046.435 3528.625 1047.435 ;
    END
  END DIG_MON_SEL[60]
  PIN DIG_MON_PMOS_NOSF[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3525.545 1046.435 3525.825 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[59]
  PIN MASKV[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3521.905 1046.435 3522.185 1047.435 ;
    END
  END MASKV[59]
  PIN Data_PMOS_NOSF[621]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3520.225 1046.435 3520.505 1047.435 ;
    END
  END Data_PMOS_NOSF[621]
  PIN Data_PMOS_NOSF[629]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3492.505 1046.435 3492.785 1047.435 ;
    END
  END Data_PMOS_NOSF[629]
  PIN Data_PMOS_NOSF[616]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3491.385 1046.435 3491.665 1047.435 ;
    END
  END Data_PMOS_NOSF[616]
  PIN DIG_MON_SEL[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18885.225 1046.435 18885.505 1047.435 ;
    END
  END DIG_MON_SEL[444]
  PIN BcidMtx[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3486.345 1046.435 3486.625 1047.435 ;
    END
  END BcidMtx[177]
  PIN Read_PMOS_NOSF[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3485.225 1046.435 3485.505 1047.435 ;
    END
  END Read_PMOS_NOSF[29]
  PIN BcidMtx[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3483.545 1046.435 3483.825 1047.435 ;
    END
  END BcidMtx[174]
  PIN Data_PMOS_NOSF[618]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3480.185 1046.435 3480.465 1047.435 ;
    END
  END Data_PMOS_NOSF[618]
  PIN Data_PMOS_NOSF[619]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3466.185 1046.435 3466.465 1047.435 ;
    END
  END Data_PMOS_NOSF[619]
  PIN Data_PMOS_NOSF[620]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3464.505 1046.435 3464.785 1047.435 ;
    END
  END Data_PMOS_NOSF[620]
  PIN MASKH[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3461.705 1046.435 3461.985 1047.435 ;
    END
  END MASKH[29]
  PIN DIG_MON_PMOS_NOSF[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3460.025 1046.435 3460.305 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[58]
  PIN DIG_MON_SEL[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3458.345 1046.435 3458.625 1047.435 ;
    END
  END DIG_MON_SEL[58]
  PIN MASKV[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3453.865 1046.435 3454.145 1047.435 ;
    END
  END MASKV[57]
  PIN Data_PMOS_NOSF[596]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3412.985 1046.435 3413.265 1047.435 ;
    END
  END Data_PMOS_NOSF[596]
  PIN Data_PMOS_NOSF[607]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3411.865 1046.435 3412.145 1047.435 ;
    END
  END Data_PMOS_NOSF[607]
  PIN Data_PMOS_NOSF[595]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3409.065 1046.435 3409.345 1047.435 ;
    END
  END Data_PMOS_NOSF[595]
  PIN INJ_IN[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3407.385 1046.435 3407.665 1047.435 ;
    END
  END INJ_IN[57]
  PIN DIG_MON_HV[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18882.425 1046.435 18882.705 1047.435 ;
    END
  END DIG_MON_HV[107]
  PIN FREEZE_PMOS_NOSF[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3403.465 1046.435 3403.745 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[28]
  PIN BcidMtx[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3402.345 1046.435 3402.625 1047.435 ;
    END
  END BcidMtx[170]
  PIN BcidMtx[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3401.225 1046.435 3401.505 1047.435 ;
    END
  END BcidMtx[168]
  PIN Data_PMOS_NOSF[603]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3388.905 1046.435 3389.185 1047.435 ;
    END
  END Data_PMOS_NOSF[603]
  PIN Data_PMOS_NOSF[592]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3387.785 1046.435 3388.065 1047.435 ;
    END
  END Data_PMOS_NOSF[592]
  PIN Data_PMOS_NOSF[599]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3386.665 1046.435 3386.945 1047.435 ;
    END
  END Data_PMOS_NOSF[599]
  PIN MASKH[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3381.905 1046.435 3382.185 1047.435 ;
    END
  END MASKH[28]
  PIN DIG_MON_PMOS_NOSF[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3380.225 1046.435 3380.505 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[56]
  PIN DIG_MON_SEL[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3378.545 1046.435 3378.825 1047.435 ;
    END
  END DIG_MON_SEL[56]
  PIN INJ_ROW[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4468.585 1046.435 4468.865 1047.435 ;
    END
  END INJ_ROW[41]
  PIN Data_PMOS_NOSF[879]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4467.465 1046.435 4467.745 1047.435 ;
    END
  END Data_PMOS_NOSF[879]
  PIN Data_PMOS_NOSF[873]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4466.345 1046.435 4466.625 1047.435 ;
    END
  END Data_PMOS_NOSF[873]
  PIN Data_PMOS_NOSF[875]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4463.545 1046.435 4463.825 1047.435 ;
    END
  END Data_PMOS_NOSF[875]
  PIN Data_PMOS_NOSF[867]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4462.425 1046.435 4462.705 1047.435 ;
    END
  END Data_PMOS_NOSF[867]
  PIN nTOK_PMOS_NOSF[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4460.185 1046.435 4460.465 1047.435 ;
    END
  END nTOK_PMOS_NOSF[41]
  PIN MASKV[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18880.745 1046.435 18881.025 1047.435 ;
    END
  END MASKV[443]
  PIN BcidMtx[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4442.825 1046.435 4443.105 1047.435 ;
    END
  END BcidMtx[248]
  PIN BcidMtx[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4441.705 1046.435 4441.985 1047.435 ;
    END
  END BcidMtx[246]
  PIN Data_PMOS_NOSF[876]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4437.785 1046.435 4438.065 1047.435 ;
    END
  END Data_PMOS_NOSF[876]
  PIN Data_PMOS_NOSF[865]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4436.665 1046.435 4436.945 1047.435 ;
    END
  END Data_PMOS_NOSF[865]
  PIN Data_PMOS_NOSF[872]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4435.545 1046.435 4435.825 1047.435 ;
    END
  END Data_PMOS_NOSF[872]
  PIN MASKH[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4394.105 1046.435 4394.385 1047.435 ;
    END
  END MASKH[41]
  PIN DIG_MON_PMOS_NOSF[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4392.425 1046.435 4392.705 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[82]
  PIN DIG_MON_SEL[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4390.745 1046.435 4391.025 1047.435 ;
    END
  END DIG_MON_SEL[82]
  PIN MASKV[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4386.265 1046.435 4386.545 1047.435 ;
    END
  END MASKV[81]
  PIN Data_PMOS_NOSF[848]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4385.145 1046.435 4385.425 1047.435 ;
    END
  END Data_PMOS_NOSF[848]
  PIN Data_PMOS_NOSF[859]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4384.025 1046.435 4384.305 1047.435 ;
    END
  END Data_PMOS_NOSF[859]
  PIN Data_PMOS_NOSF[847]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4381.225 1046.435 4381.505 1047.435 ;
    END
  END Data_PMOS_NOSF[847]
  PIN INJ_IN[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4371.145 1046.435 4371.425 1047.435 ;
    END
  END INJ_IN[81]
  PIN BcidMtx[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4368.905 1046.435 4369.185 1047.435 ;
    END
  END BcidMtx[245]
  PIN BcidMtx[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4366.105 1046.435 4366.385 1047.435 ;
    END
  END BcidMtx[242]
  PIN BcidMtx[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4364.985 1046.435 4365.265 1047.435 ;
    END
  END BcidMtx[240]
  PIN Data_PMOS_NOSF[843]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4360.785 1046.435 4361.065 1047.435 ;
    END
  END Data_PMOS_NOSF[843]
  PIN Data_PMOS_NOSF[844]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4332.505 1046.435 4332.785 1047.435 ;
    END
  END Data_PMOS_NOSF[844]
  PIN Data_PMOS_NOSF[851]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4331.385 1046.435 4331.665 1047.435 ;
    END
  END Data_PMOS_NOSF[851]
  PIN Data_PMOS_NOSF[840]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4330.265 1046.435 4330.545 1047.435 ;
    END
  END Data_PMOS_NOSF[840]
  PIN DIG_MON_PMOS_NOSF[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4326.905 1046.435 4327.185 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[80]
  PIN DIG_MON_SEL[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4325.225 1046.435 4325.505 1047.435 ;
    END
  END DIG_MON_SEL[80]
  PIN DIG_MON_PMOS_NOSF[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4322.425 1046.435 4322.705 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[79]
  PIN Data_PMOS_NOSF[827]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4319.625 1046.435 4319.905 1047.435 ;
    END
  END Data_PMOS_NOSF[827]
  PIN Data_PMOS_NOSF[838]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4305.625 1046.435 4305.905 1047.435 ;
    END
  END Data_PMOS_NOSF[838]
  PIN MASKV[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7680.745 1046.435 7681.025 1047.435 ;
    END
  END MASKV[163]
  PIN Data_PMOS[537]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7666.185 1046.435 7666.465 1047.435 ;
    END
  END Data_PMOS[537]
  PIN Data_PMOS[530]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7665.065 1046.435 7665.345 1047.435 ;
    END
  END Data_PMOS[530]
  PIN Data_PMOS[532]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7662.825 1046.435 7663.105 1047.435 ;
    END
  END Data_PMOS[532]
  PIN nTOK_PMOS[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7660.025 1046.435 7660.305 1047.435 ;
    END
  END nTOK_PMOS[25]
  PIN BcidMtx[490]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7658.345 1046.435 7658.625 1047.435 ;
    END
  END BcidMtx[490]
  PIN BcidMtx[488]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7656.105 1046.435 7656.385 1047.435 ;
    END
  END BcidMtx[488]
  PIN INJ_IN[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7653.865 1046.435 7654.145 1047.435 ;
    END
  END INJ_IN[162]
  PIN Data_PMOS[527]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7613.545 1046.435 7613.825 1047.435 ;
    END
  END Data_PMOS[527]
  PIN Data_PMOS[529]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7611.305 1046.435 7611.585 1047.435 ;
    END
  END Data_PMOS[529]
  PIN Data_PMOS[526]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7609.625 1046.435 7609.905 1047.435 ;
    END
  END Data_PMOS[526]
  PIN Data_PMOS[542]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7608.505 1046.435 7608.785 1047.435 ;
    END
  END Data_PMOS[542]
  PIN DIG_MON_PMOS[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7605.705 1046.435 7605.985 1047.435 ;
    END
  END DIG_MON_PMOS[50]
  PIN DIG_MON_SEL[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7603.465 1046.435 7603.745 1047.435 ;
    END
  END DIG_MON_SEL[161]
  PIN DIG_MON_PMOS[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7601.225 1046.435 7601.505 1047.435 ;
    END
  END DIG_MON_PMOS[49]
  PIN Data_PMOS[512]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7590.025 1046.435 7590.305 1047.435 ;
    END
  END Data_PMOS[512]
  PIN Data_PMOS[509]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7588.345 1046.435 7588.625 1047.435 ;
    END
  END Data_PMOS[509]
  PIN Data_PMOS[524]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7587.225 1046.435 7587.505 1047.435 ;
    END
  END Data_PMOS[524]
  PIN INJ_IN[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7582.465 1046.435 7582.745 1047.435 ;
    END
  END INJ_IN[161]
  PIN BcidMtx[484]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7579.665 1046.435 7579.945 1047.435 ;
    END
  END BcidMtx[484]
  PIN Read_PMOS[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7552.505 1046.435 7552.785 1047.435 ;
    END
  END Read_PMOS[24]
  PIN INJ_IN[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7549.705 1046.435 7549.985 1047.435 ;
    END
  END INJ_IN[160]
  PIN Data_PMOS[513]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7547.465 1046.435 7547.745 1047.435 ;
    END
  END Data_PMOS[513]
  PIN Data_PMOS[514]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7546.345 1046.435 7546.625 1047.435 ;
    END
  END Data_PMOS[514]
  PIN Data_PMOS[505]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7544.105 1046.435 7544.385 1047.435 ;
    END
  END Data_PMOS[505]
  PIN MASKV[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7542.425 1046.435 7542.705 1047.435 ;
    END
  END MASKV[160]
  PIN MASKD[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7541.305 1046.435 7541.585 1047.435 ;
    END
  END MASKD[160]
  PIN DIG_MON_SEL[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7525.065 1046.435 7525.345 1047.435 ;
    END
  END DIG_MON_SEL[159]
  PIN INJ_ROW[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7521.705 1046.435 7521.985 1047.435 ;
    END
  END INJ_ROW[79]
  PIN Data_PMOS[501]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7520.585 1046.435 7520.865 1047.435 ;
    END
  END Data_PMOS[501]
  PIN Data_PMOS[488]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7518.345 1046.435 7518.625 1047.435 ;
    END
  END Data_PMOS[488]
  PIN Data_PMOS[497]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7516.665 1046.435 7516.945 1047.435 ;
    END
  END Data_PMOS[497]
  PIN Data_PMOS[489]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7515.545 1046.435 7515.825 1047.435 ;
    END
  END Data_PMOS[489]
  PIN Data_HV[1075]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18664.025 1046.435 18664.305 1047.435 ;
    END
  END Data_HV[1075]
  PIN BcidMtx[478]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7472.425 1046.435 7472.705 1047.435 ;
    END
  END BcidMtx[478]
  PIN FREEZE_PMOS[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7471.305 1046.435 7471.585 1047.435 ;
    END
  END FREEZE_PMOS[23]
  PIN BcidMtx[474]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7469.065 1046.435 7469.345 1047.435 ;
    END
  END BcidMtx[474]
  PIN Data_PMOS[485]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7466.265 1046.435 7466.545 1047.435 ;
    END
  END Data_PMOS[485]
  PIN Data_PMOS[498]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7465.145 1046.435 7465.425 1047.435 ;
    END
  END Data_PMOS[498]
  PIN Data_PMOS[494]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7462.905 1046.435 7463.185 1047.435 ;
    END
  END Data_PMOS[494]
  PIN Data_PMOS[500]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7461.225 1046.435 7461.505 1047.435 ;
    END
  END Data_PMOS[500]
  PIN MASKH[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7451.705 1046.435 7451.985 1047.435 ;
    END
  END MASKH[79]
  PIN DIG_MON_SEL[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7448.345 1046.435 7448.625 1047.435 ;
    END
  END DIG_MON_SEL[158]
  PIN INJ_ROW[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7442.465 1046.435 7442.745 1047.435 ;
    END
  END INJ_ROW[78]
  PIN Data_PMOS[480]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7441.345 1046.435 7441.625 1047.435 ;
    END
  END Data_PMOS[480]
  PIN Data_PMOS[481]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7439.665 1046.435 7439.945 1047.435 ;
    END
  END Data_PMOS[481]
  PIN Data_PMOS[476]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7411.945 1046.435 7412.225 1047.435 ;
    END
  END Data_PMOS[476]
  PIN Data_PMOS[468]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7410.825 1046.435 7411.105 1047.435 ;
    END
  END Data_PMOS[468]
  PIN BcidMtx[473]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7407.465 1046.435 7407.745 1047.435 ;
    END
  END BcidMtx[473]
  PIN FREEZE_PMOS[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7405.785 1046.435 7406.065 1047.435 ;
    END
  END FREEZE_PMOS[22]
  PIN Data_HV[1114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18809.625 1046.435 18809.905 1047.435 ;
    END
  END Data_HV[1114]
  PIN BcidMtx[469]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7404.105 1046.435 7404.385 1047.435 ;
    END
  END BcidMtx[469]
  PIN Data_PMOS[464]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7400.745 1046.435 7401.025 1047.435 ;
    END
  END Data_PMOS[464]
  PIN Data_PMOS[477]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7386.745 1046.435 7387.025 1047.435 ;
    END
  END Data_PMOS[477]
  PIN Data_PMOS[478]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7385.065 1046.435 7385.345 1047.435 ;
    END
  END Data_PMOS[478]
  PIN MASKV[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7382.265 1046.435 7382.545 1047.435 ;
    END
  END MASKV[156]
  PIN DIG_MON_PMOS[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7380.025 1046.435 7380.305 1047.435 ;
    END
  END DIG_MON_PMOS[44]
  PIN DIG_MON_SEL[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7377.785 1046.435 7378.065 1047.435 ;
    END
  END DIG_MON_SEL[155]
  PIN INJ_ROW[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7374.425 1046.435 7374.705 1047.435 ;
    END
  END INJ_ROW[77]
  PIN Data_PMOS[449]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7332.985 1046.435 7333.265 1047.435 ;
    END
  END Data_PMOS[449]
  PIN Data_PMOS[446]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7331.305 1046.435 7331.585 1047.435 ;
    END
  END Data_PMOS[446]
  PIN Data_PMOS[455]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7329.625 1046.435 7329.905 1047.435 ;
    END
  END Data_PMOS[455]
  PIN INJ_IN[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7327.385 1046.435 7327.665 1047.435 ;
    END
  END INJ_IN[155]
  PIN Data_HV[1124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18810.185 1046.435 18810.465 1047.435 ;
    END
  END Data_HV[1124]
  PIN FREEZE_PMOS[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7323.465 1046.435 7323.745 1047.435 ;
    END
  END FREEZE_PMOS[21]
  PIN BcidMtx[463]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7321.785 1046.435 7322.065 1047.435 ;
    END
  END BcidMtx[463]
  PIN INJ_IN[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7311.705 1046.435 7311.985 1047.435 ;
    END
  END INJ_IN[154]
  PIN Data_PMOS[456]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7308.905 1046.435 7309.185 1047.435 ;
    END
  END Data_PMOS[456]
  PIN Data_PMOS[457]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7307.225 1046.435 7307.505 1047.435 ;
    END
  END Data_PMOS[457]
  PIN Data_PMOS[441]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7305.545 1046.435 7305.825 1047.435 ;
    END
  END Data_PMOS[441]
  PIN MASKH[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7301.905 1046.435 7302.185 1047.435 ;
    END
  END MASKH[77]
  PIN DIG_MON_PMOS[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7300.225 1046.435 7300.505 1047.435 ;
    END
  END DIG_MON_PMOS[42]
  PIN FREEZE_PMOS[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7553.065 1046.435 7553.345 1047.435 ;
    END
  END FREEZE_PMOS[24]
  PIN INJ_ROW[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8388.585 1046.435 8388.865 1047.435 ;
    END
  END INJ_ROW[90]
  PIN Data_PMOS[732]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8387.465 1046.435 8387.745 1047.435 ;
    END
  END Data_PMOS[732]
  PIN Data_PMOS[733]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8385.785 1046.435 8386.065 1047.435 ;
    END
  END Data_PMOS[733]
  PIN Data_PMOS[728]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8383.545 1046.435 8383.825 1047.435 ;
    END
  END Data_PMOS[728]
  PIN Data_PMOS[720]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8382.425 1046.435 8382.705 1047.435 ;
    END
  END Data_PMOS[720]
  PIN BcidMtx[545]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8365.625 1046.435 8365.905 1047.435 ;
    END
  END BcidMtx[545]
  PIN Read_PMOS[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8363.385 1046.435 8363.665 1047.435 ;
    END
  END Read_PMOS[34]
  PIN BcidMtx[541]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8362.265 1046.435 8362.545 1047.435 ;
    END
  END BcidMtx[541]
  PIN Data_PMOS[717]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8359.465 1046.435 8359.745 1047.435 ;
    END
  END Data_PMOS[717]
  PIN Data_PMOS[724]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8357.225 1046.435 8357.505 1047.435 ;
    END
  END Data_PMOS[724]
  PIN Data_PMOS[730]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8356.105 1046.435 8356.385 1047.435 ;
    END
  END Data_PMOS[730]
  PIN Data_PMOS[714]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8354.425 1046.435 8354.705 1047.435 ;
    END
  END Data_PMOS[714]
  PIN MASKD[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8313.545 1046.435 8313.825 1047.435 ;
    END
  END MASKD[180]
  PIN MASKD[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8309.065 1046.435 8309.345 1047.435 ;
    END
  END MASKD[179]
  PIN Data_PMOS[711]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8305.705 1046.435 8305.985 1047.435 ;
    END
  END Data_PMOS[711]
  PIN Data_PMOS[705]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8304.585 1046.435 8304.865 1047.435 ;
    END
  END Data_PMOS[705]
  PIN Data_PMOS[706]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8302.905 1046.435 8303.185 1047.435 ;
    END
  END Data_PMOS[706]
  PIN Data_PMOS[699]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8292.265 1046.435 8292.545 1047.435 ;
    END
  END Data_PMOS[699]
  PIN nTOK_PMOS[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8290.025 1046.435 8290.305 1047.435 ;
    END
  END nTOK_PMOS[33]
  PIN BcidMtx[537]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8287.785 1046.435 8288.065 1047.435 ;
    END
  END BcidMtx[537]
  PIN BcidMtx[535]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8285.545 1046.435 8285.825 1047.435 ;
    END
  END BcidMtx[535]
  PIN BcidMtx[534]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8284.985 1046.435 8285.265 1047.435 ;
    END
  END BcidMtx[534]
  PIN Data_PMOS[695]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8280.225 1046.435 8280.505 1047.435 ;
    END
  END Data_PMOS[695]
  PIN Data_PMOS[697]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8252.505 1046.435 8252.785 1047.435 ;
    END
  END Data_PMOS[697]
  PIN Data_PMOS[704]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8251.385 1046.435 8251.665 1047.435 ;
    END
  END Data_PMOS[704]
  PIN Data_PMOS[710]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8249.705 1046.435 8249.985 1047.435 ;
    END
  END Data_PMOS[710]
  PIN DIG_MON_PMOS[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8246.905 1046.435 8247.185 1047.435 ;
    END
  END DIG_MON_PMOS[66]
  PIN DIG_MON_SEL[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8245.225 1046.435 8245.505 1047.435 ;
    END
  END DIG_MON_SEL[178]
  PIN Data_PMOS[837]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8800.185 1046.435 8800.465 1047.435 ;
    END
  END Data_PMOS[837]
  PIN Data_PMOS[838]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8785.625 1046.435 8785.905 1047.435 ;
    END
  END Data_PMOS[838]
  PIN Data_PMOS[833]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8783.385 1046.435 8783.665 1047.435 ;
    END
  END Data_PMOS[833]
  PIN Data_PMOS[825]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8782.265 1046.435 8782.545 1047.435 ;
    END
  END Data_PMOS[825]
  PIN BcidMtx[575]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8778.905 1046.435 8779.185 1047.435 ;
    END
  END BcidMtx[575]
  PIN FREEZE_PMOS[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8777.225 1046.435 8777.505 1047.435 ;
    END
  END FREEZE_PMOS[39]
  PIN BcidMtx[571]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8775.545 1046.435 8775.825 1047.435 ;
    END
  END BcidMtx[571]
  PIN Data_PMOS[822]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8734.105 1046.435 8734.385 1047.435 ;
    END
  END Data_PMOS[822]
  PIN Data_PMOS[834]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8732.425 1046.435 8732.705 1047.435 ;
    END
  END Data_PMOS[834]
  PIN Data_PMOS[835]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8730.745 1046.435 8731.025 1047.435 ;
    END
  END Data_PMOS[835]
  PIN Data_PMOS[819]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8729.065 1046.435 8729.345 1047.435 ;
    END
  END Data_PMOS[819]
  PIN MASKH[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8727.385 1046.435 8727.665 1047.435 ;
    END
  END MASKH[95]
  PIN MASKD[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8722.345 1046.435 8722.625 1047.435 ;
    END
  END MASKD[189]
  PIN MASKV[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8711.145 1046.435 8711.425 1047.435 ;
    END
  END MASKV[189]
  PIN Data_PMOS[810]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8709.465 1046.435 8709.745 1047.435 ;
    END
  END Data_PMOS[810]
  PIN Data_PMOS[811]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8707.785 1046.435 8708.065 1047.435 ;
    END
  END Data_PMOS[811]
  PIN Data_PMOS[805]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8706.105 1046.435 8706.385 1047.435 ;
    END
  END Data_PMOS[805]
  PIN nTOK_PMOS[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8701.345 1046.435 8701.625 1047.435 ;
    END
  END nTOK_PMOS[38]
  PIN BcidMtx[567]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8699.105 1046.435 8699.385 1047.435 ;
    END
  END BcidMtx[567]
  PIN BcidMtx[564]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8670.825 1046.435 8671.105 1047.435 ;
    END
  END BcidMtx[564]
  PIN Data_PMOS[801]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8668.585 1046.435 8668.865 1047.435 ;
    END
  END Data_PMOS[801]
  PIN Data_PMOS[813]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8666.905 1046.435 8667.185 1047.435 ;
    END
  END Data_PMOS[813]
  PIN Data_PMOS[799]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8664.105 1046.435 8664.385 1047.435 ;
    END
  END Data_PMOS[799]
  PIN Data_PMOS[815]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8662.985 1046.435 8663.265 1047.435 ;
    END
  END Data_PMOS[815]
  PIN MASKD[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8661.305 1046.435 8661.585 1047.435 ;
    END
  END MASKD[188]
  PIN DIG_MON_SEL[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8645.065 1046.435 8645.345 1047.435 ;
    END
  END DIG_MON_SEL[187]
  PIN DIG_MON_PMOS[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8642.825 1046.435 8643.105 1047.435 ;
    END
  END DIG_MON_PMOS[75]
  PIN MASKV[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18807.945 1046.435 18808.225 1047.435 ;
    END
  END MASKV[442]
  PIN Data_PMOS[785]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8640.025 1046.435 8640.305 1047.435 ;
    END
  END Data_PMOS[785]
  PIN Data_PMOS[782]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8638.345 1046.435 8638.625 1047.435 ;
    END
  END Data_PMOS[782]
  PIN Data_PMOS[791]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8636.665 1046.435 8636.945 1047.435 ;
    END
  END Data_PMOS[791]
  PIN nTOK_PMOS[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8594.105 1046.435 8594.385 1047.435 ;
    END
  END nTOK_PMOS[37]
  PIN BcidMtx[562]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8592.425 1046.435 8592.705 1047.435 ;
    END
  END BcidMtx[562]
  PIN Read_PMOS[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8590.745 1046.435 8591.025 1047.435 ;
    END
  END Read_PMOS[37]
  PIN Data_PMOS[780]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8586.825 1046.435 8587.105 1047.435 ;
    END
  END Data_PMOS[780]
  PIN Data_PMOS[786]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8585.705 1046.435 8585.985 1047.435 ;
    END
  END Data_PMOS[786]
  PIN Data_PMOS[781]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8584.025 1046.435 8584.305 1047.435 ;
    END
  END Data_PMOS[781]
  PIN Data_PMOS[778]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8582.345 1046.435 8582.625 1047.435 ;
    END
  END Data_PMOS[778]
  PIN MASKV[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8572.265 1046.435 8572.545 1047.435 ;
    END
  END MASKV[186]
  PIN DIG_MON_PMOS[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8570.025 1046.435 8570.305 1047.435 ;
    END
  END DIG_MON_PMOS[74]
  PIN MASKD[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8566.665 1046.435 8566.945 1047.435 ;
    END
  END MASKD[185]
  PIN MASKV[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8561.905 1046.435 8562.185 1047.435 ;
    END
  END MASKV[185]
  PIN Data_PMOS[768]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8560.225 1046.435 8560.505 1047.435 ;
    END
  END Data_PMOS[768]
  PIN Data_HV[1058]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18640.785 1046.435 18641.065 1047.435 ;
    END
  END Data_HV[1058]
  PIN Data_PMOS[770]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8531.945 1046.435 8532.225 1047.435 ;
    END
  END Data_PMOS[770]
  PIN INJ_IN[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8529.705 1046.435 8529.985 1047.435 ;
    END
  END INJ_IN[185]
  PIN BcidMtx[555]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8526.345 1046.435 8526.625 1047.435 ;
    END
  END BcidMtx[555]
  PIN Read_PMOS[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8525.225 1046.435 8525.505 1047.435 ;
    END
  END Read_PMOS[36]
  PIN BcidMtx[552]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8523.545 1046.435 8523.825 1047.435 ;
    END
  END BcidMtx[552]
  PIN Data_PMOS[758]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8520.745 1046.435 8521.025 1047.435 ;
    END
  END Data_PMOS[758]
  PIN Data_PMOS[766]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8506.185 1046.435 8506.465 1047.435 ;
    END
  END Data_PMOS[766]
  PIN Data_PMOS[767]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8504.505 1046.435 8504.785 1047.435 ;
    END
  END Data_PMOS[767]
  PIN MASKV[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8502.265 1046.435 8502.545 1047.435 ;
    END
  END MASKV[184]
  PIN DIG_MON_PMOS[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8500.025 1046.435 8500.305 1047.435 ;
    END
  END DIG_MON_PMOS[72]
  PIN DIG_MON_SEL[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8498.345 1046.435 8498.625 1047.435 ;
    END
  END DIG_MON_SEL[184]
  PIN MASKV[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8493.865 1046.435 8494.145 1047.435 ;
    END
  END MASKV[183]
  PIN Data_PMOS[753]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8453.545 1046.435 8453.825 1047.435 ;
    END
  END Data_PMOS[753]
  PIN Data_PMOS[754]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8451.865 1046.435 8452.145 1047.435 ;
    END
  END Data_PMOS[754]
  PIN Data_PMOS[742]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8449.065 1046.435 8449.345 1047.435 ;
    END
  END Data_PMOS[742]
  PIN INJ_IN[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8447.385 1046.435 8447.665 1047.435 ;
    END
  END INJ_IN[183]
  PIN FREEZE_PMOS[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8443.465 1046.435 8443.745 1047.435 ;
    END
  END FREEZE_PMOS[35]
  PIN BcidMtx[548]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8442.345 1046.435 8442.625 1047.435 ;
    END
  END BcidMtx[548]
  PIN BcidMtx[546]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8441.225 1046.435 8441.505 1047.435 ;
    END
  END BcidMtx[546]
  PIN Data_PMOS[750]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8428.905 1046.435 8429.185 1047.435 ;
    END
  END Data_PMOS[750]
  PIN Data_PMOS[745]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8428.345 1046.435 8428.625 1047.435 ;
    END
  END Data_PMOS[745]
  PIN Data_PMOS[746]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8426.665 1046.435 8426.945 1047.435 ;
    END
  END Data_PMOS[746]
  PIN MASKH[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8421.905 1046.435 8422.185 1047.435 ;
    END
  END MASKH[91]
  PIN DIG_MON_SEL[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9511.945 1046.435 9512.225 1047.435 ;
    END
  END DIG_MON_SEL[209]
  PIN DIG_MON_PMOS[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9509.705 1046.435 9509.985 1047.435 ;
    END
  END DIG_MON_PMOS[97]
  PIN Data_PMOS[1026]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9507.465 1046.435 9507.745 1047.435 ;
    END
  END Data_PMOS[1026]
  PIN Data_PMOS[1020]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9506.345 1046.435 9506.625 1047.435 ;
    END
  END Data_PMOS[1020]
  PIN Data_PMOS[1028]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9504.105 1046.435 9504.385 1047.435 ;
    END
  END Data_PMOS[1028]
  PIN Data_PMOS[1015]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9502.985 1046.435 9503.265 1047.435 ;
    END
  END Data_PMOS[1015]
  PIN nTOK_PMOS[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9500.185 1046.435 9500.465 1047.435 ;
    END
  END nTOK_PMOS[48]
  PIN Read_PMOS[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9483.385 1046.435 9483.665 1047.435 ;
    END
  END Read_PMOS[48]
  PIN BcidMtx[626]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9482.825 1046.435 9483.105 1047.435 ;
    END
  END BcidMtx[626]
  PIN INJ_IN[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9480.585 1046.435 9480.865 1047.435 ;
    END
  END INJ_IN[208]
  PIN Data_PMOS[1018]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9477.225 1046.435 9477.505 1047.435 ;
    END
  END Data_PMOS[1018]
  PIN Data_PMOS[1012]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9476.665 1046.435 9476.945 1047.435 ;
    END
  END Data_PMOS[1012]
  PIN Data_PMOS[1009]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9474.985 1046.435 9475.265 1047.435 ;
    END
  END Data_PMOS[1009]
  PIN MASKH[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9434.105 1046.435 9434.385 1047.435 ;
    END
  END MASKH[104]
  PIN DIG_MON_SEL[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9430.185 1046.435 9430.465 1047.435 ;
    END
  END DIG_MON_SEL[207]
  PIN Data_PMOS[1005]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9425.705 1046.435 9425.985 1047.435 ;
    END
  END Data_PMOS[1005]
  PIN Data_PMOS[999]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9424.585 1046.435 9424.865 1047.435 ;
    END
  END Data_PMOS[999]
  PIN Data_PMOS[992]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9423.465 1046.435 9423.745 1047.435 ;
    END
  END Data_PMOS[992]
  PIN Data_PMOS[994]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9421.225 1046.435 9421.505 1047.435 ;
    END
  END Data_PMOS[994]
  PIN Data_PMOS[993]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9412.265 1046.435 9412.545 1047.435 ;
    END
  END Data_PMOS[993]
  PIN BcidMtx[623]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9408.905 1046.435 9409.185 1047.435 ;
    END
  END BcidMtx[623]
  PIN FREEZE_PMOS[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9407.225 1046.435 9407.505 1047.435 ;
    END
  END FREEZE_PMOS[47]
  PIN BcidMtx[619]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9405.545 1046.435 9405.825 1047.435 ;
    END
  END BcidMtx[619]
  PIN Data_PMOS[990]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9400.785 1046.435 9401.065 1047.435 ;
    END
  END Data_PMOS[990]
  PIN Data_PMOS[991]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9372.505 1046.435 9372.785 1047.435 ;
    END
  END Data_PMOS[991]
  PIN Data_PMOS[988]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9370.825 1046.435 9371.105 1047.435 ;
    END
  END Data_PMOS[988]
  PIN MASKV[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9369.145 1046.435 9369.425 1047.435 ;
    END
  END MASKV[206]
  PIN DIG_MON_PMOS[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9366.905 1046.435 9367.185 1047.435 ;
    END
  END DIG_MON_PMOS[94]
  PIN DIG_MON_SEL[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9364.665 1046.435 9364.945 1047.435 ;
    END
  END DIG_MON_SEL[205]
  PIN INJ_ROW[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9361.305 1046.435 9361.585 1047.435 ;
    END
  END INJ_ROW[102]
  PIN Data_PMOS[974]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9359.625 1046.435 9359.905 1047.435 ;
    END
  END Data_PMOS[974]
  PIN MASKD[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7123.545 1046.435 7123.825 1047.435 ;
    END
  END MASKD[149]
  PIN Data_PMOS[396]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7120.185 1046.435 7120.465 1047.435 ;
    END
  END Data_PMOS[396]
  PIN Data_PMOS[397]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7105.625 1046.435 7105.905 1047.435 ;
    END
  END Data_PMOS[397]
  PIN Data_PMOS[391]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7104.505 1046.435 7104.785 1047.435 ;
    END
  END Data_PMOS[391]
  PIN Data_PMOS[384]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7102.265 1046.435 7102.545 1047.435 ;
    END
  END Data_PMOS[384]
  PIN BcidMtx[449]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7098.905 1046.435 7099.185 1047.435 ;
    END
  END BcidMtx[449]
  PIN BcidMtx[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7097.785 1046.435 7098.065 1047.435 ;
    END
  END BcidMtx[447]
  PIN BcidMtx[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7095.545 1046.435 7095.825 1047.435 ;
    END
  END BcidMtx[445]
  PIN Data_PMOS[381]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7054.105 1046.435 7054.385 1047.435 ;
    END
  END Data_PMOS[381]
  PIN Data_PMOS[393]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7052.425 1046.435 7052.705 1047.435 ;
    END
  END Data_PMOS[393]
  PIN Data_PMOS[394]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7050.745 1046.435 7051.025 1047.435 ;
    END
  END Data_PMOS[394]
  PIN Data_PMOS[378]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7049.065 1046.435 7049.345 1047.435 ;
    END
  END Data_PMOS[378]
  PIN MASKV[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7047.945 1046.435 7048.225 1047.435 ;
    END
  END MASKV[148]
  PIN MASKD[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7042.345 1046.435 7042.625 1047.435 ;
    END
  END MASKD[147]
  PIN INJ_ROW[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7031.705 1046.435 7031.985 1047.435 ;
    END
  END INJ_ROW[73]
  PIN Data_PMOS[369]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7029.465 1046.435 7029.745 1047.435 ;
    END
  END Data_PMOS[369]
  PIN Data_PMOS[370]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7027.785 1046.435 7028.065 1047.435 ;
    END
  END Data_PMOS[370]
  PIN Data_PMOS[364]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7026.105 1046.435 7026.385 1047.435 ;
    END
  END Data_PMOS[364]
  PIN nTOK_PMOS[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7021.345 1046.435 7021.625 1047.435 ;
    END
  END nTOK_PMOS[17]
  PIN BcidMtx[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7019.105 1046.435 7019.385 1047.435 ;
    END
  END BcidMtx[441]
  PIN BcidMtx[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6991.945 1046.435 6992.225 1047.435 ;
    END
  END BcidMtx[440]
  PIN Data_PMOS[360]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6988.585 1046.435 6988.865 1047.435 ;
    END
  END Data_PMOS[360]
  PIN Data_PMOS[372]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6986.905 1046.435 6987.185 1047.435 ;
    END
  END Data_PMOS[372]
  PIN Data_PMOS[361]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6985.785 1046.435 6986.065 1047.435 ;
    END
  END Data_PMOS[361]
  PIN Data_PMOS[357]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6983.545 1046.435 6983.825 1047.435 ;
    END
  END Data_PMOS[357]
  PIN MASKH[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6981.865 1046.435 6982.145 1047.435 ;
    END
  END MASKH[73]
  PIN DIG_MON_PMOS[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6980.185 1046.435 6980.465 1047.435 ;
    END
  END DIG_MON_PMOS[34]
  PIN MASKD[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6963.945 1046.435 6964.225 1047.435 ;
    END
  END MASKD[145]
  PIN MASKV[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6961.145 1046.435 6961.425 1047.435 ;
    END
  END MASKV[145]
  PIN Data_PMOS[344]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6960.025 1046.435 6960.305 1047.435 ;
    END
  END Data_PMOS[344]
  PIN Data_PMOS[349]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6957.785 1046.435 6958.065 1047.435 ;
    END
  END Data_PMOS[349]
  PIN Data_PMOS[343]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6956.105 1046.435 6956.385 1047.435 ;
    END
  END Data_PMOS[343]
  PIN INJ_IN[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6954.425 1046.435 6954.705 1047.435 ;
    END
  END INJ_IN[145]
  PIN BcidMtx[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6911.865 1046.435 6912.145 1047.435 ;
    END
  END BcidMtx[435]
  PIN BcidMtx[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6910.185 1046.435 6910.465 1047.435 ;
    END
  END BcidMtx[434]
  PIN BcidMtx[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6909.625 1046.435 6909.905 1047.435 ;
    END
  END BcidMtx[433]
  PIN Data_PMOS[338]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6906.265 1046.435 6906.545 1047.435 ;
    END
  END Data_PMOS[338]
  PIN Data_PMOS[346]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6904.585 1046.435 6904.865 1047.435 ;
    END
  END Data_PMOS[346]
  PIN Data_PMOS[352]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6903.465 1046.435 6903.745 1047.435 ;
    END
  END Data_PMOS[352]
  PIN Data_PMOS[353]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6901.225 1046.435 6901.505 1047.435 ;
    END
  END Data_PMOS[353]
  PIN MASKD[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6891.145 1046.435 6891.425 1047.435 ;
    END
  END MASKD[144]
  PIN MASKV[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6881.905 1046.435 6882.185 1047.435 ;
    END
  END MASKV[143]
  PIN Data_PMOS[323]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6880.785 1046.435 6881.065 1047.435 ;
    END
  END Data_PMOS[323]
  PIN Data_PMOS[334]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6879.665 1046.435 6879.945 1047.435 ;
    END
  END Data_PMOS[334]
  PIN Data_PMOS[335]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6852.505 1046.435 6852.785 1047.435 ;
    END
  END Data_PMOS[335]
  PIN Data_PMOS[321]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6850.825 1046.435 6851.105 1047.435 ;
    END
  END Data_PMOS[321]
  PIN BcidMtx[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6846.345 1046.435 6846.625 1047.435 ;
    END
  END BcidMtx[429]
  PIN BcidMtx[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6844.665 1046.435 6844.945 1047.435 ;
    END
  END BcidMtx[428]
  PIN BcidMtx[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6843.545 1046.435 6843.825 1047.435 ;
    END
  END BcidMtx[426]
  PIN Data_PMOS[324]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6840.185 1046.435 6840.465 1047.435 ;
    END
  END Data_PMOS[324]
  PIN Data_PMOS[319]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6825.625 1046.435 6825.905 1047.435 ;
    END
  END Data_PMOS[319]
  PIN Data_PMOS[326]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6824.505 1046.435 6824.785 1047.435 ;
    END
  END Data_PMOS[326]
  PIN MASKV[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6822.265 1046.435 6822.545 1047.435 ;
    END
  END MASKV[142]
  PIN DIG_MON_PMOS[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6820.025 1046.435 6820.305 1047.435 ;
    END
  END DIG_MON_PMOS[30]
  PIN DIG_MON_SEL[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6818.345 1046.435 6818.625 1047.435 ;
    END
  END DIG_MON_SEL[142]
  PIN INJ_ROW[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6814.425 1046.435 6814.705 1047.435 ;
    END
  END INJ_ROW[70]
  PIN Data_PMOS[302]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6772.985 1046.435 6773.265 1047.435 ;
    END
  END Data_PMOS[302]
  PIN Data_PMOS[313]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6771.865 1046.435 6772.145 1047.435 ;
    END
  END Data_PMOS[313]
  PIN Data_PMOS[308]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6769.625 1046.435 6769.905 1047.435 ;
    END
  END Data_PMOS[308]
  PIN INJ_IN[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6767.385 1046.435 6767.665 1047.435 ;
    END
  END INJ_IN[141]
  PIN BcidMtx[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6765.145 1046.435 6765.425 1047.435 ;
    END
  END BcidMtx[425]
  PIN Read_PMOS[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6762.905 1046.435 6763.185 1047.435 ;
    END
  END Read_PMOS[14]
  PIN BcidMtx[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6761.225 1046.435 6761.505 1047.435 ;
    END
  END BcidMtx[420]
  PIN INJ_IN[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6751.705 1046.435 6751.985 1047.435 ;
    END
  END INJ_IN[140]
  PIN Data_PMOS[309]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6748.905 1046.435 6749.185 1047.435 ;
    END
  END Data_PMOS[309]
  PIN Data_PMOS[298]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6747.785 1046.435 6748.065 1047.435 ;
    END
  END Data_PMOS[298]
  PIN Data_PMOS[305]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6746.665 1046.435 6746.945 1047.435 ;
    END
  END Data_PMOS[305]
  PIN MASKV[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6742.465 1046.435 6742.745 1047.435 ;
    END
  END MASKV[140]
  PIN DIG_MON_PMOS[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6740.225 1046.435 6740.505 1047.435 ;
    END
  END DIG_MON_PMOS[28]
  PIN DIG_MON_SEL[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6738.545 1046.435 6738.825 1047.435 ;
    END
  END DIG_MON_SEL[140]
  PIN DIG_MON_PMOS[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7829.705 1046.435 7829.985 1047.435 ;
    END
  END DIG_MON_PMOS[55]
  PIN Data_PMOS[585]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7827.465 1046.435 7827.745 1047.435 ;
    END
  END Data_PMOS[585]
  PIN Data_PMOS[579]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7826.345 1046.435 7826.625 1047.435 ;
    END
  END Data_PMOS[579]
  PIN Data_PMOS[587]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7824.105 1046.435 7824.385 1047.435 ;
    END
  END Data_PMOS[587]
  PIN Data_PMOS[573]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7822.425 1046.435 7822.705 1047.435 ;
    END
  END Data_PMOS[573]
  PIN nTOK_PMOS[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7820.185 1046.435 7820.465 1047.435 ;
    END
  END nTOK_PMOS[27]
  PIN FREEZE_PMOS[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7803.945 1046.435 7804.225 1047.435 ;
    END
  END FREEZE_PMOS[27]
  PIN BcidMtx[499]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7802.265 1046.435 7802.545 1047.435 ;
    END
  END BcidMtx[499]
  PIN INJ_IN[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7800.585 1046.435 7800.865 1047.435 ;
    END
  END INJ_IN[166]
  PIN Data_PMOS[576]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7798.345 1046.435 7798.625 1047.435 ;
    END
  END Data_PMOS[576]
  PIN Data_PMOS[571]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7796.665 1046.435 7796.945 1047.435 ;
    END
  END Data_PMOS[571]
  PIN Data_PMOS[578]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7795.545 1046.435 7795.825 1047.435 ;
    END
  END Data_PMOS[578]
  PIN MASKV[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7754.665 1046.435 7754.945 1047.435 ;
    END
  END MASKV[166]
  PIN DIG_MON_PMOS[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7752.425 1046.435 7752.705 1047.435 ;
    END
  END DIG_MON_PMOS[54]
  PIN DIG_MON_SEL[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7750.745 1046.435 7751.025 1047.435 ;
    END
  END DIG_MON_SEL[166]
  PIN INJ_ROW[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7746.825 1046.435 7747.105 1047.435 ;
    END
  END INJ_ROW[82]
  PIN Data_PMOS[554]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7745.145 1046.435 7745.425 1047.435 ;
    END
  END Data_PMOS[554]
  PIN Data_PMOS[565]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7744.025 1046.435 7744.305 1047.435 ;
    END
  END Data_PMOS[565]
  PIN Data_PMOS[560]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7741.785 1046.435 7742.065 1047.435 ;
    END
  END Data_PMOS[560]
  PIN INJ_IN[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7731.145 1046.435 7731.425 1047.435 ;
    END
  END INJ_IN[165]
  PIN BcidMtx[497]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7728.905 1046.435 7729.185 1047.435 ;
    END
  END BcidMtx[497]
  PIN Read_PMOS[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7726.665 1046.435 7726.945 1047.435 ;
    END
  END Read_PMOS[26]
  PIN BcidMtx[492]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7724.985 1046.435 7725.265 1047.435 ;
    END
  END BcidMtx[492]
  PIN Data_PMOS[549]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7720.785 1046.435 7721.065 1047.435 ;
    END
  END Data_PMOS[549]
  PIN Data_HV[1117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18811.305 1046.435 18811.585 1047.435 ;
    END
  END Data_HV[1117]
  PIN Data_PMOS[562]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7691.945 1046.435 7692.225 1047.435 ;
    END
  END Data_PMOS[562]
  PIN Data_PMOS[547]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7690.825 1046.435 7691.105 1047.435 ;
    END
  END Data_PMOS[547]
  PIN MASKH[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7688.585 1046.435 7688.865 1047.435 ;
    END
  END MASKH[82]
  PIN DIG_MON_SEL[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7684.665 1046.435 7684.945 1047.435 ;
    END
  END DIG_MON_SEL[163]
  PIN Data_PMOS[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5985.625 1046.435 5985.905 1047.435 ;
    END
  END Data_PMOS[103]
  PIN Data_PMOS[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5984.505 1046.435 5984.785 1047.435 ;
    END
  END Data_PMOS[97]
  PIN Data_PMOS[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5982.825 1046.435 5983.105 1047.435 ;
    END
  END Data_PMOS[91]
  PIN BcidMtx[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5978.905 1046.435 5979.185 1047.435 ;
    END
  END BcidMtx[365]
  PIN BcidMtx[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5977.785 1046.435 5978.065 1047.435 ;
    END
  END BcidMtx[363]
  PIN BcidMtx[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5976.105 1046.435 5976.385 1047.435 ;
    END
  END BcidMtx[362]
  PIN Data_PMOS[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5934.105 1046.435 5934.385 1047.435 ;
    END
  END Data_PMOS[87]
  PIN Data_PMOS[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5932.985 1046.435 5933.265 1047.435 ;
    END
  END Data_PMOS[93]
  PIN Data_PMOS[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5931.305 1046.435 5931.585 1047.435 ;
    END
  END Data_PMOS[88]
  PIN Data_PMOS[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5929.065 1046.435 5929.345 1047.435 ;
    END
  END Data_PMOS[84]
  PIN MASKV[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5927.945 1046.435 5928.225 1047.435 ;
    END
  END MASKV[120]
  PIN DIG_MON_PMOS[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5925.705 1046.435 5925.985 1047.435 ;
    END
  END DIG_MON_PMOS[8]
  PIN MASKD[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5922.345 1046.435 5922.625 1047.435 ;
    END
  END MASKD[119]
  PIN INJ_ROW[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5911.705 1046.435 5911.985 1047.435 ;
    END
  END INJ_ROW[59]
  PIN Data_PMOS[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5910.025 1046.435 5910.305 1047.435 ;
    END
  END Data_PMOS[71]
  PIN Data_PMOS[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5907.785 1046.435 5908.065 1047.435 ;
    END
  END Data_PMOS[76]
  PIN Data_PMOS[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5906.665 1046.435 5906.945 1047.435 ;
    END
  END Data_PMOS[77]
  PIN INJ_IN[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5902.465 1046.435 5902.745 1047.435 ;
    END
  END INJ_IN[119]
  PIN BcidMtx[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5899.105 1046.435 5899.385 1047.435 ;
    END
  END BcidMtx[357]
  PIN BcidMtx[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5871.945 1046.435 5872.225 1047.435 ;
    END
  END BcidMtx[356]
  PIN INJ_IN[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5869.705 1046.435 5869.985 1047.435 ;
    END
  END INJ_IN[118]
  PIN Data_PMOS[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5866.905 1046.435 5867.185 1047.435 ;
    END
  END Data_PMOS[78]
  PIN Data_PMOS[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5865.225 1046.435 5865.505 1047.435 ;
    END
  END Data_PMOS[79]
  PIN Data_PMOS[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5864.105 1046.435 5864.385 1047.435 ;
    END
  END Data_PMOS[64]
  PIN MASKH[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5861.865 1046.435 5862.145 1047.435 ;
    END
  END MASKH[59]
  PIN MASKD[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5843.945 1046.435 5844.225 1047.435 ;
    END
  END MASKD[117]
  PIN MASKV[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5841.145 1046.435 5841.425 1047.435 ;
    END
  END MASKV[117]
  PIN Data_PMOS[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5839.465 1046.435 5839.745 1047.435 ;
    END
  END Data_PMOS[54]
  PIN Data_PMOS[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5837.785 1046.435 5838.065 1047.435 ;
    END
  END Data_PMOS[55]
  PIN Data_PMOS[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5836.105 1046.435 5836.385 1047.435 ;
    END
  END Data_PMOS[49]
  PIN nTOK_PMOS[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5794.105 1046.435 5794.385 1047.435 ;
    END
  END nTOK_PMOS[2]
  PIN BcidMtx[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5791.865 1046.435 5792.145 1047.435 ;
    END
  END BcidMtx[351]
  PIN BcidMtx[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5790.185 1046.435 5790.465 1047.435 ;
    END
  END BcidMtx[350]
  PIN INJ_IN[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5787.945 1046.435 5788.225 1047.435 ;
    END
  END INJ_IN[116]
  PIN Data_PMOS[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5785.705 1046.435 5785.985 1047.435 ;
    END
  END Data_PMOS[51]
  PIN Data_PMOS[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5785.145 1046.435 5785.425 1047.435 ;
    END
  END Data_PMOS[57]
  PIN Data_PMOS[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5783.465 1046.435 5783.745 1047.435 ;
    END
  END Data_PMOS[58]
  PIN Data_PMOS[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5781.785 1046.435 5782.065 1047.435 ;
    END
  END Data_PMOS[42]
  PIN MASKH[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5771.705 1046.435 5771.985 1047.435 ;
    END
  END MASKH[58]
  PIN MASKD[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5766.665 1046.435 5766.945 1047.435 ;
    END
  END MASKD[115]
  PIN INJ_ROW[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5762.465 1046.435 5762.745 1047.435 ;
    END
  END INJ_ROW[57]
  PIN Data_PMOS[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5760.225 1046.435 5760.505 1047.435 ;
    END
  END Data_PMOS[33]
  PIN Data_PMOS[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5733.065 1046.435 5733.345 1047.435 ;
    END
  END Data_PMOS[34]
  PIN Data_PMOS[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5731.385 1046.435 5731.665 1047.435 ;
    END
  END Data_PMOS[28]
  PIN INJ_IN[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5729.705 1046.435 5729.985 1047.435 ;
    END
  END INJ_IN[115]
  PIN BcidMtx[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5726.905 1046.435 5727.185 1047.435 ;
    END
  END BcidMtx[346]
  PIN FREEZE_PMOS[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5725.785 1046.435 5726.065 1047.435 ;
    END
  END FREEZE_PMOS[1]
  PIN BcidMtx[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5724.665 1046.435 5724.945 1047.435 ;
    END
  END BcidMtx[344]
  PIN INJ_IN[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5722.425 1046.435 5722.705 1047.435 ;
    END
  END INJ_IN[114]
  PIN Data_PMOS[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5706.745 1046.435 5707.025 1047.435 ;
    END
  END Data_PMOS[36]
  PIN Data_PMOS[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5705.065 1046.435 5705.345 1047.435 ;
    END
  END Data_PMOS[37]
  PIN Data_PMOS[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5703.945 1046.435 5704.225 1047.435 ;
    END
  END Data_PMOS[22]
  PIN MASKV[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5702.265 1046.435 5702.545 1047.435 ;
    END
  END MASKV[114]
  PIN DIG_MON_PMOS[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5700.025 1046.435 5700.305 1047.435 ;
    END
  END DIG_MON_PMOS[2]
  PIN MASKD[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5696.665 1046.435 5696.945 1047.435 ;
    END
  END MASKD[113]
  PIN Data_PMOS[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5653.545 1046.435 5653.825 1047.435 ;
    END
  END Data_PMOS[18]
  PIN Data_PMOS[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5652.425 1046.435 5652.705 1047.435 ;
    END
  END Data_PMOS[12]
  PIN Data_PMOS[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5650.745 1046.435 5651.025 1047.435 ;
    END
  END Data_PMOS[13]
  PIN Data_PMOS[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5649.065 1046.435 5649.345 1047.435 ;
    END
  END Data_PMOS[7]
  PIN nTOK_PMOS[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5646.265 1046.435 5646.545 1047.435 ;
    END
  END nTOK_PMOS[0]
  PIN BcidMtx[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5644.025 1046.435 5644.305 1047.435 ;
    END
  END BcidMtx[339]
  PIN BcidMtx[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5642.345 1046.435 5642.625 1047.435 ;
    END
  END BcidMtx[338]
  PIN BcidMtx[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5641.225 1046.435 5641.505 1047.435 ;
    END
  END BcidMtx[336]
  PIN Data_PMOS[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5630.585 1046.435 5630.865 1047.435 ;
    END
  END Data_PMOS[3]
  PIN Data_PMOS[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5627.785 1046.435 5628.065 1047.435 ;
    END
  END Data_PMOS[4]
  PIN Data_PMOS[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5626.665 1046.435 5626.945 1047.435 ;
    END
  END Data_PMOS[11]
  PIN MASKV[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5622.465 1046.435 5622.745 1047.435 ;
    END
  END MASKV[112]
  PIN MASKD[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5621.345 1046.435 5621.625 1047.435 ;
    END
  END MASKD[112]
  PIN DIG_MON_SEL[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5618.545 1046.435 5618.825 1047.435 ;
    END
  END DIG_MON_SEL[112]
  PIN INJ_ROW[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6708.585 1046.435 6708.865 1047.435 ;
    END
  END INJ_ROW[69]
  PIN Data_PMOS[281]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6706.905 1046.435 6707.185 1047.435 ;
    END
  END Data_PMOS[281]
  PIN Data_PMOS[285]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6706.345 1046.435 6706.625 1047.435 ;
    END
  END Data_PMOS[285]
  PIN Data_PMOS[293]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6704.105 1046.435 6704.385 1047.435 ;
    END
  END Data_PMOS[293]
  PIN Data_PMOS[279]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6702.425 1046.435 6702.705 1047.435 ;
    END
  END Data_PMOS[279]
  PIN BcidMtx[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6685.625 1046.435 6685.905 1047.435 ;
    END
  END BcidMtx[419]
  PIN FREEZE_PMOS[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6683.945 1046.435 6684.225 1047.435 ;
    END
  END FREEZE_PMOS[13]
  PIN BcidMtx[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6682.265 1046.435 6682.545 1047.435 ;
    END
  END BcidMtx[415]
  PIN Data_PMOS[276]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6679.465 1046.435 6679.745 1047.435 ;
    END
  END Data_PMOS[276]
  PIN Data_PMOS[288]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6677.785 1046.435 6678.065 1047.435 ;
    END
  END Data_PMOS[288]
  PIN Data_PMOS[289]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6676.105 1046.435 6676.385 1047.435 ;
    END
  END Data_PMOS[289]
  PIN Data_PMOS[274]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6674.985 1046.435 6675.265 1047.435 ;
    END
  END Data_PMOS[274]
  PIN MASKH[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6634.105 1046.435 6634.385 1047.435 ;
    END
  END MASKH[69]
  PIN DIG_MON_PMOS[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6632.425 1046.435 6632.705 1047.435 ;
    END
  END DIG_MON_PMOS[26]
  PIN DIG_MON_SEL[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6630.185 1046.435 6630.465 1047.435 ;
    END
  END DIG_MON_SEL[137]
  PIN INJ_ROW[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6626.825 1046.435 6627.105 1047.435 ;
    END
  END INJ_ROW[68]
  PIN Data_PMOS[260]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6625.145 1046.435 6625.425 1047.435 ;
    END
  END Data_PMOS[260]
  PIN Data_PMOS[257]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6623.465 1046.435 6623.745 1047.435 ;
    END
  END Data_PMOS[257]
  PIN Data_PMOS[266]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6621.785 1046.435 6622.065 1047.435 ;
    END
  END Data_PMOS[266]
  PIN INJ_IN[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6611.145 1046.435 6611.425 1047.435 ;
    END
  END INJ_IN[137]
  PIN BcidMtx[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6608.345 1046.435 6608.625 1047.435 ;
    END
  END BcidMtx[412]
  PIN Read_PMOS[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6606.665 1046.435 6606.945 1047.435 ;
    END
  END Read_PMOS[12]
  PIN BcidMtx[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6604.985 1046.435 6605.265 1047.435 ;
    END
  END BcidMtx[408]
  PIN Data_PMOS[255]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6600.785 1046.435 6601.065 1047.435 ;
    END
  END Data_PMOS[255]
  PIN Data_PMOS[262]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6598.545 1046.435 6598.825 1047.435 ;
    END
  END Data_PMOS[262]
  PIN Data_PMOS[263]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6571.385 1046.435 6571.665 1047.435 ;
    END
  END Data_PMOS[263]
  PIN Data_PMOS[252]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6570.265 1046.435 6570.545 1047.435 ;
    END
  END Data_PMOS[252]
  PIN MASKD[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6568.025 1046.435 6568.305 1047.435 ;
    END
  END MASKD[136]
  PIN MASKD[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18646.665 1046.435 18646.945 1047.435 ;
    END
  END MASKD[437]
  PIN MASKD[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6563.545 1046.435 6563.825 1047.435 ;
    END
  END MASKD[135]
  PIN MASKV[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6560.745 1046.435 6561.025 1047.435 ;
    END
  END MASKV[135]
  PIN Data_PMOS[243]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6546.185 1046.435 6546.465 1047.435 ;
    END
  END Data_PMOS[243]
  PIN Data_PMOS[244]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6544.505 1046.435 6544.785 1047.435 ;
    END
  END Data_PMOS[244]
  PIN Data_PMOS[238]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6542.825 1046.435 6543.105 1047.435 ;
    END
  END Data_PMOS[238]
  PIN nTOK_PMOS[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6540.025 1046.435 6540.305 1047.435 ;
    END
  END nTOK_PMOS[11]
  PIN FREEZE_PMOS[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6537.225 1046.435 6537.505 1047.435 ;
    END
  END FREEZE_PMOS[11]
  PIN BcidMtx[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6536.105 1046.435 6536.385 1047.435 ;
    END
  END BcidMtx[404]
  PIN INJ_IN[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6533.865 1046.435 6534.145 1047.435 ;
    END
  END INJ_IN[134]
  PIN Data_PMOS[240]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6492.985 1046.435 6493.265 1047.435 ;
    END
  END Data_PMOS[240]
  PIN Data_PMOS[235]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6491.305 1046.435 6491.585 1047.435 ;
    END
  END Data_PMOS[235]
  PIN Data_PMOS[232]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6489.625 1046.435 6489.905 1047.435 ;
    END
  END Data_PMOS[232]
  PIN MASKV[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6487.945 1046.435 6488.225 1047.435 ;
    END
  END MASKV[134]
  PIN DIG_MON_PMOS[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6485.705 1046.435 6485.985 1047.435 ;
    END
  END DIG_MON_PMOS[22]
  PIN DIG_MON_SEL[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6483.465 1046.435 6483.745 1047.435 ;
    END
  END DIG_MON_SEL[133]
  PIN DIG_MON_PMOS[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6481.225 1046.435 6481.505 1047.435 ;
    END
  END DIG_MON_PMOS[21]
  PIN Data_PMOS[218]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6470.025 1046.435 6470.305 1047.435 ;
    END
  END Data_PMOS[218]
  PIN Data_PMOS[215]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6468.345 1046.435 6468.625 1047.435 ;
    END
  END Data_PMOS[215]
  PIN Data_PMOS[230]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6467.225 1046.435 6467.505 1047.435 ;
    END
  END Data_PMOS[230]
  PIN INJ_IN[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6462.465 1046.435 6462.745 1047.435 ;
    END
  END INJ_IN[133]
  PIN BcidMtx[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6459.665 1046.435 6459.945 1047.435 ;
    END
  END BcidMtx[400]
  PIN Read_PMOS[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6432.505 1046.435 6432.785 1047.435 ;
    END
  END Read_PMOS[10]
  PIN INJ_IN[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6429.705 1046.435 6429.985 1047.435 ;
    END
  END INJ_IN[132]
  PIN Data_PMOS[219]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6427.465 1046.435 6427.745 1047.435 ;
    END
  END Data_PMOS[219]
  PIN Data_PMOS[214]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6425.785 1046.435 6426.065 1047.435 ;
    END
  END Data_PMOS[214]
  PIN Data_PMOS[211]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6424.105 1046.435 6424.385 1047.435 ;
    END
  END Data_PMOS[211]
  PIN MASKV[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6422.425 1046.435 6422.705 1047.435 ;
    END
  END MASKV[132]
  PIN DIG_MON_PMOS[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6420.185 1046.435 6420.465 1047.435 ;
    END
  END DIG_MON_PMOS[20]
  PIN DIG_MON_SEL[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6405.065 1046.435 6405.345 1047.435 ;
    END
  END DIG_MON_SEL[131]
  PIN INJ_ROW[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6401.705 1046.435 6401.985 1047.435 ;
    END
  END INJ_ROW[65]
  PIN Data_PMOS[207]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6400.585 1046.435 6400.865 1047.435 ;
    END
  END Data_PMOS[207]
  PIN Data_PMOS[194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6398.345 1046.435 6398.625 1047.435 ;
    END
  END Data_PMOS[194]
  PIN Data_PMOS[203]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6396.665 1046.435 6396.945 1047.435 ;
    END
  END Data_PMOS[203]
  PIN INJ_IN[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6394.425 1046.435 6394.705 1047.435 ;
    END
  END INJ_IN[131]
  PIN BcidMtx[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6352.425 1046.435 6352.705 1047.435 ;
    END
  END BcidMtx[394]
  PIN Read_PMOS[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6350.745 1046.435 6351.025 1047.435 ;
    END
  END Read_PMOS[9]
  PIN BcidMtx[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6349.065 1046.435 6349.345 1047.435 ;
    END
  END BcidMtx[390]
  PIN Data_PMOS[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6346.265 1046.435 6346.545 1047.435 ;
    END
  END Data_PMOS[191]
  PIN Data_PMOS[199]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6344.585 1046.435 6344.865 1047.435 ;
    END
  END Data_PMOS[199]
  PIN Data_PMOS[205]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6343.465 1046.435 6343.745 1047.435 ;
    END
  END Data_PMOS[205]
  PIN Data_PMOS[206]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6341.225 1046.435 6341.505 1047.435 ;
    END
  END Data_PMOS[206]
  PIN MASKD[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6331.145 1046.435 6331.425 1047.435 ;
    END
  END MASKD[130]
  PIN DIG_MON_PMOS[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6325.545 1046.435 6325.825 1047.435 ;
    END
  END DIG_MON_PMOS[17]
  PIN Data_PMOS[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6321.345 1046.435 6321.625 1047.435 ;
    END
  END Data_PMOS[186]
  PIN Data_PMOS[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6319.665 1046.435 6319.945 1047.435 ;
    END
  END Data_PMOS[187]
  PIN Data_PMOS[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6292.505 1046.435 6292.785 1047.435 ;
    END
  END Data_PMOS[188]
  PIN Data_PMOS[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6290.825 1046.435 6291.105 1047.435 ;
    END
  END Data_PMOS[174]
  PIN BcidMtx[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6287.465 1046.435 6287.745 1047.435 ;
    END
  END BcidMtx[389]
  PIN FREEZE_PMOS[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6285.785 1046.435 6286.065 1047.435 ;
    END
  END FREEZE_PMOS[8]
  PIN BcidMtx[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6284.105 1046.435 6284.385 1047.435 ;
    END
  END BcidMtx[385]
  PIN INJ_IN[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6282.425 1046.435 6282.705 1047.435 ;
    END
  END INJ_IN[128]
  PIN Data_PMOS[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6266.745 1046.435 6267.025 1047.435 ;
    END
  END Data_PMOS[183]
  PIN Data_PMOS[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6265.625 1046.435 6265.905 1047.435 ;
    END
  END Data_PMOS[172]
  PIN Data_PMOS[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6264.505 1046.435 6264.785 1047.435 ;
    END
  END Data_PMOS[179]
  PIN MASKV[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6262.265 1046.435 6262.545 1047.435 ;
    END
  END MASKV[128]
  PIN DIG_MON_PMOS[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6260.025 1046.435 6260.305 1047.435 ;
    END
  END DIG_MON_PMOS[16]
  PIN DIG_MON_SEL[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6258.345 1046.435 6258.625 1047.435 ;
    END
  END DIG_MON_SEL[128]
  PIN INJ_ROW[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6254.425 1046.435 6254.705 1047.435 ;
    END
  END INJ_ROW[63]
  PIN Data_PMOS[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6212.985 1046.435 6213.265 1047.435 ;
    END
  END Data_PMOS[155]
  PIN Data_PMOS[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6211.865 1046.435 6212.145 1047.435 ;
    END
  END Data_PMOS[166]
  PIN Data_PMOS[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6209.625 1046.435 6209.905 1047.435 ;
    END
  END Data_PMOS[161]
  PIN INJ_IN[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6207.385 1046.435 6207.665 1047.435 ;
    END
  END INJ_IN[127]
  PIN BcidMtx[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6205.145 1046.435 6205.425 1047.435 ;
    END
  END BcidMtx[383]
  PIN Read_PMOS[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6202.905 1046.435 6203.185 1047.435 ;
    END
  END Read_PMOS[7]
  PIN BcidMtx[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6201.225 1046.435 6201.505 1047.435 ;
    END
  END BcidMtx[378]
  PIN Data_PMOS[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6190.025 1046.435 6190.305 1047.435 ;
    END
  END Data_PMOS[149]
  PIN Data_PMOS[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6188.345 1046.435 6188.625 1047.435 ;
    END
  END Data_PMOS[157]
  PIN Data_PMOS[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6186.665 1046.435 6186.945 1047.435 ;
    END
  END Data_PMOS[158]
  PIN Data_PMOS[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6184.985 1046.435 6185.265 1047.435 ;
    END
  END Data_PMOS[164]
  PIN INJ_IN[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18853.865 1046.435 18854.145 1047.435 ;
    END
  END INJ_IN[442]
  PIN DIG_MON_PMOS[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6180.225 1046.435 6180.505 1047.435 ;
    END
  END DIG_MON_PMOS[14]
  PIN DIG_MON_SEL[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6178.545 1046.435 6178.825 1047.435 ;
    END
  END DIG_MON_SEL[126]
  PIN DIG_MON_PMOS[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7269.705 1046.435 7269.985 1047.435 ;
    END
  END DIG_MON_PMOS[41]
  PIN Data_PMOS[438]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7267.465 1046.435 7267.745 1047.435 ;
    END
  END Data_PMOS[438]
  PIN Data_PMOS[432]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7266.345 1046.435 7266.625 1047.435 ;
    END
  END Data_PMOS[432]
  PIN Data_PMOS[440]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7264.105 1046.435 7264.385 1047.435 ;
    END
  END Data_PMOS[440]
  PIN Data_PMOS[426]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7262.425 1046.435 7262.705 1047.435 ;
    END
  END Data_PMOS[426]
  PIN BcidMtx[461]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7245.625 1046.435 7245.905 1047.435 ;
    END
  END BcidMtx[461]
  PIN FREEZE_PMOS[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7243.945 1046.435 7244.225 1047.435 ;
    END
  END FREEZE_PMOS[20]
  PIN BcidMtx[457]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7242.265 1046.435 7242.545 1047.435 ;
    END
  END BcidMtx[457]
  PIN INJ_IN[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7240.585 1046.435 7240.865 1047.435 ;
    END
  END INJ_IN[152]
  PIN Data_PMOS[435]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7237.785 1046.435 7238.065 1047.435 ;
    END
  END Data_PMOS[435]
  PIN Data_PMOS[436]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7236.105 1046.435 7236.385 1047.435 ;
    END
  END Data_PMOS[436]
  PIN Data_PMOS[421]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7234.985 1046.435 7235.265 1047.435 ;
    END
  END Data_PMOS[421]
  PIN MASKH[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7194.105 1046.435 7194.385 1047.435 ;
    END
  END MASKH[76]
  PIN MASKD[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7189.065 1046.435 7189.345 1047.435 ;
    END
  END MASKD[151]
  PIN MASKV[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7186.265 1046.435 7186.545 1047.435 ;
    END
  END MASKV[151]
  PIN Data_PMOS[411]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7184.585 1046.435 7184.865 1047.435 ;
    END
  END Data_PMOS[411]
  PIN Data_PMOS[404]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7183.465 1046.435 7183.745 1047.435 ;
    END
  END Data_PMOS[404]
  PIN Data_PMOS[406]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7181.225 1046.435 7181.505 1047.435 ;
    END
  END Data_PMOS[406]
  PIN nTOK_PMOS[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7170.025 1046.435 7170.305 1047.435 ;
    END
  END nTOK_PMOS[19]
  PIN BcidMtx[454]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7168.345 1046.435 7168.625 1047.435 ;
    END
  END BcidMtx[454]
  PIN BcidMtx[452]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7166.105 1046.435 7166.385 1047.435 ;
    END
  END BcidMtx[452]
  PIN INJ_IN[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7161.905 1046.435 7162.185 1047.435 ;
    END
  END INJ_IN[150]
  PIN Data_PMOS[401]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7160.225 1046.435 7160.505 1047.435 ;
    END
  END Data_PMOS[401]
  PIN Data_PMOS[403]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7132.505 1046.435 7132.785 1047.435 ;
    END
  END Data_PMOS[403]
  PIN Data_PMOS[410]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7131.385 1046.435 7131.665 1047.435 ;
    END
  END Data_PMOS[410]
  PIN Data_PMOS[416]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7129.705 1046.435 7129.985 1047.435 ;
    END
  END Data_PMOS[416]
  PIN MASKD[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7128.025 1046.435 7128.305 1047.435 ;
    END
  END MASKD[150]
  PIN DIG_MON_SEL[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7125.225 1046.435 7125.505 1047.435 ;
    END
  END DIG_MON_SEL[150]
  PIN Data_PMOS_NOSF[839]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4303.945 1046.435 4304.225 1047.435 ;
    END
  END Data_PMOS_NOSF[839]
  PIN nTOK_PMOS_NOSF[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4300.025 1046.435 4300.305 1047.435 ;
    END
  END nTOK_PMOS_NOSF[39]
  PIN BcidMtx[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4298.345 1046.435 4298.625 1047.435 ;
    END
  END BcidMtx[238]
  PIN FREEZE_PMOS_NOSF[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4297.225 1046.435 4297.505 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[39]
  PIN BcidMtx[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4294.985 1046.435 4295.265 1047.435 ;
    END
  END BcidMtx[234]
  PIN Data_PMOS_NOSF[822]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4254.105 1046.435 4254.385 1047.435 ;
    END
  END Data_PMOS_NOSF[822]
  PIN Data_PMOS_NOSF[828]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4252.985 1046.435 4253.265 1047.435 ;
    END
  END Data_PMOS_NOSF[828]
  PIN Data_PMOS_NOSF[830]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4250.185 1046.435 4250.465 1047.435 ;
    END
  END Data_PMOS_NOSF[830]
  PIN Data_PMOS_NOSF[819]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4249.065 1046.435 4249.345 1047.435 ;
    END
  END Data_PMOS_NOSF[819]
  PIN MASKV[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4247.945 1046.435 4248.225 1047.435 ;
    END
  END MASKV[78]
  PIN DIG_MON_SEL[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4244.025 1046.435 4244.305 1047.435 ;
    END
  END DIG_MON_SEL[78]
  PIN MASKD[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4242.345 1046.435 4242.625 1047.435 ;
    END
  END MASKD[77]
  PIN INJ_ROW[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4231.705 1046.435 4231.985 1047.435 ;
    END
  END INJ_ROW[38]
  PIN Data_PMOS_NOSF[810]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4229.465 1046.435 4229.745 1047.435 ;
    END
  END Data_PMOS_NOSF[810]
  PIN Data_PMOS_NOSF[811]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4227.785 1046.435 4228.065 1047.435 ;
    END
  END Data_PMOS_NOSF[811]
  PIN Data_PMOS_NOSF[812]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4226.665 1046.435 4226.945 1047.435 ;
    END
  END Data_PMOS_NOSF[812]
  PIN nTOK_PMOS_NOSF[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4221.345 1046.435 4221.625 1047.435 ;
    END
  END nTOK_PMOS_NOSF[38]
  PIN BcidMtx[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4219.105 1046.435 4219.385 1047.435 ;
    END
  END BcidMtx[231]
  PIN BcidMtx[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4191.945 1046.435 4192.225 1047.435 ;
    END
  END BcidMtx[230]
  PIN Data_PMOS_NOSF[801]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4188.585 1046.435 4188.865 1047.435 ;
    END
  END Data_PMOS_NOSF[801]
  PIN Data_PMOS_NOSF[813]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4186.905 1046.435 4187.185 1047.435 ;
    END
  END Data_PMOS_NOSF[813]
  PIN Data_PMOS_NOSF[802]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4185.785 1046.435 4186.065 1047.435 ;
    END
  END Data_PMOS_NOSF[802]
  PIN Data_PMOS_NOSF[798]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4183.545 1046.435 4183.825 1047.435 ;
    END
  END Data_PMOS_NOSF[798]
  PIN MASKH[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4181.865 1046.435 4182.145 1047.435 ;
    END
  END MASKH[38]
  PIN DIG_MON_PMOS_NOSF[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4180.185 1046.435 4180.465 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[76]
  PIN DIG_MON_SEL[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4165.065 1046.435 4165.345 1047.435 ;
    END
  END DIG_MON_SEL[75]
  PIN INJ_ROW[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4161.705 1046.435 4161.985 1047.435 ;
    END
  END INJ_ROW[37]
  PIN Data_PMOS_NOSF[795]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4160.585 1046.435 4160.865 1047.435 ;
    END
  END Data_PMOS_NOSF[795]
  PIN Data_PMOS_NOSF[782]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4158.345 1046.435 4158.625 1047.435 ;
    END
  END Data_PMOS_NOSF[782]
  PIN Data_PMOS_NOSF[791]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4156.665 1046.435 4156.945 1047.435 ;
    END
  END Data_PMOS_NOSF[791]
  PIN Data_PMOS_NOSF[783]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4155.545 1046.435 4155.825 1047.435 ;
    END
  END Data_PMOS_NOSF[783]
  PIN BcidMtx[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4112.425 1046.435 4112.705 1047.435 ;
    END
  END BcidMtx[226]
  PIN Read_PMOS_NOSF[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4110.745 1046.435 4111.025 1047.435 ;
    END
  END Read_PMOS_NOSF[37]
  PIN BcidMtx[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4109.625 1046.435 4109.905 1047.435 ;
    END
  END BcidMtx[223]
  PIN Data_PMOS_NOSF[779]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4106.265 1046.435 4106.545 1047.435 ;
    END
  END Data_PMOS_NOSF[779]
  PIN Data_PMOS_NOSF[787]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4104.585 1046.435 4104.865 1047.435 ;
    END
  END Data_PMOS_NOSF[787]
  PIN Data_PMOS_NOSF[793]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4103.465 1046.435 4103.745 1047.435 ;
    END
  END Data_PMOS_NOSF[793]
  PIN Data_PMOS_NOSF[794]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4101.225 1046.435 4101.505 1047.435 ;
    END
  END Data_PMOS_NOSF[794]
  PIN MASKD[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4091.145 1046.435 4091.425 1047.435 ;
    END
  END MASKD[74]
  PIN INJ_ROW[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4082.465 1046.435 4082.745 1047.435 ;
    END
  END INJ_ROW[36]
  PIN Data_PMOS_NOSF[764]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4080.785 1046.435 4081.065 1047.435 ;
    END
  END Data_PMOS_NOSF[764]
  PIN Data_PMOS_NOSF[775]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4079.665 1046.435 4079.945 1047.435 ;
    END
  END Data_PMOS_NOSF[775]
  PIN Data_PMOS_NOSF[770]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4051.945 1046.435 4052.225 1047.435 ;
    END
  END Data_PMOS_NOSF[770]
  PIN INJ_IN[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4049.705 1046.435 4049.985 1047.435 ;
    END
  END INJ_IN[73]
  PIN BcidMtx[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4047.465 1046.435 4047.745 1047.435 ;
    END
  END BcidMtx[221]
  PIN Read_PMOS_NOSF[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4045.225 1046.435 4045.505 1047.435 ;
    END
  END Read_PMOS_NOSF[36]
  PIN BcidMtx[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4043.545 1046.435 4043.825 1047.435 ;
    END
  END BcidMtx[216]
  PIN Data_PMOS_NOSF[759]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4041.305 1046.435 4041.585 1047.435 ;
    END
  END Data_PMOS_NOSF[759]
  PIN Data_PMOS_NOSF[766]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4026.185 1046.435 4026.465 1047.435 ;
    END
  END Data_PMOS_NOSF[766]
  PIN Data_PMOS_NOSF[767]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4024.505 1046.435 4024.785 1047.435 ;
    END
  END Data_PMOS_NOSF[767]
  PIN Data_PMOS_NOSF[756]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4023.385 1046.435 4023.665 1047.435 ;
    END
  END Data_PMOS_NOSF[756]
  PIN MASKD[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4021.145 1046.435 4021.425 1047.435 ;
    END
  END MASKD[72]
  PIN DIG_MON_SEL[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4018.345 1046.435 4018.625 1047.435 ;
    END
  END DIG_MON_SEL[72]
  PIN MASKD[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4016.665 1046.435 4016.945 1047.435 ;
    END
  END MASKD[71]
  PIN Data_PMOS_NOSF[753]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3973.545 1046.435 3973.825 1047.435 ;
    END
  END Data_PMOS_NOSF[753]
  PIN Data_PMOS_NOSF[754]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3971.865 1046.435 3972.145 1047.435 ;
    END
  END Data_PMOS_NOSF[754]
  PIN Data_PMOS_NOSF[748]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3970.745 1046.435 3971.025 1047.435 ;
    END
  END Data_PMOS_NOSF[748]
  PIN Data_PMOS_NOSF[749]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3969.625 1046.435 3969.905 1047.435 ;
    END
  END Data_PMOS_NOSF[749]
  PIN Data_HV[1132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18865.625 1046.435 18865.905 1047.435 ;
    END
  END Data_HV[1132]
  PIN nTOK_PMOS_NOSF[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3966.265 1046.435 3966.545 1047.435 ;
    END
  END nTOK_PMOS_NOSF[35]
  PIN FREEZE_PMOS_NOSF[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3963.465 1046.435 3963.745 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[35]
  PIN BcidMtx[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3961.785 1046.435 3962.065 1047.435 ;
    END
  END BcidMtx[211]
  PIN BcidMtx[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3961.225 1046.435 3961.505 1047.435 ;
    END
  END BcidMtx[210]
  PIN Data_PMOS_NOSF[750]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3948.905 1046.435 3949.185 1047.435 ;
    END
  END Data_PMOS_NOSF[750]
  PIN Data_PMOS_NOSF[751]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3947.225 1046.435 3947.505 1047.435 ;
    END
  END Data_PMOS_NOSF[751]
  PIN Data_PMOS_NOSF[736]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3946.105 1046.435 3946.385 1047.435 ;
    END
  END Data_PMOS_NOSF[736]
  PIN MASKH[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3941.905 1046.435 3942.185 1047.435 ;
    END
  END MASKH[35]
  PIN FREEZE_PMOS_NOSF[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4193.065 1046.435 4193.345 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[38]
  PIN INJ_ROW[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5028.585 1046.435 5028.865 1047.435 ;
    END
  END INJ_ROW[48]
  PIN Data_PMOS_NOSF[1016]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5026.905 1046.435 5027.185 1047.435 ;
    END
  END Data_PMOS_NOSF[1016]
  PIN Data_PMOS_NOSF[1027]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5025.785 1046.435 5026.065 1047.435 ;
    END
  END Data_PMOS_NOSF[1027]
  PIN Data_PMOS_NOSF[1028]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5024.105 1046.435 5024.385 1047.435 ;
    END
  END Data_PMOS_NOSF[1028]
  PIN Data_PMOS_NOSF[1014]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5022.425 1046.435 5022.705 1047.435 ;
    END
  END Data_PMOS_NOSF[1014]
  PIN Data_HV[1118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18865.065 1046.435 18865.345 1047.435 ;
    END
  END Data_HV[1118]
  PIN BcidMtx[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5005.065 1046.435 5005.345 1047.435 ;
    END
  END BcidMtx[292]
  PIN Read_PMOS_NOSF[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5003.385 1046.435 5003.665 1047.435 ;
    END
  END Read_PMOS_NOSF[48]
  PIN BcidMtx[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5002.265 1046.435 5002.545 1047.435 ;
    END
  END BcidMtx[289]
  PIN Data_PMOS_NOSF[1010]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4998.905 1046.435 4999.185 1047.435 ;
    END
  END Data_PMOS_NOSF[1010]
  PIN Data_PMOS_NOSF[1018]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4997.225 1046.435 4997.505 1047.435 ;
    END
  END Data_PMOS_NOSF[1018]
  PIN Data_PMOS_NOSF[1024]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4996.105 1046.435 4996.385 1047.435 ;
    END
  END Data_PMOS_NOSF[1024]
  PIN Data_PMOS_NOSF[1025]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4993.865 1046.435 4994.145 1047.435 ;
    END
  END Data_PMOS_NOSF[1025]
  PIN MASKD[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4953.545 1046.435 4953.825 1047.435 ;
    END
  END MASKD[96]
  PIN DIG_MON_PMOS_NOSF[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4947.945 1046.435 4948.225 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[95]
  PIN MASKV[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4946.265 1046.435 4946.545 1047.435 ;
    END
  END MASKV[95]
  PIN Data_PMOS_NOSF[995]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4945.145 1046.435 4945.425 1047.435 ;
    END
  END Data_PMOS_NOSF[995]
  PIN Data_PMOS_NOSF[1000]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4942.905 1046.435 4943.185 1047.435 ;
    END
  END Data_PMOS_NOSF[1000]
  PIN Data_HV[1126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18864.505 1046.435 18864.785 1047.435 ;
    END
  END Data_HV[1126]
  PIN Data_PMOS_NOSF[993]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4932.265 1046.435 4932.545 1047.435 ;
    END
  END Data_PMOS_NOSF[993]
  PIN BcidMtx[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4928.345 1046.435 4928.625 1047.435 ;
    END
  END BcidMtx[286]
  PIN Read_PMOS_NOSF[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4926.665 1046.435 4926.945 1047.435 ;
    END
  END Read_PMOS_NOSF[47]
  PIN BcidMtx[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4925.545 1046.435 4925.825 1047.435 ;
    END
  END BcidMtx[283]
  PIN Data_PMOS_NOSF[989]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4920.225 1046.435 4920.505 1047.435 ;
    END
  END Data_PMOS_NOSF[989]
  PIN Data_PMOS_NOSF[997]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4918.545 1046.435 4918.825 1047.435 ;
    END
  END Data_PMOS_NOSF[997]
  PIN Data_PMOS_NOSF[1003]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4891.945 1046.435 4892.225 1047.435 ;
    END
  END Data_PMOS_NOSF[1003]
  PIN Data_PMOS_NOSF[1004]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4889.705 1046.435 4889.985 1047.435 ;
    END
  END Data_PMOS_NOSF[1004]
  PIN MASKD[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4888.025 1046.435 4888.305 1047.435 ;
    END
  END MASKD[94]
  PIN DIG_MON_PMOS_NOSF[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4882.425 1046.435 4882.705 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[93]
  PIN Data_PMOS_NOSF[984]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4880.185 1046.435 4880.465 1047.435 ;
    END
  END Data_PMOS_NOSF[984]
  PIN INJ_IN[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18861.145 1046.435 18861.425 1047.435 ;
    END
  END INJ_IN[443]
  PIN Data_PMOS_NOSF[1127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5423.385 1046.435 5423.665 1047.435 ;
    END
  END Data_PMOS_NOSF[1127]
  PIN Data_PMOS_NOSF[1119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5422.265 1046.435 5422.545 1047.435 ;
    END
  END Data_PMOS_NOSF[1119]
  PIN BcidMtx[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5418.345 1046.435 5418.625 1047.435 ;
    END
  END BcidMtx[322]
  PIN Read_PMOS_NOSF[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5416.665 1046.435 5416.945 1047.435 ;
    END
  END Read_PMOS_NOSF[53]
  PIN BcidMtx[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5415.545 1046.435 5415.825 1047.435 ;
    END
  END BcidMtx[319]
  PIN Data_PMOS_NOSF[1115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5373.545 1046.435 5373.825 1047.435 ;
    END
  END Data_PMOS_NOSF[1115]
  PIN Data_PMOS_NOSF[1123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5371.865 1046.435 5372.145 1047.435 ;
    END
  END Data_PMOS_NOSF[1123]
  PIN Data_PMOS_NOSF[1129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5370.745 1046.435 5371.025 1047.435 ;
    END
  END Data_PMOS_NOSF[1129]
  PIN Data_PMOS_NOSF[1130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5368.505 1046.435 5368.785 1047.435 ;
    END
  END Data_PMOS_NOSF[1130]
  PIN MASKD[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5366.825 1046.435 5367.105 1047.435 ;
    END
  END MASKD[106]
  PIN DIG_MON_PMOS_NOSF[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5361.225 1046.435 5361.505 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[105]
  PIN Data_PMOS_NOSF[1110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5350.585 1046.435 5350.865 1047.435 ;
    END
  END Data_PMOS_NOSF[1110]
  PIN Data_PMOS_NOSF[1104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5349.465 1046.435 5349.745 1047.435 ;
    END
  END Data_PMOS_NOSF[1104]
  PIN Data_PMOS_NOSF[1112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5347.225 1046.435 5347.505 1047.435 ;
    END
  END Data_PMOS_NOSF[1112]
  PIN Data_PMOS_NOSF[1098]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5345.545 1046.435 5345.825 1047.435 ;
    END
  END Data_PMOS_NOSF[1098]
  PIN nTOK_PMOS_NOSF[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5341.345 1046.435 5341.625 1047.435 ;
    END
  END nTOK_PMOS_NOSF[52]
  PIN Read_PMOS_NOSF[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5312.505 1046.435 5312.785 1047.435 ;
    END
  END Read_PMOS_NOSF[52]
  PIN BcidMtx[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5310.825 1046.435 5311.105 1047.435 ;
    END
  END BcidMtx[312]
  PIN Data_PMOS_NOSF[1095]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5308.585 1046.435 5308.865 1047.435 ;
    END
  END Data_PMOS_NOSF[1095]
  PIN Data_PMOS_NOSF[1102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5306.345 1046.435 5306.625 1047.435 ;
    END
  END Data_PMOS_NOSF[1102]
  PIN Data_PMOS_NOSF[1103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5304.665 1046.435 5304.945 1047.435 ;
    END
  END Data_PMOS_NOSF[1103]
  PIN Data_PMOS_NOSF[1092]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5303.545 1046.435 5303.825 1047.435 ;
    END
  END Data_PMOS_NOSF[1092]
  PIN MASKD[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5301.305 1046.435 5301.585 1047.435 ;
    END
  END MASKD[104]
  PIN DIG_MON_SEL[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5285.625 1046.435 5285.905 1047.435 ;
    END
  END DIG_MON_SEL[104]
  PIN MASKD[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5283.945 1046.435 5284.225 1047.435 ;
    END
  END MASKD[103]
  PIN Data_PMOS_NOSF[1089]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5280.585 1046.435 5280.865 1047.435 ;
    END
  END Data_PMOS_NOSF[1089]
  PIN Data_PMOS_NOSF[1090]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5278.905 1046.435 5279.185 1047.435 ;
    END
  END Data_PMOS_NOSF[1090]
  PIN Data_PMOS_NOSF[1084]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5277.785 1046.435 5278.065 1047.435 ;
    END
  END Data_PMOS_NOSF[1084]
  PIN Data_PMOS_NOSF[1077]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5275.545 1046.435 5275.825 1047.435 ;
    END
  END Data_PMOS_NOSF[1077]
  PIN BcidMtx[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5232.985 1046.435 5233.265 1047.435 ;
    END
  END BcidMtx[311]
  PIN FREEZE_PMOS_NOSF[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5231.305 1046.435 5231.585 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[51]
  PIN BcidMtx[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5229.065 1046.435 5229.345 1047.435 ;
    END
  END BcidMtx[306]
  PIN Data_PMOS_NOSF[1073]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5226.265 1046.435 5226.545 1047.435 ;
    END
  END Data_PMOS_NOSF[1073]
  PIN Data_PMOS_NOSF[1081]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5224.585 1046.435 5224.865 1047.435 ;
    END
  END Data_PMOS_NOSF[1081]
  PIN Data_PMOS_NOSF[1082]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5222.905 1046.435 5223.185 1047.435 ;
    END
  END Data_PMOS_NOSF[1082]
  PIN Data_PMOS_NOSF[1088]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5221.225 1046.435 5221.505 1047.435 ;
    END
  END Data_PMOS_NOSF[1088]
  PIN MASKD[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5211.145 1046.435 5211.425 1047.435 ;
    END
  END MASKD[102]
  PIN Data_HV[1127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18863.385 1046.435 18863.665 1047.435 ;
    END
  END Data_HV[1127]
  PIN DIG_MON_SEL[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5208.345 1046.435 5208.625 1047.435 ;
    END
  END DIG_MON_SEL[102]
  PIN DIG_MON_PMOS_NOSF[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5205.545 1046.435 5205.825 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[101]
  PIN Data_PMOS_NOSF[1068]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5201.345 1046.435 5201.625 1047.435 ;
    END
  END Data_PMOS_NOSF[1068]
  PIN Data_PMOS_NOSF[1069]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5199.665 1046.435 5199.945 1047.435 ;
    END
  END Data_PMOS_NOSF[1069]
  PIN Data_PMOS_NOSF[1070]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5172.505 1046.435 5172.785 1047.435 ;
    END
  END Data_PMOS_NOSF[1070]
  PIN Data_PMOS_NOSF[1056]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5170.825 1046.435 5171.105 1047.435 ;
    END
  END Data_PMOS_NOSF[1056]
  PIN BcidMtx[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5167.465 1046.435 5167.745 1047.435 ;
    END
  END BcidMtx[305]
  PIN FREEZE_PMOS_NOSF[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5165.785 1046.435 5166.065 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[50]
  PIN BcidMtx[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5164.105 1046.435 5164.385 1047.435 ;
    END
  END BcidMtx[301]
  PIN Data_PMOS_NOSF[1053]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5161.305 1046.435 5161.585 1047.435 ;
    END
  END Data_PMOS_NOSF[1053]
  PIN Data_PMOS_NOSF[1065]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5146.745 1046.435 5147.025 1047.435 ;
    END
  END Data_PMOS_NOSF[1065]
  PIN Data_PMOS_NOSF[1066]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5145.065 1046.435 5145.345 1047.435 ;
    END
  END Data_PMOS_NOSF[1066]
  PIN Data_PMOS_NOSF[1050]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5143.385 1046.435 5143.665 1047.435 ;
    END
  END Data_PMOS_NOSF[1050]
  PIN MASKH[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5141.705 1046.435 5141.985 1047.435 ;
    END
  END MASKH[50]
  PIN MASKD[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5136.665 1046.435 5136.945 1047.435 ;
    END
  END MASKD[99]
  PIN DIG_MON_PMOS_NOSF[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5135.545 1046.435 5135.825 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[99]
  PIN Data_PMOS_NOSF[1047]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5093.545 1046.435 5093.825 1047.435 ;
    END
  END Data_PMOS_NOSF[1047]
  PIN Data_PMOS_NOSF[1048]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5091.865 1046.435 5092.145 1047.435 ;
    END
  END Data_PMOS_NOSF[1048]
  PIN Data_PMOS_NOSF[1049]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5090.185 1046.435 5090.465 1047.435 ;
    END
  END Data_PMOS_NOSF[1049]
  PIN Data_PMOS_NOSF[1036]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5089.065 1046.435 5089.345 1047.435 ;
    END
  END Data_PMOS_NOSF[1036]
  PIN BcidMtx[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5085.145 1046.435 5085.425 1047.435 ;
    END
  END BcidMtx[299]
  PIN FREEZE_PMOS_NOSF[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5083.465 1046.435 5083.745 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[49]
  PIN BcidMtx[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5082.345 1046.435 5082.625 1047.435 ;
    END
  END BcidMtx[296]
  PIN BcidMtx[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5081.225 1046.435 5081.505 1047.435 ;
    END
  END BcidMtx[294]
  PIN Data_PMOS_NOSF[1031]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5070.025 1046.435 5070.305 1047.435 ;
    END
  END Data_PMOS_NOSF[1031]
  PIN Data_PMOS_NOSF[1045]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5067.225 1046.435 5067.505 1047.435 ;
    END
  END Data_PMOS_NOSF[1045]
  PIN Data_PMOS_NOSF[1040]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5066.665 1046.435 5066.945 1047.435 ;
    END
  END Data_PMOS_NOSF[1040]
  PIN Data_PMOS_NOSF[1046]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5064.985 1046.435 5065.265 1047.435 ;
    END
  END Data_PMOS_NOSF[1046]
  PIN DIG_MON_SEL[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5058.545 1046.435 5058.825 1047.435 ;
    END
  END DIG_MON_SEL[98]
  PIN MASKD[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6150.825 1046.435 6151.105 1047.435 ;
    END
  END MASKD[125]
  PIN Data_PMOS[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6146.905 1046.435 6147.185 1047.435 ;
    END
  END Data_PMOS[134]
  PIN Data_PMOS[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6146.345 1046.435 6146.625 1047.435 ;
    END
  END Data_PMOS[138]
  PIN Data_PMOS[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6144.665 1046.435 6144.945 1047.435 ;
    END
  END Data_PMOS[139]
  PIN INJ_IN[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6141.305 1046.435 6141.585 1047.435 ;
    END
  END INJ_IN[125]
  PIN nTOK_PMOS[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6140.185 1046.435 6140.465 1047.435 ;
    END
  END nTOK_PMOS[6]
  PIN BcidMtx[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6124.505 1046.435 6124.785 1047.435 ;
    END
  END BcidMtx[375]
  PIN BcidMtx[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6121.705 1046.435 6121.985 1047.435 ;
    END
  END BcidMtx[372]
  PIN INJ_IN[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6120.585 1046.435 6120.865 1047.435 ;
    END
  END INJ_IN[124]
  PIN Data_PMOS[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6118.345 1046.435 6118.625 1047.435 ;
    END
  END Data_PMOS[135]
  PIN Data_PMOS[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6115.545 1046.435 6115.825 1047.435 ;
    END
  END Data_PMOS[137]
  PIN Data_PMOS[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6114.425 1046.435 6114.705 1047.435 ;
    END
  END Data_PMOS[126]
  PIN MASKV[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6074.665 1046.435 6074.945 1047.435 ;
    END
  END MASKV[124]
  PIN DIG_MON_SEL[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6070.185 1046.435 6070.465 1047.435 ;
    END
  END DIG_MON_SEL[123]
  PIN INJ_ROW[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6066.825 1046.435 6067.105 1047.435 ;
    END
  END INJ_ROW[61]
  PIN Data_PMOS[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6064.585 1046.435 6064.865 1047.435 ;
    END
  END Data_PMOS[117]
  PIN Data_PMOS[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6063.465 1046.435 6063.745 1047.435 ;
    END
  END Data_PMOS[110]
  PIN Data_PMOS[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6061.785 1046.435 6062.065 1047.435 ;
    END
  END Data_PMOS[119]
  PIN nTOK_PMOS[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6050.025 1046.435 6050.305 1047.435 ;
    END
  END nTOK_PMOS[5]
  PIN BcidMtx[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6048.345 1046.435 6048.625 1047.435 ;
    END
  END BcidMtx[370]
  PIN Read_PMOS[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6046.665 1046.435 6046.945 1047.435 ;
    END
  END Read_PMOS[5]
  PIN INJ_IN[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6041.905 1046.435 6042.185 1047.435 ;
    END
  END INJ_IN[122]
  PIN Data_PMOS[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6040.225 1046.435 6040.505 1047.435 ;
    END
  END Data_PMOS[107]
  PIN Data_PMOS[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6038.545 1046.435 6038.825 1047.435 ;
    END
  END Data_PMOS[115]
  PIN Data_PMOS[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6010.825 1046.435 6011.105 1047.435 ;
    END
  END Data_PMOS[106]
  PIN Data_PMOS[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6009.705 1046.435 6009.985 1047.435 ;
    END
  END Data_PMOS[122]
  PIN MASKD[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6008.025 1046.435 6008.305 1047.435 ;
    END
  END MASKD[122]
  PIN DIG_MON_SEL[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6004.665 1046.435 6004.945 1047.435 ;
    END
  END DIG_MON_SEL[121]
  PIN DIG_MON_PMOS[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6002.425 1046.435 6002.705 1047.435 ;
    END
  END DIG_MON_PMOS[9]
  PIN MASKV[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6000.745 1046.435 6001.025 1047.435 ;
    END
  END MASKV[121]
  PIN Data_PMOS_NOSF[978]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4866.185 1046.435 4866.465 1047.435 ;
    END
  END Data_PMOS_NOSF[978]
  PIN Data_PMOS_NOSF[986]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4863.945 1046.435 4864.225 1047.435 ;
    END
  END Data_PMOS_NOSF[986]
  PIN Data_PMOS_NOSF[972]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4862.265 1046.435 4862.545 1047.435 ;
    END
  END Data_PMOS_NOSF[972]
  PIN nTOK_PMOS_NOSF[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4860.025 1046.435 4860.305 1047.435 ;
    END
  END nTOK_PMOS_NOSF[46]
  PIN FREEZE_PMOS_NOSF[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4857.225 1046.435 4857.505 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[46]
  PIN BcidMtx[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4855.545 1046.435 4855.825 1047.435 ;
    END
  END BcidMtx[277]
  PIN INJ_IN[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4853.865 1046.435 4854.145 1047.435 ;
    END
  END INJ_IN[92]
  PIN Data_PMOS_NOSF[981]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4812.425 1046.435 4812.705 1047.435 ;
    END
  END Data_PMOS_NOSF[981]
  PIN Data_PMOS_NOSF[982]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4810.745 1046.435 4811.025 1047.435 ;
    END
  END Data_PMOS_NOSF[982]
  PIN Data_PMOS_NOSF[967]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4809.625 1046.435 4809.905 1047.435 ;
    END
  END Data_PMOS_NOSF[967]
  PIN MASKV[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4807.945 1046.435 4808.225 1047.435 ;
    END
  END MASKV[92]
  PIN INJ_ROW[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4791.705 1046.435 4791.985 1047.435 ;
    END
  END INJ_ROW[45]
  PIN Data_PMOS_NOSF[953]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4790.025 1046.435 4790.305 1047.435 ;
    END
  END Data_PMOS_NOSF[953]
  PIN Data_PMOS_NOSF[964]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4788.905 1046.435 4789.185 1047.435 ;
    END
  END Data_PMOS_NOSF[964]
  PIN Data_PMOS_NOSF[959]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4786.665 1046.435 4786.945 1047.435 ;
    END
  END Data_PMOS_NOSF[959]
  PIN INJ_IN[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4782.465 1046.435 4782.745 1047.435 ;
    END
  END INJ_IN[91]
  PIN BcidMtx[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4780.225 1046.435 4780.505 1047.435 ;
    END
  END BcidMtx[275]
  PIN BcidMtx[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4751.945 1046.435 4752.225 1047.435 ;
    END
  END BcidMtx[272]
  PIN INJ_IN[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4749.705 1046.435 4749.985 1047.435 ;
    END
  END INJ_IN[90]
  PIN Data_PMOS_NOSF[947]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4748.025 1046.435 4748.305 1047.435 ;
    END
  END Data_PMOS_NOSF[947]
  PIN Data_PMOS_NOSF[949]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4745.785 1046.435 4746.065 1047.435 ;
    END
  END Data_PMOS_NOSF[949]
  PIN Data_PMOS_NOSF[946]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4744.105 1046.435 4744.385 1047.435 ;
    END
  END Data_PMOS_NOSF[946]
  PIN Data_PMOS_NOSF[962]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4742.985 1046.435 4743.265 1047.435 ;
    END
  END Data_PMOS_NOSF[962]
  PIN DIG_MON_PMOS_NOSF[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4740.185 1046.435 4740.465 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[90]
  PIN DIG_MON_SEL[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4725.065 1046.435 4725.345 1047.435 ;
    END
  END DIG_MON_SEL[89]
  PIN DIG_MON_PMOS_NOSF[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4722.825 1046.435 4723.105 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[89]
  PIN Data_PMOS_NOSF[932]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4720.025 1046.435 4720.305 1047.435 ;
    END
  END Data_PMOS_NOSF[932]
  PIN Data_PMOS_NOSF[929]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4718.345 1046.435 4718.625 1047.435 ;
    END
  END Data_PMOS_NOSF[929]
  PIN Data_PMOS_NOSF[944]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4717.225 1046.435 4717.505 1047.435 ;
    END
  END Data_PMOS_NOSF[944]
  PIN INJ_IN[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4714.425 1046.435 4714.705 1047.435 ;
    END
  END INJ_IN[89]
  PIN BcidMtx[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4672.425 1046.435 4672.705 1047.435 ;
    END
  END BcidMtx[268]
  PIN FREEZE_PMOS_NOSF[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4671.305 1046.435 4671.585 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[44]
  PIN BcidMtx[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4669.065 1046.435 4669.345 1047.435 ;
    END
  END BcidMtx[264]
  PIN Data_PMOS_NOSF[926]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4666.265 1046.435 4666.545 1047.435 ;
    END
  END Data_PMOS_NOSF[926]
  PIN Data_PMOS_NOSF[939]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4665.145 1046.435 4665.425 1047.435 ;
    END
  END Data_PMOS_NOSF[939]
  PIN Data_PMOS_NOSF[935]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4662.905 1046.435 4663.185 1047.435 ;
    END
  END Data_PMOS_NOSF[935]
  PIN Data_PMOS_NOSF[941]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4661.225 1046.435 4661.505 1047.435 ;
    END
  END Data_PMOS_NOSF[941]
  PIN MASKH[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4651.705 1046.435 4651.985 1047.435 ;
    END
  END MASKH[44]
  PIN DIG_MON_SEL[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4648.345 1046.435 4648.625 1047.435 ;
    END
  END DIG_MON_SEL[88]
  PIN DIG_MON_PMOS_NOSF[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4645.545 1046.435 4645.825 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[87]
  PIN MASKV[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4641.905 1046.435 4642.185 1047.435 ;
    END
  END MASKV[87]
  PIN Data_PMOS_NOSF[922]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4639.665 1046.435 4639.945 1047.435 ;
    END
  END Data_PMOS_NOSF[922]
  PIN Data_PMOS_NOSF[923]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4612.505 1046.435 4612.785 1047.435 ;
    END
  END Data_PMOS_NOSF[923]
  PIN Data_PMOS_NOSF[910]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4611.385 1046.435 4611.665 1047.435 ;
    END
  END Data_PMOS_NOSF[910]
  PIN BcidMtx[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4607.465 1046.435 4607.745 1047.435 ;
    END
  END BcidMtx[263]
  PIN FREEZE_PMOS_NOSF[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4605.785 1046.435 4606.065 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[43]
  PIN BcidMtx[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4604.665 1046.435 4604.945 1047.435 ;
    END
  END BcidMtx[260]
  PIN Data_PMOS_NOSF[906]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4601.305 1046.435 4601.585 1047.435 ;
    END
  END Data_PMOS_NOSF[906]
  PIN Data_PMOS_NOSF[918]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4586.745 1046.435 4587.025 1047.435 ;
    END
  END Data_PMOS_NOSF[918]
  PIN Data_PMOS_NOSF[907]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4585.625 1046.435 4585.905 1047.435 ;
    END
  END Data_PMOS_NOSF[907]
  PIN Data_PMOS_NOSF[903]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4583.385 1046.435 4583.665 1047.435 ;
    END
  END Data_PMOS_NOSF[903]
  PIN MASKH[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4581.705 1046.435 4581.985 1047.435 ;
    END
  END MASKH[43]
  PIN DIG_MON_PMOS_NOSF[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4580.025 1046.435 4580.305 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[86]
  PIN MASKD[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4576.665 1046.435 4576.945 1047.435 ;
    END
  END MASKD[85]
  PIN MASKV[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4573.865 1046.435 4574.145 1047.435 ;
    END
  END MASKV[85]
  PIN Data_PMOS_NOSF[900]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4533.545 1046.435 4533.825 1047.435 ;
    END
  END Data_PMOS_NOSF[900]
  PIN Data_HV[1120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18862.825 1046.435 18863.105 1047.435 ;
    END
  END Data_HV[1120]
  PIN Data_PMOS_NOSF[902]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4530.185 1046.435 4530.465 1047.435 ;
    END
  END Data_PMOS_NOSF[902]
  PIN Data_PMOS_NOSF[889]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4529.065 1046.435 4529.345 1047.435 ;
    END
  END Data_PMOS_NOSF[889]
  PIN BcidMtx[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4525.145 1046.435 4525.425 1047.435 ;
    END
  END BcidMtx[257]
  PIN BcidMtx[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4524.025 1046.435 4524.305 1047.435 ;
    END
  END BcidMtx[255]
  PIN Read_PMOS_NOSF[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4522.905 1046.435 4523.185 1047.435 ;
    END
  END Read_PMOS_NOSF[42]
  PIN INJ_IN[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4511.705 1046.435 4511.985 1047.435 ;
    END
  END INJ_IN[84]
  PIN Data_PMOS_NOSF[891]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4509.465 1046.435 4509.745 1047.435 ;
    END
  END Data_PMOS_NOSF[891]
  PIN Data_PMOS_NOSF[892]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4508.345 1046.435 4508.625 1047.435 ;
    END
  END Data_PMOS_NOSF[892]
  PIN Data_PMOS_NOSF[883]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4506.105 1046.435 4506.385 1047.435 ;
    END
  END Data_PMOS_NOSF[883]
  PIN MASKV[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4502.465 1046.435 4502.745 1047.435 ;
    END
  END MASKV[84]
  PIN MASKD[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4501.345 1046.435 4501.625 1047.435 ;
    END
  END MASKD[84]
  PIN FREEZE_PMOS_NOSF[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4753.065 1046.435 4753.345 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[45]
  PIN DIG_MON_PMOS_NOSF[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5589.705 1046.435 5589.985 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[111]
  PIN MASKV[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5588.025 1046.435 5588.305 1047.435 ;
    END
  END MASKV[111]
  PIN Data_PMOS_NOSF[1174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5585.785 1046.435 5586.065 1047.435 ;
    END
  END Data_PMOS_NOSF[1174]
  PIN Data_PMOS_NOSF[1168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5584.665 1046.435 5584.945 1047.435 ;
    END
  END Data_PMOS_NOSF[1168]
  PIN Data_PMOS_NOSF[1169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5583.545 1046.435 5583.825 1047.435 ;
    END
  END Data_PMOS_NOSF[1169]
  PIN nTOK_PMOS_NOSF[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5580.185 1046.435 5580.465 1047.435 ;
    END
  END nTOK_PMOS_NOSF[55]
  PIN BcidMtx[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5564.505 1046.435 5564.785 1047.435 ;
    END
  END BcidMtx[333]
  PIN Read_PMOS_NOSF[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5563.385 1046.435 5563.665 1047.435 ;
    END
  END Read_PMOS_NOSF[55]
  PIN INJ_IN[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5560.585 1046.435 5560.865 1047.435 ;
    END
  END INJ_IN[110]
  PIN Data_PMOS_NOSF[1164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5558.345 1046.435 5558.625 1047.435 ;
    END
  END Data_PMOS_NOSF[1164]
  PIN Data_PMOS_NOSF[1165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5557.225 1046.435 5557.505 1047.435 ;
    END
  END Data_PMOS_NOSF[1165]
  PIN Data_PMOS_NOSF[1156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5554.985 1046.435 5555.265 1047.435 ;
    END
  END Data_PMOS_NOSF[1156]
  PIN MASKV[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5514.665 1046.435 5514.945 1047.435 ;
    END
  END MASKV[110]
  PIN MASKD[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5513.545 1046.435 5513.825 1047.435 ;
    END
  END MASKD[110]
  PIN DIG_MON_SEL[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5510.185 1046.435 5510.465 1047.435 ;
    END
  END DIG_MON_SEL[109]
  PIN INJ_ROW[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5506.825 1046.435 5507.105 1047.435 ;
    END
  END INJ_ROW[54]
  PIN Data_PMOS_NOSF[1152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5505.705 1046.435 5505.985 1047.435 ;
    END
  END Data_PMOS_NOSF[1152]
  PIN Data_PMOS_NOSF[1139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5503.465 1046.435 5503.745 1047.435 ;
    END
  END Data_PMOS_NOSF[1139]
  PIN Data_PMOS_NOSF[1148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5501.785 1046.435 5502.065 1047.435 ;
    END
  END Data_PMOS_NOSF[1148]
  PIN Data_PMOS_NOSF[1140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5492.265 1046.435 5492.545 1047.435 ;
    END
  END Data_PMOS_NOSF[1140]
  PIN BcidMtx[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5488.345 1046.435 5488.625 1047.435 ;
    END
  END BcidMtx[328]
  PIN Read_PMOS_NOSF[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5486.665 1046.435 5486.945 1047.435 ;
    END
  END Read_PMOS_NOSF[54]
  PIN BcidMtx[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5485.545 1046.435 5485.825 1047.435 ;
    END
  END BcidMtx[325]
  PIN Data_PMOS_NOSF[1136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5480.225 1046.435 5480.505 1047.435 ;
    END
  END Data_PMOS_NOSF[1136]
  PIN Data_PMOS_NOSF[1144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5478.545 1046.435 5478.825 1047.435 ;
    END
  END Data_PMOS_NOSF[1144]
  PIN Data_PMOS_NOSF[1150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5451.945 1046.435 5452.225 1047.435 ;
    END
  END Data_PMOS_NOSF[1150]
  PIN Data_PMOS_NOSF[1151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5449.705 1046.435 5449.985 1047.435 ;
    END
  END Data_PMOS_NOSF[1151]
  PIN MASKD[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5448.025 1046.435 5448.305 1047.435 ;
    END
  END MASKD[108]
  PIN DIG_MON_PMOS_NOSF[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5442.425 1046.435 5442.705 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[107]
  PIN Data_PMOS_NOSF[1131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5440.185 1046.435 5440.465 1047.435 ;
    END
  END Data_PMOS_NOSF[1131]
  PIN Data_PMOS_NOSF[1125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5426.185 1046.435 5426.465 1047.435 ;
    END
  END Data_PMOS_NOSF[1125]
  PIN DIG_MON_PMOS[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8242.425 1046.435 8242.705 1047.435 ;
    END
  END DIG_MON_PMOS[65]
  PIN Data_PMOS[680]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8239.625 1046.435 8239.905 1047.435 ;
    END
  END Data_PMOS[680]
  PIN Data_PMOS[691]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8225.625 1046.435 8225.905 1047.435 ;
    END
  END Data_PMOS[691]
  PIN Data_PMOS[692]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8223.945 1046.435 8224.225 1047.435 ;
    END
  END Data_PMOS[692]
  PIN INJ_IN[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8221.145 1046.435 8221.425 1047.435 ;
    END
  END INJ_IN[177]
  PIN BcidMtx[533]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8218.905 1046.435 8219.185 1047.435 ;
    END
  END BcidMtx[533]
  PIN FREEZE_PMOS[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8217.225 1046.435 8217.505 1047.435 ;
    END
  END FREEZE_PMOS[32]
  PIN BcidMtx[530]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8216.105 1046.435 8216.385 1047.435 ;
    END
  END BcidMtx[530]
  PIN INJ_IN[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8213.865 1046.435 8214.145 1047.435 ;
    END
  END INJ_IN[176]
  PIN Data_PMOS[674]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8173.545 1046.435 8173.825 1047.435 ;
    END
  END Data_PMOS[674]
  PIN Data_PMOS[682]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8171.865 1046.435 8172.145 1047.435 ;
    END
  END Data_PMOS[682]
  PIN Data_PMOS[673]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8169.625 1046.435 8169.905 1047.435 ;
    END
  END Data_PMOS[673]
  PIN Data_PMOS[689]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8168.505 1046.435 8168.785 1047.435 ;
    END
  END Data_PMOS[689]
  PIN MASKD[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8166.825 1046.435 8167.105 1047.435 ;
    END
  END MASKD[176]
  PIN DIG_MON_SEL[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8163.465 1046.435 8163.745 1047.435 ;
    END
  END DIG_MON_SEL[175]
  PIN DIG_MON_PMOS[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8161.225 1046.435 8161.505 1047.435 ;
    END
  END DIG_MON_PMOS[63]
  PIN Data_PMOS[669]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8150.585 1046.435 8150.865 1047.435 ;
    END
  END Data_PMOS[669]
  PIN Data_PMOS[656]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8148.345 1046.435 8148.625 1047.435 ;
    END
  END Data_PMOS[656]
  PIN Data_PMOS[671]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8147.225 1046.435 8147.505 1047.435 ;
    END
  END Data_PMOS[671]
  PIN Data_PMOS[657]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8145.545 1046.435 8145.825 1047.435 ;
    END
  END Data_PMOS[657]
  PIN BcidMtx[526]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8139.665 1046.435 8139.945 1047.435 ;
    END
  END BcidMtx[526]
  PIN Read_PMOS[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8112.505 1046.435 8112.785 1047.435 ;
    END
  END Read_PMOS[31]
  PIN INJ_IN[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8109.705 1046.435 8109.985 1047.435 ;
    END
  END INJ_IN[174]
  PIN Data_PMOS[660]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8107.465 1046.435 8107.745 1047.435 ;
    END
  END Data_PMOS[660]
  PIN Data_PMOS[661]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8106.345 1046.435 8106.625 1047.435 ;
    END
  END Data_PMOS[661]
  PIN Data_PMOS[662]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8104.665 1046.435 8104.945 1047.435 ;
    END
  END Data_PMOS[662]
  PIN MASKV[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8102.425 1046.435 8102.705 1047.435 ;
    END
  END MASKV[174]
  PIN MASKD[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8101.305 1046.435 8101.585 1047.435 ;
    END
  END MASKD[174]
  PIN DIG_MON_SEL[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8085.625 1046.435 8085.905 1047.435 ;
    END
  END DIG_MON_SEL[174]
  PIN INJ_ROW[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8081.705 1046.435 8081.985 1047.435 ;
    END
  END INJ_ROW[86]
  PIN Data_PMOS[648]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8080.585 1046.435 8080.865 1047.435 ;
    END
  END Data_PMOS[648]
  PIN Data_PMOS[649]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8078.905 1046.435 8079.185 1047.435 ;
    END
  END Data_PMOS[649]
  PIN Data_PMOS[644]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8076.665 1046.435 8076.945 1047.435 ;
    END
  END Data_PMOS[644]
  PIN Data_PMOS[636]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8075.545 1046.435 8075.825 1047.435 ;
    END
  END Data_PMOS[636]
  PIN BcidMtx[521]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8032.985 1046.435 8033.265 1047.435 ;
    END
  END BcidMtx[521]
  PIN Read_PMOS[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8030.745 1046.435 8031.025 1047.435 ;
    END
  END Read_PMOS[30]
  PIN BcidMtx[517]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8029.625 1046.435 8029.905 1047.435 ;
    END
  END BcidMtx[517]
  PIN Data_PMOS[633]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8026.825 1046.435 8027.105 1047.435 ;
    END
  END Data_PMOS[633]
  PIN Data_PMOS[640]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8024.585 1046.435 8024.865 1047.435 ;
    END
  END Data_PMOS[640]
  PIN Data_PMOS[646]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8023.465 1046.435 8023.745 1047.435 ;
    END
  END Data_PMOS[646]
  PIN Data_PMOS[630]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8021.785 1046.435 8022.065 1047.435 ;
    END
  END Data_PMOS[630]
  PIN MASKD[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8011.145 1046.435 8011.425 1047.435 ;
    END
  END MASKD[172]
  PIN MASKD[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8006.665 1046.435 8006.945 1047.435 ;
    END
  END MASKD[171]
  PIN Data_PMOS[617]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8000.785 1046.435 8001.065 1047.435 ;
    END
  END Data_PMOS[617]
  PIN Data_PMOS[628]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7999.665 1046.435 7999.945 1047.435 ;
    END
  END Data_PMOS[628]
  PIN Data_PMOS[622]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7973.065 1046.435 7973.345 1047.435 ;
    END
  END Data_PMOS[622]
  PIN INJ_IN[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7969.705 1046.435 7969.985 1047.435 ;
    END
  END INJ_IN[171]
  PIN BcidMtx[515]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7967.465 1046.435 7967.745 1047.435 ;
    END
  END BcidMtx[515]
  PIN BcidMtx[513]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7966.345 1046.435 7966.625 1047.435 ;
    END
  END BcidMtx[513]
  PIN BcidMtx[511]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7964.105 1046.435 7964.385 1047.435 ;
    END
  END BcidMtx[511]
  PIN Data_PMOS[612]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7961.305 1046.435 7961.585 1047.435 ;
    END
  END Data_PMOS[612]
  PIN Data_PMOS[624]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7946.745 1046.435 7947.025 1047.435 ;
    END
  END Data_PMOS[624]
  PIN Data_PMOS[625]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7945.065 1046.435 7945.345 1047.435 ;
    END
  END Data_PMOS[625]
  PIN Data_PMOS[609]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7943.385 1046.435 7943.665 1047.435 ;
    END
  END Data_PMOS[609]
  PIN MASKH[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7941.705 1046.435 7941.985 1047.435 ;
    END
  END MASKH[85]
  PIN DIG_MON_SEL[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7938.345 1046.435 7938.625 1047.435 ;
    END
  END DIG_MON_SEL[170]
  PIN MASKD[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7936.665 1046.435 7936.945 1047.435 ;
    END
  END MASKD[169]
  PIN MASKV[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7933.865 1046.435 7934.145 1047.435 ;
    END
  END MASKV[169]
  PIN Data_PMOS[607]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7891.865 1046.435 7892.145 1047.435 ;
    END
  END Data_PMOS[607]
  PIN Data_PMOS[608]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7890.185 1046.435 7890.465 1047.435 ;
    END
  END Data_PMOS[608]
  PIN Data_PMOS[595]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7889.065 1046.435 7889.345 1047.435 ;
    END
  END Data_PMOS[595]
  PIN BcidMtx[509]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7885.145 1046.435 7885.425 1047.435 ;
    END
  END BcidMtx[509]
  PIN BcidMtx[507]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7884.025 1046.435 7884.305 1047.435 ;
    END
  END BcidMtx[507]
  PIN Read_PMOS[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7882.905 1046.435 7883.185 1047.435 ;
    END
  END Read_PMOS[28]
  PIN INJ_IN[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7871.705 1046.435 7871.985 1047.435 ;
    END
  END INJ_IN[168]
  PIN Data_PMOS[597]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7869.465 1046.435 7869.745 1047.435 ;
    END
  END Data_PMOS[597]
  PIN Data_PMOS[592]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7867.785 1046.435 7868.065 1047.435 ;
    END
  END Data_PMOS[592]
  PIN Data_PMOS[589]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7866.105 1046.435 7866.385 1047.435 ;
    END
  END Data_PMOS[589]
  PIN MASKV[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7862.465 1046.435 7862.745 1047.435 ;
    END
  END MASKV[168]
  PIN DIG_MON_PMOS[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7860.225 1046.435 7860.505 1047.435 ;
    END
  END DIG_MON_PMOS[56]
  PIN DIG_MON_SEL[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8951.945 1046.435 8952.225 1047.435 ;
    END
  END DIG_MON_SEL[195]
  PIN DIG_MON_PMOS[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8949.705 1046.435 8949.985 1047.435 ;
    END
  END DIG_MON_PMOS[83]
  PIN Data_PMOS[879]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8947.465 1046.435 8947.745 1047.435 ;
    END
  END Data_PMOS[879]
  PIN Data_PMOS[880]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8945.785 1046.435 8946.065 1047.435 ;
    END
  END Data_PMOS[880]
  PIN Data_PMOS[881]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8944.105 1046.435 8944.385 1047.435 ;
    END
  END Data_PMOS[881]
  PIN Data_PMOS[867]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8942.425 1046.435 8942.705 1047.435 ;
    END
  END Data_PMOS[867]
  PIN BcidMtx[586]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8925.065 1046.435 8925.345 1047.435 ;
    END
  END BcidMtx[586]
  PIN FREEZE_PMOS[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8923.945 1046.435 8924.225 1047.435 ;
    END
  END FREEZE_PMOS[41]
  PIN BcidMtx[583]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8922.265 1046.435 8922.545 1047.435 ;
    END
  END BcidMtx[583]
  PIN Data_PMOS[863]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8918.905 1046.435 8919.185 1047.435 ;
    END
  END Data_PMOS[863]
  PIN Data_PMOS[876]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8917.785 1046.435 8918.065 1047.435 ;
    END
  END Data_PMOS[876]
  PIN Data_PMOS[877]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8916.105 1046.435 8916.385 1047.435 ;
    END
  END Data_PMOS[877]
  PIN Data_PMOS[861]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8914.425 1046.435 8914.705 1047.435 ;
    END
  END Data_PMOS[861]
  PIN MASKH[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8874.105 1046.435 8874.385 1047.435 ;
    END
  END MASKH[97]
  PIN MASKD[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8869.065 1046.435 8869.345 1047.435 ;
    END
  END MASKD[193]
  PIN MASKV[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8866.265 1046.435 8866.545 1047.435 ;
    END
  END MASKV[193]
  PIN Data_PMOS[852]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8864.585 1046.435 8864.865 1047.435 ;
    END
  END Data_PMOS[852]
  PIN Data_PMOS[860]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8862.345 1046.435 8862.625 1047.435 ;
    END
  END Data_PMOS[860]
  PIN Data_PMOS[847]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8861.225 1046.435 8861.505 1047.435 ;
    END
  END Data_PMOS[847]
  PIN nTOK_PMOS[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8850.025 1046.435 8850.305 1047.435 ;
    END
  END nTOK_PMOS[40]
  PIN BcidMtx[580]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8848.345 1046.435 8848.625 1047.435 ;
    END
  END BcidMtx[580]
  PIN Read_PMOS[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8846.665 1046.435 8846.945 1047.435 ;
    END
  END Read_PMOS[40]
  PIN BcidMtx[576]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8844.985 1046.435 8845.265 1047.435 ;
    END
  END BcidMtx[576]
  PIN Data_PMOS[842]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8840.225 1046.435 8840.505 1047.435 ;
    END
  END Data_PMOS[842]
  PIN Data_PMOS[850]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8838.545 1046.435 8838.825 1047.435 ;
    END
  END Data_PMOS[850]
  PIN Data_PMOS[851]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8811.385 1046.435 8811.665 1047.435 ;
    END
  END Data_PMOS[851]
  PIN Data_PMOS[857]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8809.705 1046.435 8809.985 1047.435 ;
    END
  END Data_PMOS[857]
  PIN MASKD[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8808.025 1046.435 8808.305 1047.435 ;
    END
  END MASKD[192]
  PIN DIG_MON_SEL[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8805.225 1046.435 8805.505 1047.435 ;
    END
  END DIG_MON_SEL[192]
  PIN INJ_ROW[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8801.305 1046.435 8801.585 1047.435 ;
    END
  END INJ_ROW[95]
  PIN Data_PMOS[971]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9345.065 1046.435 9345.345 1047.435 ;
    END
  END Data_PMOS[971]
  PIN Data_PMOS[980]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9343.385 1046.435 9343.665 1047.435 ;
    END
  END Data_PMOS[980]
  PIN nTOK_PMOS[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9340.025 1046.435 9340.305 1047.435 ;
    END
  END nTOK_PMOS[46]
  PIN BcidMtx[616]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9338.345 1046.435 9338.625 1047.435 ;
    END
  END BcidMtx[616]
  PIN Read_PMOS[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9336.665 1046.435 9336.945 1047.435 ;
    END
  END Read_PMOS[46]
  PIN INJ_IN[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9333.865 1046.435 9334.145 1047.435 ;
    END
  END INJ_IN[204]
  PIN Data_PMOS[968]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9293.545 1046.435 9293.825 1047.435 ;
    END
  END Data_PMOS[968]
  PIN Data_PMOS[976]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9291.865 1046.435 9292.145 1047.435 ;
    END
  END Data_PMOS[976]
  PIN Data_PMOS[967]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9289.625 1046.435 9289.905 1047.435 ;
    END
  END Data_PMOS[967]
  PIN Data_PMOS[983]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9288.505 1046.435 9288.785 1047.435 ;
    END
  END Data_PMOS[983]
  PIN MASKD[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9286.825 1046.435 9287.105 1047.435 ;
    END
  END MASKD[204]
  PIN DIG_MON_SEL[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9284.025 1046.435 9284.305 1047.435 ;
    END
  END DIG_MON_SEL[204]
  PIN DIG_MON_PMOS[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9281.225 1046.435 9281.505 1047.435 ;
    END
  END DIG_MON_PMOS[91]
  PIN Data_PMOS[963]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9270.585 1046.435 9270.865 1047.435 ;
    END
  END Data_PMOS[963]
  PIN Data_PMOS[964]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9268.905 1046.435 9269.185 1047.435 ;
    END
  END Data_PMOS[964]
  PIN Data_PMOS[965]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9267.225 1046.435 9267.505 1047.435 ;
    END
  END Data_PMOS[965]
  PIN Data_PMOS[951]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9265.545 1046.435 9265.825 1047.435 ;
    END
  END Data_PMOS[951]
  PIN BcidMtx[610]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9259.665 1046.435 9259.945 1047.435 ;
    END
  END BcidMtx[610]
  PIN Read_PMOS[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9232.505 1046.435 9232.785 1047.435 ;
    END
  END Read_PMOS[45]
  PIN BcidMtx[606]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9230.825 1046.435 9231.105 1047.435 ;
    END
  END BcidMtx[606]
  PIN Data_PMOS[947]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9228.025 1046.435 9228.305 1047.435 ;
    END
  END Data_PMOS[947]
  PIN Data_PMOS[955]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9226.345 1046.435 9226.625 1047.435 ;
    END
  END Data_PMOS[955]
  PIN Data_PMOS[956]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9224.665 1046.435 9224.945 1047.435 ;
    END
  END Data_PMOS[956]
  PIN Data_PMOS[962]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9222.985 1046.435 9223.265 1047.435 ;
    END
  END Data_PMOS[962]
  PIN MASKD[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9221.305 1046.435 9221.585 1047.435 ;
    END
  END MASKD[202]
  PIN DIG_MON_SEL[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9205.625 1046.435 9205.905 1047.435 ;
    END
  END DIG_MON_SEL[202]
  PIN DIG_MON_PMOS[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9202.825 1046.435 9203.105 1047.435 ;
    END
  END DIG_MON_PMOS[89]
  PIN MASKV[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9201.145 1046.435 9201.425 1047.435 ;
    END
  END MASKV[201]
  PIN Data_PMOS[936]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9199.465 1046.435 9199.745 1047.435 ;
    END
  END Data_PMOS[936]
  PIN Data_PMOS[944]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9197.225 1046.435 9197.505 1047.435 ;
    END
  END Data_PMOS[944]
  PIN Data_PMOS[931]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9196.105 1046.435 9196.385 1047.435 ;
    END
  END Data_PMOS[931]
  PIN nTOK_PMOS[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9154.105 1046.435 9154.385 1047.435 ;
    END
  END nTOK_PMOS[44]
  PIN BcidMtx[603]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9151.865 1046.435 9152.145 1047.435 ;
    END
  END BcidMtx[603]
  PIN BcidMtx[602]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9150.185 1046.435 9150.465 1047.435 ;
    END
  END BcidMtx[602]
  PIN INJ_IN[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9147.945 1046.435 9148.225 1047.435 ;
    END
  END INJ_IN[200]
  PIN Data_PMOS[933]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9145.705 1046.435 9145.985 1047.435 ;
    END
  END Data_PMOS[933]
  PIN Data_PMOS[928]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9144.025 1046.435 9144.305 1047.435 ;
    END
  END Data_PMOS[928]
  PIN Data_PMOS[925]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9142.345 1046.435 9142.625 1047.435 ;
    END
  END Data_PMOS[925]
  PIN MASKH[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9131.705 1046.435 9131.985 1047.435 ;
    END
  END MASKH[100]
  PIN DIG_MON_PMOS[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9130.025 1046.435 9130.305 1047.435 ;
    END
  END DIG_MON_PMOS[88]
  PIN DIG_MON_SEL[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9127.785 1046.435 9128.065 1047.435 ;
    END
  END DIG_MON_SEL[199]
  PIN INJ_ROW[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9122.465 1046.435 9122.745 1047.435 ;
    END
  END INJ_ROW[99]
  PIN MASKV[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9121.905 1046.435 9122.185 1047.435 ;
    END
  END MASKV[199]
  PIN Data_PMOS[915]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9120.225 1046.435 9120.505 1047.435 ;
    END
  END Data_PMOS[915]
  PIN Data_PMOS[923]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9092.505 1046.435 9092.785 1047.435 ;
    END
  END Data_PMOS[923]
  PIN Data_PMOS[910]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9091.385 1046.435 9091.665 1047.435 ;
    END
  END Data_PMOS[910]
  PIN nTOK_PMOS[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9088.585 1046.435 9088.865 1047.435 ;
    END
  END nTOK_PMOS[43]
  PIN FREEZE_PMOS[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9085.785 1046.435 9086.065 1047.435 ;
    END
  END FREEZE_PMOS[43]
  PIN BcidMtx[596]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9084.665 1046.435 9084.945 1047.435 ;
    END
  END BcidMtx[596]
  PIN INJ_IN[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9082.425 1046.435 9082.705 1047.435 ;
    END
  END INJ_IN[198]
  PIN Data_PMOS[918]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9066.745 1046.435 9067.025 1047.435 ;
    END
  END Data_PMOS[918]
  PIN Data_PMOS[907]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9065.625 1046.435 9065.905 1047.435 ;
    END
  END Data_PMOS[907]
  PIN Data_PMOS[904]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9063.945 1046.435 9064.225 1047.435 ;
    END
  END Data_PMOS[904]
  PIN MASKV[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9062.265 1046.435 9062.545 1047.435 ;
    END
  END MASKV[198]
  PIN DIG_MON_PMOS[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9060.025 1046.435 9060.305 1047.435 ;
    END
  END DIG_MON_PMOS[86]
  PIN DIG_MON_SEL[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9057.785 1046.435 9058.065 1047.435 ;
    END
  END DIG_MON_SEL[197]
  PIN INJ_ROW[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9054.425 1046.435 9054.705 1047.435 ;
    END
  END INJ_ROW[98]
  PIN Data_PMOS[890]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9012.985 1046.435 9013.265 1047.435 ;
    END
  END Data_PMOS[890]
  PIN Data_PMOS[887]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9011.305 1046.435 9011.585 1047.435 ;
    END
  END Data_PMOS[887]
  PIN Data_PMOS[896]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9009.625 1046.435 9009.905 1047.435 ;
    END
  END Data_PMOS[896]
  PIN Data_PMOS[888]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9008.505 1046.435 9008.785 1047.435 ;
    END
  END Data_PMOS[888]
  PIN BcidMtx[592]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9004.585 1046.435 9004.865 1047.435 ;
    END
  END BcidMtx[592]
  PIN Read_PMOS[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9002.905 1046.435 9003.185 1047.435 ;
    END
  END Read_PMOS[42]
  PIN BcidMtx[589]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9001.785 1046.435 9002.065 1047.435 ;
    END
  END BcidMtx[589]
  PIN Data_PMOS[884]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8990.025 1046.435 8990.305 1047.435 ;
    END
  END Data_PMOS[884]
  PIN Data_PMOS[892]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8988.345 1046.435 8988.625 1047.435 ;
    END
  END Data_PMOS[892]
  PIN Data_PMOS[886]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8987.785 1046.435 8988.065 1047.435 ;
    END
  END Data_PMOS[886]
  PIN Data_PMOS[899]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8984.985 1046.435 8985.265 1047.435 ;
    END
  END Data_PMOS[899]
  PIN MASKD[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8981.345 1046.435 8981.625 1047.435 ;
    END
  END MASKD[196]
  PIN MASKD[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10070.825 1046.435 10071.105 1047.435 ;
    END
  END MASKD[223]
  PIN INJ_ROW[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10068.585 1046.435 10068.865 1047.435 ;
    END
  END INJ_ROW[111]
  PIN Data_PMOS[1173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10067.465 1046.435 10067.745 1047.435 ;
    END
  END Data_PMOS[1173]
  PIN Data_PMOS[1160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10065.225 1046.435 10065.505 1047.435 ;
    END
  END Data_PMOS[1160]
  PIN Data_PMOS[1169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10063.545 1046.435 10063.825 1047.435 ;
    END
  END Data_PMOS[1169]
  PIN INJ_IN[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10061.305 1046.435 10061.585 1047.435 ;
    END
  END INJ_IN[223]
  PIN BcidMtx[670]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10045.065 1046.435 10045.345 1047.435 ;
    END
  END BcidMtx[670]
  PIN Read_PMOS[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10043.385 1046.435 10043.665 1047.435 ;
    END
  END Read_PMOS[55]
  PIN BcidMtx[667]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10042.265 1046.435 10042.545 1047.435 ;
    END
  END BcidMtx[667]
  PIN Data_PMOS[1157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10038.905 1046.435 10039.185 1047.435 ;
    END
  END Data_PMOS[1157]
  PIN Data_PMOS[1165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10037.225 1046.435 10037.505 1047.435 ;
    END
  END Data_PMOS[1165]
  PIN Data_PMOS[1166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10035.545 1046.435 10035.825 1047.435 ;
    END
  END Data_PMOS[1166]
  PIN Data_PMOS[1172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10033.865 1046.435 10034.145 1047.435 ;
    END
  END Data_PMOS[1172]
  PIN MASKD[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9993.545 1046.435 9993.825 1047.435 ;
    END
  END MASKD[222]
  PIN DIG_MON_SEL[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9990.745 1046.435 9991.025 1047.435 ;
    END
  END DIG_MON_SEL[222]
  PIN DIG_MON_PMOS[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9987.945 1046.435 9988.225 1047.435 ;
    END
  END DIG_MON_PMOS[109]
  PIN Data_HV[1069]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18639.665 1046.435 18639.945 1047.435 ;
    END
  END Data_HV[1069]
  PIN Data_PMOS[1146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9984.585 1046.435 9984.865 1047.435 ;
    END
  END Data_PMOS[1146]
  PIN Data_PMOS[1147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9982.905 1046.435 9983.185 1047.435 ;
    END
  END Data_PMOS[1147]
  PIN Data_PMOS[1141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9981.225 1046.435 9981.505 1047.435 ;
    END
  END Data_PMOS[1141]
  PIN INJ_IN[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9971.145 1046.435 9971.425 1047.435 ;
    END
  END INJ_IN[221]
  PIN BcidMtx[663]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9967.785 1046.435 9968.065 1047.435 ;
    END
  END BcidMtx[663]
  PIN BcidMtx[662]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9966.105 1046.435 9966.385 1047.435 ;
    END
  END BcidMtx[662]
  PIN BcidMtx[660]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9964.985 1046.435 9965.265 1047.435 ;
    END
  END BcidMtx[660]
  PIN Data_PMOS[1143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9959.665 1046.435 9959.945 1047.435 ;
    END
  END Data_PMOS[1143]
  PIN Data_PMOS[1138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9932.505 1046.435 9932.785 1047.435 ;
    END
  END Data_PMOS[1138]
  PIN Data_PMOS[1145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9931.385 1046.435 9931.665 1047.435 ;
    END
  END Data_PMOS[1145]
  PIN MASKV[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9929.145 1046.435 9929.425 1047.435 ;
    END
  END MASKV[220]
  PIN DIG_MON_PMOS[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9926.905 1046.435 9927.185 1047.435 ;
    END
  END DIG_MON_PMOS[108]
  PIN INJ_ROW[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9921.305 1046.435 9921.585 1047.435 ;
    END
  END INJ_ROW[109]
  PIN Data_PMOS[1121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9919.625 1046.435 9919.905 1047.435 ;
    END
  END Data_PMOS[1121]
  PIN DIG_MON_COMP[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13286.905 1046.435 13287.185 1047.435 ;
    END
  END DIG_MON_COMP[80]
  PIN DIG_MON_SEL[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13284.665 1046.435 13284.945 1047.435 ;
    END
  END DIG_MON_SEL[303]
  PIN INJ_ROW[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13281.305 1046.435 13281.585 1047.435 ;
    END
  END INJ_ROW[151]
  PIN Data_COMP[837]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13280.185 1046.435 13280.465 1047.435 ;
    END
  END Data_COMP[837]
  PIN Data_COMP[824]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13265.065 1046.435 13265.345 1047.435 ;
    END
  END Data_COMP[824]
  PIN Data_COMP[833]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13263.385 1046.435 13263.665 1047.435 ;
    END
  END Data_COMP[833]
  PIN Data_COMP[825]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13262.265 1046.435 13262.545 1047.435 ;
    END
  END Data_COMP[825]
  PIN BcidMtx[910]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13258.345 1046.435 13258.625 1047.435 ;
    END
  END BcidMtx[910]
  PIN Read_COMP[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13256.665 1046.435 13256.945 1047.435 ;
    END
  END Read_COMP[39]
  PIN BcidMtx[906]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13254.985 1046.435 13255.265 1047.435 ;
    END
  END BcidMtx[906]
  PIN Data_COMP[821]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13213.545 1046.435 13213.825 1047.435 ;
    END
  END Data_COMP[821]
  PIN Data_COMP[829]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13211.865 1046.435 13212.145 1047.435 ;
    END
  END Data_COMP[829]
  PIN Data_COMP[835]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13210.745 1046.435 13211.025 1047.435 ;
    END
  END Data_COMP[835]
  PIN Data_COMP[836]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13208.505 1046.435 13208.785 1047.435 ;
    END
  END Data_COMP[836]
  PIN MASKD[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13206.825 1046.435 13207.105 1047.435 ;
    END
  END MASKD[302]
  PIN INJ_IN[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18609.705 1046.435 18609.985 1047.435 ;
    END
  END INJ_IN[437]
  PIN INJ_ROW[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13191.705 1046.435 13191.985 1047.435 ;
    END
  END INJ_ROW[150]
  PIN Data_COMP[816]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13190.585 1046.435 13190.865 1047.435 ;
    END
  END Data_COMP[816]
  PIN Data_COMP[803]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13188.345 1046.435 13188.625 1047.435 ;
    END
  END Data_COMP[803]
  PIN Data_COMP[812]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13186.665 1046.435 13186.945 1047.435 ;
    END
  END Data_COMP[812]
  PIN Data_COMP[804]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13185.545 1046.435 13185.825 1047.435 ;
    END
  END Data_COMP[804]
  PIN BcidMtx[904]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13179.665 1046.435 13179.945 1047.435 ;
    END
  END BcidMtx[904]
  PIN BcidMtx[902]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13151.945 1046.435 13152.225 1047.435 ;
    END
  END BcidMtx[902]
  PIN BcidMtx[900]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13150.825 1046.435 13151.105 1047.435 ;
    END
  END BcidMtx[900]
  PIN Data_COMP[807]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13147.465 1046.435 13147.745 1047.435 ;
    END
  END Data_COMP[807]
  PIN Data_COMP[802]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13145.785 1046.435 13146.065 1047.435 ;
    END
  END Data_COMP[802]
  PIN Data_COMP[809]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13144.665 1046.435 13144.945 1047.435 ;
    END
  END Data_COMP[809]
  PIN MASKV[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13142.425 1046.435 13142.705 1047.435 ;
    END
  END MASKV[300]
  PIN DIG_MON_COMP[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13140.185 1046.435 13140.465 1047.435 ;
    END
  END DIG_MON_COMP[76]
  PIN DIG_MON_SEL[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13125.625 1046.435 13125.905 1047.435 ;
    END
  END DIG_MON_SEL[300]
  PIN DIG_MON_COMP[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13122.825 1046.435 13123.105 1047.435 ;
    END
  END DIG_MON_COMP[75]
  PIN Data_HV[1108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18745.225 1046.435 18745.505 1047.435 ;
    END
  END Data_HV[1108]
  PIN Data_COMP[785]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13120.025 1046.435 13120.305 1047.435 ;
    END
  END Data_COMP[785]
  PIN Data_COMP[782]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13118.345 1046.435 13118.625 1047.435 ;
    END
  END Data_COMP[782]
  PIN Data_COMP[791]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13116.665 1046.435 13116.945 1047.435 ;
    END
  END Data_COMP[791]
  PIN Data_COMP[783]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13115.545 1046.435 13115.825 1047.435 ;
    END
  END Data_COMP[783]
  PIN BcidMtx[898]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13072.425 1046.435 13072.705 1047.435 ;
    END
  END BcidMtx[898]
  PIN Read_COMP[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13070.745 1046.435 13071.025 1047.435 ;
    END
  END Read_COMP[37]
  PIN BcidMtx[895]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13069.625 1046.435 13069.905 1047.435 ;
    END
  END BcidMtx[895]
  PIN Data_COMP[779]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13066.265 1046.435 13066.545 1047.435 ;
    END
  END Data_COMP[779]
  PIN Data_COMP[787]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13064.585 1046.435 13064.865 1047.435 ;
    END
  END Data_COMP[787]
  PIN Data_COMP[788]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13062.905 1046.435 13063.185 1047.435 ;
    END
  END Data_COMP[788]
  PIN Data_COMP[794]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13061.225 1046.435 13061.505 1047.435 ;
    END
  END Data_COMP[794]
  PIN MASKD[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13051.145 1046.435 13051.425 1047.435 ;
    END
  END MASKD[298]
  PIN DIG_MON_SEL[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13047.785 1046.435 13048.065 1047.435 ;
    END
  END DIG_MON_SEL[297]
  PIN Data_COMP[774]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13041.345 1046.435 13041.625 1047.435 ;
    END
  END Data_COMP[774]
  PIN Data_COMP[768]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13040.225 1046.435 13040.505 1047.435 ;
    END
  END Data_COMP[768]
  PIN Data_HV[1066]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18585.065 1046.435 18585.345 1047.435 ;
    END
  END Data_HV[1066]
  PIN Data_COMP[776]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13012.505 1046.435 13012.785 1047.435 ;
    END
  END Data_COMP[776]
  PIN Data_COMP[763]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13011.385 1046.435 13011.665 1047.435 ;
    END
  END Data_COMP[763]
  PIN BcidMtx[893]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13007.465 1046.435 13007.745 1047.435 ;
    END
  END BcidMtx[893]
  PIN FREEZE_COMP[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13005.785 1046.435 13006.065 1047.435 ;
    END
  END FREEZE_COMP[36]
  PIN BcidMtx[890]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13004.665 1046.435 13004.945 1047.435 ;
    END
  END BcidMtx[890]
  PIN Data_COMP[759]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13001.305 1046.435 13001.585 1047.435 ;
    END
  END Data_COMP[759]
  PIN Data_COMP[771]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12986.745 1046.435 12987.025 1047.435 ;
    END
  END Data_COMP[771]
  PIN Data_COMP[760]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12985.625 1046.435 12985.905 1047.435 ;
    END
  END Data_COMP[760]
  PIN Data_COMP[756]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12983.385 1046.435 12983.665 1047.435 ;
    END
  END Data_COMP[756]
  PIN MASKH[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12981.705 1046.435 12981.985 1047.435 ;
    END
  END MASKH[148]
  PIN DIG_MON_COMP[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12980.025 1046.435 12980.305 1047.435 ;
    END
  END DIG_MON_COMP[72]
  PIN MASKD[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12976.665 1046.435 12976.945 1047.435 ;
    END
  END MASKD[295]
  PIN MASKV[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12973.865 1046.435 12974.145 1047.435 ;
    END
  END MASKV[295]
  PIN Data_COMP[743]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12932.985 1046.435 12933.265 1047.435 ;
    END
  END Data_COMP[743]
  PIN Data_COMP[748]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12930.745 1046.435 12931.025 1047.435 ;
    END
  END Data_COMP[748]
  PIN Data_COMP[742]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12929.065 1046.435 12929.345 1047.435 ;
    END
  END Data_COMP[742]
  PIN INJ_IN[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12927.385 1046.435 12927.665 1047.435 ;
    END
  END INJ_IN[295]
  PIN BcidMtx[885]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12924.025 1046.435 12924.305 1047.435 ;
    END
  END BcidMtx[885]
  PIN BcidMtx[884]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12922.345 1046.435 12922.625 1047.435 ;
    END
  END BcidMtx[884]
  PIN BcidMtx[882]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12921.225 1046.435 12921.505 1047.435 ;
    END
  END BcidMtx[882]
  PIN Data_COMP[744]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12909.465 1046.435 12909.745 1047.435 ;
    END
  END Data_COMP[744]
  PIN Data_COMP[739]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12907.785 1046.435 12908.065 1047.435 ;
    END
  END Data_COMP[739]
  PIN Data_COMP[746]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12906.665 1046.435 12906.945 1047.435 ;
    END
  END Data_COMP[746]
  PIN MASKV[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12902.465 1046.435 12902.745 1047.435 ;
    END
  END MASKV[294]
  PIN DIG_MON_COMP[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12900.225 1046.435 12900.505 1047.435 ;
    END
  END DIG_MON_COMP[70]
  PIN DIG_MON_SEL[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12898.545 1046.435 12898.825 1047.435 ;
    END
  END DIG_MON_SEL[294]
  PIN DIG_MON_COMP[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13989.705 1046.435 13989.985 1047.435 ;
    END
  END DIG_MON_COMP[97]
  PIN Data_COMP[1026]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13987.465 1046.435 13987.745 1047.435 ;
    END
  END Data_COMP[1026]
  PIN Data_HV[1093]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18744.105 1046.435 18744.385 1047.435 ;
    END
  END Data_HV[1093]
  PIN Data_COMP[1021]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13984.665 1046.435 13984.945 1047.435 ;
    END
  END Data_COMP[1021]
  PIN Data_COMP[1015]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13982.985 1046.435 13983.265 1047.435 ;
    END
  END Data_COMP[1015]
  PIN INJ_IN[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13981.305 1046.435 13981.585 1047.435 ;
    END
  END INJ_IN[321]
  PIN BcidMtx[963]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13964.505 1046.435 13964.785 1047.435 ;
    END
  END BcidMtx[963]
  PIN BcidMtx[962]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13962.825 1046.435 13963.105 1047.435 ;
    END
  END BcidMtx[962]
  PIN BcidMtx[960]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13961.705 1046.435 13961.985 1047.435 ;
    END
  END BcidMtx[960]
  PIN Data_COMP[1017]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13958.345 1046.435 13958.625 1047.435 ;
    END
  END Data_COMP[1017]
  PIN Data_COMP[1012]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13956.665 1046.435 13956.945 1047.435 ;
    END
  END Data_COMP[1012]
  PIN Data_COMP[1019]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13955.545 1046.435 13955.825 1047.435 ;
    END
  END Data_COMP[1019]
  PIN MASKV[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13914.665 1046.435 13914.945 1047.435 ;
    END
  END MASKV[320]
  PIN DIG_MON_COMP[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13912.425 1046.435 13912.705 1047.435 ;
    END
  END DIG_MON_COMP[96]
  PIN DIG_MON_SEL[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13910.745 1046.435 13911.025 1047.435 ;
    END
  END DIG_MON_SEL[320]
  PIN INJ_ROW[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13906.825 1046.435 13907.105 1047.435 ;
    END
  END INJ_ROW[159]
  PIN Data_COMP[995]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13905.145 1046.435 13905.425 1047.435 ;
    END
  END Data_COMP[995]
  PIN Data_COMP[1006]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13904.025 1046.435 13904.305 1047.435 ;
    END
  END Data_COMP[1006]
  PIN Data_COMP[1001]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13901.785 1046.435 13902.065 1047.435 ;
    END
  END Data_COMP[1001]
  PIN INJ_IN[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13891.145 1046.435 13891.425 1047.435 ;
    END
  END INJ_IN[319]
  PIN BcidMtx[959]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13888.905 1046.435 13889.185 1047.435 ;
    END
  END BcidMtx[959]
  PIN Read_COMP[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13886.665 1046.435 13886.945 1047.435 ;
    END
  END Read_COMP[47]
  PIN BcidMtx[954]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13884.985 1046.435 13885.265 1047.435 ;
    END
  END BcidMtx[954]
  PIN Data_COMP[990]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13880.785 1046.435 13881.065 1047.435 ;
    END
  END Data_COMP[990]
  PIN Data_COMP[997]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13878.545 1046.435 13878.825 1047.435 ;
    END
  END Data_COMP[997]
  PIN Data_COMP[998]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13851.385 1046.435 13851.665 1047.435 ;
    END
  END Data_COMP[998]
  PIN Data_COMP[1134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14410.265 1046.435 14410.545 1047.435 ;
    END
  END Data_COMP[1134]
  PIN MASKH[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14408.585 1046.435 14408.865 1047.435 ;
    END
  END MASKH[166]
  PIN DIG_MON_SEL[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14405.225 1046.435 14405.505 1047.435 ;
    END
  END DIG_MON_SEL[332]
  PIN MASKD[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14403.545 1046.435 14403.825 1047.435 ;
    END
  END MASKD[331]
  PIN MASKV[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14400.745 1046.435 14401.025 1047.435 ;
    END
  END MASKV[331]
  PIN Data_COMP[1132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14385.625 1046.435 14385.905 1047.435 ;
    END
  END Data_COMP[1132]
  PIN Data_COMP[1126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14384.505 1046.435 14384.785 1047.435 ;
    END
  END Data_COMP[1126]
  PIN Data_COMP[1120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14382.825 1046.435 14383.105 1047.435 ;
    END
  END Data_COMP[1120]
  PIN BcidMtx[995]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14378.905 1046.435 14379.185 1047.435 ;
    END
  END BcidMtx[995]
  PIN BcidMtx[993]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14377.785 1046.435 14378.065 1047.435 ;
    END
  END BcidMtx[993]
  PIN BcidMtx[992]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14376.105 1046.435 14376.385 1047.435 ;
    END
  END BcidMtx[992]
  PIN Data_COMP[1116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14334.105 1046.435 14334.385 1047.435 ;
    END
  END Data_COMP[1116]
  PIN Data_COMP[1122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14332.985 1046.435 14333.265 1047.435 ;
    END
  END Data_COMP[1122]
  PIN Data_COMP[1117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14331.305 1046.435 14331.585 1047.435 ;
    END
  END Data_COMP[1117]
  PIN Data_COMP[1113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14329.065 1046.435 14329.345 1047.435 ;
    END
  END Data_COMP[1113]
  PIN MASKV[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14327.945 1046.435 14328.225 1047.435 ;
    END
  END MASKV[330]
  PIN DIG_MON_COMP[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14325.705 1046.435 14325.985 1047.435 ;
    END
  END DIG_MON_COMP[106]
  PIN MASKD[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14322.345 1046.435 14322.625 1047.435 ;
    END
  END MASKD[329]
  PIN INJ_ROW[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14311.705 1046.435 14311.985 1047.435 ;
    END
  END INJ_ROW[164]
  PIN Data_COMP[1100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14310.025 1046.435 14310.305 1047.435 ;
    END
  END Data_COMP[1100]
  PIN Data_COMP[1105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14307.785 1046.435 14308.065 1047.435 ;
    END
  END Data_COMP[1105]
  PIN Data_COMP[1106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14306.665 1046.435 14306.945 1047.435 ;
    END
  END Data_COMP[1106]
  PIN INJ_IN[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14302.465 1046.435 14302.745 1047.435 ;
    END
  END INJ_IN[329]
  PIN BcidMtx[987]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14299.105 1046.435 14299.385 1047.435 ;
    END
  END BcidMtx[987]
  PIN BcidMtx[986]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14271.945 1046.435 14272.225 1047.435 ;
    END
  END BcidMtx[986]
  PIN Data_COMP[1095]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14268.585 1046.435 14268.865 1047.435 ;
    END
  END Data_COMP[1095]
  PIN Data_COMP[1107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14266.905 1046.435 14267.185 1047.435 ;
    END
  END Data_COMP[1107]
  PIN Data_COMP[1096]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14265.785 1046.435 14266.065 1047.435 ;
    END
  END Data_COMP[1096]
  PIN Data_COMP[1093]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14264.105 1046.435 14264.385 1047.435 ;
    END
  END Data_COMP[1093]
  PIN MASKH[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14261.865 1046.435 14262.145 1047.435 ;
    END
  END MASKH[164]
  PIN MASKD[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14261.305 1046.435 14261.585 1047.435 ;
    END
  END MASKD[328]
  PIN DIG_MON_SEL[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14245.625 1046.435 14245.905 1047.435 ;
    END
  END DIG_MON_SEL[328]
  PIN INJ_ROW[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14241.705 1046.435 14241.985 1047.435 ;
    END
  END INJ_ROW[163]
  PIN Data_COMP[1089]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14240.585 1046.435 14240.865 1047.435 ;
    END
  END Data_COMP[1089]
  PIN Data_COMP[1090]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14238.905 1046.435 14239.185 1047.435 ;
    END
  END Data_COMP[1090]
  PIN Data_COMP[1085]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14236.665 1046.435 14236.945 1047.435 ;
    END
  END Data_COMP[1085]
  PIN Data_COMP[1077]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14235.545 1046.435 14235.825 1047.435 ;
    END
  END Data_COMP[1077]
  PIN BcidMtx[983]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14192.985 1046.435 14193.265 1047.435 ;
    END
  END BcidMtx[983]
  PIN Read_COMP[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14190.745 1046.435 14191.025 1047.435 ;
    END
  END Read_COMP[51]
  PIN BcidMtx[979]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14189.625 1046.435 14189.905 1047.435 ;
    END
  END BcidMtx[979]
  PIN Data_COMP[1074]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14186.825 1046.435 14187.105 1047.435 ;
    END
  END Data_COMP[1074]
  PIN Data_COMP[1081]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14184.585 1046.435 14184.865 1047.435 ;
    END
  END Data_COMP[1081]
  PIN Data_COMP[1087]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14183.465 1046.435 14183.745 1047.435 ;
    END
  END Data_COMP[1087]
  PIN Data_COMP[1071]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14181.785 1046.435 14182.065 1047.435 ;
    END
  END Data_COMP[1071]
  PIN MASKD[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14171.145 1046.435 14171.425 1047.435 ;
    END
  END MASKD[326]
  PIN DIG_MON_SEL[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14167.785 1046.435 14168.065 1047.435 ;
    END
  END DIG_MON_SEL[325]
  PIN MASKV[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14161.905 1046.435 14162.185 1047.435 ;
    END
  END MASKV[325]
  PIN Data_COMP[1058]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14160.785 1046.435 14161.065 1047.435 ;
    END
  END Data_COMP[1058]
  PIN Data_COMP[1055]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14159.105 1046.435 14159.385 1047.435 ;
    END
  END Data_COMP[1055]
  PIN Data_COMP[1057]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14131.385 1046.435 14131.665 1047.435 ;
    END
  END Data_COMP[1057]
  PIN INJ_IN[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14129.705 1046.435 14129.985 1047.435 ;
    END
  END INJ_IN[325]
  PIN BcidMtx[976]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14126.905 1046.435 14127.185 1047.435 ;
    END
  END BcidMtx[976]
  PIN BcidMtx[974]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14124.665 1046.435 14124.945 1047.435 ;
    END
  END BcidMtx[974]
  PIN BcidMtx[972]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14123.545 1046.435 14123.825 1047.435 ;
    END
  END BcidMtx[972]
  PIN Data_COMP[1052]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14120.745 1046.435 14121.025 1047.435 ;
    END
  END Data_COMP[1052]
  PIN Data_COMP[1054]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14105.625 1046.435 14105.905 1047.435 ;
    END
  END Data_COMP[1054]
  PIN Data_COMP[1061]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14104.505 1046.435 14104.785 1047.435 ;
    END
  END Data_COMP[1061]
  PIN Data_COMP[1067]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14102.825 1046.435 14103.105 1047.435 ;
    END
  END Data_COMP[1067]
  PIN MASKD[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14101.145 1046.435 14101.425 1047.435 ;
    END
  END MASKD[324]
  PIN MASKD[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14096.665 1046.435 14096.945 1047.435 ;
    END
  END MASKD[323]
  PIN Data_COMP[1047]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14053.545 1046.435 14053.825 1047.435 ;
    END
  END Data_COMP[1047]
  PIN Data_COMP[1041]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14052.425 1046.435 14052.705 1047.435 ;
    END
  END Data_COMP[1041]
  PIN Data_COMP[1042]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14050.745 1046.435 14051.025 1047.435 ;
    END
  END Data_COMP[1042]
  PIN Data_COMP[1035]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14048.505 1046.435 14048.785 1047.435 ;
    END
  END Data_COMP[1035]
  PIN nTOK_COMP[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14046.265 1046.435 14046.545 1047.435 ;
    END
  END nTOK_COMP[49]
  PIN BcidMtx[969]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14044.025 1046.435 14044.305 1047.435 ;
    END
  END BcidMtx[969]
  PIN BcidMtx[966]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14041.225 1046.435 14041.505 1047.435 ;
    END
  END BcidMtx[966]
  PIN Data_COMP[1032]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14030.585 1046.435 14030.865 1047.435 ;
    END
  END Data_COMP[1032]
  PIN Data_COMP[1038]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14029.465 1046.435 14029.745 1047.435 ;
    END
  END Data_COMP[1038]
  PIN Data_COMP[1040]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14026.665 1046.435 14026.945 1047.435 ;
    END
  END Data_COMP[1040]
  PIN Data_COMP[1046]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14024.985 1046.435 14025.265 1047.435 ;
    END
  END Data_COMP[1046]
  PIN MASKH[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14021.905 1046.435 14022.185 1047.435 ;
    END
  END MASKH[161]
  PIN DIG_MON_SEL[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15111.945 1046.435 15112.225 1047.435 ;
    END
  END DIG_MON_SEL[349]
  PIN INJ_ROW[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15108.585 1046.435 15108.865 1047.435 ;
    END
  END INJ_ROW[174]
  PIN Data_HV[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15106.905 1046.435 15107.185 1047.435 ;
    END
  END Data_HV[134]
  PIN Data_HV[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15105.225 1046.435 15105.505 1047.435 ;
    END
  END Data_HV[131]
  PIN Data_HV[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15103.545 1046.435 15103.825 1047.435 ;
    END
  END Data_HV[140]
  PIN nTOK_HV[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15100.185 1046.435 15100.465 1047.435 ;
    END
  END nTOK_HV[6]
  PIN BcidMtx[1048]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15085.065 1046.435 15085.345 1047.435 ;
    END
  END BcidMtx[1048]
  PIN Read_HV[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15083.385 1046.435 15083.665 1047.435 ;
    END
  END Read_HV[6]
  PIN INJ_IN[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15080.585 1046.435 15080.865 1047.435 ;
    END
  END INJ_IN[348]
  PIN Data_HV[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15078.345 1046.435 15078.625 1047.435 ;
    END
  END Data_HV[135]
  PIN Data_HV[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15077.225 1046.435 15077.505 1047.435 ;
    END
  END Data_HV[136]
  PIN Data_HV[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15074.985 1046.435 15075.265 1047.435 ;
    END
  END Data_HV[127]
  PIN MASKV[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15034.665 1046.435 15034.945 1047.435 ;
    END
  END MASKV[348]
  PIN MASKD[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15033.545 1046.435 15033.825 1047.435 ;
    END
  END MASKD[348]
  PIN DIG_MON_SEL[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15030.185 1046.435 15030.465 1047.435 ;
    END
  END DIG_MON_SEL[347]
  PIN INJ_ROW[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15026.825 1046.435 15027.105 1047.435 ;
    END
  END INJ_ROW[173]
  PIN Data_HV[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15025.145 1046.435 15025.425 1047.435 ;
    END
  END Data_HV[113]
  PIN Data_HV[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15023.465 1046.435 15023.745 1047.435 ;
    END
  END Data_HV[110]
  PIN Data_HV[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15021.785 1046.435 15022.065 1047.435 ;
    END
  END Data_HV[119]
  PIN INJ_IN[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15011.145 1046.435 15011.425 1047.435 ;
    END
  END INJ_IN[347]
  PIN BcidMtx[1041]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15007.785 1046.435 15008.065 1047.435 ;
    END
  END BcidMtx[1041]
  PIN Read_HV[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15006.665 1046.435 15006.945 1047.435 ;
    END
  END Read_HV[5]
  PIN BcidMtx[1038]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15004.985 1046.435 15005.265 1047.435 ;
    END
  END BcidMtx[1038]
  PIN Data_HV[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15000.225 1046.435 15000.505 1047.435 ;
    END
  END Data_HV[107]
  PIN Data_HV[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14998.545 1046.435 14998.825 1047.435 ;
    END
  END Data_HV[115]
  PIN Data_HV[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14971.385 1046.435 14971.665 1047.435 ;
    END
  END Data_HV[116]
  PIN MASKV[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14969.145 1046.435 14969.425 1047.435 ;
    END
  END MASKV[346]
  PIN DIG_MON_COMP[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12726.905 1046.435 12727.185 1047.435 ;
    END
  END DIG_MON_COMP[66]
  PIN DIG_MON_SEL[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12724.665 1046.435 12724.945 1047.435 ;
    END
  END DIG_MON_SEL[289]
  PIN INJ_ROW[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12721.305 1046.435 12721.585 1047.435 ;
    END
  END INJ_ROW[144]
  PIN Data_COMP[680]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12719.625 1046.435 12719.905 1047.435 ;
    END
  END Data_COMP[680]
  PIN Data_COMP[677]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12705.065 1046.435 12705.345 1047.435 ;
    END
  END Data_COMP[677]
  PIN Data_COMP[686]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12703.385 1046.435 12703.665 1047.435 ;
    END
  END Data_COMP[686]
  PIN Data_COMP[678]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12702.265 1046.435 12702.545 1047.435 ;
    END
  END Data_COMP[678]
  PIN BcidMtx[868]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12698.345 1046.435 12698.625 1047.435 ;
    END
  END BcidMtx[868]
  PIN Read_COMP[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12696.665 1046.435 12696.945 1047.435 ;
    END
  END Read_COMP[32]
  PIN INJ_IN[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12693.865 1046.435 12694.145 1047.435 ;
    END
  END INJ_IN[288]
  PIN Data_COMP[674]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12653.545 1046.435 12653.825 1047.435 ;
    END
  END Data_COMP[674]
  PIN Data_COMP[682]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12651.865 1046.435 12652.145 1047.435 ;
    END
  END Data_COMP[682]
  PIN Data_COMP[683]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12650.185 1046.435 12650.465 1047.435 ;
    END
  END Data_COMP[683]
  PIN Data_COMP[689]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12648.505 1046.435 12648.785 1047.435 ;
    END
  END Data_COMP[689]
  PIN MASKD[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12646.825 1046.435 12647.105 1047.435 ;
    END
  END MASKD[288]
  PIN DIG_MON_SEL[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12644.025 1046.435 12644.305 1047.435 ;
    END
  END DIG_MON_SEL[288]
  PIN DIG_MON_COMP[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12641.225 1046.435 12641.505 1047.435 ;
    END
  END DIG_MON_COMP[63]
  PIN Data_COMP[669]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12630.585 1046.435 12630.865 1047.435 ;
    END
  END Data_COMP[669]
  PIN Data_COMP[659]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12630.025 1046.435 12630.305 1047.435 ;
    END
  END Data_COMP[659]
  PIN Data_COMP[664]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12627.785 1046.435 12628.065 1047.435 ;
    END
  END Data_COMP[664]
  PIN Data_COMP[658]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12626.105 1046.435 12626.385 1047.435 ;
    END
  END Data_COMP[658]
  PIN INJ_IN[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12622.465 1046.435 12622.745 1047.435 ;
    END
  END INJ_IN[287]
  PIN BcidMtx[861]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12619.105 1046.435 12619.385 1047.435 ;
    END
  END BcidMtx[861]
  PIN BcidMtx[859]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12591.385 1046.435 12591.665 1047.435 ;
    END
  END BcidMtx[859]
  PIN Data_COMP[654]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12588.585 1046.435 12588.865 1047.435 ;
    END
  END Data_COMP[654]
  PIN Data_COMP[666]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12586.905 1046.435 12587.185 1047.435 ;
    END
  END Data_COMP[666]
  PIN Data_COMP[667]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12585.225 1046.435 12585.505 1047.435 ;
    END
  END Data_COMP[667]
  PIN Data_COMP[651]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12583.545 1046.435 12583.825 1047.435 ;
    END
  END Data_COMP[651]
  PIN MASKH[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12581.865 1046.435 12582.145 1047.435 ;
    END
  END MASKH[143]
  PIN MASKD[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12563.945 1046.435 12564.225 1047.435 ;
    END
  END MASKD[285]
  PIN MASKV[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12561.145 1046.435 12561.425 1047.435 ;
    END
  END MASKV[285]
  PIN Data_COMP[642]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12559.465 1046.435 12559.745 1047.435 ;
    END
  END Data_COMP[642]
  PIN Data_COMP[643]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12557.785 1046.435 12558.065 1047.435 ;
    END
  END Data_COMP[643]
  PIN Data_HV[1094]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18748.025 1046.435 18748.305 1047.435 ;
    END
  END Data_HV[1094]
  PIN INJ_IN[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12554.425 1046.435 12554.705 1047.435 ;
    END
  END INJ_IN[285]
  PIN BcidMtx[856]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12512.425 1046.435 12512.705 1047.435 ;
    END
  END BcidMtx[856]
  PIN Read_COMP[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12510.745 1046.435 12511.025 1047.435 ;
    END
  END Read_COMP[30]
  PIN BcidMtx[852]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12509.065 1046.435 12509.345 1047.435 ;
    END
  END BcidMtx[852]
  PIN Data_COMP[633]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12506.825 1046.435 12507.105 1047.435 ;
    END
  END Data_COMP[633]
  PIN Data_COMP[640]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12504.585 1046.435 12504.865 1047.435 ;
    END
  END Data_COMP[640]
  PIN Data_COMP[641]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12502.905 1046.435 12503.185 1047.435 ;
    END
  END Data_COMP[641]
  PIN Data_COMP[630]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12501.785 1046.435 12502.065 1047.435 ;
    END
  END Data_COMP[630]
  PIN MASKD[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12491.145 1046.435 12491.425 1047.435 ;
    END
  END MASKD[284]
  PIN DIG_MON_SEL[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12488.345 1046.435 12488.625 1047.435 ;
    END
  END DIG_MON_SEL[284]
  PIN MASKD[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12486.665 1046.435 12486.945 1047.435 ;
    END
  END MASKD[283]
  PIN Data_COMP[627]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12481.345 1046.435 12481.625 1047.435 ;
    END
  END Data_COMP[627]
  PIN Data_COMP[628]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12479.665 1046.435 12479.945 1047.435 ;
    END
  END Data_COMP[628]
  PIN Data_COMP[622]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12453.065 1046.435 12453.345 1047.435 ;
    END
  END Data_COMP[622]
  PIN Data_COMP[616]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12451.385 1046.435 12451.665 1047.435 ;
    END
  END Data_COMP[616]
  PIN nTOK_COMP[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12448.585 1046.435 12448.865 1047.435 ;
    END
  END nTOK_COMP[29]
  PIN BcidMtx[849]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12446.345 1046.435 12446.625 1047.435 ;
    END
  END BcidMtx[849]
  PIN BcidMtx[848]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12444.665 1046.435 12444.945 1047.435 ;
    END
  END BcidMtx[848]
  PIN INJ_IN[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12442.425 1046.435 12442.705 1047.435 ;
    END
  END INJ_IN[282]
  PIN Data_COMP[611]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12440.745 1046.435 12441.025 1047.435 ;
    END
  END Data_COMP[611]
  PIN Data_COMP[613]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12425.625 1046.435 12425.905 1047.435 ;
    END
  END Data_COMP[613]
  PIN Data_COMP[610]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12423.945 1046.435 12424.225 1047.435 ;
    END
  END Data_COMP[610]
  PIN MASKV[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12422.265 1046.435 12422.545 1047.435 ;
    END
  END MASKV[282]
  PIN DIG_MON_COMP[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12420.025 1046.435 12420.305 1047.435 ;
    END
  END DIG_MON_COMP[58]
  PIN DIG_MON_SEL[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12417.785 1046.435 12418.065 1047.435 ;
    END
  END DIG_MON_SEL[281]
  PIN INJ_ROW[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12414.425 1046.435 12414.705 1047.435 ;
    END
  END INJ_ROW[140]
  PIN Data_COMP[596]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12372.985 1046.435 12373.265 1047.435 ;
    END
  END Data_COMP[596]
  PIN Data_COMP[593]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12371.305 1046.435 12371.585 1047.435 ;
    END
  END Data_COMP[593]
  PIN Data_COMP[608]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12370.185 1046.435 12370.465 1047.435 ;
    END
  END Data_COMP[608]
  PIN Data_COMP[594]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12368.505 1046.435 12368.785 1047.435 ;
    END
  END Data_COMP[594]
  PIN BcidMtx[845]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12365.145 1046.435 12365.425 1047.435 ;
    END
  END BcidMtx[845]
  PIN BcidMtx[843]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12364.025 1046.435 12364.305 1047.435 ;
    END
  END BcidMtx[843]
  PIN BcidMtx[841]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12361.785 1046.435 12362.065 1047.435 ;
    END
  END BcidMtx[841]
  PIN Data_COMP[591]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12350.585 1046.435 12350.865 1047.435 ;
    END
  END Data_COMP[591]
  PIN Data_COMP[603]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12348.905 1046.435 12349.185 1047.435 ;
    END
  END Data_COMP[603]
  PIN Data_COMP[604]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12347.225 1046.435 12347.505 1047.435 ;
    END
  END Data_COMP[604]
  PIN Data_COMP[588]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12345.545 1046.435 12345.825 1047.435 ;
    END
  END Data_COMP[588]
  PIN MASKH[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12341.905 1046.435 12342.185 1047.435 ;
    END
  END MASKH[140]
  PIN DIG_MON_SEL[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13431.945 1046.435 13432.225 1047.435 ;
    END
  END DIG_MON_SEL[307]
  PIN DIG_MON_COMP[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13429.705 1046.435 13429.985 1047.435 ;
    END
  END DIG_MON_COMP[83]
  PIN Data_COMP[869]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13426.905 1046.435 13427.185 1047.435 ;
    END
  END Data_COMP[869]
  PIN Data_COMP[866]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13425.225 1046.435 13425.505 1047.435 ;
    END
  END Data_COMP[866]
  PIN Data_COMP[881]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13424.105 1046.435 13424.385 1047.435 ;
    END
  END Data_COMP[881]
  PIN Data_COMP[867]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13422.425 1046.435 13422.705 1047.435 ;
    END
  END Data_COMP[867]
  PIN BcidMtx[923]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13405.625 1046.435 13405.905 1047.435 ;
    END
  END BcidMtx[923]
  PIN BcidMtx[921]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13404.505 1046.435 13404.785 1047.435 ;
    END
  END BcidMtx[921]
  PIN BcidMtx[919]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13402.265 1046.435 13402.545 1047.435 ;
    END
  END BcidMtx[919]
  PIN Data_COMP[864]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13399.465 1046.435 13399.745 1047.435 ;
    END
  END Data_COMP[864]
  PIN Data_COMP[870]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13398.345 1046.435 13398.625 1047.435 ;
    END
  END Data_COMP[870]
  PIN Data_COMP[877]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13396.105 1046.435 13396.385 1047.435 ;
    END
  END Data_COMP[877]
  PIN Data_COMP[861]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13394.425 1046.435 13394.705 1047.435 ;
    END
  END Data_COMP[861]
  PIN MASKV[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13354.665 1046.435 13354.945 1047.435 ;
    END
  END MASKV[306]
  PIN MASKD[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13349.065 1046.435 13349.345 1047.435 ;
    END
  END MASKD[305]
  PIN MASKV[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13346.265 1046.435 13346.545 1047.435 ;
    END
  END MASKV[305]
  PIN Data_COMP[852]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13344.585 1046.435 13344.865 1047.435 ;
    END
  END Data_COMP[852]
  PIN Data_COMP[853]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13342.905 1046.435 13343.185 1047.435 ;
    END
  END Data_COMP[853]
  PIN Data_COMP[847]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13341.225 1046.435 13341.505 1047.435 ;
    END
  END Data_COMP[847]
  PIN nTOK_COMP[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13330.025 1046.435 13330.305 1047.435 ;
    END
  END nTOK_COMP[40]
  PIN BcidMtx[915]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13327.785 1046.435 13328.065 1047.435 ;
    END
  END BcidMtx[915]
  PIN Read_COMP[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13326.665 1046.435 13326.945 1047.435 ;
    END
  END Read_COMP[40]
  PIN INJ_IN[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13321.905 1046.435 13322.185 1047.435 ;
    END
  END INJ_IN[304]
  PIN Data_COMP[849]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13319.665 1046.435 13319.945 1047.435 ;
    END
  END Data_COMP[849]
  PIN Data_COMP[850]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13318.545 1046.435 13318.825 1047.435 ;
    END
  END Data_COMP[850]
  PIN Data_COMP[841]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13290.825 1046.435 13291.105 1047.435 ;
    END
  END Data_COMP[841]
  PIN Data_COMP[857]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13289.705 1046.435 13289.985 1047.435 ;
    END
  END Data_COMP[857]
  PIN DIG_MON_COMP[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11602.425 1046.435 11602.705 1047.435 ;
    END
  END DIG_MON_COMP[37]
  PIN Data_COMP[396]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11600.185 1046.435 11600.465 1047.435 ;
    END
  END Data_COMP[396]
  PIN Data_COMP[390]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11586.185 1046.435 11586.465 1047.435 ;
    END
  END Data_COMP[390]
  PIN Data_COMP[398]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11583.945 1046.435 11584.225 1047.435 ;
    END
  END Data_COMP[398]
  PIN Data_COMP[384]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11582.265 1046.435 11582.545 1047.435 ;
    END
  END Data_COMP[384]
  PIN nTOK_COMP[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11580.025 1046.435 11580.305 1047.435 ;
    END
  END nTOK_COMP[18]
  PIN FREEZE_COMP[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11577.225 1046.435 11577.505 1047.435 ;
    END
  END FREEZE_COMP[18]
  PIN BcidMtx[781]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11575.545 1046.435 11575.825 1047.435 ;
    END
  END BcidMtx[781]
  PIN INJ_IN[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11573.865 1046.435 11574.145 1047.435 ;
    END
  END INJ_IN[260]
  PIN Data_COMP[393]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11532.425 1046.435 11532.705 1047.435 ;
    END
  END Data_COMP[393]
  PIN Data_COMP[394]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11530.745 1046.435 11531.025 1047.435 ;
    END
  END Data_COMP[394]
  PIN Data_COMP[379]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11529.625 1046.435 11529.905 1047.435 ;
    END
  END Data_COMP[379]
  PIN MASKH[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11527.385 1046.435 11527.665 1047.435 ;
    END
  END MASKH[130]
  PIN DIG_MON_SEL[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11523.465 1046.435 11523.745 1047.435 ;
    END
  END DIG_MON_SEL[259]
  PIN MASKV[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11511.145 1046.435 11511.425 1047.435 ;
    END
  END MASKV[259]
  PIN Data_COMP[369]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11509.465 1046.435 11509.745 1047.435 ;
    END
  END Data_COMP[369]
  PIN Data_COMP[362]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11508.345 1046.435 11508.625 1047.435 ;
    END
  END Data_COMP[362]
  PIN Data_COMP[364]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11506.105 1046.435 11506.385 1047.435 ;
    END
  END Data_COMP[364]
  PIN nTOK_COMP[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11501.345 1046.435 11501.625 1047.435 ;
    END
  END nTOK_COMP[17]
  PIN BcidMtx[778]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11499.665 1046.435 11499.945 1047.435 ;
    END
  END BcidMtx[778]
  PIN BcidMtx[775]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11471.385 1046.435 11471.665 1047.435 ;
    END
  END BcidMtx[775]
  PIN Data_COMP[360]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11468.585 1046.435 11468.865 1047.435 ;
    END
  END Data_COMP[360]
  PIN Data_COMP[366]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11467.465 1046.435 11467.745 1047.435 ;
    END
  END Data_COMP[366]
  PIN Data_COMP[373]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11465.225 1046.435 11465.505 1047.435 ;
    END
  END Data_COMP[373]
  PIN Data_COMP[357]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11463.545 1046.435 11463.825 1047.435 ;
    END
  END Data_COMP[357]
  PIN MASKV[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11462.425 1046.435 11462.705 1047.435 ;
    END
  END MASKV[258]
  PIN MASKD[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11443.945 1046.435 11444.225 1047.435 ;
    END
  END MASKD[257]
  PIN INJ_ROW[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11441.705 1046.435 11441.985 1047.435 ;
    END
  END INJ_ROW[128]
  PIN Data_COMP[348]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11439.465 1046.435 11439.745 1047.435 ;
    END
  END Data_COMP[348]
  PIN Data_COMP[349]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11437.785 1046.435 11438.065 1047.435 ;
    END
  END Data_COMP[349]
  PIN Data_COMP[350]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11436.665 1046.435 11436.945 1047.435 ;
    END
  END Data_COMP[350]
  PIN nTOK_COMP[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11394.105 1046.435 11394.385 1047.435 ;
    END
  END nTOK_COMP[16]
  PIN BcidMtx[771]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11391.865 1046.435 11392.145 1047.435 ;
    END
  END BcidMtx[771]
  PIN nTOK_HV[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18781.345 1046.435 18781.625 1047.435 ;
    END
  END nTOK_HV[52]
  PIN BcidMtx[1325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18780.225 1046.435 18780.505 1047.435 ;
    END
  END BcidMtx[1325]
  PIN Data_COMP[339]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11386.825 1046.435 11387.105 1047.435 ;
    END
  END Data_COMP[339]
  PIN Data_COMP[345]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11385.705 1046.435 11385.985 1047.435 ;
    END
  END Data_COMP[345]
  PIN Data_COMP[352]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11383.465 1046.435 11383.745 1047.435 ;
    END
  END Data_COMP[352]
  PIN Data_COMP[336]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11381.785 1046.435 11382.065 1047.435 ;
    END
  END Data_COMP[336]
  PIN MASKV[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11372.265 1046.435 11372.545 1047.435 ;
    END
  END MASKV[256]
  PIN MASKD[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11366.665 1046.435 11366.945 1047.435 ;
    END
  END MASKD[255]
  PIN INJ_ROW[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11362.465 1046.435 11362.745 1047.435 ;
    END
  END INJ_ROW[127]
  PIN Data_COMP[327]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11360.225 1046.435 11360.505 1047.435 ;
    END
  END Data_COMP[327]
  PIN Data_COMP[328]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11333.065 1046.435 11333.345 1047.435 ;
    END
  END Data_COMP[328]
  PIN Data_COMP[329]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11331.945 1046.435 11332.225 1047.435 ;
    END
  END Data_COMP[329]
  PIN nTOK_COMP[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11328.585 1046.435 11328.865 1047.435 ;
    END
  END nTOK_COMP[15]
  PIN BcidMtx[765]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11326.345 1046.435 11326.625 1047.435 ;
    END
  END BcidMtx[765]
  PIN Read_COMP[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11325.225 1046.435 11325.505 1047.435 ;
    END
  END Read_COMP[15]
  PIN INJ_IN[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11322.425 1046.435 11322.705 1047.435 ;
    END
  END INJ_IN[254]
  PIN Data_COMP[317]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11320.745 1046.435 11321.025 1047.435 ;
    END
  END Data_COMP[317]
  PIN Data_COMP[330]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11306.745 1046.435 11307.025 1047.435 ;
    END
  END Data_COMP[330]
  PIN Data_COMP[326]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11304.505 1046.435 11304.785 1047.435 ;
    END
  END Data_COMP[326]
  PIN Data_COMP[332]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11302.825 1046.435 11303.105 1047.435 ;
    END
  END Data_COMP[332]
  PIN MASKD[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11301.145 1046.435 11301.425 1047.435 ;
    END
  END MASKD[254]
  PIN DIG_MON_SEL[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11298.345 1046.435 11298.625 1047.435 ;
    END
  END DIG_MON_SEL[254]
  PIN DIG_MON_COMP[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11295.545 1046.435 11295.825 1047.435 ;
    END
  END DIG_MON_COMP[29]
  PIN Data_COMP[312]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11253.545 1046.435 11253.825 1047.435 ;
    END
  END Data_COMP[312]
  PIN Data_COMP[313]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11251.865 1046.435 11252.145 1047.435 ;
    END
  END Data_COMP[313]
  PIN Data_COMP[314]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11250.185 1046.435 11250.465 1047.435 ;
    END
  END Data_COMP[314]
  PIN Data_COMP[300]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11248.505 1046.435 11248.785 1047.435 ;
    END
  END Data_COMP[300]
  PIN BcidMtx[761]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11245.145 1046.435 11245.425 1047.435 ;
    END
  END BcidMtx[761]
  PIN FREEZE_COMP[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11243.465 1046.435 11243.745 1047.435 ;
    END
  END FREEZE_COMP[14]
  PIN BcidMtx[757]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11241.785 1046.435 11242.065 1047.435 ;
    END
  END BcidMtx[757]
  PIN INJ_IN[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11231.705 1046.435 11231.985 1047.435 ;
    END
  END INJ_IN[252]
  PIN Data_COMP[303]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11229.465 1046.435 11229.745 1047.435 ;
    END
  END Data_COMP[303]
  PIN Data_COMP[298]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11227.785 1046.435 11228.065 1047.435 ;
    END
  END Data_COMP[298]
  PIN Data_COMP[295]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11226.105 1046.435 11226.385 1047.435 ;
    END
  END Data_COMP[295]
  PIN MASKV[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11222.465 1046.435 11222.745 1047.435 ;
    END
  END MASKV[252]
  PIN DIG_MON_COMP[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11220.225 1046.435 11220.505 1047.435 ;
    END
  END DIG_MON_COMP[28]
  PIN FREEZE_COMP[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11473.065 1046.435 11473.345 1047.435 ;
    END
  END FREEZE_COMP[17]
  PIN DIG_MON_COMP[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12309.705 1046.435 12309.985 1047.435 ;
    END
  END DIG_MON_COMP[55]
  PIN Data_COMP[585]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12307.465 1046.435 12307.745 1047.435 ;
    END
  END Data_COMP[585]
  PIN Data_COMP[586]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12305.785 1046.435 12306.065 1047.435 ;
    END
  END Data_COMP[586]
  PIN Data_COMP[587]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12304.105 1046.435 12304.385 1047.435 ;
    END
  END Data_COMP[587]
  PIN Data_COMP[573]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12302.425 1046.435 12302.705 1047.435 ;
    END
  END Data_COMP[573]
  PIN BcidMtx[839]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12285.625 1046.435 12285.905 1047.435 ;
    END
  END BcidMtx[839]
  PIN FREEZE_COMP[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12283.945 1046.435 12284.225 1047.435 ;
    END
  END FREEZE_COMP[27]
  PIN BcidMtx[835]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12282.265 1046.435 12282.545 1047.435 ;
    END
  END BcidMtx[835]
  PIN Data_HV[1056]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18610.825 1046.435 18611.105 1047.435 ;
    END
  END Data_HV[1056]
  PIN Data_COMP[569]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12278.905 1046.435 12279.185 1047.435 ;
    END
  END Data_COMP[569]
  PIN Data_COMP[577]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12277.225 1046.435 12277.505 1047.435 ;
    END
  END Data_COMP[577]
  PIN Data_COMP[583]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12276.105 1046.435 12276.385 1047.435 ;
    END
  END Data_COMP[583]
  PIN Data_COMP[584]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12273.865 1046.435 12274.145 1047.435 ;
    END
  END Data_COMP[584]
  PIN MASKD[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12233.545 1046.435 12233.825 1047.435 ;
    END
  END MASKD[278]
  PIN DIG_MON_SEL[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12230.185 1046.435 12230.465 1047.435 ;
    END
  END DIG_MON_SEL[277]
  PIN INJ_ROW[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12226.825 1046.435 12227.105 1047.435 ;
    END
  END INJ_ROW[138]
  PIN Data_COMP[565]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12224.025 1046.435 12224.305 1047.435 ;
    END
  END Data_COMP[565]
  PIN Data_COMP[551]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12223.465 1046.435 12223.745 1047.435 ;
    END
  END Data_COMP[551]
  PIN Data_COMP[560]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12221.785 1046.435 12222.065 1047.435 ;
    END
  END Data_COMP[560]
  PIN BcidMtx[833]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12208.905 1046.435 12209.185 1047.435 ;
    END
  END BcidMtx[833]
  PIN BcidMtx[832]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12208.345 1046.435 12208.625 1047.435 ;
    END
  END BcidMtx[832]
  PIN Read_COMP[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12206.665 1046.435 12206.945 1047.435 ;
    END
  END Read_COMP[26]
  PIN Data_COMP[549]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12200.785 1046.435 12201.065 1047.435 ;
    END
  END Data_COMP[549]
  PIN Data_COMP[548]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12200.225 1046.435 12200.505 1047.435 ;
    END
  END Data_COMP[548]
  PIN Data_COMP[556]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12198.545 1046.435 12198.825 1047.435 ;
    END
  END Data_COMP[556]
  PIN Data_COMP[546]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12170.265 1046.435 12170.545 1047.435 ;
    END
  END Data_COMP[546]
  PIN Data_COMP[563]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12169.705 1046.435 12169.985 1047.435 ;
    END
  END Data_COMP[563]
  PIN MASKD[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12168.025 1046.435 12168.305 1047.435 ;
    END
  END MASKD[276]
  PIN MASKD[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12163.545 1046.435 12163.825 1047.435 ;
    END
  END MASKD[275]
  PIN DIG_MON_COMP[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12162.425 1046.435 12162.705 1047.435 ;
    END
  END DIG_MON_COMP[51]
  PIN Data_COMP[543]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12160.185 1046.435 12160.465 1047.435 ;
    END
  END Data_COMP[543]
  PIN Data_COMP[538]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12144.505 1046.435 12144.785 1047.435 ;
    END
  END Data_COMP[538]
  PIN Data_COMP[539]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12143.385 1046.435 12143.665 1047.435 ;
    END
  END Data_COMP[539]
  PIN Data_COMP[531]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12142.265 1046.435 12142.545 1047.435 ;
    END
  END Data_COMP[531]
  PIN BcidMtx[826]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12138.345 1046.435 12138.625 1047.435 ;
    END
  END BcidMtx[826]
  PIN FREEZE_COMP[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12137.225 1046.435 12137.505 1047.435 ;
    END
  END FREEZE_COMP[25]
  PIN BcidMtx[823]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12135.545 1046.435 12135.825 1047.435 ;
    END
  END BcidMtx[823]
  PIN Data_COMP[527]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12093.545 1046.435 12093.825 1047.435 ;
    END
  END Data_COMP[527]
  PIN Data_COMP[540]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12092.425 1046.435 12092.705 1047.435 ;
    END
  END Data_COMP[540]
  PIN Data_COMP[541]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12090.745 1046.435 12091.025 1047.435 ;
    END
  END Data_COMP[541]
  PIN Data_COMP[542]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12088.505 1046.435 12088.785 1047.435 ;
    END
  END Data_COMP[542]
  PIN MASKH[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12087.385 1046.435 12087.665 1047.435 ;
    END
  END MASKH[137]
  PIN DIG_MON_COMP[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12081.225 1046.435 12081.505 1047.435 ;
    END
  END DIG_MON_COMP[49]
  PIN MASKV[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12071.145 1046.435 12071.425 1047.435 ;
    END
  END MASKV[273]
  PIN Data_COMP[516]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12069.465 1046.435 12069.745 1047.435 ;
    END
  END Data_COMP[516]
  PIN Data_COMP[524]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12067.225 1046.435 12067.505 1047.435 ;
    END
  END Data_COMP[524]
  PIN Data_COMP[511]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12066.105 1046.435 12066.385 1047.435 ;
    END
  END Data_COMP[511]
  PIN INJ_IN[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12062.465 1046.435 12062.745 1047.435 ;
    END
  END INJ_IN[273]
  PIN BcidMtx[819]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12059.105 1046.435 12059.385 1047.435 ;
    END
  END BcidMtx[819]
  PIN BcidMtx[818]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12031.945 1046.435 12032.225 1047.435 ;
    END
  END BcidMtx[818]
  PIN INJ_IN[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12029.705 1046.435 12029.985 1047.435 ;
    END
  END INJ_IN[272]
  PIN Data_COMP[519]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12026.905 1046.435 12027.185 1047.435 ;
    END
  END Data_COMP[519]
  PIN Data_COMP[508]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12025.785 1046.435 12026.065 1047.435 ;
    END
  END Data_COMP[508]
  PIN Data_COMP[505]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12024.105 1046.435 12024.385 1047.435 ;
    END
  END Data_COMP[505]
  PIN MASKD[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12021.305 1046.435 12021.585 1047.435 ;
    END
  END MASKD[272]
  PIN MASKD[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12003.945 1046.435 12004.225 1047.435 ;
    END
  END MASKD[271]
  PIN Data_COMP[501]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12000.585 1046.435 12000.865 1047.435 ;
    END
  END Data_COMP[501]
  PIN Data_COMP[495]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11999.465 1046.435 11999.745 1047.435 ;
    END
  END Data_COMP[495]
  PIN Data_COMP[496]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11997.785 1046.435 11998.065 1047.435 ;
    END
  END Data_COMP[496]
  PIN Data_COMP[489]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11995.545 1046.435 11995.825 1047.435 ;
    END
  END Data_COMP[489]
  PIN nTOK_COMP[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11954.105 1046.435 11954.385 1047.435 ;
    END
  END nTOK_COMP[23]
  PIN BcidMtx[814]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11952.425 1046.435 11952.705 1047.435 ;
    END
  END BcidMtx[814]
  PIN BcidMtx[812]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11950.185 1046.435 11950.465 1047.435 ;
    END
  END BcidMtx[812]
  PIN BcidMtx[810]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11949.065 1046.435 11949.345 1047.435 ;
    END
  END BcidMtx[810]
  PIN Data_COMP[485]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11946.265 1046.435 11946.545 1047.435 ;
    END
  END Data_COMP[485]
  PIN Data_COMP[487]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11944.025 1046.435 11944.305 1047.435 ;
    END
  END Data_COMP[487]
  PIN Data_COMP[494]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11942.905 1046.435 11943.185 1047.435 ;
    END
  END Data_COMP[494]
  PIN Data_COMP[500]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11941.225 1046.435 11941.505 1047.435 ;
    END
  END Data_COMP[500]
  PIN DIG_MON_COMP[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11930.025 1046.435 11930.305 1047.435 ;
    END
  END DIG_MON_COMP[46]
  PIN DIG_MON_SEL[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11928.345 1046.435 11928.625 1047.435 ;
    END
  END DIG_MON_SEL[270]
  PIN DIG_MON_COMP[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11925.545 1046.435 11925.825 1047.435 ;
    END
  END DIG_MON_COMP[45]
  PIN Data_COMP[470]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11920.785 1046.435 11921.065 1047.435 ;
    END
  END Data_COMP[470]
  PIN Data_COMP[467]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11919.105 1046.435 11919.385 1047.435 ;
    END
  END Data_COMP[467]
  PIN Data_COMP[482]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11892.505 1046.435 11892.785 1047.435 ;
    END
  END Data_COMP[482]
  PIN nTOK_COMP[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11888.585 1046.435 11888.865 1047.435 ;
    END
  END nTOK_COMP[22]
  PIN BcidMtx[808]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11886.905 1046.435 11887.185 1047.435 ;
    END
  END BcidMtx[808]
  PIN BcidMtx[1320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18750.825 1046.435 18751.105 1047.435 ;
    END
  END BcidMtx[1320]
  PIN BcidMtx[805]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11884.105 1046.435 11884.385 1047.435 ;
    END
  END BcidMtx[805]
  PIN Data_COMP[465]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11881.305 1046.435 11881.585 1047.435 ;
    END
  END Data_COMP[465]
  PIN Data_COMP[477]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11866.745 1046.435 11867.025 1047.435 ;
    END
  END Data_COMP[477]
  PIN Data_COMP[478]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11865.065 1046.435 11865.345 1047.435 ;
    END
  END Data_COMP[478]
  PIN Data_COMP[462]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11863.385 1046.435 11863.665 1047.435 ;
    END
  END Data_COMP[462]
  PIN MASKH[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11861.705 1046.435 11861.985 1047.435 ;
    END
  END MASKH[134]
  PIN MASKD[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11856.665 1046.435 11856.945 1047.435 ;
    END
  END MASKD[267]
  PIN MASKV[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11853.865 1046.435 11854.145 1047.435 ;
    END
  END MASKV[267]
  PIN Data_COMP[449]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11812.985 1046.435 11813.265 1047.435 ;
    END
  END Data_COMP[449]
  PIN Data_COMP[460]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11811.865 1046.435 11812.145 1047.435 ;
    END
  END Data_COMP[460]
  PIN Data_COMP[461]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11810.185 1046.435 11810.465 1047.435 ;
    END
  END Data_COMP[461]
  PIN INJ_IN[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11807.385 1046.435 11807.665 1047.435 ;
    END
  END INJ_IN[267]
  PIN BcidMtx[803]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11805.145 1046.435 11805.425 1047.435 ;
    END
  END BcidMtx[803]
  PIN FREEZE_COMP[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11803.465 1046.435 11803.745 1047.435 ;
    END
  END FREEZE_COMP[21]
  PIN BcidMtx[800]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11802.345 1046.435 11802.625 1047.435 ;
    END
  END BcidMtx[800]
  PIN Data_COMP[444]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11790.585 1046.435 11790.865 1047.435 ;
    END
  END Data_COMP[444]
  PIN Data_COMP[456]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11788.905 1046.435 11789.185 1047.435 ;
    END
  END Data_COMP[456]
  PIN Data_COMP[457]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11787.225 1046.435 11787.505 1047.435 ;
    END
  END Data_COMP[457]
  PIN Data_COMP[442]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11786.105 1046.435 11786.385 1047.435 ;
    END
  END Data_COMP[442]
  PIN MASKH[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11781.905 1046.435 11782.185 1047.435 ;
    END
  END MASKH[133]
  PIN DIG_MON_COMP[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11780.225 1046.435 11780.505 1047.435 ;
    END
  END DIG_MON_COMP[42]
  PIN FREEZE_COMP[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12033.065 1046.435 12033.345 1047.435 ;
    END
  END FREEZE_COMP[24]
  PIN MASKD[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12870.825 1046.435 12871.105 1047.435 ;
    END
  END MASKD[293]
  PIN Data_COMP[732]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12867.465 1046.435 12867.745 1047.435 ;
    END
  END Data_COMP[732]
  PIN Data_COMP[733]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12865.785 1046.435 12866.065 1047.435 ;
    END
  END Data_COMP[733]
  PIN Data_COMP[727]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12864.665 1046.435 12864.945 1047.435 ;
    END
  END Data_COMP[727]
  PIN Data_COMP[721]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12862.985 1046.435 12863.265 1047.435 ;
    END
  END Data_COMP[721]
  PIN BcidMtx[881]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12845.625 1046.435 12845.905 1047.435 ;
    END
  END BcidMtx[881]
  PIN INJ_IN[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18749.705 1046.435 18749.985 1047.435 ;
    END
  END INJ_IN[440]
  PIN Read_COMP[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12843.385 1046.435 12843.665 1047.435 ;
    END
  END Read_COMP[34]
  PIN INJ_IN[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12840.585 1046.435 12840.865 1047.435 ;
    END
  END INJ_IN[292]
  PIN Data_COMP[716]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12838.905 1046.435 12839.185 1047.435 ;
    END
  END Data_COMP[716]
  PIN Data_COMP[724]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12837.225 1046.435 12837.505 1047.435 ;
    END
  END Data_COMP[724]
  PIN Data_COMP[725]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12835.545 1046.435 12835.825 1047.435 ;
    END
  END Data_COMP[725]
  PIN Data_COMP[731]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12833.865 1046.435 12834.145 1047.435 ;
    END
  END Data_COMP[731]
  PIN MASKD[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12793.545 1046.435 12793.825 1047.435 ;
    END
  END MASKD[292]
  PIN DIG_MON_SEL[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12790.745 1046.435 12791.025 1047.435 ;
    END
  END DIG_MON_SEL[292]
  PIN MASKD[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12789.065 1046.435 12789.345 1047.435 ;
    END
  END MASKD[291]
  PIN INJ_ROW[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12786.825 1046.435 12787.105 1047.435 ;
    END
  END INJ_ROW[145]
  PIN Data_COMP[712]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12784.025 1046.435 12784.305 1047.435 ;
    END
  END Data_COMP[712]
  PIN Data_COMP[706]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12782.905 1046.435 12783.185 1047.435 ;
    END
  END Data_COMP[706]
  PIN Data_COMP[699]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12772.265 1046.435 12772.545 1047.435 ;
    END
  END Data_COMP[699]
  PIN BcidMtx[875]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12768.905 1046.435 12769.185 1047.435 ;
    END
  END BcidMtx[875]
  PIN BcidMtx[873]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12767.785 1046.435 12768.065 1047.435 ;
    END
  END BcidMtx[873]
  PIN Read_COMP[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12766.665 1046.435 12766.945 1047.435 ;
    END
  END Read_COMP[33]
  PIN Data_COMP[696]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12760.785 1046.435 12761.065 1047.435 ;
    END
  END Data_COMP[696]
  PIN Data_COMP[708]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12759.105 1046.435 12759.385 1047.435 ;
    END
  END Data_COMP[708]
  PIN Data_COMP[703]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12758.545 1046.435 12758.825 1047.435 ;
    END
  END Data_COMP[703]
  PIN Data_COMP[694]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12730.825 1046.435 12731.105 1047.435 ;
    END
  END Data_COMP[694]
  PIN MASKV[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12729.145 1046.435 12729.425 1047.435 ;
    END
  END MASKV[290]
  PIN Data_PMOS[1132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9905.625 1046.435 9905.905 1047.435 ;
    END
  END Data_PMOS[1132]
  PIN Data_PMOS[1127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9903.385 1046.435 9903.665 1047.435 ;
    END
  END Data_PMOS[1127]
  PIN INJ_IN[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9901.145 1046.435 9901.425 1047.435 ;
    END
  END INJ_IN[219]
  PIN BcidMtx[659]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9898.905 1046.435 9899.185 1047.435 ;
    END
  END BcidMtx[659]
  PIN BcidMtx[657]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9897.785 1046.435 9898.065 1047.435 ;
    END
  END BcidMtx[657]
  PIN BcidMtx[654]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9894.985 1046.435 9895.265 1047.435 ;
    END
  END BcidMtx[654]
  PIN Data_PMOS[1115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9853.545 1046.435 9853.825 1047.435 ;
    END
  END Data_PMOS[1115]
  PIN Data_PMOS[1123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9851.865 1046.435 9852.145 1047.435 ;
    END
  END Data_PMOS[1123]
  PIN Data_PMOS[1124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9850.185 1046.435 9850.465 1047.435 ;
    END
  END Data_PMOS[1124]
  PIN Data_PMOS[1130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9848.505 1046.435 9848.785 1047.435 ;
    END
  END Data_PMOS[1130]
  PIN MASKD[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9846.825 1046.435 9847.105 1047.435 ;
    END
  END MASKD[218]
  PIN DIG_MON_SEL[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9843.465 1046.435 9843.745 1047.435 ;
    END
  END DIG_MON_SEL[217]
  PIN DIG_MON_PMOS[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9841.225 1046.435 9841.505 1047.435 ;
    END
  END DIG_MON_PMOS[105]
  PIN Data_PMOS[1110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9830.585 1046.435 9830.865 1047.435 ;
    END
  END Data_PMOS[1110]
  PIN Data_PMOS[1097]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9828.345 1046.435 9828.625 1047.435 ;
    END
  END Data_PMOS[1097]
  PIN Data_PMOS[1106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9826.665 1046.435 9826.945 1047.435 ;
    END
  END Data_PMOS[1106]
  PIN Data_PMOS[1098]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9825.545 1046.435 9825.825 1047.435 ;
    END
  END Data_PMOS[1098]
  PIN BcidMtx[652]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9819.665 1046.435 9819.945 1047.435 ;
    END
  END BcidMtx[652]
  PIN Read_PMOS[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9792.505 1046.435 9792.785 1047.435 ;
    END
  END Read_PMOS[52]
  PIN BcidMtx[648]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9790.825 1046.435 9791.105 1047.435 ;
    END
  END BcidMtx[648]
  PIN Data_PMOS[1101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9787.465 1046.435 9787.745 1047.435 ;
    END
  END Data_PMOS[1101]
  PIN Data_PMOS[1102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9786.345 1046.435 9786.625 1047.435 ;
    END
  END Data_PMOS[1102]
  PIN Data_PMOS[1103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9784.665 1046.435 9784.945 1047.435 ;
    END
  END Data_PMOS[1103]
  PIN MASKV[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9782.425 1046.435 9782.705 1047.435 ;
    END
  END MASKV[216]
  PIN Data_HV[1087]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18663.465 1046.435 18663.745 1047.435 ;
    END
  END Data_HV[1087]
  PIN DIG_MON_PMOS[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9780.185 1046.435 9780.465 1047.435 ;
    END
  END DIG_MON_PMOS[104]
  PIN MASKD[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9763.945 1046.435 9764.225 1047.435 ;
    END
  END MASKD[215]
  PIN INJ_ROW[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9761.705 1046.435 9761.985 1047.435 ;
    END
  END INJ_ROW[107]
  PIN Data_PMOS[1079]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9760.025 1046.435 9760.305 1047.435 ;
    END
  END Data_PMOS[1079]
  PIN Data_PMOS[1084]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9757.785 1046.435 9758.065 1047.435 ;
    END
  END Data_PMOS[1084]
  PIN Data_PMOS[1085]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9756.665 1046.435 9756.945 1047.435 ;
    END
  END Data_PMOS[1085]
  PIN INJ_IN[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9754.425 1046.435 9754.705 1047.435 ;
    END
  END INJ_IN[215]
  PIN BcidMtx[645]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9711.865 1046.435 9712.145 1047.435 ;
    END
  END BcidMtx[645]
  PIN Read_PMOS[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9710.745 1046.435 9711.025 1047.435 ;
    END
  END Read_PMOS[51]
  PIN BcidMtx[642]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9709.065 1046.435 9709.345 1047.435 ;
    END
  END BcidMtx[642]
  PIN Data_PMOS[1080]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9705.705 1046.435 9705.985 1047.435 ;
    END
  END Data_PMOS[1080]
  PIN Data_PMOS[1081]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9704.585 1046.435 9704.865 1047.435 ;
    END
  END Data_PMOS[1081]
  PIN Data_PMOS[1082]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9702.905 1046.435 9703.185 1047.435 ;
    END
  END Data_PMOS[1082]
  PIN MASKV[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9692.265 1046.435 9692.545 1047.435 ;
    END
  END MASKV[214]
  PIN MASKD[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9691.145 1046.435 9691.425 1047.435 ;
    END
  END MASKD[214]
  PIN Data_HV[1055]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18639.105 1046.435 18639.385 1047.435 ;
    END
  END Data_HV[1055]
  PIN MASKD[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9686.665 1046.435 9686.945 1047.435 ;
    END
  END MASKD[213]
  PIN INJ_ROW[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9682.465 1046.435 9682.745 1047.435 ;
    END
  END INJ_ROW[106]
  PIN Data_PMOS[1068]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9681.345 1046.435 9681.625 1047.435 ;
    END
  END Data_PMOS[1068]
  PIN Data_PMOS[1069]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9679.665 1046.435 9679.945 1047.435 ;
    END
  END Data_PMOS[1069]
  PIN Data_PMOS[1064]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9651.945 1046.435 9652.225 1047.435 ;
    END
  END Data_PMOS[1064]
  PIN Data_PMOS[1056]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9650.825 1046.435 9651.105 1047.435 ;
    END
  END Data_PMOS[1056]
  PIN nTOK_PMOS[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9648.585 1046.435 9648.865 1047.435 ;
    END
  END nTOK_PMOS[50]
  PIN Read_PMOS[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9645.225 1046.435 9645.505 1047.435 ;
    END
  END Read_PMOS[50]
  PIN BcidMtx[637]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9644.105 1046.435 9644.385 1047.435 ;
    END
  END BcidMtx[637]
  PIN INJ_IN[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9642.425 1046.435 9642.705 1047.435 ;
    END
  END INJ_IN[212]
  PIN Data_PMOS[1060]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9626.185 1046.435 9626.465 1047.435 ;
    END
  END Data_PMOS[1060]
  PIN Data_PMOS[1066]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9625.065 1046.435 9625.345 1047.435 ;
    END
  END Data_PMOS[1066]
  PIN Data_PMOS[1051]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9623.945 1046.435 9624.225 1047.435 ;
    END
  END Data_PMOS[1051]
  PIN MASKD[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9621.145 1046.435 9621.425 1047.435 ;
    END
  END MASKD[212]
  PIN DIG_MON_PMOS[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9620.025 1046.435 9620.305 1047.435 ;
    END
  END DIG_MON_PMOS[100]
  PIN DIG_MON_SEL[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9618.345 1046.435 9618.625 1047.435 ;
    END
  END DIG_MON_SEL[212]
  PIN INJ_ROW[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9614.425 1046.435 9614.705 1047.435 ;
    END
  END INJ_ROW[105]
  PIN Data_PMOS[1047]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9573.545 1046.435 9573.825 1047.435 ;
    END
  END Data_PMOS[1047]
  PIN Data_PMOS[1041]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9572.425 1046.435 9572.705 1047.435 ;
    END
  END Data_PMOS[1041]
  PIN Data_PMOS[1049]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9570.185 1046.435 9570.465 1047.435 ;
    END
  END Data_PMOS[1049]
  PIN Data_PMOS[1036]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9569.065 1046.435 9569.345 1047.435 ;
    END
  END Data_PMOS[1036]
  PIN nTOK_PMOS[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9566.265 1046.435 9566.545 1047.435 ;
    END
  END nTOK_PMOS[49]
  PIN FREEZE_PMOS[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9563.465 1046.435 9563.745 1047.435 ;
    END
  END FREEZE_PMOS[49]
  PIN BcidMtx[632]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9562.345 1046.435 9562.625 1047.435 ;
    END
  END BcidMtx[632]
  PIN INJ_IN[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9551.705 1046.435 9551.985 1047.435 ;
    END
  END INJ_IN[210]
  PIN Data_PMOS[1044]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9548.905 1046.435 9549.185 1047.435 ;
    END
  END Data_PMOS[1044]
  PIN Data_PMOS[1033]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9547.785 1046.435 9548.065 1047.435 ;
    END
  END Data_PMOS[1033]
  PIN Data_PMOS[1030]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9546.105 1046.435 9546.385 1047.435 ;
    END
  END Data_PMOS[1030]
  PIN MASKH[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9541.905 1046.435 9542.185 1047.435 ;
    END
  END MASKH[105]
  PIN DIG_MON_PMOS[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9540.225 1046.435 9540.505 1047.435 ;
    END
  END DIG_MON_PMOS[98]
  PIN DIG_MON_SEL[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9538.545 1046.435 9538.825 1047.435 ;
    END
  END DIG_MON_SEL[210]
  PIN DIG_MON_COMP[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10629.705 1046.435 10629.985 1047.435 ;
    END
  END DIG_MON_COMP[13]
  PIN MASKV[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10628.025 1046.435 10628.305 1047.435 ;
    END
  END MASKV[237]
  PIN Data_COMP[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10626.345 1046.435 10626.625 1047.435 ;
    END
  END Data_COMP[138]
  PIN Data_COMP[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10623.545 1046.435 10623.825 1047.435 ;
    END
  END Data_COMP[140]
  PIN Data_COMP[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10622.425 1046.435 10622.705 1047.435 ;
    END
  END Data_COMP[132]
  PIN nTOK_COMP[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10620.185 1046.435 10620.465 1047.435 ;
    END
  END nTOK_COMP[6]
  PIN Read_COMP[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10603.385 1046.435 10603.665 1047.435 ;
    END
  END Read_COMP[6]
  PIN BcidMtx[709]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10602.265 1046.435 10602.545 1047.435 ;
    END
  END BcidMtx[709]
  PIN INJ_IN[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10600.585 1046.435 10600.865 1047.435 ;
    END
  END INJ_IN[236]
  PIN Data_COMP[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10597.225 1046.435 10597.505 1047.435 ;
    END
  END Data_COMP[136]
  PIN Data_COMP[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10596.105 1046.435 10596.385 1047.435 ;
    END
  END Data_COMP[142]
  PIN Data_COMP[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10594.985 1046.435 10595.265 1047.435 ;
    END
  END Data_COMP[127]
  PIN MASKD[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10553.545 1046.435 10553.825 1047.435 ;
    END
  END MASKD[236]
  PIN DIG_MON_SEL[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10550.185 1046.435 10550.465 1047.435 ;
    END
  END DIG_MON_SEL[235]
  PIN MASKV[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10546.265 1046.435 10546.545 1047.435 ;
    END
  END MASKV[235]
  PIN Data_COMP[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10545.145 1046.435 10545.425 1047.435 ;
    END
  END Data_COMP[113]
  PIN Data_COMP[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10544.025 1046.435 10544.305 1047.435 ;
    END
  END Data_COMP[124]
  PIN Data_COMP[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10541.225 1046.435 10541.505 1047.435 ;
    END
  END Data_COMP[112]
  PIN INJ_IN[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10531.145 1046.435 10531.425 1047.435 ;
    END
  END INJ_IN[235]
  PIN BcidMtx[707]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10528.905 1046.435 10529.185 1047.435 ;
    END
  END BcidMtx[707]
  PIN BcidMtx[704]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10526.105 1046.435 10526.385 1047.435 ;
    END
  END BcidMtx[704]
  PIN BcidMtx[702]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10524.985 1046.435 10525.265 1047.435 ;
    END
  END BcidMtx[702]
  PIN Data_COMP[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10520.785 1046.435 10521.065 1047.435 ;
    END
  END Data_COMP[108]
  PIN Data_COMP[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10492.505 1046.435 10492.785 1047.435 ;
    END
  END Data_COMP[109]
  PIN Data_COMP[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10491.385 1046.435 10491.665 1047.435 ;
    END
  END Data_COMP[116]
  PIN Data_COMP[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10490.265 1046.435 10490.545 1047.435 ;
    END
  END Data_COMP[105]
  PIN DIG_MON_COMP[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10486.905 1046.435 10487.185 1047.435 ;
    END
  END DIG_MON_COMP[10]
  PIN DIG_MON_SEL[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10485.225 1046.435 10485.505 1047.435 ;
    END
  END DIG_MON_SEL[234]
  PIN DIG_MON_COMP[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10482.425 1046.435 10482.705 1047.435 ;
    END
  END DIG_MON_COMP[9]
  PIN MASKV[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11040.745 1046.435 11041.025 1047.435 ;
    END
  END MASKV[247]
  PIN Data_COMP[243]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11026.185 1046.435 11026.465 1047.435 ;
    END
  END Data_COMP[243]
  PIN Data_COMP[236]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11025.065 1046.435 11025.345 1047.435 ;
    END
  END Data_COMP[236]
  PIN Data_COMP[238]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11022.825 1046.435 11023.105 1047.435 ;
    END
  END Data_COMP[238]
  PIN nTOK_COMP[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11020.025 1046.435 11020.305 1047.435 ;
    END
  END nTOK_COMP[11]
  PIN BcidMtx[742]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11018.345 1046.435 11018.625 1047.435 ;
    END
  END BcidMtx[742]
  PIN BcidMtx[740]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11016.105 1046.435 11016.385 1047.435 ;
    END
  END BcidMtx[740]
  PIN INJ_IN[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11013.865 1046.435 11014.145 1047.435 ;
    END
  END INJ_IN[246]
  PIN Data_COMP[233]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10973.545 1046.435 10973.825 1047.435 ;
    END
  END Data_COMP[233]
  PIN Data_COMP[235]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10971.305 1046.435 10971.585 1047.435 ;
    END
  END Data_COMP[235]
  PIN Data_COMP[232]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10969.625 1046.435 10969.905 1047.435 ;
    END
  END Data_COMP[232]
  PIN Data_COMP[248]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10968.505 1046.435 10968.785 1047.435 ;
    END
  END Data_COMP[248]
  PIN MASKD[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10966.825 1046.435 10967.105 1047.435 ;
    END
  END MASKD[246]
  PIN DIG_MON_SEL[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10963.465 1046.435 10963.745 1047.435 ;
    END
  END DIG_MON_SEL[245]
  PIN DIG_MON_COMP[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10961.225 1046.435 10961.505 1047.435 ;
    END
  END DIG_MON_COMP[21]
  PIN Data_COMP[218]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10950.025 1046.435 10950.305 1047.435 ;
    END
  END Data_COMP[218]
  PIN Data_COMP[215]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10948.345 1046.435 10948.625 1047.435 ;
    END
  END Data_COMP[215]
  PIN Data_COMP[230]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10947.225 1046.435 10947.505 1047.435 ;
    END
  END Data_COMP[230]
  PIN INJ_IN[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10942.465 1046.435 10942.745 1047.435 ;
    END
  END INJ_IN[245]
  PIN BcidMtx[736]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10939.665 1046.435 10939.945 1047.435 ;
    END
  END BcidMtx[736]
  PIN Read_COMP[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10912.505 1046.435 10912.785 1047.435 ;
    END
  END Read_COMP[10]
  PIN Data_HV[1082]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18662.905 1046.435 18663.185 1047.435 ;
    END
  END Data_HV[1082]
  PIN Data_COMP[213]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10908.585 1046.435 10908.865 1047.435 ;
    END
  END Data_COMP[213]
  PIN Data_COMP[219]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10907.465 1046.435 10907.745 1047.435 ;
    END
  END Data_COMP[219]
  PIN Data_COMP[226]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10905.225 1046.435 10905.505 1047.435 ;
    END
  END Data_COMP[226]
  PIN Data_COMP[210]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10903.545 1046.435 10903.825 1047.435 ;
    END
  END Data_COMP[210]
  PIN MASKV[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10902.425 1046.435 10902.705 1047.435 ;
    END
  END MASKV[244]
  PIN MASKD[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10883.945 1046.435 10884.225 1047.435 ;
    END
  END MASKD[243]
  PIN INJ_ROW[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10881.705 1046.435 10881.985 1047.435 ;
    END
  END INJ_ROW[121]
  PIN Data_COMP[201]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10879.465 1046.435 10879.745 1047.435 ;
    END
  END Data_COMP[201]
  PIN Data_COMP[202]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10877.785 1046.435 10878.065 1047.435 ;
    END
  END Data_COMP[202]
  PIN Data_COMP[203]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10876.665 1046.435 10876.945 1047.435 ;
    END
  END Data_COMP[203]
  PIN nTOK_COMP[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10834.105 1046.435 10834.385 1047.435 ;
    END
  END nTOK_COMP[9]
  PIN BcidMtx[729]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10831.865 1046.435 10832.145 1047.435 ;
    END
  END BcidMtx[729]
  PIN Read_COMP[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10830.745 1046.435 10831.025 1047.435 ;
    END
  END Read_COMP[9]
  PIN INJ_IN[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10827.945 1046.435 10828.225 1047.435 ;
    END
  END INJ_IN[242]
  PIN Data_COMP[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10826.265 1046.435 10826.545 1047.435 ;
    END
  END Data_COMP[191]
  PIN Data_HV[1064]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18611.945 1046.435 18612.225 1047.435 ;
    END
  END Data_HV[1064]
  PIN Data_COMP[205]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10823.465 1046.435 10823.745 1047.435 ;
    END
  END Data_COMP[205]
  PIN Data_COMP[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10821.785 1046.435 10822.065 1047.435 ;
    END
  END Data_COMP[189]
  PIN MASKV[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10812.265 1046.435 10812.545 1047.435 ;
    END
  END MASKV[242]
  PIN MASKD[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10806.665 1046.435 10806.945 1047.435 ;
    END
  END MASKD[241]
  PIN INJ_ROW[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10802.465 1046.435 10802.745 1047.435 ;
    END
  END INJ_ROW[120]
  PIN Data_COMP[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10800.225 1046.435 10800.505 1047.435 ;
    END
  END Data_COMP[180]
  PIN Data_COMP[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10773.065 1046.435 10773.345 1047.435 ;
    END
  END Data_COMP[181]
  PIN Data_COMP[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10771.945 1046.435 10772.225 1047.435 ;
    END
  END Data_COMP[182]
  PIN nTOK_COMP[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10768.585 1046.435 10768.865 1047.435 ;
    END
  END nTOK_COMP[8]
  PIN BcidMtx[723]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10766.345 1046.435 10766.625 1047.435 ;
    END
  END BcidMtx[723]
  PIN Read_COMP[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10765.225 1046.435 10765.505 1047.435 ;
    END
  END Read_COMP[8]
  PIN INJ_IN[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10762.425 1046.435 10762.705 1047.435 ;
    END
  END INJ_IN[240]
  PIN Data_COMP[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10760.745 1046.435 10761.025 1047.435 ;
    END
  END Data_COMP[170]
  PIN Data_COMP[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10746.745 1046.435 10747.025 1047.435 ;
    END
  END Data_COMP[183]
  PIN INJ_IN[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18782.465 1046.435 18782.745 1047.435 ;
    END
  END INJ_IN[441]
  PIN Data_COMP[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10743.945 1046.435 10744.225 1047.435 ;
    END
  END Data_COMP[169]
  PIN Data_COMP[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10742.825 1046.435 10743.105 1047.435 ;
    END
  END Data_COMP[185]
  PIN DIG_MON_COMP[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10740.025 1046.435 10740.305 1047.435 ;
    END
  END DIG_MON_COMP[16]
  PIN DIG_MON_SEL[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10737.785 1046.435 10738.065 1047.435 ;
    END
  END DIG_MON_SEL[239]
  PIN DIG_MON_COMP[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10735.545 1046.435 10735.825 1047.435 ;
    END
  END DIG_MON_COMP[15]
  PIN Data_COMP[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10692.985 1046.435 10693.265 1047.435 ;
    END
  END Data_COMP[155]
  PIN Data_COMP[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10691.305 1046.435 10691.585 1047.435 ;
    END
  END Data_COMP[152]
  PIN Data_COMP[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10690.185 1046.435 10690.465 1047.435 ;
    END
  END Data_COMP[167]
  PIN INJ_IN[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10687.385 1046.435 10687.665 1047.435 ;
    END
  END INJ_IN[239]
  PIN BcidMtx[718]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10684.585 1046.435 10684.865 1047.435 ;
    END
  END BcidMtx[718]
  PIN FREEZE_COMP[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10683.465 1046.435 10683.745 1047.435 ;
    END
  END FREEZE_COMP[7]
  PIN BcidMtx[714]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10681.225 1046.435 10681.505 1047.435 ;
    END
  END BcidMtx[714]
  PIN Data_COMP[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10670.025 1046.435 10670.305 1047.435 ;
    END
  END Data_COMP[149]
  PIN Data_COMP[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10668.905 1046.435 10669.185 1047.435 ;
    END
  END Data_COMP[162]
  PIN Data_COMP[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10666.665 1046.435 10666.945 1047.435 ;
    END
  END Data_COMP[158]
  PIN Data_COMP[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10664.985 1046.435 10665.265 1047.435 ;
    END
  END Data_COMP[164]
  PIN MASKH[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10661.905 1046.435 10662.185 1047.435 ;
    END
  END MASKH[119]
  PIN DIG_MON_SEL[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10658.545 1046.435 10658.825 1047.435 ;
    END
  END DIG_MON_SEL[238]
  PIN MASKD[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11750.825 1046.435 11751.105 1047.435 ;
    END
  END MASKD[265]
  PIN INJ_ROW[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11748.585 1046.435 11748.865 1047.435 ;
    END
  END INJ_ROW[132]
  PIN Data_COMP[432]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11746.345 1046.435 11746.625 1047.435 ;
    END
  END Data_COMP[432]
  PIN Data_COMP[433]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11744.665 1046.435 11744.945 1047.435 ;
    END
  END Data_COMP[433]
  PIN Data_COMP[434]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11743.545 1046.435 11743.825 1047.435 ;
    END
  END Data_COMP[434]
  PIN nTOK_COMP[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11740.185 1046.435 11740.465 1047.435 ;
    END
  END nTOK_COMP[20]
  PIN BcidMtx[795]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11724.505 1046.435 11724.785 1047.435 ;
    END
  END BcidMtx[795]
  PIN Read_COMP[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11723.385 1046.435 11723.665 1047.435 ;
    END
  END Read_COMP[20]
  PIN INJ_IN[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11720.585 1046.435 11720.865 1047.435 ;
    END
  END INJ_IN[264]
  PIN Data_COMP[429]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11718.345 1046.435 11718.625 1047.435 ;
    END
  END Data_COMP[429]
  PIN Data_COMP[430]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11717.225 1046.435 11717.505 1047.435 ;
    END
  END Data_COMP[430]
  PIN Data_COMP[421]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11714.985 1046.435 11715.265 1047.435 ;
    END
  END Data_COMP[421]
  PIN MASKV[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11674.665 1046.435 11674.945 1047.435 ;
    END
  END MASKV[264]
  PIN MASKD[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11673.545 1046.435 11673.825 1047.435 ;
    END
  END MASKD[264]
  PIN DIG_MON_SEL[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11670.185 1046.435 11670.465 1047.435 ;
    END
  END DIG_MON_SEL[263]
  PIN INJ_ROW[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11666.825 1046.435 11667.105 1047.435 ;
    END
  END INJ_ROW[131]
  PIN Data_COMP[417]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11665.705 1046.435 11665.985 1047.435 ;
    END
  END Data_COMP[417]
  PIN Data_COMP[404]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11663.465 1046.435 11663.745 1047.435 ;
    END
  END Data_COMP[404]
  PIN Data_COMP[413]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11661.785 1046.435 11662.065 1047.435 ;
    END
  END Data_COMP[413]
  PIN Data_COMP[405]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11652.265 1046.435 11652.545 1047.435 ;
    END
  END Data_COMP[405]
  PIN BcidMtx[790]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11648.345 1046.435 11648.625 1047.435 ;
    END
  END BcidMtx[790]
  PIN Read_COMP[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11646.665 1046.435 11646.945 1047.435 ;
    END
  END Read_COMP[19]
  PIN BcidMtx[787]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11645.545 1046.435 11645.825 1047.435 ;
    END
  END BcidMtx[787]
  PIN Data_COMP[401]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11640.225 1046.435 11640.505 1047.435 ;
    END
  END Data_COMP[401]
  PIN Data_COMP[409]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11638.545 1046.435 11638.825 1047.435 ;
    END
  END Data_COMP[409]
  PIN Data_COMP[415]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11611.945 1046.435 11612.225 1047.435 ;
    END
  END Data_COMP[415]
  PIN Data_COMP[416]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11609.705 1046.435 11609.985 1047.435 ;
    END
  END Data_COMP[416]
  PIN MASKD[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11608.025 1046.435 11608.305 1047.435 ;
    END
  END MASKD[262]
  PIN Data_COMP[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10466.185 1046.435 10466.465 1047.435 ;
    END
  END Data_COMP[96]
  PIN Data_COMP[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10465.625 1046.435 10465.905 1047.435 ;
    END
  END Data_COMP[103]
  PIN Data_COMP[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10463.945 1046.435 10464.225 1047.435 ;
    END
  END Data_COMP[104]
  PIN nTOK_COMP[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10460.025 1046.435 10460.305 1047.435 ;
    END
  END nTOK_COMP[4]
  PIN BcidMtx[700]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10458.345 1046.435 10458.625 1047.435 ;
    END
  END BcidMtx[700]
  PIN FREEZE_COMP[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10457.225 1046.435 10457.505 1047.435 ;
    END
  END FREEZE_COMP[4]
  PIN INJ_IN[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10453.865 1046.435 10454.145 1047.435 ;
    END
  END INJ_IN[232]
  PIN Data_COMP[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10413.545 1046.435 10413.825 1047.435 ;
    END
  END Data_COMP[86]
  PIN Data_COMP[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10412.425 1046.435 10412.705 1047.435 ;
    END
  END Data_COMP[99]
  PIN Data_COMP[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10409.625 1046.435 10409.905 1047.435 ;
    END
  END Data_COMP[85]
  PIN Data_COMP[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10408.505 1046.435 10408.785 1047.435 ;
    END
  END Data_COMP[101]
  PIN MASKH[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10407.385 1046.435 10407.665 1047.435 ;
    END
  END MASKH[116]
  PIN DIG_MON_SEL[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10403.465 1046.435 10403.745 1047.435 ;
    END
  END DIG_MON_SEL[231]
  PIN DIG_MON_COMP[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10401.225 1046.435 10401.505 1047.435 ;
    END
  END DIG_MON_COMP[7]
  PIN MASKV[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10391.145 1046.435 10391.425 1047.435 ;
    END
  END MASKV[231]
  PIN Data_COMP[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10388.345 1046.435 10388.625 1047.435 ;
    END
  END Data_COMP[68]
  PIN Data_COMP[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10387.225 1046.435 10387.505 1047.435 ;
    END
  END Data_COMP[83]
  PIN Data_COMP[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10386.105 1046.435 10386.385 1047.435 ;
    END
  END Data_COMP[70]
  PIN BcidMtx[694]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10379.665 1046.435 10379.945 1047.435 ;
    END
  END BcidMtx[694]
  PIN Read_COMP[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10352.505 1046.435 10352.785 1047.435 ;
    END
  END Read_COMP[3]
  PIN BcidMtx[691]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10351.385 1046.435 10351.665 1047.435 ;
    END
  END BcidMtx[691]
  PIN Data_COMP[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10347.465 1046.435 10347.745 1047.435 ;
    END
  END Data_COMP[72]
  PIN Data_COMP[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10346.345 1046.435 10346.625 1047.435 ;
    END
  END Data_COMP[73]
  PIN Data_COMP[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10345.785 1046.435 10346.065 1047.435 ;
    END
  END Data_COMP[67]
  PIN Data_COMP[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10342.985 1046.435 10343.265 1047.435 ;
    END
  END Data_COMP[80]
  PIN MASKH[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10341.865 1046.435 10342.145 1047.435 ;
    END
  END MASKH[115]
  PIN DIG_MON_COMP[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10340.185 1046.435 10340.465 1047.435 ;
    END
  END DIG_MON_COMP[6]
  PIN DIG_MON_COMP[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10322.825 1046.435 10323.105 1047.435 ;
    END
  END DIG_MON_COMP[5]
  PIN MASKV[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10321.145 1046.435 10321.425 1047.435 ;
    END
  END MASKV[229]
  PIN Data_COMP[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10320.025 1046.435 10320.305 1047.435 ;
    END
  END Data_COMP[50]
  PIN Data_COMP[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10317.225 1046.435 10317.505 1047.435 ;
    END
  END Data_COMP[62]
  PIN Data_COMP[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10316.105 1046.435 10316.385 1047.435 ;
    END
  END Data_COMP[49]
  PIN INJ_IN[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10314.425 1046.435 10314.705 1047.435 ;
    END
  END INJ_IN[229]
  PIN FREEZE_COMP[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10271.305 1046.435 10271.585 1047.435 ;
    END
  END FREEZE_COMP[2]
  PIN BcidMtx[686]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10270.185 1046.435 10270.465 1047.435 ;
    END
  END BcidMtx[686]
  PIN BcidMtx[684]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10269.065 1046.435 10269.345 1047.435 ;
    END
  END BcidMtx[684]
  PIN Data_COMP[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10265.705 1046.435 10265.985 1047.435 ;
    END
  END Data_COMP[51]
  PIN Data_COMP[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10264.025 1046.435 10264.305 1047.435 ;
    END
  END Data_COMP[46]
  PIN Data_HV[1111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18788.905 1046.435 18789.185 1047.435 ;
    END
  END Data_HV[1111]
  PIN Data_COMP[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10261.225 1046.435 10261.505 1047.435 ;
    END
  END Data_COMP[59]
  PIN MASKH[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10251.705 1046.435 10251.985 1047.435 ;
    END
  END MASKH[114]
  PIN DIG_MON_COMP[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10250.025 1046.435 10250.305 1047.435 ;
    END
  END DIG_MON_COMP[4]
  PIN MASKD[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10246.665 1046.435 10246.945 1047.435 ;
    END
  END MASKD[227]
  PIN MASKV[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10241.905 1046.435 10242.185 1047.435 ;
    END
  END MASKV[227]
  PIN Data_COMP[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10240.785 1046.435 10241.065 1047.435 ;
    END
  END Data_COMP[29]
  PIN Data_COMP[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10213.065 1046.435 10213.345 1047.435 ;
    END
  END Data_COMP[34]
  PIN Data_COMP[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10211.385 1046.435 10211.665 1047.435 ;
    END
  END Data_COMP[28]
  PIN INJ_IN[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10209.705 1046.435 10209.985 1047.435 ;
    END
  END INJ_IN[227]
  PIN BcidMtx[682]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10206.905 1046.435 10207.185 1047.435 ;
    END
  END BcidMtx[682]
  PIN Read_COMP[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10205.225 1046.435 10205.505 1047.435 ;
    END
  END Read_COMP[1]
  PIN BcidMtx[679]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10204.105 1046.435 10204.385 1047.435 ;
    END
  END BcidMtx[679]
  PIN Data_COMP[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10200.745 1046.435 10201.025 1047.435 ;
    END
  END Data_COMP[23]
  PIN Data_COMP[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10186.185 1046.435 10186.465 1047.435 ;
    END
  END Data_COMP[31]
  PIN Data_COMP[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10185.065 1046.435 10185.345 1047.435 ;
    END
  END Data_COMP[37]
  PIN Data_COMP[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10183.385 1046.435 10183.665 1047.435 ;
    END
  END Data_COMP[21]
  PIN MASKH[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10181.705 1046.435 10181.985 1047.435 ;
    END
  END MASKH[113]
  PIN Data_HV[1112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18787.225 1046.435 18787.505 1047.435 ;
    END
  END Data_HV[1112]
  PIN DIG_MON_SEL[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10177.785 1046.435 10178.065 1047.435 ;
    END
  END DIG_MON_SEL[225]
  PIN INJ_ROW[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10174.425 1046.435 10174.705 1047.435 ;
    END
  END INJ_ROW[112]
  PIN Data_COMP[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10133.545 1046.435 10133.825 1047.435 ;
    END
  END Data_COMP[18]
  PIN Data_COMP[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10131.305 1046.435 10131.585 1047.435 ;
    END
  END Data_COMP[5]
  PIN Data_COMP[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10129.625 1046.435 10129.905 1047.435 ;
    END
  END Data_COMP[14]
  PIN Data_COMP[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10128.505 1046.435 10128.785 1047.435 ;
    END
  END Data_COMP[6]
  PIN BcidMtx[675]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10124.025 1046.435 10124.305 1047.435 ;
    END
  END BcidMtx[675]
  PIN BcidMtx[674]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10122.345 1046.435 10122.625 1047.435 ;
    END
  END BcidMtx[674]
  PIN BcidMtx[672]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10121.225 1046.435 10121.505 1047.435 ;
    END
  END BcidMtx[672]
  PIN Data_COMP[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10109.465 1046.435 10109.745 1047.435 ;
    END
  END Data_COMP[9]
  PIN Data_COMP[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10107.785 1046.435 10108.065 1047.435 ;
    END
  END Data_COMP[4]
  PIN Data_COMP[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10106.665 1046.435 10106.945 1047.435 ;
    END
  END Data_COMP[11]
  PIN MASKV[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10102.465 1046.435 10102.745 1047.435 ;
    END
  END MASKV[224]
  PIN DIG_MON_COMP[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10100.225 1046.435 10100.505 1047.435 ;
    END
  END DIG_MON_COMP[0]
  PIN DIG_MON_SEL[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10098.545 1046.435 10098.825 1047.435 ;
    END
  END DIG_MON_SEL[224]
  PIN DIG_MON_COMP[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11189.705 1046.435 11189.985 1047.435 ;
    END
  END DIG_MON_COMP[27]
  PIN Data_COMP[291]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11187.465 1046.435 11187.745 1047.435 ;
    END
  END Data_COMP[291]
  PIN Data_COMP[285]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11186.345 1046.435 11186.625 1047.435 ;
    END
  END Data_COMP[285]
  PIN Data_COMP[293]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11184.105 1046.435 11184.385 1047.435 ;
    END
  END Data_COMP[293]
  PIN Data_COMP[279]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11182.425 1046.435 11182.705 1047.435 ;
    END
  END Data_COMP[279]
  PIN nTOK_COMP[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11180.185 1046.435 11180.465 1047.435 ;
    END
  END nTOK_COMP[13]
  PIN FREEZE_COMP[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11163.945 1046.435 11164.225 1047.435 ;
    END
  END FREEZE_COMP[13]
  PIN BcidMtx[751]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11162.265 1046.435 11162.545 1047.435 ;
    END
  END BcidMtx[751]
  PIN INJ_IN[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11160.585 1046.435 11160.865 1047.435 ;
    END
  END INJ_IN[250]
  PIN Data_COMP[288]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11157.785 1046.435 11158.065 1047.435 ;
    END
  END Data_COMP[288]
  PIN Data_COMP[289]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11156.105 1046.435 11156.385 1047.435 ;
    END
  END Data_COMP[289]
  PIN Data_COMP[274]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11154.985 1046.435 11155.265 1047.435 ;
    END
  END Data_COMP[274]
  PIN Data_HV[1106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18786.665 1046.435 18786.945 1047.435 ;
    END
  END Data_HV[1106]
  PIN MASKD[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11113.545 1046.435 11113.825 1047.435 ;
    END
  END MASKD[250]
  PIN DIG_MON_COMP[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11107.945 1046.435 11108.225 1047.435 ;
    END
  END DIG_MON_COMP[25]
  PIN MASKV[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11106.265 1046.435 11106.545 1047.435 ;
    END
  END MASKV[249]
  PIN Data_COMP[260]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11105.145 1046.435 11105.425 1047.435 ;
    END
  END Data_COMP[260]
  PIN Data_COMP[272]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11102.345 1046.435 11102.625 1047.435 ;
    END
  END Data_COMP[272]
  PIN Data_COMP[258]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11092.265 1046.435 11092.545 1047.435 ;
    END
  END Data_COMP[258]
  PIN nTOK_COMP[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11090.025 1046.435 11090.305 1047.435 ;
    END
  END nTOK_COMP[12]
  PIN FREEZE_COMP[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11087.225 1046.435 11087.505 1047.435 ;
    END
  END FREEZE_COMP[12]
  PIN BcidMtx[745]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11085.545 1046.435 11085.825 1047.435 ;
    END
  END BcidMtx[745]
  PIN INJ_IN[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11081.905 1046.435 11082.185 1047.435 ;
    END
  END INJ_IN[248]
  PIN Data_COMP[267]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11079.105 1046.435 11079.385 1047.435 ;
    END
  END Data_COMP[267]
  PIN Data_COMP[268]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11051.945 1046.435 11052.225 1047.435 ;
    END
  END Data_COMP[268]
  PIN Data_COMP[253]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11050.825 1046.435 11051.105 1047.435 ;
    END
  END Data_COMP[253]
  PIN MASKH[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11048.585 1046.435 11048.865 1047.435 ;
    END
  END MASKH[124]
  PIN DIG_MON_SEL[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11044.665 1046.435 11044.945 1047.435 ;
    END
  END DIG_MON_SEL[247]
  PIN Data_COMP[987]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13850.265 1046.435 13850.545 1047.435 ;
    END
  END Data_COMP[987]
  PIN MASKD[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13848.025 1046.435 13848.305 1047.435 ;
    END
  END MASKD[318]
  PIN DIG_MON_SEL[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13845.225 1046.435 13845.505 1047.435 ;
    END
  END DIG_MON_SEL[318]
  PIN MASKD[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13843.545 1046.435 13843.825 1047.435 ;
    END
  END MASKD[317]
  PIN Data_COMP[984]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13840.185 1046.435 13840.465 1047.435 ;
    END
  END Data_COMP[984]
  PIN Data_COMP[985]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13825.625 1046.435 13825.905 1047.435 ;
    END
  END Data_COMP[985]
  PIN Data_COMP[979]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13824.505 1046.435 13824.785 1047.435 ;
    END
  END Data_COMP[979]
  PIN Data_COMP[972]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13822.265 1046.435 13822.545 1047.435 ;
    END
  END Data_COMP[972]
  PIN BcidMtx[953]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13818.905 1046.435 13819.185 1047.435 ;
    END
  END BcidMtx[953]
  PIN BcidMtx[951]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13817.785 1046.435 13818.065 1047.435 ;
    END
  END BcidMtx[951]
  PIN BcidMtx[949]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13815.545 1046.435 13815.825 1047.435 ;
    END
  END BcidMtx[949]
  PIN Data_COMP[969]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13774.105 1046.435 13774.385 1047.435 ;
    END
  END Data_COMP[969]
  PIN Data_COMP[975]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13772.985 1046.435 13773.265 1047.435 ;
    END
  END Data_COMP[975]
  PIN Data_COMP[982]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13770.745 1046.435 13771.025 1047.435 ;
    END
  END Data_COMP[982]
  PIN Data_COMP[966]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13769.065 1046.435 13769.345 1047.435 ;
    END
  END Data_COMP[966]
  PIN MASKV[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13767.945 1046.435 13768.225 1047.435 ;
    END
  END MASKV[316]
  PIN MASKD[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13762.345 1046.435 13762.625 1047.435 ;
    END
  END MASKD[315]
  PIN INJ_ROW[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13751.705 1046.435 13751.985 1047.435 ;
    END
  END INJ_ROW[157]
  PIN Data_COMP[957]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13749.465 1046.435 13749.745 1047.435 ;
    END
  END Data_COMP[957]
  PIN Data_COMP[958]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13747.785 1046.435 13748.065 1047.435 ;
    END
  END Data_COMP[958]
  PIN Data_COMP[959]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13746.665 1046.435 13746.945 1047.435 ;
    END
  END Data_COMP[959]
  PIN nTOK_COMP[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13741.345 1046.435 13741.625 1047.435 ;
    END
  END nTOK_COMP[45]
  PIN BcidMtx[945]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13739.105 1046.435 13739.385 1047.435 ;
    END
  END BcidMtx[945]
  PIN BcidMtx[944]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13711.945 1046.435 13712.225 1047.435 ;
    END
  END BcidMtx[944]
  PIN Data_COMP[948]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13708.585 1046.435 13708.865 1047.435 ;
    END
  END Data_COMP[948]
  PIN Data_COMP[960]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13706.905 1046.435 13707.185 1047.435 ;
    END
  END Data_COMP[960]
  PIN Data_COMP[949]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13705.785 1046.435 13706.065 1047.435 ;
    END
  END Data_COMP[949]
  PIN Data_COMP[945]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13703.545 1046.435 13703.825 1047.435 ;
    END
  END Data_COMP[945]
  PIN MASKH[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13701.865 1046.435 13702.145 1047.435 ;
    END
  END MASKH[157]
  PIN DIG_MON_COMP[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13700.185 1046.435 13700.465 1047.435 ;
    END
  END DIG_MON_COMP[90]
  PIN DIG_MON_SEL[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13685.065 1046.435 13685.345 1047.435 ;
    END
  END DIG_MON_SEL[313]
  PIN DIG_MON_COMP[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13682.825 1046.435 13683.105 1047.435 ;
    END
  END DIG_MON_COMP[89]
  PIN MASKV[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13681.145 1046.435 13681.425 1047.435 ;
    END
  END MASKV[313]
  PIN Data_COMP[943]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13678.905 1046.435 13679.185 1047.435 ;
    END
  END Data_COMP[943]
  PIN Data_COMP[944]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13677.225 1046.435 13677.505 1047.435 ;
    END
  END Data_COMP[944]
  PIN Data_COMP[931]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13676.105 1046.435 13676.385 1047.435 ;
    END
  END Data_COMP[931]
  PIN BcidMtx[941]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13632.985 1046.435 13633.265 1047.435 ;
    END
  END BcidMtx[941]
  PIN FREEZE_COMP[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13631.305 1046.435 13631.585 1047.435 ;
    END
  END FREEZE_COMP[44]
  PIN BcidMtx[938]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13630.185 1046.435 13630.465 1047.435 ;
    END
  END BcidMtx[938]
  PIN Data_COMP[927]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13626.825 1046.435 13627.105 1047.435 ;
    END
  END Data_COMP[927]
  PIN Data_COMP[939]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13625.145 1046.435 13625.425 1047.435 ;
    END
  END Data_COMP[939]
  PIN Data_COMP[928]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13624.025 1046.435 13624.305 1047.435 ;
    END
  END Data_COMP[928]
  PIN Data_COMP[924]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13621.785 1046.435 13622.065 1047.435 ;
    END
  END Data_COMP[924]
  PIN MASKH[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13611.705 1046.435 13611.985 1047.435 ;
    END
  END MASKH[156]
  PIN DIG_MON_COMP[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13610.025 1046.435 13610.305 1047.435 ;
    END
  END DIG_MON_COMP[88]
  PIN DIG_MON_SEL[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13607.785 1046.435 13608.065 1047.435 ;
    END
  END DIG_MON_SEL[311]
  PIN DIG_MON_COMP[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13605.545 1046.435 13605.825 1047.435 ;
    END
  END DIG_MON_COMP[87]
  PIN MASKV[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13601.905 1046.435 13602.185 1047.435 ;
    END
  END MASKV[311]
  PIN Data_COMP[922]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13599.665 1046.435 13599.945 1047.435 ;
    END
  END Data_COMP[922]
  PIN Data_COMP[923]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13572.505 1046.435 13572.785 1047.435 ;
    END
  END Data_COMP[923]
  PIN Data_COMP[910]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13571.385 1046.435 13571.665 1047.435 ;
    END
  END Data_COMP[910]
  PIN BcidMtx[935]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13567.465 1046.435 13567.745 1047.435 ;
    END
  END BcidMtx[935]
  PIN FREEZE_COMP[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13565.785 1046.435 13566.065 1047.435 ;
    END
  END FREEZE_COMP[43]
  PIN BcidMtx[932]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13564.665 1046.435 13564.945 1047.435 ;
    END
  END BcidMtx[932]
  PIN Data_COMP[906]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13561.305 1046.435 13561.585 1047.435 ;
    END
  END Data_COMP[906]
  PIN Data_COMP[918]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13546.745 1046.435 13547.025 1047.435 ;
    END
  END Data_COMP[918]
  PIN Data_COMP[907]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13545.625 1046.435 13545.905 1047.435 ;
    END
  END Data_COMP[907]
  PIN Data_COMP[903]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13543.385 1046.435 13543.665 1047.435 ;
    END
  END Data_COMP[903]
  PIN MASKH[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13541.705 1046.435 13541.985 1047.435 ;
    END
  END MASKH[155]
  PIN DIG_MON_COMP[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13540.025 1046.435 13540.305 1047.435 ;
    END
  END DIG_MON_COMP[86]
  PIN MASKD[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18741.305 1046.435 18741.585 1047.435 ;
    END
  END MASKD[440]
  PIN INJ_ROW[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13534.425 1046.435 13534.705 1047.435 ;
    END
  END INJ_ROW[154]
  PIN Data_COMP[900]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13493.545 1046.435 13493.825 1047.435 ;
    END
  END Data_COMP[900]
  PIN Data_COMP[887]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13491.305 1046.435 13491.585 1047.435 ;
    END
  END Data_COMP[887]
  PIN Data_COMP[896]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13489.625 1046.435 13489.905 1047.435 ;
    END
  END Data_COMP[896]
  PIN Data_COMP[888]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13488.505 1046.435 13488.785 1047.435 ;
    END
  END Data_COMP[888]
  PIN BcidMtx[928]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13484.585 1046.435 13484.865 1047.435 ;
    END
  END BcidMtx[928]
  PIN BcidMtx[926]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13482.345 1046.435 13482.625 1047.435 ;
    END
  END BcidMtx[926]
  PIN BcidMtx[924]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13481.225 1046.435 13481.505 1047.435 ;
    END
  END BcidMtx[924]
  PIN Data_COMP[885]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13470.585 1046.435 13470.865 1047.435 ;
    END
  END Data_COMP[885]
  PIN Data_COMP[886]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13467.785 1046.435 13468.065 1047.435 ;
    END
  END Data_COMP[886]
  PIN Data_COMP[898]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13467.225 1046.435 13467.505 1047.435 ;
    END
  END Data_COMP[898]
  PIN Data_COMP[882]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13465.545 1046.435 13465.825 1047.435 ;
    END
  END Data_COMP[882]
  PIN MASKD[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13461.345 1046.435 13461.625 1047.435 ;
    END
  END MASKD[308]
  PIN DIG_MON_SEL[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14551.945 1046.435 14552.225 1047.435 ;
    END
  END DIG_MON_SEL[335]
  PIN INJ_ROW[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14548.585 1046.435 14548.865 1047.435 ;
    END
  END INJ_ROW[167]
  PIN Data_COMP[1173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14547.465 1046.435 14547.745 1047.435 ;
    END
  END Data_COMP[1173]
  PIN Data_COMP[1174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14545.785 1046.435 14546.065 1047.435 ;
    END
  END Data_COMP[1174]
  PIN Data_COMP[1162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14542.985 1046.435 14543.265 1047.435 ;
    END
  END Data_COMP[1162]
  PIN nTOK_COMP[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14540.185 1046.435 14540.465 1047.435 ;
    END
  END nTOK_COMP[55]
  PIN BcidMtx[1005]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14524.505 1046.435 14524.785 1047.435 ;
    END
  END BcidMtx[1005]
  PIN BcidMtx[1004]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14522.825 1046.435 14523.105 1047.435 ;
    END
  END BcidMtx[1004]
  PIN INJ_IN[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14520.585 1046.435 14520.865 1047.435 ;
    END
  END INJ_IN[334]
  PIN Data_COMP[1164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14518.345 1046.435 14518.625 1047.435 ;
    END
  END Data_COMP[1164]
  PIN Data_COMP[1159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14516.665 1046.435 14516.945 1047.435 ;
    END
  END Data_COMP[1159]
  PIN Data_COMP[1156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14514.985 1046.435 14515.265 1047.435 ;
    END
  END Data_COMP[1156]
  PIN MASKV[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14474.665 1046.435 14474.945 1047.435 ;
    END
  END MASKV[334]
  PIN DIG_MON_COMP[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14472.425 1046.435 14472.705 1047.435 ;
    END
  END DIG_MON_COMP[110]
  PIN DIG_MON_SEL[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14470.185 1046.435 14470.465 1047.435 ;
    END
  END DIG_MON_SEL[333]
  PIN INJ_ROW[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14466.825 1046.435 14467.105 1047.435 ;
    END
  END INJ_ROW[166]
  PIN Data_COMP[1142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14465.145 1046.435 14465.425 1047.435 ;
    END
  END Data_COMP[1142]
  PIN Data_COMP[1139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14463.465 1046.435 14463.745 1047.435 ;
    END
  END Data_COMP[1139]
  PIN Data_COMP[1148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14461.785 1046.435 14462.065 1047.435 ;
    END
  END Data_COMP[1148]
  PIN INJ_IN[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14451.145 1046.435 14451.425 1047.435 ;
    END
  END INJ_IN[333]
  PIN BcidMtx[1001]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14448.905 1046.435 14449.185 1047.435 ;
    END
  END BcidMtx[1001]
  PIN FREEZE_COMP[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14447.225 1046.435 14447.505 1047.435 ;
    END
  END FREEZE_COMP[54]
  PIN BcidMtx[996]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14444.985 1046.435 14445.265 1047.435 ;
    END
  END BcidMtx[996]
  PIN Data_COMP[1137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14440.785 1046.435 14441.065 1047.435 ;
    END
  END Data_COMP[1137]
  PIN Data_COMP[1149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14439.105 1046.435 14439.385 1047.435 ;
    END
  END Data_COMP[1149]
  PIN Data_COMP[1145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14411.385 1046.435 14411.665 1047.435 ;
    END
  END Data_COMP[1145]
  PIN MASKD[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14968.025 1046.435 14968.305 1047.435 ;
    END
  END MASKD[346]
  PIN DIG_MON_SEL[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14965.225 1046.435 14965.505 1047.435 ;
    END
  END DIG_MON_SEL[346]
  PIN INJ_ROW[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14961.305 1046.435 14961.585 1047.435 ;
    END
  END INJ_ROW[172]
  PIN Data_HV[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14960.185 1046.435 14960.465 1047.435 ;
    END
  END Data_HV[102]
  PIN Data_HV[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14945.625 1046.435 14945.905 1047.435 ;
    END
  END Data_HV[103]
  PIN Data_HV[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14943.945 1046.435 14944.225 1047.435 ;
    END
  END Data_HV[104]
  PIN Data_HV[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14942.265 1046.435 14942.545 1047.435 ;
    END
  END Data_HV[90]
  PIN BcidMtx[1037]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14938.905 1046.435 14939.185 1047.435 ;
    END
  END BcidMtx[1037]
  PIN FREEZE_HV[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14937.225 1046.435 14937.505 1047.435 ;
    END
  END FREEZE_HV[4]
  PIN BcidMtx[1033]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14935.545 1046.435 14935.825 1047.435 ;
    END
  END BcidMtx[1033]
  PIN Data_HV[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14894.105 1046.435 14894.385 1047.435 ;
    END
  END Data_HV[87]
  PIN Data_HV[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14892.425 1046.435 14892.705 1047.435 ;
    END
  END Data_HV[99]
  PIN Data_HV[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14891.305 1046.435 14891.585 1047.435 ;
    END
  END Data_HV[88]
  PIN Data_HV[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14889.625 1046.435 14889.905 1047.435 ;
    END
  END Data_HV[85]
  PIN MASKV[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14887.945 1046.435 14888.225 1047.435 ;
    END
  END MASKV[344]
  PIN DIG_MON_HV[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14885.705 1046.435 14885.985 1047.435 ;
    END
  END DIG_MON_HV[8]
  PIN DIG_MON_SEL[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14883.465 1046.435 14883.745 1047.435 ;
    END
  END DIG_MON_SEL[343]
  PIN INJ_ROW[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14871.705 1046.435 14871.985 1047.435 ;
    END
  END INJ_ROW[171]
  PIN Data_HV[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14870.025 1046.435 14870.305 1047.435 ;
    END
  END Data_HV[71]
  PIN Data_HV[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14868.345 1046.435 14868.625 1047.435 ;
    END
  END Data_HV[68]
  PIN Data_HV[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14866.665 1046.435 14866.945 1047.435 ;
    END
  END Data_HV[77]
  PIN INJ_IN[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14862.465 1046.435 14862.745 1047.435 ;
    END
  END INJ_IN[343]
  PIN BcidMtx[1030]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14859.665 1046.435 14859.945 1047.435 ;
    END
  END BcidMtx[1030]
  PIN BcidMtx[1027]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14831.385 1046.435 14831.665 1047.435 ;
    END
  END BcidMtx[1027]
  PIN INJ_IN[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14829.705 1046.435 14829.985 1047.435 ;
    END
  END INJ_IN[342]
  PIN Data_HV[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14827.465 1046.435 14827.745 1047.435 ;
    END
  END Data_HV[72]
  PIN Data_HV[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14825.225 1046.435 14825.505 1047.435 ;
    END
  END Data_HV[79]
  PIN Data_HV[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14824.105 1046.435 14824.385 1047.435 ;
    END
  END Data_HV[64]
  PIN MASKV[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14822.425 1046.435 14822.705 1047.435 ;
    END
  END MASKV[342]
  PIN DIG_MON_HV[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14820.185 1046.435 14820.465 1047.435 ;
    END
  END DIG_MON_HV[6]
  PIN DIG_MON_SEL[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14805.065 1046.435 14805.345 1047.435 ;
    END
  END DIG_MON_SEL[341]
  PIN INJ_ROW[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14801.705 1046.435 14801.985 1047.435 ;
    END
  END INJ_ROW[170]
  PIN Data_HV[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14800.025 1046.435 14800.305 1047.435 ;
    END
  END Data_HV[50]
  PIN Data_HV[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14798.345 1046.435 14798.625 1047.435 ;
    END
  END Data_HV[47]
  PIN Data_HV[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14796.665 1046.435 14796.945 1047.435 ;
    END
  END Data_HV[56]
  PIN INJ_IN[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14794.425 1046.435 14794.705 1047.435 ;
    END
  END INJ_IN[341]
  PIN BcidMtx[1024]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14752.425 1046.435 14752.705 1047.435 ;
    END
  END BcidMtx[1024]
  PIN Read_HV[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14750.745 1046.435 14751.025 1047.435 ;
    END
  END Read_HV[2]
  PIN BcidMtx[1020]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14749.065 1046.435 14749.345 1047.435 ;
    END
  END BcidMtx[1020]
  PIN MASKD[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18723.945 1046.435 18724.225 1047.435 ;
    END
  END MASKD[439]
  PIN Data_HV[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14745.145 1046.435 14745.425 1047.435 ;
    END
  END Data_HV[57]
  PIN Data_HV[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14742.905 1046.435 14743.185 1047.435 ;
    END
  END Data_HV[53]
  PIN Data_HV[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14741.225 1046.435 14741.505 1047.435 ;
    END
  END Data_HV[59]
  PIN MASKD[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14731.145 1046.435 14731.425 1047.435 ;
    END
  END MASKD[340]
  PIN DIG_MON_SEL[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14728.345 1046.435 14728.625 1047.435 ;
    END
  END DIG_MON_SEL[340]
  PIN MASKD[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14726.665 1046.435 14726.945 1047.435 ;
    END
  END MASKD[339]
  PIN MASKV[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14721.905 1046.435 14722.185 1047.435 ;
    END
  END MASKV[339]
  PIN Data_HV[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14719.665 1046.435 14719.945 1047.435 ;
    END
  END Data_HV[40]
  PIN Data_HV[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14693.065 1046.435 14693.345 1047.435 ;
    END
  END Data_HV[34]
  PIN Data_HV[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14691.385 1046.435 14691.665 1047.435 ;
    END
  END Data_HV[28]
  PIN BcidMtx[1018]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14686.905 1046.435 14687.185 1047.435 ;
    END
  END BcidMtx[1018]
  PIN FREEZE_HV[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14685.785 1046.435 14686.065 1047.435 ;
    END
  END FREEZE_HV[1]
  PIN BcidMtx[1015]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14684.105 1046.435 14684.385 1047.435 ;
    END
  END BcidMtx[1015]
  PIN Data_HV[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14681.305 1046.435 14681.585 1047.435 ;
    END
  END Data_HV[24]
  PIN Data_HV[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14666.745 1046.435 14667.025 1047.435 ;
    END
  END Data_HV[36]
  PIN Data_HV[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14665.625 1046.435 14665.905 1047.435 ;
    END
  END Data_HV[25]
  PIN Data_HV[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14663.945 1046.435 14664.225 1047.435 ;
    END
  END Data_HV[22]
  PIN MASKV[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14662.265 1046.435 14662.545 1047.435 ;
    END
  END MASKV[338]
  PIN DIG_MON_HV[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14660.025 1046.435 14660.305 1047.435 ;
    END
  END DIG_MON_HV[2]
  PIN DIG_MON_HV[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14655.545 1046.435 14655.825 1047.435 ;
    END
  END DIG_MON_HV[1]
  PIN INJ_ROW[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14654.425 1046.435 14654.705 1047.435 ;
    END
  END INJ_ROW[168]
  PIN Data_HV[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14612.985 1046.435 14613.265 1047.435 ;
    END
  END Data_HV[8]
  PIN Data_HV[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14610.745 1046.435 14611.025 1047.435 ;
    END
  END Data_HV[13]
  PIN Data_HV[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14609.065 1046.435 14609.345 1047.435 ;
    END
  END Data_HV[7]
  PIN INJ_IN[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14607.385 1046.435 14607.665 1047.435 ;
    END
  END INJ_IN[337]
  PIN BcidMtx[1011]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14604.025 1046.435 14604.305 1047.435 ;
    END
  END BcidMtx[1011]
  PIN BcidMtx[1010]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14602.345 1046.435 14602.625 1047.435 ;
    END
  END BcidMtx[1010]
  PIN INJ_IN[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14591.705 1046.435 14591.985 1047.435 ;
    END
  END INJ_IN[336]
  PIN Data_HV[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14588.905 1046.435 14589.185 1047.435 ;
    END
  END Data_HV[15]
  PIN Data_HV[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14587.785 1046.435 14588.065 1047.435 ;
    END
  END Data_HV[4]
  PIN Data_HV[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14586.105 1046.435 14586.385 1047.435 ;
    END
  END Data_HV[1]
  PIN Data_HV[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14585.545 1046.435 14585.825 1047.435 ;
    END
  END Data_HV[0]
  PIN MASKD[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14581.345 1046.435 14581.625 1047.435 ;
    END
  END MASKD[336]
  PIN DIG_MON_SEL[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14578.545 1046.435 14578.825 1047.435 ;
    END
  END DIG_MON_SEL[336]
  PIN MASKD[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15670.825 1046.435 15671.105 1047.435 ;
    END
  END MASKD[363]
  PIN MASKV[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15668.025 1046.435 15668.305 1047.435 ;
    END
  END MASKV[363]
  PIN Data_HV[285]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15666.345 1046.435 15666.625 1047.435 ;
    END
  END Data_HV[285]
  PIN Data_HV[293]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15664.105 1046.435 15664.385 1047.435 ;
    END
  END Data_HV[293]
  PIN Data_HV[279]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15662.425 1046.435 15662.705 1047.435 ;
    END
  END Data_HV[279]
  PIN nTOK_HV[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15660.185 1046.435 15660.465 1047.435 ;
    END
  END nTOK_HV[13]
  PIN Read_HV[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15643.385 1046.435 15643.665 1047.435 ;
    END
  END Read_HV[13]
  PIN BcidMtx[1088]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15642.825 1046.435 15643.105 1047.435 ;
    END
  END BcidMtx[1088]
  PIN INJ_IN[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15640.585 1046.435 15640.865 1047.435 ;
    END
  END INJ_IN[362]
  PIN Data_HV[283]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15637.225 1046.435 15637.505 1047.435 ;
    END
  END Data_HV[283]
  PIN Data_HV[289]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15636.105 1046.435 15636.385 1047.435 ;
    END
  END Data_HV[289]
  PIN Data_HV[274]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15634.985 1046.435 15635.265 1047.435 ;
    END
  END Data_HV[274]
  PIN MASKD[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15593.545 1046.435 15593.825 1047.435 ;
    END
  END MASKD[362]
  PIN DIG_MON_SEL[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15590.185 1046.435 15590.465 1047.435 ;
    END
  END DIG_MON_SEL[361]
  PIN Data_HV[270]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15585.705 1046.435 15585.985 1047.435 ;
    END
  END Data_HV[270]
  PIN Data_HV[260]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15585.145 1046.435 15585.425 1047.435 ;
    END
  END Data_HV[260]
  PIN Data_HV[257]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15583.465 1046.435 15583.745 1047.435 ;
    END
  END Data_HV[257]
  PIN Data_HV[258]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15572.265 1046.435 15572.545 1047.435 ;
    END
  END Data_HV[258]
  PIN INJ_IN[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15571.145 1046.435 15571.425 1047.435 ;
    END
  END INJ_IN[361]
  PIN BcidMtx[1084]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15568.345 1046.435 15568.625 1047.435 ;
    END
  END BcidMtx[1084]
  PIN Read_HV[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15566.665 1046.435 15566.945 1047.435 ;
    END
  END Read_HV[12]
  PIN BcidMtx[1081]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15565.545 1046.435 15565.825 1047.435 ;
    END
  END BcidMtx[1081]
  PIN Data_HV[254]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15560.225 1046.435 15560.505 1047.435 ;
    END
  END Data_HV[254]
  PIN Data_HV[262]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15558.545 1046.435 15558.825 1047.435 ;
    END
  END Data_HV[262]
  PIN Data_HV[263]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15531.385 1046.435 15531.665 1047.435 ;
    END
  END Data_HV[263]
  PIN Data_HV[269]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15529.705 1046.435 15529.985 1047.435 ;
    END
  END Data_HV[269]
  PIN MASKD[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15528.025 1046.435 15528.305 1047.435 ;
    END
  END MASKD[360]
  PIN DIG_MON_SEL[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15525.225 1046.435 15525.505 1047.435 ;
    END
  END DIG_MON_SEL[360]
  PIN DIG_MON_HV[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15522.425 1046.435 15522.705 1047.435 ;
    END
  END DIG_MON_HV[23]
  PIN Data_HV[249]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15520.185 1046.435 15520.465 1047.435 ;
    END
  END Data_HV[249]
  PIN Data_HV[250]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15505.625 1046.435 15505.905 1047.435 ;
    END
  END Data_HV[250]
  PIN Data_HV[251]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15503.945 1046.435 15504.225 1047.435 ;
    END
  END Data_HV[251]
  PIN Data_HV[237]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15502.265 1046.435 15502.545 1047.435 ;
    END
  END Data_HV[237]
  PIN BcidMtx[1078]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15498.345 1046.435 15498.625 1047.435 ;
    END
  END BcidMtx[1078]
  PIN FREEZE_HV[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15497.225 1046.435 15497.505 1047.435 ;
    END
  END FREEZE_HV[11]
  PIN Data_HV[1071]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18661.785 1046.435 18662.065 1047.435 ;
    END
  END Data_HV[1071]
  PIN INJ_IN[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15493.865 1046.435 15494.145 1047.435 ;
    END
  END INJ_IN[358]
  PIN Data_HV[233]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15453.545 1046.435 15453.825 1047.435 ;
    END
  END Data_HV[233]
  PIN Data_HV[241]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15451.865 1046.435 15452.145 1047.435 ;
    END
  END Data_HV[241]
  PIN Data_HV[242]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15450.185 1046.435 15450.465 1047.435 ;
    END
  END Data_HV[242]
  PIN Data_HV[248]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15448.505 1046.435 15448.785 1047.435 ;
    END
  END Data_HV[248]
  PIN MASKD[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15446.825 1046.435 15447.105 1047.435 ;
    END
  END MASKD[358]
  PIN DIG_MON_SEL[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15444.025 1046.435 15444.305 1047.435 ;
    END
  END DIG_MON_SEL[358]
  PIN DIG_MON_HV[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15441.225 1046.435 15441.505 1047.435 ;
    END
  END DIG_MON_HV[21]
  PIN Data_HV[228]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15430.585 1046.435 15430.865 1047.435 ;
    END
  END Data_HV[228]
  PIN Data_HV[229]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15428.905 1046.435 15429.185 1047.435 ;
    END
  END Data_HV[229]
  PIN Data_HV[230]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15427.225 1046.435 15427.505 1047.435 ;
    END
  END Data_HV[230]
  PIN Data_HV[216]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15425.545 1046.435 15425.825 1047.435 ;
    END
  END Data_HV[216]
  PIN BcidMtx[1073]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15420.225 1046.435 15420.505 1047.435 ;
    END
  END BcidMtx[1073]
  PIN Read_HV[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15392.505 1046.435 15392.785 1047.435 ;
    END
  END Read_HV[10]
  PIN BcidMtx[1069]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15391.385 1046.435 15391.665 1047.435 ;
    END
  END BcidMtx[1069]
  PIN Read_HV[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18605.225 1046.435 18605.505 1047.435 ;
    END
  END Read_HV[50]
  PIN Data_HV[212]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15388.025 1046.435 15388.305 1047.435 ;
    END
  END Data_HV[212]
  PIN Data_HV[220]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15386.345 1046.435 15386.625 1047.435 ;
    END
  END Data_HV[220]
  PIN Data_HV[211]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15384.105 1046.435 15384.385 1047.435 ;
    END
  END Data_HV[211]
  PIN Data_HV[227]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15382.985 1046.435 15383.265 1047.435 ;
    END
  END Data_HV[227]
  PIN MASKD[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15381.305 1046.435 15381.585 1047.435 ;
    END
  END MASKD[356]
  PIN DIG_MON_SEL[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15365.065 1046.435 15365.345 1047.435 ;
    END
  END DIG_MON_SEL[355]
  PIN DIG_MON_HV[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15362.825 1046.435 15363.105 1047.435 ;
    END
  END DIG_MON_HV[19]
  PIN Data_HV[207]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15360.585 1046.435 15360.865 1047.435 ;
    END
  END Data_HV[207]
  PIN Data_HV[194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15358.345 1046.435 15358.625 1047.435 ;
    END
  END Data_HV[194]
  PIN Data_HV[209]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15357.225 1046.435 15357.505 1047.435 ;
    END
  END Data_HV[209]
  PIN Data_HV[195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15355.545 1046.435 15355.825 1047.435 ;
    END
  END Data_HV[195]
  PIN BcidMtx[1067]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15312.985 1046.435 15313.265 1047.435 ;
    END
  END BcidMtx[1067]
  PIN FREEZE_HV[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15311.305 1046.435 15311.585 1047.435 ;
    END
  END FREEZE_HV[9]
  PIN BcidMtx[1064]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15310.185 1046.435 15310.465 1047.435 ;
    END
  END BcidMtx[1064]
  PIN INJ_IN[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15307.945 1046.435 15308.225 1047.435 ;
    END
  END INJ_IN[354]
  PIN Data_HV[1061]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18584.505 1046.435 18584.785 1047.435 ;
    END
  END Data_HV[1061]
  PIN Data_HV[204]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15305.145 1046.435 15305.425 1047.435 ;
    END
  END Data_HV[204]
  PIN Data_HV[200]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15302.905 1046.435 15303.185 1047.435 ;
    END
  END Data_HV[200]
  PIN Data_HV[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15301.785 1046.435 15302.065 1047.435 ;
    END
  END Data_HV[189]
  PIN MASKH[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15291.705 1046.435 15291.985 1047.435 ;
    END
  END MASKH[177]
  PIN MASKD[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15286.665 1046.435 15286.945 1047.435 ;
    END
  END MASKD[353]
  PIN MASKV[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15281.905 1046.435 15282.185 1047.435 ;
    END
  END MASKV[353]
  PIN Data_HV[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15280.225 1046.435 15280.505 1047.435 ;
    END
  END Data_HV[180]
  PIN Data_HV[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15253.065 1046.435 15253.345 1047.435 ;
    END
  END Data_HV[181]
  PIN Data_HV[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15251.385 1046.435 15251.665 1047.435 ;
    END
  END Data_HV[175]
  PIN BcidMtx[1061]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15247.465 1046.435 15247.745 1047.435 ;
    END
  END BcidMtx[1061]
  PIN BcidMtx[1059]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15246.345 1046.435 15246.625 1047.435 ;
    END
  END BcidMtx[1059]
  PIN BcidMtx[1058]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15244.665 1046.435 15244.945 1047.435 ;
    END
  END BcidMtx[1058]
  PIN Data_HV[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15241.305 1046.435 15241.585 1047.435 ;
    END
  END Data_HV[171]
  PIN Data_HV[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15240.185 1046.435 15240.465 1047.435 ;
    END
  END Data_HV[177]
  PIN Data_HV[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15225.625 1046.435 15225.905 1047.435 ;
    END
  END Data_HV[172]
  PIN Data_HV[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15223.945 1046.435 15224.225 1047.435 ;
    END
  END Data_HV[169]
  PIN MASKV[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15222.265 1046.435 15222.545 1047.435 ;
    END
  END MASKV[352]
  PIN DIG_MON_HV[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15220.025 1046.435 15220.305 1047.435 ;
    END
  END DIG_MON_HV[16]
  PIN DIG_MON_SEL[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15217.785 1046.435 15218.065 1047.435 ;
    END
  END DIG_MON_SEL[351]
  PIN INJ_ROW[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15214.425 1046.435 15214.705 1047.435 ;
    END
  END INJ_ROW[175]
  PIN Data_HV[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15172.985 1046.435 15173.265 1047.435 ;
    END
  END Data_HV[155]
  PIN Data_HV[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15170.745 1046.435 15171.025 1047.435 ;
    END
  END Data_HV[160]
  PIN Data_HV[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15169.625 1046.435 15169.905 1047.435 ;
    END
  END Data_HV[161]
  PIN INJ_IN[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15167.385 1046.435 15167.665 1047.435 ;
    END
  END INJ_IN[351]
  PIN BcidMtx[1053]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15164.025 1046.435 15164.305 1047.435 ;
    END
  END BcidMtx[1053]
  PIN Read_HV[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15162.905 1046.435 15163.185 1047.435 ;
    END
  END Read_HV[7]
  PIN BcidMtx[1050]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15161.225 1046.435 15161.505 1047.435 ;
    END
  END BcidMtx[1050]
  PIN Data_HV[1083]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18719.465 1046.435 18719.745 1047.435 ;
    END
  END Data_HV[1083]
  PIN Data_HV[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15148.905 1046.435 15149.185 1047.435 ;
    END
  END Data_HV[162]
  PIN Data_HV[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15147.225 1046.435 15147.505 1047.435 ;
    END
  END Data_HV[163]
  PIN Data_HV[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15144.985 1046.435 15145.265 1047.435 ;
    END
  END Data_HV[164]
  PIN MASKH[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15141.905 1046.435 15142.185 1047.435 ;
    END
  END MASKH[175]
  PIN MASKD[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16230.825 1046.435 16231.105 1047.435 ;
    END
  END MASKD[377]
  PIN INJ_ROW[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16228.585 1046.435 16228.865 1047.435 ;
    END
  END INJ_ROW[188]
  PIN Data_HV[428]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16226.905 1046.435 16227.185 1047.435 ;
    END
  END Data_HV[428]
  PIN Data_HV[425]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16225.225 1046.435 16225.505 1047.435 ;
    END
  END Data_HV[425]
  PIN Data_HV[434]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16223.545 1046.435 16223.825 1047.435 ;
    END
  END Data_HV[434]
  PIN INJ_IN[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16221.305 1046.435 16221.585 1047.435 ;
    END
  END INJ_IN[377]
  PIN BcidMtx[1132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16205.065 1046.435 16205.345 1047.435 ;
    END
  END BcidMtx[1132]
  PIN Read_HV[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16203.385 1046.435 16203.665 1047.435 ;
    END
  END Read_HV[20]
  PIN BcidMtx[1128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16201.705 1046.435 16201.985 1047.435 ;
    END
  END BcidMtx[1128]
  PIN Data_HV[422]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16198.905 1046.435 16199.185 1047.435 ;
    END
  END Data_HV[422]
  PIN Data_HV[435]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16197.785 1046.435 16198.065 1047.435 ;
    END
  END Data_HV[435]
  PIN Data_HV[431]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16195.545 1046.435 16195.825 1047.435 ;
    END
  END Data_HV[431]
  PIN Data_HV[437]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16193.865 1046.435 16194.145 1047.435 ;
    END
  END Data_HV[437]
  PIN MASKH[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16154.105 1046.435 16154.385 1047.435 ;
    END
  END MASKH[188]
  PIN DIG_MON_SEL[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16150.745 1046.435 16151.025 1047.435 ;
    END
  END DIG_MON_SEL[376]
  PIN DIG_MON_HV[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16147.945 1046.435 16148.225 1047.435 ;
    END
  END DIG_MON_HV[39]
  PIN INJ_ROW[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16146.825 1046.435 16147.105 1047.435 ;
    END
  END INJ_ROW[187]
  PIN Data_HV[418]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16144.025 1046.435 16144.305 1047.435 ;
    END
  END Data_HV[418]
  PIN Data_HV[419]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16142.345 1046.435 16142.625 1047.435 ;
    END
  END Data_HV[419]
  PIN Data_HV[406]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16141.225 1046.435 16141.505 1047.435 ;
    END
  END Data_HV[406]
  PIN BcidMtx[1127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16128.905 1046.435 16129.185 1047.435 ;
    END
  END BcidMtx[1127]
  PIN FREEZE_HV[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16127.225 1046.435 16127.505 1047.435 ;
    END
  END FREEZE_HV[19]
  PIN BcidMtx[1124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16126.105 1046.435 16126.385 1047.435 ;
    END
  END BcidMtx[1124]
  PIN Data_HV[402]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16120.785 1046.435 16121.065 1047.435 ;
    END
  END Data_HV[402]
  PIN Data_HV[414]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16119.105 1046.435 16119.385 1047.435 ;
    END
  END Data_HV[414]
  PIN Data_HV[415]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16091.945 1046.435 16092.225 1047.435 ;
    END
  END Data_HV[415]
  PIN Data_HV[399]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16090.265 1046.435 16090.545 1047.435 ;
    END
  END Data_HV[399]
  PIN Data_HV[998]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18331.385 1046.435 18331.665 1047.435 ;
    END
  END Data_HV[998]
  PIN Data_HV[1004]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18329.705 1046.435 18329.985 1047.435 ;
    END
  END Data_HV[1004]
  PIN MASKD[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18328.025 1046.435 18328.305 1047.435 ;
    END
  END MASKD[430]
  PIN DIG_MON_SEL[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18325.225 1046.435 18325.505 1047.435 ;
    END
  END DIG_MON_SEL[430]
  PIN DIG_MON_HV[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18322.425 1046.435 18322.705 1047.435 ;
    END
  END DIG_MON_HV[93]
  PIN Data_HV[984]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18320.185 1046.435 18320.465 1047.435 ;
    END
  END Data_HV[984]
  PIN Data_HV[978]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18306.185 1046.435 18306.465 1047.435 ;
    END
  END Data_HV[978]
  PIN Data_HV[986]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18303.945 1046.435 18304.225 1047.435 ;
    END
  END Data_HV[986]
  PIN Data_HV[972]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18302.265 1046.435 18302.545 1047.435 ;
    END
  END Data_HV[972]
  PIN nTOK_HV[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18300.025 1046.435 18300.305 1047.435 ;
    END
  END nTOK_HV[46]
  PIN BcidMtx[1288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18298.345 1046.435 18298.625 1047.435 ;
    END
  END BcidMtx[1288]
  PIN Read_HV[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18296.665 1046.435 18296.945 1047.435 ;
    END
  END Read_HV[46]
  PIN Data_HV[969]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18254.105 1046.435 18254.385 1047.435 ;
    END
  END Data_HV[969]
  PIN Data_HV[968]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18253.545 1046.435 18253.825 1047.435 ;
    END
  END Data_HV[968]
  PIN Data_HV[976]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18251.865 1046.435 18252.145 1047.435 ;
    END
  END Data_HV[976]
  PIN Data_HV[966]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18249.065 1046.435 18249.345 1047.435 ;
    END
  END Data_HV[966]
  PIN Data_HV[983]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18248.505 1046.435 18248.785 1047.435 ;
    END
  END Data_HV[983]
  PIN MASKH[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18247.385 1046.435 18247.665 1047.435 ;
    END
  END MASKH[214]
  PIN DIG_MON_SEL[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18244.025 1046.435 18244.305 1047.435 ;
    END
  END DIG_MON_SEL[428]
  PIN DIG_MON_SEL[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18243.465 1046.435 18243.745 1047.435 ;
    END
  END DIG_MON_SEL[427]
  PIN INJ_ROW[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18231.705 1046.435 18231.985 1047.435 ;
    END
  END INJ_ROW[213]
  PIN Data_HV[964]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18228.905 1046.435 18229.185 1047.435 ;
    END
  END Data_HV[964]
  PIN Data_HV[950]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18228.345 1046.435 18228.625 1047.435 ;
    END
  END Data_HV[950]
  PIN Data_HV[959]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18226.665 1046.435 18226.945 1047.435 ;
    END
  END Data_HV[959]
  PIN BcidMtx[1283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18220.225 1046.435 18220.505 1047.435 ;
    END
  END BcidMtx[1283]
  PIN BcidMtx[1282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18219.665 1046.435 18219.945 1047.435 ;
    END
  END BcidMtx[1282]
  PIN BcidMtx[1280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18191.945 1046.435 18192.225 1047.435 ;
    END
  END BcidMtx[1280]
  PIN Data_HV[947]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18188.025 1046.435 18188.305 1047.435 ;
    END
  END Data_HV[947]
  PIN Data_HV[960]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18186.905 1046.435 18187.185 1047.435 ;
    END
  END Data_HV[960]
  PIN Data_HV[961]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18185.225 1046.435 18185.505 1047.435 ;
    END
  END Data_HV[961]
  PIN MASKV[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18182.425 1046.435 18182.705 1047.435 ;
    END
  END MASKV[426]
  PIN MASKD[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18181.305 1046.435 18181.585 1047.435 ;
    END
  END MASKD[426]
  PIN MASKD[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18163.945 1046.435 18164.225 1047.435 ;
    END
  END MASKD[425]
  PIN INJ_ROW[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18161.705 1046.435 18161.985 1047.435 ;
    END
  END INJ_ROW[212]
  PIN Data_HV[932]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18160.025 1046.435 18160.305 1047.435 ;
    END
  END Data_HV[932]
  PIN Data_HV[937]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18157.785 1046.435 18158.065 1047.435 ;
    END
  END Data_HV[937]
  PIN Data_HV[938]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18156.665 1046.435 18156.945 1047.435 ;
    END
  END Data_HV[938]
  PIN INJ_IN[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18154.425 1046.435 18154.705 1047.435 ;
    END
  END INJ_IN[425]
  PIN BcidMtx[1275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18111.865 1046.435 18112.145 1047.435 ;
    END
  END BcidMtx[1275]
  PIN Read_HV[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18110.745 1046.435 18111.025 1047.435 ;
    END
  END Read_HV[44]
  PIN BcidMtx[1272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18109.065 1046.435 18109.345 1047.435 ;
    END
  END BcidMtx[1272]
  PIN Data_HV[933]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18105.705 1046.435 18105.985 1047.435 ;
    END
  END Data_HV[933]
  PIN Data_HV[934]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18104.585 1046.435 18104.865 1047.435 ;
    END
  END Data_HV[934]
  PIN Data_HV[935]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18102.905 1046.435 18103.185 1047.435 ;
    END
  END Data_HV[935]
  PIN MASKV[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18092.265 1046.435 18092.545 1047.435 ;
    END
  END MASKV[424]
  PIN MASKD[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18091.145 1046.435 18091.425 1047.435 ;
    END
  END MASKD[424]
  PIN DIG_MON_HV[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18085.545 1046.435 18085.825 1047.435 ;
    END
  END DIG_MON_HV[87]
  PIN INJ_ROW[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18082.465 1046.435 18082.745 1047.435 ;
    END
  END INJ_ROW[211]
  PIN Data_HV[911]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18080.785 1046.435 18081.065 1047.435 ;
    END
  END Data_HV[911]
  PIN Data_HV[923]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18052.505 1046.435 18052.785 1047.435 ;
    END
  END Data_HV[923]
  PIN Data_HV[910]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18051.385 1046.435 18051.665 1047.435 ;
    END
  END Data_HV[910]
  PIN INJ_IN[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18049.705 1046.435 18049.985 1047.435 ;
    END
  END INJ_IN[423]
  PIN FREEZE_HV[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18045.785 1046.435 18046.065 1047.435 ;
    END
  END FREEZE_HV[43]
  PIN BcidMtx[1268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18044.665 1046.435 18044.945 1047.435 ;
    END
  END BcidMtx[1268]
  PIN INJ_IN[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18042.425 1046.435 18042.705 1047.435 ;
    END
  END INJ_IN[422]
  PIN Data_HV[918]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18026.745 1046.435 18027.025 1047.435 ;
    END
  END Data_HV[918]
  PIN Data_HV[907]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18025.625 1046.435 18025.905 1047.435 ;
    END
  END Data_HV[907]
  PIN Data_HV[904]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18023.945 1046.435 18024.225 1047.435 ;
    END
  END Data_HV[904]
  PIN MASKH[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18021.705 1046.435 18021.985 1047.435 ;
    END
  END MASKH[211]
  PIN DIG_MON_HV[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18020.025 1046.435 18020.305 1047.435 ;
    END
  END DIG_MON_HV[86]
  PIN Data_HV[1052]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18600.745 1046.435 18601.025 1047.435 ;
    END
  END Data_HV[1052]
  PIN INJ_ROW[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18014.425 1046.435 18014.705 1047.435 ;
    END
  END INJ_ROW[210]
  PIN Data_HV[900]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17973.545 1046.435 17973.825 1047.435 ;
    END
  END Data_HV[900]
  PIN Data_HV[901]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17971.865 1046.435 17972.145 1047.435 ;
    END
  END Data_HV[901]
  PIN Data_HV[896]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17969.625 1046.435 17969.905 1047.435 ;
    END
  END Data_HV[896]
  PIN Data_HV[888]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17968.505 1046.435 17968.785 1047.435 ;
    END
  END Data_HV[888]
  PIN BcidMtx[1265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17965.145 1046.435 17965.425 1047.435 ;
    END
  END BcidMtx[1265]
  PIN Read_HV[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17962.905 1046.435 17963.185 1047.435 ;
    END
  END Read_HV[42]
  PIN BcidMtx[1260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17961.225 1046.435 17961.505 1047.435 ;
    END
  END BcidMtx[1260]
  PIN Data_HV[885]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17950.585 1046.435 17950.865 1047.435 ;
    END
  END Data_HV[885]
  PIN Data_HV[892]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17948.345 1046.435 17948.625 1047.435 ;
    END
  END Data_HV[892]
  PIN Data_HV[893]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17946.665 1046.435 17946.945 1047.435 ;
    END
  END Data_HV[893]
  PIN Data_HV[899]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17944.985 1046.435 17945.265 1047.435 ;
    END
  END Data_HV[899]
  PIN MASKD[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17941.345 1046.435 17941.625 1047.435 ;
    END
  END MASKD[420]
  PIN DIG_MON_SEL[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17938.545 1046.435 17938.825 1047.435 ;
    END
  END DIG_MON_SEL[420]
  PIN MASKD[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 19030.825 1046.435 19031.105 1047.435 ;
    END
  END MASKD[447]
  PIN MASKV[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 19028.025 1046.435 19028.305 1047.435 ;
    END
  END MASKV[447]
  PIN Data_HV[1167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 19026.345 1046.435 19026.625 1047.435 ;
    END
  END Data_HV[1167]
  PIN Data_HV[1168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 19024.665 1046.435 19024.945 1047.435 ;
    END
  END Data_HV[1168]
  PIN Data_HV[1162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 19022.985 1046.435 19023.265 1047.435 ;
    END
  END Data_HV[1162]
  PIN nTOK_HV[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 19020.185 1046.435 19020.465 1047.435 ;
    END
  END nTOK_HV[55]
  PIN BcidMtx[1341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 19004.505 1046.435 19004.785 1047.435 ;
    END
  END BcidMtx[1341]
  PIN Read_HV[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 19003.385 1046.435 19003.665 1047.435 ;
    END
  END Read_HV[55]
  PIN BcidMtx[1339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 19002.265 1046.435 19002.545 1047.435 ;
    END
  END BcidMtx[1339]
  PIN Data_HV[1158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18999.465 1046.435 18999.745 1047.435 ;
    END
  END Data_HV[1158]
  PIN Data_HV[1165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18997.225 1046.435 18997.505 1047.435 ;
    END
  END Data_HV[1165]
  PIN Data_HV[1171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18996.105 1046.435 18996.385 1047.435 ;
    END
  END Data_HV[1171]
  PIN Data_HV[1155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18994.425 1046.435 18994.705 1047.435 ;
    END
  END Data_HV[1155]
  PIN MASKV[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18954.665 1046.435 18954.945 1047.435 ;
    END
  END MASKV[446]
  PIN MASKD[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18949.065 1046.435 18949.345 1047.435 ;
    END
  END MASKD[445]
  PIN MASKV[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18946.265 1046.435 18946.545 1047.435 ;
    END
  END MASKV[445]
  PIN Data_HV[1142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18945.145 1046.435 18945.425 1047.435 ;
    END
  END Data_HV[1142]
  PIN Data_HV[1147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18942.905 1046.435 18943.185 1047.435 ;
    END
  END Data_HV[1147]
  PIN Data_HV[1148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18941.785 1046.435 18942.065 1047.435 ;
    END
  END Data_HV[1148]
  PIN INJ_IN[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18931.145 1046.435 18931.425 1047.435 ;
    END
  END INJ_IN[445]
  PIN BcidMtx[1337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18928.905 1046.435 18929.185 1047.435 ;
    END
  END BcidMtx[1337]
  PIN Read_HV[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18926.665 1046.435 18926.945 1047.435 ;
    END
  END Read_HV[54]
  PIN BcidMtx[1332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18924.985 1046.435 18925.265 1047.435 ;
    END
  END BcidMtx[1332]
  PIN DIG_MON_PMOS_NOSF[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1669.705 1046.435 1669.985 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[13]
  PIN MASKH[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16088.585 1046.435 16088.865 1047.435 ;
    END
  END MASKH[187]
  PIN DIG_MON_HV[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16086.905 1046.435 16087.185 1047.435 ;
    END
  END DIG_MON_HV[38]
  PIN MASKD[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16083.545 1046.435 16083.825 1047.435 ;
    END
  END MASKD[373]
  PIN MASKV[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16080.745 1046.435 16081.025 1047.435 ;
    END
  END MASKV[373]
  PIN Data_HV[397]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16065.625 1046.435 16065.905 1047.435 ;
    END
  END Data_HV[397]
  PIN Data_HV[391]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16064.505 1046.435 16064.785 1047.435 ;
    END
  END Data_HV[391]
  PIN Data_HV[385]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16062.825 1046.435 16063.105 1047.435 ;
    END
  END Data_HV[385]
  PIN nTOK_HV[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16060.025 1046.435 16060.305 1047.435 ;
    END
  END nTOK_HV[18]
  PIN BcidMtx[1119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16057.785 1046.435 16058.065 1047.435 ;
    END
  END BcidMtx[1119]
  PIN BcidMtx[1118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16056.105 1046.435 16056.385 1047.435 ;
    END
  END BcidMtx[1118]
  PIN INJ_IN[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16053.865 1046.435 16054.145 1047.435 ;
    END
  END INJ_IN[372]
  PIN Data_HV[387]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16012.985 1046.435 16013.265 1047.435 ;
    END
  END Data_HV[387]
  PIN Data_HV[382]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16011.305 1046.435 16011.585 1047.435 ;
    END
  END Data_HV[382]
  PIN Data_HV[389]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16010.185 1046.435 16010.465 1047.435 ;
    END
  END Data_HV[389]
  PIN MASKV[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16007.945 1046.435 16008.225 1047.435 ;
    END
  END MASKV[372]
  PIN DIG_MON_HV[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16005.705 1046.435 16005.985 1047.435 ;
    END
  END DIG_MON_HV[36]
  PIN DIG_MON_SEL[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16004.025 1046.435 16004.305 1047.435 ;
    END
  END DIG_MON_SEL[372]
  PIN INJ_ROW[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15991.705 1046.435 15991.985 1047.435 ;
    END
  END INJ_ROW[185]
  PIN Data_HV[365]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15990.025 1046.435 15990.305 1047.435 ;
    END
  END Data_HV[365]
  PIN Data_HV[369]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15989.465 1046.435 15989.745 1047.435 ;
    END
  END Data_HV[369]
  PIN Data_HV[377]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15987.225 1046.435 15987.505 1047.435 ;
    END
  END Data_HV[377]
  PIN Data_HV[363]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15985.545 1046.435 15985.825 1047.435 ;
    END
  END Data_HV[363]
  PIN Data_HV[1090]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18718.905 1046.435 18719.185 1047.435 ;
    END
  END Data_HV[1090]
  PIN BcidMtx[1114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15979.665 1046.435 15979.945 1047.435 ;
    END
  END BcidMtx[1114]
  PIN BcidMtx[1112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15951.945 1046.435 15952.225 1047.435 ;
    END
  END BcidMtx[1112]
  PIN BcidMtx[1110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15950.825 1046.435 15951.105 1047.435 ;
    END
  END BcidMtx[1110]
  PIN Data_HV[366]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15947.465 1046.435 15947.745 1047.435 ;
    END
  END Data_HV[366]
  PIN Data_HV[361]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15945.785 1046.435 15946.065 1047.435 ;
    END
  END Data_HV[361]
  PIN Data_HV[373]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15945.225 1046.435 15945.505 1047.435 ;
    END
  END Data_HV[373]
  PIN Data_HV[357]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15943.545 1046.435 15943.825 1047.435 ;
    END
  END Data_HV[357]
  PIN DIG_MON_HV[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15940.185 1046.435 15940.465 1047.435 ;
    END
  END DIG_MON_HV[34]
  PIN DIG_MON_SEL[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15925.065 1046.435 15925.345 1047.435 ;
    END
  END DIG_MON_SEL[369]
  PIN INJ_ROW[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15921.705 1046.435 15921.985 1047.435 ;
    END
  END INJ_ROW[184]
  PIN Data_HV[348]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15919.465 1046.435 15919.745 1047.435 ;
    END
  END Data_HV[348]
  PIN Data_HV[341]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15918.345 1046.435 15918.625 1047.435 ;
    END
  END Data_HV[341]
  PIN Data_HV[350]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15916.665 1046.435 15916.945 1047.435 ;
    END
  END Data_HV[350]
  PIN INJ_IN[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15914.425 1046.435 15914.705 1047.435 ;
    END
  END INJ_IN[369]
  PIN BcidMtx[1109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15872.985 1046.435 15873.265 1047.435 ;
    END
  END BcidMtx[1109]
  PIN FREEZE_HV[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15871.305 1046.435 15871.585 1047.435 ;
    END
  END FREEZE_HV[16]
  PIN BcidMtx[1105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15869.625 1046.435 15869.905 1047.435 ;
    END
  END BcidMtx[1105]
  PIN INJ_IN[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15867.945 1046.435 15868.225 1047.435 ;
    END
  END INJ_IN[368]
  PIN Data_HV[345]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15865.705 1046.435 15865.985 1047.435 ;
    END
  END Data_HV[345]
  PIN Data_HV[352]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15863.465 1046.435 15863.745 1047.435 ;
    END
  END Data_HV[352]
  PIN Data_HV[337]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15862.345 1046.435 15862.625 1047.435 ;
    END
  END Data_HV[337]
  PIN MASKD[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15851.145 1046.435 15851.425 1047.435 ;
    END
  END MASKD[368]
  PIN DIG_MON_SEL[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15847.785 1046.435 15848.065 1047.435 ;
    END
  END DIG_MON_SEL[367]
  PIN INJ_ROW[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15842.465 1046.435 15842.745 1047.435 ;
    END
  END INJ_ROW[183]
  PIN Data_HV[327]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15840.225 1046.435 15840.505 1047.435 ;
    END
  END Data_HV[327]
  PIN Data_HV[320]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15839.105 1046.435 15839.385 1047.435 ;
    END
  END Data_HV[320]
  PIN Data_HV[329]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15811.945 1046.435 15812.225 1047.435 ;
    END
  END Data_HV[329]
  PIN nTOK_HV[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15808.585 1046.435 15808.865 1047.435 ;
    END
  END nTOK_HV[15]
  PIN BcidMtx[1102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15806.905 1046.435 15807.185 1047.435 ;
    END
  END BcidMtx[1102]
  PIN FREEZE_HV[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15805.785 1046.435 15806.065 1047.435 ;
    END
  END FREEZE_HV[15]
  PIN BcidMtx[1098]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15803.545 1046.435 15803.825 1047.435 ;
    END
  END BcidMtx[1098]
  PIN Data_HV[318]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15801.305 1046.435 15801.585 1047.435 ;
    END
  END Data_HV[318]
  PIN Data_HV[330]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15786.745 1046.435 15787.025 1047.435 ;
    END
  END Data_HV[330]
  PIN Data_HV[326]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15784.505 1046.435 15784.785 1047.435 ;
    END
  END Data_HV[326]
  PIN Data_HV[315]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15783.385 1046.435 15783.665 1047.435 ;
    END
  END Data_HV[315]
  PIN MASKH[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15781.705 1046.435 15781.985 1047.435 ;
    END
  END MASKH[183]
  PIN DIG_MON_SEL[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15778.345 1046.435 15778.625 1047.435 ;
    END
  END DIG_MON_SEL[366]
  PIN MASKD[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15776.665 1046.435 15776.945 1047.435 ;
    END
  END MASKD[365]
  PIN MASKV[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15773.865 1046.435 15774.145 1047.435 ;
    END
  END MASKV[365]
  PIN Data_HV[313]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15731.865 1046.435 15732.145 1047.435 ;
    END
  END Data_HV[313]
  PIN Data_HV[307]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15730.745 1046.435 15731.025 1047.435 ;
    END
  END Data_HV[307]
  PIN Data_HV[301]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15729.065 1046.435 15729.345 1047.435 ;
    END
  END Data_HV[301]
  PIN BcidMtx[1097]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15725.145 1046.435 15725.425 1047.435 ;
    END
  END BcidMtx[1097]
  PIN BcidMtx[1095]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15724.025 1046.435 15724.305 1047.435 ;
    END
  END BcidMtx[1095]
  PIN BcidMtx[1094]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15722.345 1046.435 15722.625 1047.435 ;
    END
  END BcidMtx[1094]
  PIN INJ_IN[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15711.705 1046.435 15711.985 1047.435 ;
    END
  END INJ_IN[364]
  PIN Data_HV[296]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15710.025 1046.435 15710.305 1047.435 ;
    END
  END Data_HV[296]
  PIN Data_HV[309]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15708.905 1046.435 15709.185 1047.435 ;
    END
  END Data_HV[309]
  PIN Data_HV[295]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15706.105 1046.435 15706.385 1047.435 ;
    END
  END Data_HV[295]
  PIN Data_HV[311]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15704.985 1046.435 15705.265 1047.435 ;
    END
  END Data_HV[311]
  PIN MASKH[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15701.905 1046.435 15702.185 1047.435 ;
    END
  END MASKH[182]
  PIN FREEZE_HV[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15953.065 1046.435 15953.345 1047.435 ;
    END
  END FREEZE_HV[17]
  PIN MASKD[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16790.825 1046.435 16791.105 1047.435 ;
    END
  END MASKD[391]
  PIN INJ_ROW[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16788.585 1046.435 16788.865 1047.435 ;
    END
  END INJ_ROW[195]
  PIN Data_HV[586]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16785.785 1046.435 16786.065 1047.435 ;
    END
  END Data_HV[586]
  PIN Data_HV[580]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16784.665 1046.435 16784.945 1047.435 ;
    END
  END Data_HV[580]
  PIN Data_HV[581]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16783.545 1046.435 16783.825 1047.435 ;
    END
  END Data_HV[581]
  PIN BcidMtx[1175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16765.625 1046.435 16765.905 1047.435 ;
    END
  END BcidMtx[1175]
  PIN BcidMtx[1173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16764.505 1046.435 16764.785 1047.435 ;
    END
  END BcidMtx[1173]
  PIN Read_HV[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16763.385 1046.435 16763.665 1047.435 ;
    END
  END Read_HV[27]
  PIN INJ_IN[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16760.585 1046.435 16760.865 1047.435 ;
    END
  END INJ_IN[390]
  PIN Data_HV[569]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16758.905 1046.435 16759.185 1047.435 ;
    END
  END Data_HV[569]
  PIN Data_HV[577]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16757.225 1046.435 16757.505 1047.435 ;
    END
  END Data_HV[577]
  PIN Data_HV[568]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16754.985 1046.435 16755.265 1047.435 ;
    END
  END Data_HV[568]
  PIN Data_HV[584]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16753.865 1046.435 16754.145 1047.435 ;
    END
  END Data_HV[584]
  PIN MASKD[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16713.545 1046.435 16713.825 1047.435 ;
    END
  END MASKD[390]
  PIN DIG_MON_SEL[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16710.185 1046.435 16710.465 1047.435 ;
    END
  END DIG_MON_SEL[389]
  PIN DIG_MON_HV[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16707.945 1046.435 16708.225 1047.435 ;
    END
  END DIG_MON_HV[53]
  PIN Data_HV[564]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16705.705 1046.435 16705.985 1047.435 ;
    END
  END Data_HV[564]
  PIN Data_HV[551]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16703.465 1046.435 16703.745 1047.435 ;
    END
  END Data_HV[551]
  PIN Data_HV[566]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16702.345 1046.435 16702.625 1047.435 ;
    END
  END Data_HV[566]
  PIN Data_HV[552]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16692.265 1046.435 16692.545 1047.435 ;
    END
  END Data_HV[552]
  PIN BcidMtx[1168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16688.345 1046.435 16688.625 1047.435 ;
    END
  END BcidMtx[1168]
  PIN FREEZE_HV[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16687.225 1046.435 16687.505 1047.435 ;
    END
  END FREEZE_HV[26]
  PIN BcidMtx[1165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16685.545 1046.435 16685.825 1047.435 ;
    END
  END BcidMtx[1165]
  PIN Data_HV[555]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16679.665 1046.435 16679.945 1047.435 ;
    END
  END Data_HV[555]
  PIN Data_HV[556]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16678.545 1046.435 16678.825 1047.435 ;
    END
  END Data_HV[556]
  PIN Data_HV[562]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16651.945 1046.435 16652.225 1047.435 ;
    END
  END Data_HV[562]
  PIN Data_HV[693]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17210.265 1046.435 17210.545 1047.435 ;
    END
  END Data_HV[693]
  PIN MASKH[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17208.585 1046.435 17208.865 1047.435 ;
    END
  END MASKH[201]
  PIN DIG_MON_HV[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17206.905 1046.435 17207.185 1047.435 ;
    END
  END DIG_MON_HV[66]
  PIN MASKD[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17203.545 1046.435 17203.825 1047.435 ;
    END
  END MASKD[401]
  PIN Data_HV[1077]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18715.545 1046.435 18715.825 1047.435 ;
    END
  END Data_HV[1077]
  PIN Data_HV[690]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17200.185 1046.435 17200.465 1047.435 ;
    END
  END Data_HV[690]
  PIN Data_HV[677]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17185.065 1046.435 17185.345 1047.435 ;
    END
  END Data_HV[677]
  PIN Data_HV[686]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17183.385 1046.435 17183.665 1047.435 ;
    END
  END Data_HV[686]
  PIN Data_HV[678]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17182.265 1046.435 17182.545 1047.435 ;
    END
  END Data_HV[678]
  PIN BcidMtx[1204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17178.345 1046.435 17178.625 1047.435 ;
    END
  END BcidMtx[1204]
  PIN Read_HV[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17176.665 1046.435 17176.945 1047.435 ;
    END
  END Read_HV[32]
  PIN BcidMtx[1201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17175.545 1046.435 17175.825 1047.435 ;
    END
  END BcidMtx[1201]
  PIN Data_HV[674]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17133.545 1046.435 17133.825 1047.435 ;
    END
  END Data_HV[674]
  PIN Data_HV[682]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17131.865 1046.435 17132.145 1047.435 ;
    END
  END Data_HV[682]
  PIN Data_HV[688]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17130.745 1046.435 17131.025 1047.435 ;
    END
  END Data_HV[688]
  PIN Data_HV[672]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17129.065 1046.435 17129.345 1047.435 ;
    END
  END Data_HV[672]
  PIN MASKD[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17126.825 1046.435 17127.105 1047.435 ;
    END
  END MASKD[400]
  PIN DIG_MON_HV[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17121.225 1046.435 17121.505 1047.435 ;
    END
  END DIG_MON_HV[63]
  PIN Data_HV[669]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17110.585 1046.435 17110.865 1047.435 ;
    END
  END Data_HV[669]
  PIN Data_HV[663]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17109.465 1046.435 17109.745 1047.435 ;
    END
  END Data_HV[663]
  PIN Data_HV[671]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17107.225 1046.435 17107.505 1047.435 ;
    END
  END Data_HV[671]
  PIN Data_HV[657]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17105.545 1046.435 17105.825 1047.435 ;
    END
  END Data_HV[657]
  PIN nTOK_HV[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17101.345 1046.435 17101.625 1047.435 ;
    END
  END nTOK_HV[31]
  PIN Read_HV[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17072.505 1046.435 17072.785 1047.435 ;
    END
  END Read_HV[31]
  PIN BcidMtx[1194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17070.825 1046.435 17071.105 1047.435 ;
    END
  END BcidMtx[1194]
  PIN Data_HV[654]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17068.585 1046.435 17068.865 1047.435 ;
    END
  END Data_HV[654]
  PIN Data_HV[661]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17066.345 1046.435 17066.625 1047.435 ;
    END
  END Data_HV[661]
  PIN Data_HV[662]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17064.665 1046.435 17064.945 1047.435 ;
    END
  END Data_HV[662]
  PIN Data_HV[651]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17063.545 1046.435 17063.825 1047.435 ;
    END
  END Data_HV[651]
  PIN MASKD[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17061.305 1046.435 17061.585 1047.435 ;
    END
  END MASKD[398]
  PIN DIG_MON_SEL[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17045.625 1046.435 17045.905 1047.435 ;
    END
  END DIG_MON_SEL[398]
  PIN MASKD[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17043.945 1046.435 17044.225 1047.435 ;
    END
  END MASKD[397]
  PIN MASKV[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17041.145 1046.435 17041.425 1047.435 ;
    END
  END MASKV[397]
  PIN Data_HV[642]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17039.465 1046.435 17039.745 1047.435 ;
    END
  END Data_HV[642]
  PIN Data_HV[635]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17038.345 1046.435 17038.625 1047.435 ;
    END
  END Data_HV[635]
  PIN Data_HV[644]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17036.665 1046.435 17036.945 1047.435 ;
    END
  END Data_HV[644]
  PIN INJ_IN[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17034.425 1046.435 17034.705 1047.435 ;
    END
  END INJ_IN[397]
  PIN BcidMtx[1193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16992.985 1046.435 16993.265 1047.435 ;
    END
  END BcidMtx[1193]
  PIN Read_HV[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16990.745 1046.435 16991.025 1047.435 ;
    END
  END Read_HV[30]
  PIN BcidMtx[1188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16989.065 1046.435 16989.345 1047.435 ;
    END
  END BcidMtx[1188]
  PIN Data_HV[633]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16986.825 1046.435 16987.105 1047.435 ;
    END
  END Data_HV[633]
  PIN Data_HV[640]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16984.585 1046.435 16984.865 1047.435 ;
    END
  END Data_HV[640]
  PIN Data_HV[641]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16982.905 1046.435 16983.185 1047.435 ;
    END
  END Data_HV[641]
  PIN Data_HV[630]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16981.785 1046.435 16982.065 1047.435 ;
    END
  END Data_HV[630]
  PIN MASKD[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16971.145 1046.435 16971.425 1047.435 ;
    END
  END MASKD[396]
  PIN DIG_MON_SEL[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16968.345 1046.435 16968.625 1047.435 ;
    END
  END DIG_MON_SEL[396]
  PIN MASKD[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16966.665 1046.435 16966.945 1047.435 ;
    END
  END MASKD[395]
  PIN Data_HV[627]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16961.345 1046.435 16961.625 1047.435 ;
    END
  END Data_HV[627]
  PIN Data_HV[621]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16960.225 1046.435 16960.505 1047.435 ;
    END
  END Data_HV[621]
  PIN Data_HV[614]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16959.105 1046.435 16959.385 1047.435 ;
    END
  END Data_HV[614]
  PIN Data_HV[616]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16931.385 1046.435 16931.665 1047.435 ;
    END
  END Data_HV[616]
  PIN nTOK_HV[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16928.585 1046.435 16928.865 1047.435 ;
    END
  END nTOK_HV[29]
  PIN BcidMtx[1186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16926.905 1046.435 16927.185 1047.435 ;
    END
  END BcidMtx[1186]
  PIN BcidMtx[1184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16924.665 1046.435 16924.945 1047.435 ;
    END
  END BcidMtx[1184]
  PIN INJ_IN[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16922.425 1046.435 16922.705 1047.435 ;
    END
  END INJ_IN[394]
  PIN Data_HV[611]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16920.745 1046.435 16921.025 1047.435 ;
    END
  END Data_HV[611]
  PIN Data_HV[613]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16905.625 1046.435 16905.905 1047.435 ;
    END
  END Data_HV[613]
  PIN Data_HV[610]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16903.945 1046.435 16904.225 1047.435 ;
    END
  END Data_HV[610]
  PIN Data_HV[626]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16902.825 1046.435 16903.105 1047.435 ;
    END
  END Data_HV[626]
  PIN DIG_MON_HV[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16900.025 1046.435 16900.305 1047.435 ;
    END
  END DIG_MON_HV[58]
  PIN DIG_MON_SEL[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16897.785 1046.435 16898.065 1047.435 ;
    END
  END DIG_MON_SEL[393]
  PIN DIG_MON_HV[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16895.545 1046.435 16895.825 1047.435 ;
    END
  END DIG_MON_HV[57]
  PIN Data_HV[596]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16852.985 1046.435 16853.265 1047.435 ;
    END
  END Data_HV[596]
  PIN Data_HV[593]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16851.305 1046.435 16851.585 1047.435 ;
    END
  END Data_HV[593]
  PIN INJ_IN[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18602.425 1046.435 18602.705 1047.435 ;
    END
  END INJ_IN[436]
  PIN Data_HV[594]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16848.505 1046.435 16848.785 1047.435 ;
    END
  END Data_HV[594]
  PIN BcidMtx[1181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16845.145 1046.435 16845.425 1047.435 ;
    END
  END BcidMtx[1181]
  PIN BcidMtx[1179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16844.025 1046.435 16844.305 1047.435 ;
    END
  END BcidMtx[1179]
  PIN BcidMtx[1177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16841.785 1046.435 16842.065 1047.435 ;
    END
  END BcidMtx[1177]
  PIN Data_HV[591]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16830.585 1046.435 16830.865 1047.435 ;
    END
  END Data_HV[591]
  PIN Data_HV[597]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16829.465 1046.435 16829.745 1047.435 ;
    END
  END Data_HV[597]
  PIN Data_HV[604]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16827.225 1046.435 16827.505 1047.435 ;
    END
  END Data_HV[604]
  PIN Data_HV[588]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16825.545 1046.435 16825.825 1047.435 ;
    END
  END Data_HV[588]
  PIN MASKV[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16822.465 1046.435 16822.745 1047.435 ;
    END
  END MASKV[392]
  PIN DIG_MON_SEL[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17911.945 1046.435 17912.225 1047.435 ;
    END
  END DIG_MON_SEL[419]
  PIN DIG_MON_HV[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17909.705 1046.435 17909.985 1047.435 ;
    END
  END DIG_MON_HV[83]
  PIN Data_HV[869]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17906.905 1046.435 17907.185 1047.435 ;
    END
  END Data_HV[869]
  PIN Data_HV[866]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17905.225 1046.435 17905.505 1047.435 ;
    END
  END Data_HV[866]
  PIN Data_HV[881]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17904.105 1046.435 17904.385 1047.435 ;
    END
  END Data_HV[881]
  PIN Data_HV[867]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17902.425 1046.435 17902.705 1047.435 ;
    END
  END Data_HV[867]
  PIN BcidMtx[1259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17885.625 1046.435 17885.905 1047.435 ;
    END
  END BcidMtx[1259]
  PIN BcidMtx[1257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17884.505 1046.435 17884.785 1047.435 ;
    END
  END BcidMtx[1257]
  PIN BcidMtx[1255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17882.265 1046.435 17882.545 1047.435 ;
    END
  END BcidMtx[1255]
  PIN Data_HV[864]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17879.465 1046.435 17879.745 1047.435 ;
    END
  END Data_HV[864]
  PIN Data_HV[870]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17878.345 1046.435 17878.625 1047.435 ;
    END
  END Data_HV[870]
  PIN Data_HV[877]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17876.105 1046.435 17876.385 1047.435 ;
    END
  END Data_HV[877]
  PIN Data_HV[861]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17874.425 1046.435 17874.705 1047.435 ;
    END
  END Data_HV[861]
  PIN MASKV[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17834.665 1046.435 17834.945 1047.435 ;
    END
  END MASKV[418]
  PIN MASKD[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17829.065 1046.435 17829.345 1047.435 ;
    END
  END MASKD[417]
  PIN INJ_ROW[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17826.825 1046.435 17827.105 1047.435 ;
    END
  END INJ_ROW[208]
  PIN Data_HV[852]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17824.585 1046.435 17824.865 1047.435 ;
    END
  END Data_HV[852]
  PIN Data_HV[853]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17822.905 1046.435 17823.185 1047.435 ;
    END
  END Data_HV[853]
  PIN Data_HV[854]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17821.785 1046.435 17822.065 1047.435 ;
    END
  END Data_HV[854]
  PIN nTOK_HV[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17810.025 1046.435 17810.305 1047.435 ;
    END
  END nTOK_HV[40]
  PIN BcidMtx[1251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17807.785 1046.435 17808.065 1047.435 ;
    END
  END BcidMtx[1251]
  PIN Read_HV[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17806.665 1046.435 17806.945 1047.435 ;
    END
  END Read_HV[40]
  PIN INJ_IN[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17801.905 1046.435 17802.185 1047.435 ;
    END
  END INJ_IN[416]
  PIN Data_HV[849]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17799.665 1046.435 17799.945 1047.435 ;
    END
  END Data_HV[849]
  PIN Data_HV[850]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17798.545 1046.435 17798.825 1047.435 ;
    END
  END Data_HV[850]
  PIN Data_HV[563]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16649.705 1046.435 16649.985 1047.435 ;
    END
  END Data_HV[563]
  PIN MASKH[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16648.585 1046.435 16648.865 1047.435 ;
    END
  END MASKH[194]
  PIN DIG_MON_HV[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16642.425 1046.435 16642.705 1047.435 ;
    END
  END DIG_MON_HV[51]
  PIN INJ_ROW[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16641.305 1046.435 16641.585 1047.435 ;
    END
  END INJ_ROW[193]
  PIN Data_HV[543]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16640.185 1046.435 16640.465 1047.435 ;
    END
  END Data_HV[543]
  PIN Data_HV[538]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16624.505 1046.435 16624.785 1047.435 ;
    END
  END Data_HV[538]
  PIN BcidMtx[1310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18604.665 1046.435 18604.945 1047.435 ;
    END
  END BcidMtx[1310]
  PIN Data_HV[532]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16622.825 1046.435 16623.105 1047.435 ;
    END
  END Data_HV[532]
  PIN BcidMtx[1162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16618.345 1046.435 16618.625 1047.435 ;
    END
  END BcidMtx[1162]
  PIN FREEZE_HV[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16617.225 1046.435 16617.505 1047.435 ;
    END
  END FREEZE_HV[25]
  PIN BcidMtx[1160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16616.105 1046.435 16616.385 1047.435 ;
    END
  END BcidMtx[1160]
  PIN Data_HV[527]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16573.545 1046.435 16573.825 1047.435 ;
    END
  END Data_HV[527]
  PIN Data_HV[540]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16572.425 1046.435 16572.705 1047.435 ;
    END
  END Data_HV[540]
  PIN Data_HV[529]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16571.305 1046.435 16571.585 1047.435 ;
    END
  END Data_HV[529]
  PIN Data_HV[542]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16568.505 1046.435 16568.785 1047.435 ;
    END
  END Data_HV[542]
  PIN MASKH[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16567.385 1046.435 16567.665 1047.435 ;
    END
  END MASKH[193]
  PIN DIG_MON_HV[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16565.705 1046.435 16565.985 1047.435 ;
    END
  END DIG_MON_HV[50]
  PIN DIG_MON_HV[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16561.225 1046.435 16561.505 1047.435 ;
    END
  END DIG_MON_HV[49]
  PIN MASKV[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16551.145 1046.435 16551.425 1047.435 ;
    END
  END MASKV[385]
  PIN Data_HV[512]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16550.025 1046.435 16550.305 1047.435 ;
    END
  END Data_HV[512]
  PIN Data_HV[517]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16547.785 1046.435 16548.065 1047.435 ;
    END
  END Data_HV[517]
  PIN Data_HV[518]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16546.665 1046.435 16546.945 1047.435 ;
    END
  END Data_HV[518]
  PIN BcidMtx[1308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18603.545 1046.435 18603.825 1047.435 ;
    END
  END BcidMtx[1308]
  PIN BcidMtx[1156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16539.665 1046.435 16539.945 1047.435 ;
    END
  END BcidMtx[1156]
  PIN Read_HV[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16512.505 1046.435 16512.785 1047.435 ;
    END
  END Read_HV[24]
  PIN BcidMtx[1153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16511.385 1046.435 16511.665 1047.435 ;
    END
  END BcidMtx[1153]
  PIN Data_HV[513]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16507.465 1046.435 16507.745 1047.435 ;
    END
  END Data_HV[513]
  PIN Data_HV[514]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16506.345 1046.435 16506.625 1047.435 ;
    END
  END Data_HV[514]
  PIN Data_HV[520]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16505.225 1046.435 16505.505 1047.435 ;
    END
  END Data_HV[520]
  PIN MASKV[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16502.425 1046.435 16502.705 1047.435 ;
    END
  END MASKV[384]
  PIN MASKD[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16501.305 1046.435 16501.585 1047.435 ;
    END
  END MASKD[384]
  PIN INJ_ROW[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16481.705 1046.435 16481.985 1047.435 ;
    END
  END INJ_ROW[191]
  PIN Data_HV[501]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16480.585 1046.435 16480.865 1047.435 ;
    END
  END Data_HV[501]
  PIN Data_HV[495]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16479.465 1046.435 16479.745 1047.435 ;
    END
  END Data_HV[495]
  PIN Data_HV[497]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16476.665 1046.435 16476.945 1047.435 ;
    END
  END Data_HV[497]
  PIN Data_HV[489]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16475.545 1046.435 16475.825 1047.435 ;
    END
  END Data_HV[489]
  PIN INJ_IN[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18714.425 1046.435 18714.705 1047.435 ;
    END
  END INJ_IN[439]
  PIN FREEZE_HV[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16431.305 1046.435 16431.585 1047.435 ;
    END
  END FREEZE_HV[23]
  PIN BcidMtx[1148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16430.185 1046.435 16430.465 1047.435 ;
    END
  END BcidMtx[1148]
  PIN BcidMtx[1146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16429.065 1046.435 16429.345 1047.435 ;
    END
  END BcidMtx[1146]
  PIN Data_HV[498]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16425.145 1046.435 16425.425 1047.435 ;
    END
  END Data_HV[498]
  PIN Data_HV[487]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16424.025 1046.435 16424.305 1047.435 ;
    END
  END Data_HV[487]
  PIN Data_HV[494]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16422.905 1046.435 16423.185 1047.435 ;
    END
  END Data_HV[494]
  PIN MASKH[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16411.705 1046.435 16411.985 1047.435 ;
    END
  END MASKH[191]
  PIN DIG_MON_HV[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16410.025 1046.435 16410.305 1047.435 ;
    END
  END DIG_MON_HV[46]
  PIN DIG_MON_SEL[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16408.345 1046.435 16408.625 1047.435 ;
    END
  END DIG_MON_SEL[382]
  PIN MASKV[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16401.905 1046.435 16402.185 1047.435 ;
    END
  END MASKV[381]
  PIN Data_HV[470]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16400.785 1046.435 16401.065 1047.435 ;
    END
  END Data_HV[470]
  PIN Data_HV[481]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16399.665 1046.435 16399.945 1047.435 ;
    END
  END Data_HV[481]
  PIN Data_HV[469]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16371.385 1046.435 16371.665 1047.435 ;
    END
  END Data_HV[469]
  PIN INJ_IN[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16369.705 1046.435 16369.985 1047.435 ;
    END
  END INJ_IN[381]
  PIN BcidMtx[1145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16367.465 1046.435 16367.745 1047.435 ;
    END
  END BcidMtx[1145]
  PIN BcidMtx[1142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16364.665 1046.435 16364.945 1047.435 ;
    END
  END BcidMtx[1142]
  PIN BcidMtx[1140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16363.545 1046.435 16363.825 1047.435 ;
    END
  END BcidMtx[1140]
  PIN Data_HV[465]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16361.305 1046.435 16361.585 1047.435 ;
    END
  END Data_HV[465]
  PIN Data_HV[466]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16345.625 1046.435 16345.905 1047.435 ;
    END
  END Data_HV[466]
  PIN Data_HV[473]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16344.505 1046.435 16344.785 1047.435 ;
    END
  END Data_HV[473]
  PIN Data_HV[462]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16343.385 1046.435 16343.665 1047.435 ;
    END
  END Data_HV[462]
  PIN MASKD[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16341.145 1046.435 16341.425 1047.435 ;
    END
  END MASKD[380]
  PIN DIG_MON_SEL[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16338.345 1046.435 16338.625 1047.435 ;
    END
  END DIG_MON_SEL[380]
  PIN MASKD[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16336.665 1046.435 16336.945 1047.435 ;
    END
  END MASKD[379]
  PIN Data_HV[459]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16293.545 1046.435 16293.825 1047.435 ;
    END
  END Data_HV[459]
  PIN Data_HV[460]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16291.865 1046.435 16292.145 1047.435 ;
    END
  END Data_HV[460]
  PIN Data_HV[454]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16290.745 1046.435 16291.025 1047.435 ;
    END
  END Data_HV[454]
  PIN INJ_IN[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16287.385 1046.435 16287.665 1047.435 ;
    END
  END INJ_IN[379]
  PIN nTOK_HV[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18674.105 1046.435 18674.385 1047.435 ;
    END
  END nTOK_HV[51]
  PIN BcidMtx[1138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16284.585 1046.435 16284.865 1047.435 ;
    END
  END BcidMtx[1138]
  PIN BcidMtx[1135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16281.785 1046.435 16282.065 1047.435 ;
    END
  END BcidMtx[1135]
  PIN Data_HV[444]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16270.585 1046.435 16270.865 1047.435 ;
    END
  END Data_HV[444]
  PIN Data_HV[450]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16269.465 1046.435 16269.745 1047.435 ;
    END
  END Data_HV[450]
  PIN Data_HV[457]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16267.225 1046.435 16267.505 1047.435 ;
    END
  END Data_HV[457]
  PIN Data_HV[441]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16265.545 1046.435 16265.825 1047.435 ;
    END
  END Data_HV[441]
  PIN MASKV[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16262.465 1046.435 16262.745 1047.435 ;
    END
  END MASKV[378]
  PIN DIG_MON_HV[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16260.225 1046.435 16260.505 1047.435 ;
    END
  END DIG_MON_HV[42]
  PIN FREEZE_HV[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16513.065 1046.435 16513.345 1047.435 ;
    END
  END FREEZE_HV[24]
  PIN MASKD[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17350.825 1046.435 17351.105 1047.435 ;
    END
  END MASKD[405]
  PIN Data_HV[732]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17347.465 1046.435 17347.745 1047.435 ;
    END
  END Data_HV[732]
  PIN Data_HV[733]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17345.785 1046.435 17346.065 1047.435 ;
    END
  END Data_HV[733]
  PIN Data_HV[727]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17344.665 1046.435 17344.945 1047.435 ;
    END
  END Data_HV[727]
  PIN Data_HV[720]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17342.425 1046.435 17342.705 1047.435 ;
    END
  END Data_HV[720]
  PIN BcidMtx[1217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17325.625 1046.435 17325.905 1047.435 ;
    END
  END BcidMtx[1217]
  PIN BcidMtx[1215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17324.505 1046.435 17324.785 1047.435 ;
    END
  END BcidMtx[1215]
  PIN BcidMtx[1213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17322.265 1046.435 17322.545 1047.435 ;
    END
  END BcidMtx[1213]
  PIN Data_HV[717]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17319.465 1046.435 17319.745 1047.435 ;
    END
  END Data_HV[717]
  PIN Data_HV[723]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17318.345 1046.435 17318.625 1047.435 ;
    END
  END Data_HV[723]
  PIN Data_HV[730]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17316.105 1046.435 17316.385 1047.435 ;
    END
  END Data_HV[730]
  PIN Data_HV[714]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17314.425 1046.435 17314.705 1047.435 ;
    END
  END Data_HV[714]
  PIN MASKV[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17274.665 1046.435 17274.945 1047.435 ;
    END
  END MASKV[404]
  PIN DIG_MON_SEL[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17270.745 1046.435 17271.025 1047.435 ;
    END
  END DIG_MON_SEL[404]
  PIN DIG_MON_HV[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17267.945 1046.435 17268.225 1047.435 ;
    END
  END DIG_MON_HV[67]
  PIN MASKV[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17266.265 1046.435 17266.545 1047.435 ;
    END
  END MASKV[403]
  PIN Data_HV[712]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17264.025 1046.435 17264.305 1047.435 ;
    END
  END Data_HV[712]
  PIN Data_HV[713]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17262.345 1046.435 17262.625 1047.435 ;
    END
  END Data_HV[713]
  PIN Data_HV[700]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17261.225 1046.435 17261.505 1047.435 ;
    END
  END Data_HV[700]
  PIN BcidMtx[1211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17248.905 1046.435 17249.185 1047.435 ;
    END
  END BcidMtx[1211]
  PIN FREEZE_HV[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17247.225 1046.435 17247.505 1047.435 ;
    END
  END FREEZE_HV[33]
  PIN BcidMtx[1208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17246.105 1046.435 17246.385 1047.435 ;
    END
  END BcidMtx[1208]
  PIN Data_HV[696]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17240.785 1046.435 17241.065 1047.435 ;
    END
  END Data_HV[696]
  PIN Data_HV[708]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17239.105 1046.435 17239.385 1047.435 ;
    END
  END Data_HV[708]
  PIN Data_HV[697]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17212.505 1046.435 17212.785 1047.435 ;
    END
  END Data_HV[697]
  PIN DIG_MON_PMOS_NOSF[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2229.705 1046.435 2229.985 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[27]
  PIN INJ_ROW[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2228.585 1046.435 2228.865 1047.435 ;
    END
  END INJ_ROW[13]
  PIN Data_PMOS_NOSF[292]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2225.785 1046.435 2226.065 1047.435 ;
    END
  END Data_PMOS_NOSF[292]
  PIN Data_PMOS_NOSF[293]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2224.105 1046.435 2224.385 1047.435 ;
    END
  END Data_PMOS_NOSF[293]
  PIN Data_PMOS_NOSF[287]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2223.545 1046.435 2223.825 1047.435 ;
    END
  END Data_PMOS_NOSF[287]
  PIN BcidMtx[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2205.625 1046.435 2205.905 1047.435 ;
    END
  END BcidMtx[83]
  PIN FREEZE_PMOS_NOSF[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2203.945 1046.435 2204.225 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[13]
  PIN Read_PMOS_NOSF[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2203.385 1046.435 2203.665 1047.435 ;
    END
  END Read_PMOS_NOSF[13]
  PIN Data_PMOS_NOSF[276]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2199.465 1046.435 2199.745 1047.435 ;
    END
  END Data_PMOS_NOSF[276]
  PIN Data_PMOS_NOSF[288]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2197.785 1046.435 2198.065 1047.435 ;
    END
  END Data_PMOS_NOSF[288]
  PIN Data_PMOS_NOSF[283]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2197.225 1046.435 2197.505 1047.435 ;
    END
  END Data_PMOS_NOSF[283]
  PIN Data_PMOS_NOSF[273]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2194.425 1046.435 2194.705 1047.435 ;
    END
  END Data_PMOS_NOSF[273]
  PIN MASKH[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2154.105 1046.435 2154.385 1047.435 ;
    END
  END MASKH[13]
  PIN MASKD[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2153.545 1046.435 2153.825 1047.435 ;
    END
  END MASKD[26]
  PIN DIG_MON_SEL[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2150.185 1046.435 2150.465 1047.435 ;
    END
  END DIG_MON_SEL[25]
  PIN DIG_MON_PMOS_NOSF[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2147.945 1046.435 2148.225 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[25]
  PIN INJ_ROW[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2146.825 1046.435 2147.105 1047.435 ;
    END
  END INJ_ROW[12]
  PIN Data_PMOS_NOSF[257]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2143.465 1046.435 2143.745 1047.435 ;
    END
  END Data_PMOS_NOSF[257]
  PIN Data_PMOS_NOSF[272]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2142.345 1046.435 2142.625 1047.435 ;
    END
  END Data_PMOS_NOSF[272]
  PIN Data_PMOS_NOSF[266]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2141.785 1046.435 2142.065 1047.435 ;
    END
  END Data_PMOS_NOSF[266]
  PIN BcidMtx[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2128.905 1046.435 2129.185 1047.435 ;
    END
  END BcidMtx[77]
  PIN FREEZE_PMOS_NOSF[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2127.225 1046.435 2127.505 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[12]
  PIN Read_PMOS_NOSF[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2126.665 1046.435 2126.945 1047.435 ;
    END
  END Read_PMOS_NOSF[12]
  PIN MASKD[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1941.305 1046.435 1941.585 1047.435 ;
    END
  END MASKD[20]
  PIN Data_PMOS_NOSF[261]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2119.665 1046.435 2119.945 1047.435 ;
    END
  END Data_PMOS_NOSF[261]
  PIN Data_PMOS_NOSF[267]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2119.105 1046.435 2119.385 1047.435 ;
    END
  END Data_PMOS_NOSF[267]
  PIN Data_PMOS_NOSF[253]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2090.825 1046.435 2091.105 1047.435 ;
    END
  END Data_PMOS_NOSF[253]
  PIN MASKV[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2089.145 1046.435 2089.425 1047.435 ;
    END
  END MASKV[24]
  PIN MASKH[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2088.585 1046.435 2088.865 1047.435 ;
    END
  END MASKH[12]
  PIN DIG_MON_SEL[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2084.665 1046.435 2084.945 1047.435 ;
    END
  END DIG_MON_SEL[23]
  PIN INJ_ROW[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2081.305 1046.435 2081.585 1047.435 ;
    END
  END INJ_ROW[11]
  PIN MASKV[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2080.745 1046.435 2081.025 1047.435 ;
    END
  END MASKV[23]
  PIN Data_PMOS_NOSF[236]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2065.065 1046.435 2065.345 1047.435 ;
    END
  END Data_PMOS_NOSF[236]
  PIN Data_PMOS_NOSF[245]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2063.385 1046.435 2063.665 1047.435 ;
    END
  END Data_PMOS_NOSF[245]
  PIN Data_PMOS_NOSF[238]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2062.825 1046.435 2063.105 1047.435 ;
    END
  END Data_PMOS_NOSF[238]
  PIN BcidMtx[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2058.345 1046.435 2058.625 1047.435 ;
    END
  END BcidMtx[70]
  PIN Read_PMOS_NOSF[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2056.665 1046.435 2056.945 1047.435 ;
    END
  END Read_PMOS_NOSF[11]
  PIN BcidMtx[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2055.545 1046.435 2055.825 1047.435 ;
    END
  END BcidMtx[67]
  PIN Data_PMOS_NOSF[240]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2012.985 1046.435 2013.265 1047.435 ;
    END
  END Data_PMOS_NOSF[240]
  PIN Data_PMOS_NOSF[235]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2011.305 1046.435 2011.585 1047.435 ;
    END
  END Data_PMOS_NOSF[235]
  PIN Data_PMOS_NOSF[247]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2010.745 1046.435 2011.025 1047.435 ;
    END
  END Data_PMOS_NOSF[247]
  PIN MASKV[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2007.945 1046.435 2008.225 1047.435 ;
    END
  END MASKV[22]
  PIN DIG_MON_PMOS_NOSF[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2005.705 1046.435 2005.985 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[22]
  PIN DIG_MON_PMOS_NOSF[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2001.225 1046.435 2001.505 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[21]
  PIN Data_PMOS_NOSF[228]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1990.585 1046.435 1990.865 1047.435 ;
    END
  END Data_PMOS_NOSF[228]
  PIN Data_PMOS_NOSF[218]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1990.025 1046.435 1990.305 1047.435 ;
    END
  END Data_PMOS_NOSF[218]
  PIN Data_PMOS_NOSF[230]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1987.225 1046.435 1987.505 1047.435 ;
    END
  END Data_PMOS_NOSF[230]
  PIN Data_PMOS_NOSF[216]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1985.545 1046.435 1985.825 1047.435 ;
    END
  END Data_PMOS_NOSF[216]
  PIN INJ_IN[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1982.465 1046.435 1982.745 1047.435 ;
    END
  END INJ_IN[21]
  PIN Read_PMOS_NOSF[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1952.505 1046.435 1952.785 1047.435 ;
    END
  END Read_PMOS_NOSF[10]
  PIN BcidMtx[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1950.825 1046.435 1951.105 1047.435 ;
    END
  END BcidMtx[60]
  PIN Data_PMOS_NOSF[213]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1948.585 1046.435 1948.865 1047.435 ;
    END
  END Data_PMOS_NOSF[213]
  PIN Data_PMOS_NOSF[220]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1946.345 1046.435 1946.625 1047.435 ;
    END
  END Data_PMOS_NOSF[220]
  PIN Data_PMOS_NOSF[226]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1945.225 1046.435 1945.505 1047.435 ;
    END
  END Data_PMOS_NOSF[226]
  PIN Data_PMOS_NOSF[211]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1944.105 1046.435 1944.385 1047.435 ;
    END
  END Data_PMOS_NOSF[211]
  PIN MASKV[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1942.425 1046.435 1942.705 1047.435 ;
    END
  END MASKV[20]
  PIN DIG_MON_SEL[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1925.065 1046.435 1925.345 1047.435 ;
    END
  END DIG_MON_SEL[19]
  PIN MASKD[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1923.945 1046.435 1924.225 1047.435 ;
    END
  END MASKD[19]
  PIN MASKV[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1921.145 1046.435 1921.425 1047.435 ;
    END
  END MASKV[19]
  PIN Data_PMOS_NOSF[201]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1919.465 1046.435 1919.745 1047.435 ;
    END
  END Data_PMOS_NOSF[201]
  PIN Data_PMOS_NOSF[202]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1917.785 1046.435 1918.065 1047.435 ;
    END
  END Data_PMOS_NOSF[202]
  PIN Data_PMOS_NOSF[196]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1916.105 1046.435 1916.385 1047.435 ;
    END
  END Data_PMOS_NOSF[196]
  PIN nTOK_PMOS_NOSF[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1874.105 1046.435 1874.385 1047.435 ;
    END
  END nTOK_PMOS_NOSF[9]
  PIN BcidMtx[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1871.865 1046.435 1872.145 1047.435 ;
    END
  END BcidMtx[57]
  PIN BcidMtx[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1869.625 1046.435 1869.905 1047.435 ;
    END
  END BcidMtx[55]
  PIN INJ_IN[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1867.945 1046.435 1868.225 1047.435 ;
    END
  END INJ_IN[18]
  PIN Data_PMOS_NOSF[198]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1865.705 1046.435 1865.985 1047.435 ;
    END
  END Data_PMOS_NOSF[198]
  PIN Data_PMOS_NOSF[205]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1863.465 1046.435 1863.745 1047.435 ;
    END
  END Data_PMOS_NOSF[205]
  PIN Data_PMOS_NOSF[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1861.785 1046.435 1862.065 1047.435 ;
    END
  END Data_PMOS_NOSF[189]
  PIN MASKH[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1851.705 1046.435 1851.985 1047.435 ;
    END
  END MASKH[9]
  PIN MASKD[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1846.665 1046.435 1846.945 1047.435 ;
    END
  END MASKD[17]
  PIN INJ_ROW[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1842.465 1046.435 1842.745 1047.435 ;
    END
  END INJ_ROW[8]
  PIN Data_PMOS_NOSF[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1840.225 1046.435 1840.505 1047.435 ;
    END
  END Data_PMOS_NOSF[180]
  PIN Data_PMOS_NOSF[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1813.065 1046.435 1813.345 1047.435 ;
    END
  END Data_PMOS_NOSF[181]
  PIN Data_PMOS_NOSF[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1811.385 1046.435 1811.665 1047.435 ;
    END
  END Data_PMOS_NOSF[175]
  PIN nTOK_PMOS_NOSF[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1808.585 1046.435 1808.865 1047.435 ;
    END
  END nTOK_PMOS_NOSF[8]
  PIN BcidMtx[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1806.345 1046.435 1806.625 1047.435 ;
    END
  END BcidMtx[51]
  PIN BcidMtx[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1804.105 1046.435 1804.385 1047.435 ;
    END
  END BcidMtx[49]
  PIN Data_PMOS_NOSF[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1801.305 1046.435 1801.585 1047.435 ;
    END
  END Data_PMOS_NOSF[171]
  PIN Data_PMOS_NOSF[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1786.745 1046.435 1787.025 1047.435 ;
    END
  END Data_PMOS_NOSF[183]
  PIN Data_PMOS_NOSF[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1785.625 1046.435 1785.905 1047.435 ;
    END
  END Data_PMOS_NOSF[172]
  PIN Data_PMOS_NOSF[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1784.505 1046.435 1784.785 1047.435 ;
    END
  END Data_PMOS_NOSF[179]
  PIN Data_PMOS_NOSF[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1782.825 1046.435 1783.105 1047.435 ;
    END
  END Data_PMOS_NOSF[185]
  PIN MASKD[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1781.145 1046.435 1781.425 1047.435 ;
    END
  END MASKD[16]
  PIN MASKD[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1776.665 1046.435 1776.945 1047.435 ;
    END
  END MASKD[15]
  PIN INJ_ROW[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1774.425 1046.435 1774.705 1047.435 ;
    END
  END INJ_ROW[7]
  PIN Data_PMOS_NOSF[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1732.985 1046.435 1733.265 1047.435 ;
    END
  END Data_PMOS_NOSF[155]
  PIN Data_PMOS_NOSF[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1730.745 1046.435 1731.025 1047.435 ;
    END
  END Data_PMOS_NOSF[160]
  PIN Data_PMOS_NOSF[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1729.625 1046.435 1729.905 1047.435 ;
    END
  END Data_PMOS_NOSF[161]
  PIN INJ_IN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1727.385 1046.435 1727.665 1047.435 ;
    END
  END INJ_IN[15]
  PIN BcidMtx[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1724.585 1046.435 1724.865 1047.435 ;
    END
  END BcidMtx[46]
  PIN Read_PMOS_NOSF[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1722.905 1046.435 1723.185 1047.435 ;
    END
  END Read_PMOS_NOSF[7]
  PIN BcidMtx[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1721.225 1046.435 1721.505 1047.435 ;
    END
  END BcidMtx[42]
  PIN Data_PMOS_NOSF[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1710.025 1046.435 1710.305 1047.435 ;
    END
  END Data_PMOS_NOSF[149]
  PIN Data_PMOS_NOSF[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1708.345 1046.435 1708.625 1047.435 ;
    END
  END Data_PMOS_NOSF[157]
  PIN Data_PMOS_NOSF[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1706.665 1046.435 1706.945 1047.435 ;
    END
  END Data_PMOS_NOSF[158]
  PIN MASKV[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1702.465 1046.435 1702.745 1047.435 ;
    END
  END MASKV[14]
  PIN DIG_MON_SEL[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18577.785 1046.435 18578.065 1047.435 ;
    END
  END DIG_MON_SEL[435]
  PIN DIG_MON_SEL[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2791.945 1046.435 2792.225 1047.435 ;
    END
  END DIG_MON_SEL[41]
  PIN INJ_ROW[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2788.585 1046.435 2788.865 1047.435 ;
    END
  END INJ_ROW[20]
  PIN Data_PMOS_NOSF[428]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2786.905 1046.435 2787.185 1047.435 ;
    END
  END Data_PMOS_NOSF[428]
  PIN Data_PMOS_NOSF[425]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2785.225 1046.435 2785.505 1047.435 ;
    END
  END Data_PMOS_NOSF[425]
  PIN Data_PMOS_NOSF[434]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2783.545 1046.435 2783.825 1047.435 ;
    END
  END Data_PMOS_NOSF[434]
  PIN INJ_IN[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2781.305 1046.435 2781.585 1047.435 ;
    END
  END INJ_IN[41]
  PIN BcidMtx[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2765.065 1046.435 2765.345 1047.435 ;
    END
  END BcidMtx[124]
  PIN Read_PMOS_NOSF[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2763.385 1046.435 2763.665 1047.435 ;
    END
  END Read_PMOS_NOSF[20]
  PIN BcidMtx[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2761.705 1046.435 2761.985 1047.435 ;
    END
  END BcidMtx[120]
  PIN Data_PMOS_NOSF[429]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2758.345 1046.435 2758.625 1047.435 ;
    END
  END Data_PMOS_NOSF[429]
  PIN Data_PMOS_NOSF[430]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2757.225 1046.435 2757.505 1047.435 ;
    END
  END Data_PMOS_NOSF[430]
  PIN DIG_MON_SEL[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18578.345 1046.435 18578.625 1047.435 ;
    END
  END DIG_MON_SEL[436]
  PIN Data_PMOS_NOSF[420]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2754.425 1046.435 2754.705 1047.435 ;
    END
  END Data_PMOS_NOSF[420]
  PIN MASKH[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2714.105 1046.435 2714.385 1047.435 ;
    END
  END MASKH[20]
  PIN MASKD[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2709.065 1046.435 2709.345 1047.435 ;
    END
  END MASKD[39]
  PIN MASKV[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2706.265 1046.435 2706.545 1047.435 ;
    END
  END MASKV[39]
  PIN Data_PMOS_NOSF[407]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2705.145 1046.435 2705.425 1047.435 ;
    END
  END Data_PMOS_NOSF[407]
  PIN Data_PMOS_NOSF[419]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2702.345 1046.435 2702.625 1047.435 ;
    END
  END Data_PMOS_NOSF[419]
  PIN Data_PMOS_NOSF[413]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2701.785 1046.435 2702.065 1047.435 ;
    END
  END Data_PMOS_NOSF[413]
  PIN nTOK_PMOS_NOSF[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2690.025 1046.435 2690.305 1047.435 ;
    END
  END nTOK_PMOS_NOSF[19]
  PIN BcidMtx[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2687.785 1046.435 2688.065 1047.435 ;
    END
  END BcidMtx[117]
  PIN BcidMtx[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2686.105 1046.435 2686.385 1047.435 ;
    END
  END BcidMtx[116]
  PIN INJ_IN[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2681.905 1046.435 2682.185 1047.435 ;
    END
  END INJ_IN[38]
  PIN Data_PMOS_NOSF[401]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2680.225 1046.435 2680.505 1047.435 ;
    END
  END Data_PMOS_NOSF[401]
  PIN Data_PMOS_NOSF[409]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2678.545 1046.435 2678.825 1047.435 ;
    END
  END Data_PMOS_NOSF[409]
  PIN Data_PMOS_NOSF[410]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2651.385 1046.435 2651.665 1047.435 ;
    END
  END Data_PMOS_NOSF[410]
  PIN MASKD[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18576.665 1046.435 18576.945 1047.435 ;
    END
  END MASKD[435]
  PIN MASKH[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2648.585 1046.435 2648.865 1047.435 ;
    END
  END MASKH[19]
  PIN DIG_MON_PMOS_NOSF[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2642.425 1046.435 2642.705 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[37]
  PIN MASKV[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2640.745 1046.435 2641.025 1047.435 ;
    END
  END MASKV[37]
  PIN Data_PMOS_NOSF[390]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2626.185 1046.435 2626.465 1047.435 ;
    END
  END Data_PMOS_NOSF[390]
  PIN Data_PMOS_NOSF[383]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2625.065 1046.435 2625.345 1047.435 ;
    END
  END Data_PMOS_NOSF[383]
  PIN Data_PMOS_NOSF[392]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2623.385 1046.435 2623.665 1047.435 ;
    END
  END Data_PMOS_NOSF[392]
  PIN Data_PMOS_NOSF[384]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2622.265 1046.435 2622.545 1047.435 ;
    END
  END Data_PMOS_NOSF[384]
  PIN BcidMtx[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2618.345 1046.435 2618.625 1047.435 ;
    END
  END BcidMtx[112]
  PIN Read_PMOS_NOSF[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2616.665 1046.435 2616.945 1047.435 ;
    END
  END Read_PMOS_NOSF[18]
  PIN BcidMtx[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2615.545 1046.435 2615.825 1047.435 ;
    END
  END BcidMtx[109]
  PIN Data_PMOS_NOSF[381]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2574.105 1046.435 2574.385 1047.435 ;
    END
  END Data_PMOS_NOSF[381]
  PIN Data_PMOS_NOSF[393]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2572.425 1046.435 2572.705 1047.435 ;
    END
  END Data_PMOS_NOSF[393]
  PIN Data_PMOS_NOSF[394]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2570.745 1046.435 2571.025 1047.435 ;
    END
  END Data_PMOS_NOSF[394]
  PIN Data_PMOS_NOSF[378]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2569.065 1046.435 2569.345 1047.435 ;
    END
  END Data_PMOS_NOSF[378]
  PIN MASKV[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2567.945 1046.435 2568.225 1047.435 ;
    END
  END MASKV[36]
  PIN MASKD[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2562.345 1046.435 2562.625 1047.435 ;
    END
  END MASKD[35]
  PIN INJ_ROW[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2551.705 1046.435 2551.985 1047.435 ;
    END
  END INJ_ROW[17]
  PIN Data_PMOS_NOSF[365]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2550.025 1046.435 2550.305 1047.435 ;
    END
  END Data_PMOS_NOSF[365]
  PIN Data_PMOS_NOSF[370]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2547.785 1046.435 2548.065 1047.435 ;
    END
  END Data_PMOS_NOSF[370]
  PIN Data_PMOS_NOSF[371]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2546.665 1046.435 2546.945 1047.435 ;
    END
  END Data_PMOS_NOSF[371]
  PIN Data_PMOS_NOSF[363]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2545.545 1046.435 2545.825 1047.435 ;
    END
  END Data_PMOS_NOSF[363]
  PIN BcidMtx[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2540.225 1046.435 2540.505 1047.435 ;
    END
  END BcidMtx[107]
  PIN BcidMtx[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2511.945 1046.435 2512.225 1047.435 ;
    END
  END BcidMtx[104]
  PIN BcidMtx[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2510.825 1046.435 2511.105 1047.435 ;
    END
  END BcidMtx[102]
  PIN Data_PMOS_NOSF[359]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2508.025 1046.435 2508.305 1047.435 ;
    END
  END Data_PMOS_NOSF[359]
  PIN Data_PMOS_NOSF[361]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2505.785 1046.435 2506.065 1047.435 ;
    END
  END Data_PMOS_NOSF[361]
  PIN Data_PMOS_NOSF[358]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2504.105 1046.435 2504.385 1047.435 ;
    END
  END Data_PMOS_NOSF[358]
  PIN Data_PMOS_NOSF[374]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2502.985 1046.435 2503.265 1047.435 ;
    END
  END Data_PMOS_NOSF[374]
  PIN MASKD[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2501.305 1046.435 2501.585 1047.435 ;
    END
  END MASKD[34]
  PIN DIG_MON_SEL[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2485.065 1046.435 2485.345 1047.435 ;
    END
  END DIG_MON_SEL[33]
  PIN DIG_MON_PMOS_NOSF[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2482.825 1046.435 2483.105 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[33]
  PIN Data_PMOS_NOSF[354]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2480.585 1046.435 2480.865 1047.435 ;
    END
  END Data_PMOS_NOSF[354]
  PIN Data_PMOS_NOSF[348]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2479.465 1046.435 2479.745 1047.435 ;
    END
  END Data_PMOS_NOSF[348]
  PIN Data_PMOS_NOSF[349]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2477.785 1046.435 2478.065 1047.435 ;
    END
  END Data_PMOS_NOSF[349]
  PIN INJ_IN[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2474.425 1046.435 2474.705 1047.435 ;
    END
  END INJ_IN[33]
  PIN BcidMtx[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2432.985 1046.435 2433.265 1047.435 ;
    END
  END BcidMtx[101]
  PIN Read_PMOS_NOSF[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2430.745 1046.435 2431.025 1047.435 ;
    END
  END Read_PMOS_NOSF[16]
  PIN BcidMtx[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2429.065 1046.435 2429.345 1047.435 ;
    END
  END BcidMtx[96]
  PIN Data_PMOS_NOSF[339]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2426.825 1046.435 2427.105 1047.435 ;
    END
  END Data_PMOS_NOSF[339]
  PIN Data_PMOS_NOSF[351]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2425.145 1046.435 2425.425 1047.435 ;
    END
  END Data_PMOS_NOSF[351]
  PIN Data_PMOS_NOSF[347]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2422.905 1046.435 2423.185 1047.435 ;
    END
  END Data_PMOS_NOSF[347]
  PIN Data_PMOS_NOSF[337]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2422.345 1046.435 2422.625 1047.435 ;
    END
  END Data_PMOS_NOSF[337]
  PIN MASKH[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2411.705 1046.435 2411.985 1047.435 ;
    END
  END MASKH[16]
  PIN DIG_MON_SEL[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2408.345 1046.435 2408.625 1047.435 ;
    END
  END DIG_MON_SEL[32]
  PIN MASKV[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2401.905 1046.435 2402.185 1047.435 ;
    END
  END MASKV[31]
  PIN Data_PMOS_NOSF[323]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2400.785 1046.435 2401.065 1047.435 ;
    END
  END Data_PMOS_NOSF[323]
  PIN Data_PMOS_NOSF[328]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2373.065 1046.435 2373.345 1047.435 ;
    END
  END Data_PMOS_NOSF[328]
  PIN Data_PMOS_NOSF[321]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2370.825 1046.435 2371.105 1047.435 ;
    END
  END Data_PMOS_NOSF[321]
  PIN nTOK_PMOS_NOSF[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2368.585 1046.435 2368.865 1047.435 ;
    END
  END nTOK_PMOS_NOSF[15]
  PIN FREEZE_PMOS_NOSF[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2365.785 1046.435 2366.065 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[15]
  PIN BcidMtx[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2364.105 1046.435 2364.385 1047.435 ;
    END
  END BcidMtx[91]
  PIN INJ_IN[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2362.425 1046.435 2362.705 1047.435 ;
    END
  END INJ_IN[30]
  PIN Data_PMOS_NOSF[318]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2361.305 1046.435 2361.585 1047.435 ;
    END
  END Data_PMOS_NOSF[318]
  PIN Data_PMOS_NOSF[319]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2345.625 1046.435 2345.905 1047.435 ;
    END
  END Data_PMOS_NOSF[319]
  PIN Data_PMOS_NOSF[326]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2344.505 1046.435 2344.785 1047.435 ;
    END
  END Data_PMOS_NOSF[326]
  PIN MASKV[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2342.265 1046.435 2342.545 1047.435 ;
    END
  END MASKV[30]
  PIN DIG_MON_PMOS_NOSF[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2340.025 1046.435 2340.305 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[30]
  PIN DIG_MON_SEL[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2338.345 1046.435 2338.625 1047.435 ;
    END
  END DIG_MON_SEL[30]
  PIN INJ_ROW[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2334.425 1046.435 2334.705 1047.435 ;
    END
  END INJ_ROW[14]
  PIN Data_PMOS_NOSF[306]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2292.425 1046.435 2292.705 1047.435 ;
    END
  END Data_PMOS_NOSF[306]
  PIN Data_PMOS_NOSF[299]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2291.305 1046.435 2291.585 1047.435 ;
    END
  END Data_PMOS_NOSF[299]
  PIN Data_PMOS_NOSF[301]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2289.065 1046.435 2289.345 1047.435 ;
    END
  END Data_PMOS_NOSF[301]
  PIN nTOK_PMOS_NOSF[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2286.265 1046.435 2286.545 1047.435 ;
    END
  END nTOK_PMOS_NOSF[14]
  PIN BcidMtx[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2284.585 1046.435 2284.865 1047.435 ;
    END
  END BcidMtx[88]
  PIN FREEZE_PMOS_NOSF[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2283.465 1046.435 2283.745 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[14]
  PIN INJ_IN[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2271.705 1046.435 2271.985 1047.435 ;
    END
  END INJ_IN[28]
  PIN Data_PMOS_NOSF[296]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2270.025 1046.435 2270.305 1047.435 ;
    END
  END Data_PMOS_NOSF[296]
  PIN Data_PMOS_NOSF[309]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2268.905 1046.435 2269.185 1047.435 ;
    END
  END Data_PMOS_NOSF[309]
  PIN Data_PMOS_NOSF[305]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2266.665 1046.435 2266.945 1047.435 ;
    END
  END Data_PMOS_NOSF[305]
  PIN Data_PMOS_NOSF[294]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2265.545 1046.435 2265.825 1047.435 ;
    END
  END Data_PMOS_NOSF[294]
  PIN MASKD[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2261.345 1046.435 2261.625 1047.435 ;
    END
  END MASKD[28]
  PIN DIG_MON_SEL[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2258.545 1046.435 2258.825 1047.435 ;
    END
  END DIG_MON_SEL[28]
  PIN MASKD[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3350.825 1046.435 3351.105 1047.435 ;
    END
  END MASKD[55]
  PIN Data_PMOS_NOSF[585]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3347.465 1046.435 3347.745 1047.435 ;
    END
  END Data_PMOS_NOSF[585]
  PIN Data_PMOS_NOSF[579]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3346.345 1046.435 3346.625 1047.435 ;
    END
  END Data_PMOS_NOSF[579]
  PIN Data_PMOS_NOSF[580]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3344.665 1046.435 3344.945 1047.435 ;
    END
  END Data_PMOS_NOSF[580]
  PIN Data_PMOS_NOSF[573]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3342.425 1046.435 3342.705 1047.435 ;
    END
  END Data_PMOS_NOSF[573]
  PIN BcidMtx[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3325.625 1046.435 3325.905 1047.435 ;
    END
  END BcidMtx[167]
  PIN BcidMtx[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3324.505 1046.435 3324.785 1047.435 ;
    END
  END BcidMtx[165]
  PIN BcidMtx[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3322.265 1046.435 3322.545 1047.435 ;
    END
  END BcidMtx[163]
  PIN Data_PMOS_NOSF[570]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3319.465 1046.435 3319.745 1047.435 ;
    END
  END Data_PMOS_NOSF[570]
  PIN Data_PMOS_NOSF[569]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3318.905 1046.435 3319.185 1047.435 ;
    END
  END Data_PMOS_NOSF[569]
  PIN Data_PMOS_NOSF[571]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3316.665 1046.435 3316.945 1047.435 ;
    END
  END Data_PMOS_NOSF[571]
  PIN DIG_MON_HV[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18886.905 1046.435 18887.185 1047.435 ;
    END
  END DIG_MON_HV[108]
  PIN Data_PMOS_NOSF[567]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3314.425 1046.435 3314.705 1047.435 ;
    END
  END Data_PMOS_NOSF[567]
  PIN MASKH[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3274.105 1046.435 3274.385 1047.435 ;
    END
  END MASKH[27]
  PIN DIG_MON_SEL[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3270.745 1046.435 3271.025 1047.435 ;
    END
  END DIG_MON_SEL[54]
  PIN MASKD[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3269.065 1046.435 3269.345 1047.435 ;
    END
  END MASKD[53]
  PIN MASKV[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3266.265 1046.435 3266.545 1047.435 ;
    END
  END MASKV[53]
  PIN Data_PMOS_NOSF[565]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3264.025 1046.435 3264.305 1047.435 ;
    END
  END Data_PMOS_NOSF[565]
  PIN Data_PMOS_NOSF[559]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3262.905 1046.435 3263.185 1047.435 ;
    END
  END Data_PMOS_NOSF[559]
  PIN Data_PMOS_NOSF[553]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3261.225 1046.435 3261.505 1047.435 ;
    END
  END Data_PMOS_NOSF[553]
  PIN BcidMtx[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3248.905 1046.435 3249.185 1047.435 ;
    END
  END BcidMtx[161]
  PIN BcidMtx[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3247.785 1046.435 3248.065 1047.435 ;
    END
  END BcidMtx[159]
  PIN BcidMtx[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3246.105 1046.435 3246.385 1047.435 ;
    END
  END BcidMtx[158]
  PIN INJ_IN[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3241.905 1046.435 3242.185 1047.435 ;
    END
  END INJ_IN[52]
  PIN Data_PMOS_NOSF[555]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3239.665 1046.435 3239.945 1047.435 ;
    END
  END Data_PMOS_NOSF[555]
  PIN Data_PMOS_NOSF[562]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3211.945 1046.435 3212.225 1047.435 ;
    END
  END Data_PMOS_NOSF[562]
  PIN Data_PMOS_NOSF[546]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3210.265 1046.435 3210.545 1047.435 ;
    END
  END Data_PMOS_NOSF[546]
  PIN MASKV[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3209.145 1046.435 3209.425 1047.435 ;
    END
  END MASKV[52]
  PIN DIG_MON_PMOS_NOSF[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3206.905 1046.435 3207.185 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[52]
  PIN MASKD[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3203.545 1046.435 3203.825 1047.435 ;
    END
  END MASKD[51]
  PIN MASKV[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3200.745 1046.435 3201.025 1047.435 ;
    END
  END MASKV[51]
  PIN Data_PMOS_NOSF[537]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3186.185 1046.435 3186.465 1047.435 ;
    END
  END Data_PMOS_NOSF[537]
  PIN Data_PMOS_NOSF[538]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3184.505 1046.435 3184.785 1047.435 ;
    END
  END Data_PMOS_NOSF[538]
  PIN Data_PMOS_NOSF[532]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3182.825 1046.435 3183.105 1047.435 ;
    END
  END Data_PMOS_NOSF[532]
  PIN nTOK_PMOS_NOSF[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3180.025 1046.435 3180.305 1047.435 ;
    END
  END nTOK_PMOS_NOSF[25]
  PIN BcidMtx[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3177.785 1046.435 3178.065 1047.435 ;
    END
  END BcidMtx[153]
  PIN BcidMtx[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3176.105 1046.435 3176.385 1047.435 ;
    END
  END BcidMtx[152]
  PIN BcidMtx[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3174.985 1046.435 3175.265 1047.435 ;
    END
  END BcidMtx[150]
  PIN Data_PMOS_NOSF[534]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3132.985 1046.435 3133.265 1047.435 ;
    END
  END Data_PMOS_NOSF[534]
  PIN Data_PMOS_NOSF[529]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3131.305 1046.435 3131.585 1047.435 ;
    END
  END Data_PMOS_NOSF[529]
  PIN Data_PMOS_NOSF[536]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3130.185 1046.435 3130.465 1047.435 ;
    END
  END Data_PMOS_NOSF[536]
  PIN Data_PMOS_NOSF[542]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3128.505 1046.435 3128.785 1047.435 ;
    END
  END Data_PMOS_NOSF[542]
  PIN MASKD[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3126.825 1046.435 3127.105 1047.435 ;
    END
  END MASKD[50]
  PIN DIG_MON_SEL[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3124.025 1046.435 3124.305 1047.435 ;
    END
  END DIG_MON_SEL[50]
  PIN DIG_MON_PMOS_NOSF[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3121.225 1046.435 3121.505 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[49]
  PIN Data_PMOS_NOSF[522]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3110.585 1046.435 3110.865 1047.435 ;
    END
  END Data_PMOS_NOSF[522]
  PIN Data_PMOS_NOSF[523]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3108.905 1046.435 3109.185 1047.435 ;
    END
  END Data_PMOS_NOSF[523]
  PIN Data_PMOS_NOSF[524]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3107.225 1046.435 3107.505 1047.435 ;
    END
  END Data_PMOS_NOSF[524]
  PIN Data_PMOS_NOSF[510]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3105.545 1046.435 3105.825 1047.435 ;
    END
  END Data_PMOS_NOSF[510]
  PIN nTOK_PMOS_NOSF[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3101.345 1046.435 3101.625 1047.435 ;
    END
  END nTOK_PMOS_NOSF[24]
  PIN Read_PMOS_NOSF[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3072.505 1046.435 3072.785 1047.435 ;
    END
  END Read_PMOS_NOSF[24]
  PIN BcidMtx[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3070.825 1046.435 3071.105 1047.435 ;
    END
  END BcidMtx[144]
  PIN Data_PMOS_NOSF[507]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3068.585 1046.435 3068.865 1047.435 ;
    END
  END Data_PMOS_NOSF[507]
  PIN Data_PMOS_NOSF[514]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3066.345 1046.435 3066.625 1047.435 ;
    END
  END Data_PMOS_NOSF[514]
  PIN Data_PMOS_NOSF[515]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3064.665 1046.435 3064.945 1047.435 ;
    END
  END Data_PMOS_NOSF[515]
  PIN Data_PMOS_NOSF[504]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3063.545 1046.435 3063.825 1047.435 ;
    END
  END Data_PMOS_NOSF[504]
  PIN MASKD[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3061.305 1046.435 3061.585 1047.435 ;
    END
  END MASKD[48]
  PIN DIG_MON_SEL[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3045.625 1046.435 3045.905 1047.435 ;
    END
  END DIG_MON_SEL[48]
  PIN MASKD[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3043.945 1046.435 3044.225 1047.435 ;
    END
  END MASKD[47]
  PIN Data_PMOS_NOSF[501]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3040.585 1046.435 3040.865 1047.435 ;
    END
  END Data_PMOS_NOSF[501]
  PIN Data_PMOS_NOSF[502]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3038.905 1046.435 3039.185 1047.435 ;
    END
  END Data_PMOS_NOSF[502]
  PIN Data_PMOS_NOSF[496]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3037.785 1046.435 3038.065 1047.435 ;
    END
  END Data_PMOS_NOSF[496]
  PIN Data_PMOS_NOSF[489]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3035.545 1046.435 3035.825 1047.435 ;
    END
  END Data_PMOS_NOSF[489]
  PIN BcidMtx[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2992.985 1046.435 2993.265 1047.435 ;
    END
  END BcidMtx[143]
  PIN FREEZE_PMOS_NOSF[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2991.305 1046.435 2991.585 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[23]
  PIN BcidMtx[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2989.625 1046.435 2989.905 1047.435 ;
    END
  END BcidMtx[139]
  PIN Data_PMOS_NOSF[486]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2986.825 1046.435 2987.105 1047.435 ;
    END
  END Data_PMOS_NOSF[486]
  PIN Data_PMOS_NOSF[498]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2985.145 1046.435 2985.425 1047.435 ;
    END
  END Data_PMOS_NOSF[498]
  PIN Data_PMOS_NOSF[499]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2983.465 1046.435 2983.745 1047.435 ;
    END
  END Data_PMOS_NOSF[499]
  PIN Data_PMOS_NOSF[483]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2981.785 1046.435 2982.065 1047.435 ;
    END
  END Data_PMOS_NOSF[483]
  PIN MASKH[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2971.705 1046.435 2971.985 1047.435 ;
    END
  END MASKH[23]
  PIN MASKD[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2966.665 1046.435 2966.945 1047.435 ;
    END
  END MASKD[45]
  PIN MASKV[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2961.905 1046.435 2962.185 1047.435 ;
    END
  END MASKV[45]
  PIN Data_PMOS_NOSF[474]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2960.225 1046.435 2960.505 1047.435 ;
    END
  END Data_PMOS_NOSF[474]
  PIN Data_PMOS_NOSF[475]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2933.065 1046.435 2933.345 1047.435 ;
    END
  END Data_PMOS_NOSF[475]
  PIN Data_PMOS_NOSF[468]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2930.825 1046.435 2931.105 1047.435 ;
    END
  END Data_PMOS_NOSF[468]
  PIN nTOK_PMOS_NOSF[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2928.585 1046.435 2928.865 1047.435 ;
    END
  END nTOK_PMOS_NOSF[22]
  PIN BcidMtx[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2926.345 1046.435 2926.625 1047.435 ;
    END
  END BcidMtx[135]
  PIN MASKD[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18888.025 1046.435 18888.305 1047.435 ;
    END
  END MASKD[444]
  PIN BcidMtx[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2924.105 1046.435 2924.385 1047.435 ;
    END
  END BcidMtx[133]
  PIN Data_PMOS_NOSF[465]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2921.305 1046.435 2921.585 1047.435 ;
    END
  END Data_PMOS_NOSF[465]
  PIN Data_PMOS_NOSF[477]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2906.745 1046.435 2907.025 1047.435 ;
    END
  END Data_PMOS_NOSF[477]
  PIN Data_PMOS_NOSF[478]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2905.065 1046.435 2905.345 1047.435 ;
    END
  END Data_PMOS_NOSF[478]
  PIN Data_PMOS_NOSF[462]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2903.385 1046.435 2903.665 1047.435 ;
    END
  END Data_PMOS_NOSF[462]
  PIN MASKH[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2901.705 1046.435 2901.985 1047.435 ;
    END
  END MASKH[22]
  PIN MASKD[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2896.665 1046.435 2896.945 1047.435 ;
    END
  END MASKD[43]
  PIN MASKV[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2893.865 1046.435 2894.145 1047.435 ;
    END
  END MASKV[43]
  PIN Data_PMOS_NOSF[453]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2852.425 1046.435 2852.705 1047.435 ;
    END
  END Data_PMOS_NOSF[453]
  PIN Data_PMOS_NOSF[454]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2850.745 1046.435 2851.025 1047.435 ;
    END
  END Data_PMOS_NOSF[454]
  PIN Data_PMOS_NOSF[448]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2849.065 1046.435 2849.345 1047.435 ;
    END
  END Data_PMOS_NOSF[448]
  PIN nTOK_PMOS_NOSF[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2846.265 1046.435 2846.545 1047.435 ;
    END
  END nTOK_PMOS_NOSF[21]
  PIN BcidMtx[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2844.025 1046.435 2844.305 1047.435 ;
    END
  END BcidMtx[129]
  PIN BcidMtx[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2842.345 1046.435 2842.625 1047.435 ;
    END
  END BcidMtx[128]
  PIN BcidMtx[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2841.225 1046.435 2841.505 1047.435 ;
    END
  END BcidMtx[126]
  PIN Data_PMOS_NOSF[443]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2830.025 1046.435 2830.305 1047.435 ;
    END
  END Data_PMOS_NOSF[443]
  PIN Data_PMOS_NOSF[451]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2828.345 1046.435 2828.625 1047.435 ;
    END
  END Data_PMOS_NOSF[451]
  PIN Data_PMOS_NOSF[452]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2826.665 1046.435 2826.945 1047.435 ;
    END
  END Data_PMOS_NOSF[452]
  PIN Data_PMOS_NOSF[458]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2824.985 1046.435 2825.265 1047.435 ;
    END
  END Data_PMOS_NOSF[458]
  PIN MASKD[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2821.345 1046.435 2821.625 1047.435 ;
    END
  END MASKD[42]
  PIN DIG_MON_SEL[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2818.545 1046.435 2818.825 1047.435 ;
    END
  END DIG_MON_SEL[42]
  PIN MASKD[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3910.825 1046.435 3911.105 1047.435 ;
    END
  END MASKD[69]
  PIN MASKV[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3908.025 1046.435 3908.305 1047.435 ;
    END
  END MASKV[69]
  PIN Data_PMOS_NOSF[726]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3906.345 1046.435 3906.625 1047.435 ;
    END
  END Data_PMOS_NOSF[726]
  PIN Data_PMOS_NOSF[727]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3904.665 1046.435 3904.945 1047.435 ;
    END
  END Data_PMOS_NOSF[727]
  PIN Data_PMOS_NOSF[721]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3902.985 1046.435 3903.265 1047.435 ;
    END
  END Data_PMOS_NOSF[721]
  PIN nTOK_PMOS_NOSF[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3900.185 1046.435 3900.465 1047.435 ;
    END
  END nTOK_PMOS_NOSF[34]
  PIN BcidMtx[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3884.505 1046.435 3884.785 1047.435 ;
    END
  END BcidMtx[207]
  PIN BcidMtx[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3882.825 1046.435 3883.105 1047.435 ;
    END
  END BcidMtx[206]
  PIN BcidMtx[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3881.705 1046.435 3881.985 1047.435 ;
    END
  END BcidMtx[204]
  PIN Data_PMOS_NOSF[716]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3878.905 1046.435 3879.185 1047.435 ;
    END
  END Data_PMOS_NOSF[716]
  PIN Data_PMOS_NOSF[724]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3877.225 1046.435 3877.505 1047.435 ;
    END
  END Data_PMOS_NOSF[724]
  PIN Data_PMOS_NOSF[725]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3875.545 1046.435 3875.825 1047.435 ;
    END
  END Data_PMOS_NOSF[725]
  PIN Data_PMOS_NOSF[731]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3873.865 1046.435 3874.145 1047.435 ;
    END
  END Data_PMOS_NOSF[731]
  PIN MASKD[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3833.545 1046.435 3833.825 1047.435 ;
    END
  END MASKD[68]
  PIN DIG_MON_SEL[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3830.185 1046.435 3830.465 1047.435 ;
    END
  END DIG_MON_SEL[67]
  PIN DIG_MON_PMOS_NOSF[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3827.945 1046.435 3828.225 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[67]
  PIN Data_PMOS_NOSF[711]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3825.705 1046.435 3825.985 1047.435 ;
    END
  END Data_PMOS_NOSF[711]
  PIN Data_PMOS_NOSF[712]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3824.025 1046.435 3824.305 1047.435 ;
    END
  END Data_PMOS_NOSF[712]
  PIN Data_PMOS_NOSF[713]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3822.345 1046.435 3822.625 1047.435 ;
    END
  END Data_PMOS_NOSF[713]
  PIN Data_PMOS_NOSF[700]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3821.225 1046.435 3821.505 1047.435 ;
    END
  END Data_PMOS_NOSF[700]
  PIN BcidMtx[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3808.905 1046.435 3809.185 1047.435 ;
    END
  END BcidMtx[203]
  PIN FREEZE_PMOS_NOSF[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3807.225 1046.435 3807.505 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[33]
  PIN BcidMtx[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3806.105 1046.435 3806.385 1047.435 ;
    END
  END BcidMtx[200]
  PIN MASKD[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18651.145 1046.435 18651.425 1047.435 ;
    END
  END MASKD[438]
  PIN Data_PMOS_NOSF[695]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3800.225 1046.435 3800.505 1047.435 ;
    END
  END Data_PMOS_NOSF[695]
  PIN Data_PMOS_NOSF[708]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3799.105 1046.435 3799.385 1047.435 ;
    END
  END Data_PMOS_NOSF[708]
  PIN Data_PMOS_NOSF[704]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3771.385 1046.435 3771.665 1047.435 ;
    END
  END Data_PMOS_NOSF[704]
  PIN Data_PMOS_NOSF[710]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3769.705 1046.435 3769.985 1047.435 ;
    END
  END Data_PMOS_NOSF[710]
  PIN MASKH[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3768.585 1046.435 3768.865 1047.435 ;
    END
  END MASKH[33]
  PIN DIG_MON_SEL[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3765.225 1046.435 3765.505 1047.435 ;
    END
  END DIG_MON_SEL[66]
  PIN DIG_MON_PMOS_NOSF[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3762.425 1046.435 3762.705 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[65]
  PIN MASKV[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3760.745 1046.435 3761.025 1047.435 ;
    END
  END MASKV[65]
  PIN Data_PMOS_NOSF[680]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3759.625 1046.435 3759.905 1047.435 ;
    END
  END Data_PMOS_NOSF[680]
  PIN Data_PMOS_NOSF[677]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3745.065 1046.435 3745.345 1047.435 ;
    END
  END Data_PMOS_NOSF[677]
  PIN Data_PMOS_NOSF[679]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3742.825 1046.435 3743.105 1047.435 ;
    END
  END Data_PMOS_NOSF[679]
  PIN BcidMtx[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3738.905 1046.435 3739.185 1047.435 ;
    END
  END BcidMtx[197]
  PIN FREEZE_PMOS_NOSF[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3737.225 1046.435 3737.505 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[32]
  PIN BcidMtx[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3736.105 1046.435 3736.385 1047.435 ;
    END
  END BcidMtx[194]
  PIN Data_PMOS_NOSF[675]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3694.105 1046.435 3694.385 1047.435 ;
    END
  END Data_PMOS_NOSF[675]
  PIN Data_PMOS_NOSF[687]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3692.425 1046.435 3692.705 1047.435 ;
    END
  END Data_PMOS_NOSF[687]
  PIN Data_PMOS_NOSF[676]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3691.305 1046.435 3691.585 1047.435 ;
    END
  END Data_PMOS_NOSF[676]
  PIN Data_PMOS_NOSF[672]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3689.065 1046.435 3689.345 1047.435 ;
    END
  END Data_PMOS_NOSF[672]
  PIN MASKH[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3687.385 1046.435 3687.665 1047.435 ;
    END
  END MASKH[32]
  PIN DIG_MON_PMOS_NOSF[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3685.705 1046.435 3685.985 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[64]
  PIN MASKD[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3682.345 1046.435 3682.625 1047.435 ;
    END
  END MASKD[63]
  PIN MASKV[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3671.145 1046.435 3671.425 1047.435 ;
    END
  END MASKV[63]
  PIN Data_PMOS_NOSF[659]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3670.025 1046.435 3670.305 1047.435 ;
    END
  END Data_PMOS_NOSF[659]
  PIN Data_PMOS_NOSF[665]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3666.665 1046.435 3666.945 1047.435 ;
    END
  END Data_PMOS_NOSF[665]
  PIN Data_PMOS_NOSF[657]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3665.545 1046.435 3665.825 1047.435 ;
    END
  END Data_PMOS_NOSF[657]
  PIN BcidMtx[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3659.665 1046.435 3659.945 1047.435 ;
    END
  END BcidMtx[190]
  PIN BcidMtx[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3631.945 1046.435 3632.225 1047.435 ;
    END
  END BcidMtx[188]
  PIN BcidMtx[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3630.825 1046.435 3631.105 1047.435 ;
    END
  END BcidMtx[186]
  PIN Data_PMOS_NOSF[660]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3627.465 1046.435 3627.745 1047.435 ;
    END
  END Data_PMOS_NOSF[660]
  PIN Data_PMOS_NOSF[655]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3625.785 1046.435 3626.065 1047.435 ;
    END
  END Data_PMOS_NOSF[655]
  PIN Data_PMOS_NOSF[662]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3624.665 1046.435 3624.945 1047.435 ;
    END
  END Data_PMOS_NOSF[662]
  PIN MASKV[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3622.425 1046.435 3622.705 1047.435 ;
    END
  END MASKV[62]
  PIN MASKD[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3621.305 1046.435 3621.585 1047.435 ;
    END
  END MASKD[62]
  PIN INJ_ROW[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3601.705 1046.435 3601.985 1047.435 ;
    END
  END INJ_ROW[30]
  PIN Data_PMOS_NOSF[648]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3600.585 1046.435 3600.865 1047.435 ;
    END
  END Data_PMOS_NOSF[648]
  PIN Data_PMOS_NOSF[642]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3599.465 1046.435 3599.745 1047.435 ;
    END
  END Data_PMOS_NOSF[642]
  PIN Data_PMOS_NOSF[644]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3596.665 1046.435 3596.945 1047.435 ;
    END
  END Data_PMOS_NOSF[644]
  PIN Data_PMOS_NOSF[636]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3595.545 1046.435 3595.825 1047.435 ;
    END
  END Data_PMOS_NOSF[636]
  PIN nTOK_PMOS_NOSF[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3554.105 1046.435 3554.385 1047.435 ;
    END
  END nTOK_PMOS_NOSF[30]
  PIN Read_PMOS_NOSF[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3550.745 1046.435 3551.025 1047.435 ;
    END
  END Read_PMOS_NOSF[30]
  PIN BcidMtx[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3549.625 1046.435 3549.905 1047.435 ;
    END
  END BcidMtx[181]
  PIN INJ_IN[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3547.945 1046.435 3548.225 1047.435 ;
    END
  END INJ_IN[60]
  PIN Data_PMOS_NOSF[640]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3544.585 1046.435 3544.865 1047.435 ;
    END
  END Data_PMOS_NOSF[640]
  PIN Data_PMOS_NOSF[646]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3543.465 1046.435 3543.745 1047.435 ;
    END
  END Data_PMOS_NOSF[646]
  PIN Data_PMOS_NOSF[641]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3542.905 1046.435 3543.185 1047.435 ;
    END
  END Data_PMOS_NOSF[641]
  PIN MASKH[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3531.705 1046.435 3531.985 1047.435 ;
    END
  END MASKH[30]
  PIN DIG_MON_SEL[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3527.785 1046.435 3528.065 1047.435 ;
    END
  END DIG_MON_SEL[59]
  PIN Data_PMOS_NOSF[627]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3521.345 1046.435 3521.625 1047.435 ;
    END
  END Data_PMOS_NOSF[627]
  PIN Data_PMOS_NOSF[628]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3519.665 1046.435 3519.945 1047.435 ;
    END
  END Data_PMOS_NOSF[628]
  PIN Data_PMOS_NOSF[614]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3519.105 1046.435 3519.385 1047.435 ;
    END
  END Data_PMOS_NOSF[614]
  PIN Data_PMOS_NOSF[615]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3490.825 1046.435 3491.105 1047.435 ;
    END
  END Data_PMOS_NOSF[615]
  PIN nTOK_PMOS_NOSF[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3488.585 1046.435 3488.865 1047.435 ;
    END
  END nTOK_PMOS_NOSF[29]
  PIN BcidMtx[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3487.465 1046.435 3487.745 1047.435 ;
    END
  END BcidMtx[179]
  PIN BcidMtx[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3484.665 1046.435 3484.945 1047.435 ;
    END
  END BcidMtx[176]
  PIN INJ_IN[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3482.425 1046.435 3482.705 1047.435 ;
    END
  END INJ_IN[58]
  PIN Data_PMOS_NOSF[612]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3481.305 1046.435 3481.585 1047.435 ;
    END
  END Data_PMOS_NOSF[612]
  PIN Data_PMOS_NOSF[613]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3465.625 1046.435 3465.905 1047.435 ;
    END
  END Data_PMOS_NOSF[613]
  PIN Data_PMOS_NOSF[610]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3463.945 1046.435 3464.225 1047.435 ;
    END
  END Data_PMOS_NOSF[610]
  PIN Data_PMOS_NOSF[626]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3462.825 1046.435 3463.105 1047.435 ;
    END
  END Data_PMOS_NOSF[626]
  PIN DIG_MON_SEL[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3457.785 1046.435 3458.065 1047.435 ;
    END
  END DIG_MON_SEL[57]
  PIN DIG_MON_PMOS_NOSF[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3455.545 1046.435 3455.825 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[57]
  PIN Data_PMOS_NOSF[600]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3412.425 1046.435 3412.705 1047.435 ;
    END
  END Data_PMOS_NOSF[600]
  PIN Data_PMOS_NOSF[593]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3411.305 1046.435 3411.585 1047.435 ;
    END
  END Data_PMOS_NOSF[593]
  PIN Data_PMOS_NOSF[608]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3410.185 1046.435 3410.465 1047.435 ;
    END
  END Data_PMOS_NOSF[608]
  PIN nTOK_PMOS_NOSF[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3406.265 1046.435 3406.545 1047.435 ;
    END
  END nTOK_PMOS_NOSF[28]
  PIN BcidMtx[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3405.145 1046.435 3405.425 1047.435 ;
    END
  END BcidMtx[173]
  PIN BcidMtx[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3404.025 1046.435 3404.305 1047.435 ;
    END
  END BcidMtx[171]
  PIN BcidMtx[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3401.785 1046.435 3402.065 1047.435 ;
    END
  END BcidMtx[169]
  PIN INJ_IN[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3391.705 1046.435 3391.985 1047.435 ;
    END
  END INJ_IN[56]
  PIN Data_PMOS_NOSF[590]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3390.025 1046.435 3390.305 1047.435 ;
    END
  END Data_PMOS_NOSF[590]
  PIN Data_PMOS_NOSF[604]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3387.225 1046.435 3387.505 1047.435 ;
    END
  END Data_PMOS_NOSF[604]
  PIN Data_PMOS_NOSF[589]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3386.105 1046.435 3386.385 1047.435 ;
    END
  END Data_PMOS_NOSF[589]
  PIN Data_PMOS_NOSF[605]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3384.985 1046.435 3385.265 1047.435 ;
    END
  END Data_PMOS_NOSF[605]
  PIN FREEZE_PMOS_NOSF[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3633.065 1046.435 3633.345 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[31]
  PIN MASKD[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4470.825 1046.435 4471.105 1047.435 ;
    END
  END MASKD[83]
  PIN nRST[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17765.785 1046.435 17766.065 1047.435 ;
    END
  END nRST[208]
  PIN nRST[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18325.785 1046.435 18326.065 1047.435 ;
    END
  END nRST[215]
  PIN nRST[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1591.305 1046.435 1591.585 1047.435 ;
    END
  END nRST[6]
  PIN nRST[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2151.305 1046.435 2151.585 1047.435 ;
    END
  END nRST[13]
  PIN nRST[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16085.785 1046.435 16086.065 1047.435 ;
    END
  END nRST[187]
  PIN nRST[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16645.785 1046.435 16646.065 1047.435 ;
    END
  END nRST[194]
  PIN nRST[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17205.785 1046.435 17206.065 1047.435 ;
    END
  END nRST[201]
  PIN nRST[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13845.785 1046.435 13846.065 1047.435 ;
    END
  END nRST[159]
  PIN nRST[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14405.785 1046.435 14406.065 1047.435 ;
    END
  END nRST[166]
  PIN nRST[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14965.785 1046.435 14966.065 1047.435 ;
    END
  END nRST[173]
  PIN nRST[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15525.785 1046.435 15526.065 1047.435 ;
    END
  END nRST[180]
  PIN nRST[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12165.785 1046.435 12166.065 1047.435 ;
    END
  END nRST[138]
  PIN nRST[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12725.785 1046.435 12726.065 1047.435 ;
    END
  END nRST[145]
  PIN nRST[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13285.785 1046.435 13286.065 1047.435 ;
    END
  END nRST[152]
  PIN nRST[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11605.785 1046.435 11606.065 1047.435 ;
    END
  END nRST[131]
  PIN nRST[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18885.785 1046.435 18886.065 1047.435 ;
    END
  END nRST[222]
  PIN nRST[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2711.305 1046.435 2711.585 1047.435 ;
    END
  END nRST[20]
  PIN nRST[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3271.305 1046.435 3271.585 1047.435 ;
    END
  END nRST[27]
  PIN nRST[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13351.305 1046.435 13351.585 1047.435 ;
    END
  END nRST[153]
  PIN nRST[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13911.305 1046.435 13911.585 1047.435 ;
    END
  END nRST[160]
  PIN nRST[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14471.305 1046.435 14471.585 1047.435 ;
    END
  END nRST[167]
  PIN nRST[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15031.305 1046.435 15031.585 1047.435 ;
    END
  END nRST[174]
  PIN nRST[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16151.305 1046.435 16151.585 1047.435 ;
    END
  END nRST[188]
  PIN nRST[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16711.305 1046.435 16711.585 1047.435 ;
    END
  END nRST[195]
  PIN nRST[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17271.305 1046.435 17271.585 1047.435 ;
    END
  END nRST[202]
  PIN nRST[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17831.305 1046.435 17831.585 1047.435 ;
    END
  END nRST[209]
  PIN nRST[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10551.305 1046.435 10551.585 1047.435 ;
    END
  END nRST[118]
  PIN nRST[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11111.305 1046.435 11111.585 1047.435 ;
    END
  END nRST[125]
  PIN nRST[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11671.305 1046.435 11671.585 1047.435 ;
    END
  END nRST[132]
  PIN nRST[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12231.305 1046.435 12231.585 1047.435 ;
    END
  END nRST[139]
  PIN nRST[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12791.305 1046.435 12791.585 1047.435 ;
    END
  END nRST[146]
  PIN nRST[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8311.305 1046.435 8311.585 1047.435 ;
    END
  END nRST[90]
  PIN nRST[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8871.305 1046.435 8871.585 1047.435 ;
    END
  END nRST[97]
  PIN nRST[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9431.305 1046.435 9431.585 1047.435 ;
    END
  END nRST[104]
  PIN nRST[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9991.305 1046.435 9991.585 1047.435 ;
    END
  END nRST[111]
  PIN nRST[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3831.305 1046.435 3831.585 1047.435 ;
    END
  END nRST[34]
  PIN nRST[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4391.305 1046.435 4391.585 1047.435 ;
    END
  END nRST[41]
  PIN nRST[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4951.305 1046.435 4951.585 1047.435 ;
    END
  END nRST[48]
  PIN nRST[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7191.305 1046.435 7191.585 1047.435 ;
    END
  END nRST[76]
  PIN nRST[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7751.305 1046.435 7751.585 1047.435 ;
    END
  END nRST[83]
  PIN nRST[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5511.305 1046.435 5511.585 1047.435 ;
    END
  END nRST[55]
  PIN nRST[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6071.305 1046.435 6071.585 1047.435 ;
    END
  END nRST[62]
  PIN nRST[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6631.305 1046.435 6631.585 1047.435 ;
    END
  END nRST[69]
  PIN nRST[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15591.305 1046.435 15591.585 1047.435 ;
    END
  END nRST[181]
  PIN nRST[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18391.305 1046.435 18391.585 1047.435 ;
    END
  END nRST[216]
  PIN FREEZE_PMOS_NOSF[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4111.305 1046.435 4111.585 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[37]
  PIN INJ_IN[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4107.945 1046.435 4108.225 1047.435 ;
    END
  END INJ_IN[74]
  PIN Data_PMOS_NOSF[780]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4106.825 1046.435 4107.105 1047.435 ;
    END
  END Data_PMOS_NOSF[780]
  PIN Data_PMOS_NOSF[792]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4105.145 1046.435 4105.425 1047.435 ;
    END
  END Data_PMOS_NOSF[792]
  PIN Data_PMOS_NOSF[778]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4102.345 1046.435 4102.625 1047.435 ;
    END
  END Data_PMOS_NOSF[778]
  PIN Data_PMOS_NOSF[777]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4101.785 1046.435 4102.065 1047.435 ;
    END
  END Data_PMOS_NOSF[777]
  PIN MASKH[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4091.705 1046.435 4091.985 1047.435 ;
    END
  END MASKH[37]
  PIN DIG_MON_SEL[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4087.785 1046.435 4088.065 1047.435 ;
    END
  END DIG_MON_SEL[73]
  PIN DIG_MON_PMOS_NOSF[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4085.545 1046.435 4085.825 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[73]
  PIN Data_PMOS_NOSF[774]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4081.345 1046.435 4081.625 1047.435 ;
    END
  END Data_PMOS_NOSF[774]
  PIN Data_PMOS_NOSF[761]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4079.105 1046.435 4079.385 1047.435 ;
    END
  END Data_PMOS_NOSF[761]
  PIN Data_PMOS_NOSF[776]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4052.505 1046.435 4052.785 1047.435 ;
    END
  END Data_PMOS_NOSF[776]
  PIN Data_PMOS_NOSF[762]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4050.825 1046.435 4051.105 1047.435 ;
    END
  END Data_PMOS_NOSF[762]
  PIN BcidMtx[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4046.905 1046.435 4047.185 1047.435 ;
    END
  END BcidMtx[220]
  PIN FREEZE_PMOS_NOSF[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4045.785 1046.435 4046.065 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[36]
  PIN BcidMtx[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4044.105 1046.435 4044.385 1047.435 ;
    END
  END BcidMtx[217]
  PIN Data_PMOS_NOSF[758]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4040.745 1046.435 4041.025 1047.435 ;
    END
  END Data_PMOS_NOSF[758]
  PIN Data_PMOS_NOSF[771]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4026.745 1046.435 4027.025 1047.435 ;
    END
  END Data_PMOS_NOSF[771]
  PIN Data_PMOS_NOSF[772]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4025.065 1046.435 4025.345 1047.435 ;
    END
  END Data_PMOS_NOSF[772]
  PIN Data_PMOS_NOSF[773]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4022.825 1046.435 4023.105 1047.435 ;
    END
  END Data_PMOS_NOSF[773]
  PIN MASKH[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4021.705 1046.435 4021.985 1047.435 ;
    END
  END MASKH[36]
  PIN DIG_MON_PMOS_NOSF[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4015.545 1046.435 4015.825 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[71]
  PIN MASKV[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4013.865 1046.435 4014.145 1047.435 ;
    END
  END MASKV[71]
  PIN Data_PMOS_NOSF[747]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3972.425 1046.435 3972.705 1047.435 ;
    END
  END Data_PMOS_NOSF[747]
  PIN Data_PMOS_NOSF[755]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3970.185 1046.435 3970.465 1047.435 ;
    END
  END Data_PMOS_NOSF[755]
  PIN Data_HV[1121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18879.625 1046.435 18879.905 1047.435 ;
    END
  END Data_HV[1121]
  PIN Data_PMOS_NOSF[741]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3968.505 1046.435 3968.785 1047.435 ;
    END
  END Data_PMOS_NOSF[741]
  PIN BcidMtx[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3965.145 1046.435 3965.425 1047.435 ;
    END
  END BcidMtx[215]
  PIN BcidMtx[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3964.025 1046.435 3964.305 1047.435 ;
    END
  END BcidMtx[213]
  PIN BcidMtx[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3962.345 1046.435 3962.625 1047.435 ;
    END
  END BcidMtx[212]
  PIN Data_PMOS_NOSF[738]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3950.585 1046.435 3950.865 1047.435 ;
    END
  END Data_PMOS_NOSF[738]
  PIN Data_PMOS_NOSF[744]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3949.465 1046.435 3949.745 1047.435 ;
    END
  END Data_PMOS_NOSF[744]
  PIN Data_PMOS_NOSF[739]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3947.785 1046.435 3948.065 1047.435 ;
    END
  END Data_PMOS_NOSF[739]
  PIN Data_PMOS_NOSF[735]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3945.545 1046.435 3945.825 1047.435 ;
    END
  END Data_PMOS_NOSF[735]
  PIN MASKV[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3942.465 1046.435 3942.745 1047.435 ;
    END
  END MASKV[70]
  PIN DIG_MON_PMOS_NOSF[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3940.225 1046.435 3940.505 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[70]
  PIN DIG_MON_SEL[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5031.945 1046.435 5032.225 1047.435 ;
    END
  END DIG_MON_SEL[97]
  PIN DIG_MON_PMOS_NOSF[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5029.705 1046.435 5029.985 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[97]
  PIN Data_PMOS_NOSF[1026]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5027.465 1046.435 5027.745 1047.435 ;
    END
  END Data_PMOS_NOSF[1026]
  PIN Data_PMOS_NOSF[1013]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5025.225 1046.435 5025.505 1047.435 ;
    END
  END Data_PMOS_NOSF[1013]
  PIN Data_PMOS_NOSF[1021]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5024.665 1046.435 5024.945 1047.435 ;
    END
  END Data_PMOS_NOSF[1021]
  PIN Data_PMOS_NOSF[1015]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5022.985 1046.435 5023.265 1047.435 ;
    END
  END Data_PMOS_NOSF[1015]
  PIN Data_HV[1059]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18600.185 1046.435 18600.465 1047.435 ;
    END
  END Data_HV[1059]
  PIN BcidMtx[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5005.625 1046.435 5005.905 1047.435 ;
    END
  END BcidMtx[293]
  PIN FREEZE_PMOS_NOSF[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5003.945 1046.435 5004.225 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[48]
  PIN BcidMtx[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5001.705 1046.435 5001.985 1047.435 ;
    END
  END BcidMtx[288]
  PIN Data_PMOS_NOSF[1011]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4999.465 1046.435 4999.745 1047.435 ;
    END
  END Data_PMOS_NOSF[1011]
  PIN Data_PMOS_NOSF[1023]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4997.785 1046.435 4998.065 1047.435 ;
    END
  END Data_PMOS_NOSF[1023]
  PIN Data_PMOS_NOSF[1019]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4995.545 1046.435 4995.825 1047.435 ;
    END
  END Data_PMOS_NOSF[1019]
  PIN Data_PMOS_NOSF[1008]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4994.425 1046.435 4994.705 1047.435 ;
    END
  END Data_PMOS_NOSF[1008]
  PIN MASKH[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4954.105 1046.435 4954.385 1047.435 ;
    END
  END MASKH[48]
  PIN DIG_MON_SEL[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4950.185 1046.435 4950.465 1047.435 ;
    END
  END DIG_MON_SEL[95]
  PIN MASKD[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4949.065 1046.435 4949.345 1047.435 ;
    END
  END MASKD[95]
  PIN INJ_ROW[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4946.825 1046.435 4947.105 1047.435 ;
    END
  END INJ_ROW[47]
  PIN Data_PMOS_NOSF[999]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4944.585 1046.435 4944.865 1047.435 ;
    END
  END Data_PMOS_NOSF[999]
  PIN Data_PMOS_NOSF[992]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4943.465 1046.435 4943.745 1047.435 ;
    END
  END Data_PMOS_NOSF[992]
  PIN Data_PMOS_NOSF[1001]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4941.785 1046.435 4942.065 1047.435 ;
    END
  END Data_PMOS_NOSF[1001]
  PIN nTOK_PMOS_NOSF[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4930.025 1046.435 4930.305 1047.435 ;
    END
  END nTOK_PMOS_NOSF[47]
  PIN BcidMtx[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4928.905 1046.435 4929.185 1047.435 ;
    END
  END BcidMtx[287]
  PIN FREEZE_PMOS_NOSF[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4927.225 1046.435 4927.505 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[47]
  PIN INJ_IN[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4921.905 1046.435 4922.185 1047.435 ;
    END
  END INJ_IN[94]
  PIN Data_PMOS_NOSF[990]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4920.785 1046.435 4921.065 1047.435 ;
    END
  END Data_PMOS_NOSF[990]
  PIN Data_PMOS_NOSF[1002]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4919.105 1046.435 4919.385 1047.435 ;
    END
  END Data_PMOS_NOSF[1002]
  PIN Data_PMOS_NOSF[988]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4890.825 1046.435 4891.105 1047.435 ;
    END
  END Data_PMOS_NOSF[988]
  PIN Data_PMOS_NOSF[987]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4890.265 1046.435 4890.545 1047.435 ;
    END
  END Data_PMOS_NOSF[987]
  PIN MASKH[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4888.585 1046.435 4888.865 1047.435 ;
    END
  END MASKH[47]
  PIN DIG_MON_SEL[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4884.665 1046.435 4884.945 1047.435 ;
    END
  END DIG_MON_SEL[93]
  PIN MASKD[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4883.545 1046.435 4883.825 1047.435 ;
    END
  END MASKD[93]
  PIN MASKV[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4880.745 1046.435 4881.025 1047.435 ;
    END
  END MASKV[93]
  PIN Data_PMOS_NOSF[971]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4865.065 1046.435 4865.345 1047.435 ;
    END
  END Data_PMOS_NOSF[971]
  PIN Data_PMOS_NOSF[979]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4864.505 1046.435 4864.785 1047.435 ;
    END
  END Data_PMOS_NOSF[979]
  PIN Data_PMOS_NOSF[973]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4862.825 1046.435 4863.105 1047.435 ;
    END
  END Data_PMOS_NOSF[973]
  PIN BcidMtx[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4858.345 1046.435 4858.625 1047.435 ;
    END
  END BcidMtx[280]
  PIN BcidMtx[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4857.785 1046.435 4858.065 1047.435 ;
    END
  END BcidMtx[279]
  PIN BcidMtx[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4856.105 1046.435 4856.385 1047.435 ;
    END
  END BcidMtx[278]
  PIN Data_PMOS_NOSF[968]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4813.545 1046.435 4813.825 1047.435 ;
    END
  END Data_PMOS_NOSF[968]
  PIN Data_PMOS_NOSF[975]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4812.985 1046.435 4813.265 1047.435 ;
    END
  END Data_PMOS_NOSF[975]
  PIN Data_PMOS_NOSF[970]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4811.305 1046.435 4811.585 1047.435 ;
    END
  END Data_PMOS_NOSF[970]
  PIN Data_PMOS_NOSF[983]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4808.505 1046.435 4808.785 1047.435 ;
    END
  END Data_PMOS_NOSF[983]
  PIN MASKH[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4807.385 1046.435 4807.665 1047.435 ;
    END
  END MASKH[46]
  PIN DIG_MON_PMOS_NOSF[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4805.705 1046.435 4805.985 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[92]
  PIN MASKD[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4802.345 1046.435 4802.625 1047.435 ;
    END
  END MASKD[91]
  PIN DIG_MON_PMOS_NOSF[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4801.225 1046.435 4801.505 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[91]
  PIN Data_PMOS_NOSF[963]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4790.585 1046.435 4790.865 1047.435 ;
    END
  END Data_PMOS_NOSF[963]
  PIN Data_PMOS_NOSF[958]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4787.785 1046.435 4788.065 1047.435 ;
    END
  END Data_PMOS_NOSF[958]
  PIN Data_PMOS_NOSF[965]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4787.225 1046.435 4787.505 1047.435 ;
    END
  END Data_PMOS_NOSF[965]
  PIN Data_PMOS_NOSF[951]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4785.545 1046.435 4785.825 1047.435 ;
    END
  END Data_PMOS_NOSF[951]
  PIN BcidMtx[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4779.105 1046.435 4779.385 1047.435 ;
    END
  END BcidMtx[273]
  PIN Read_PMOS_NOSF[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4752.505 1046.435 4752.785 1047.435 ;
    END
  END Read_PMOS_NOSF[45]
  PIN BcidMtx[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4750.825 1046.435 4751.105 1047.435 ;
    END
  END BcidMtx[270]
  PIN Data_PMOS_NOSF[960]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4746.905 1046.435 4747.185 1047.435 ;
    END
  END Data_PMOS_NOSF[960]
  PIN Data_PMOS_NOSF[955]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4746.345 1046.435 4746.625 1047.435 ;
    END
  END Data_PMOS_NOSF[955]
  PIN Data_PMOS_NOSF[956]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4744.665 1046.435 4744.945 1047.435 ;
    END
  END Data_PMOS_NOSF[956]
  PIN MASKH[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4741.865 1046.435 4742.145 1047.435 ;
    END
  END MASKH[45]
  PIN MASKD[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4741.305 1046.435 4741.585 1047.435 ;
    END
  END MASKD[90]
  PIN DIG_MON_SEL[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4725.625 1046.435 4725.905 1047.435 ;
    END
  END DIG_MON_SEL[90]
  PIN MASKV[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4721.145 1046.435 4721.425 1047.435 ;
    END
  END MASKV[89]
  PIN Data_PMOS_NOSF[942]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4720.585 1046.435 4720.865 1047.435 ;
    END
  END Data_PMOS_NOSF[942]
  PIN Data_PMOS_NOSF[943]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4718.905 1046.435 4719.185 1047.435 ;
    END
  END Data_PMOS_NOSF[943]
  PIN Data_PMOS_NOSF[931]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4716.105 1046.435 4716.385 1047.435 ;
    END
  END Data_PMOS_NOSF[931]
  PIN Data_PMOS_NOSF[930]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4715.545 1046.435 4715.825 1047.435 ;
    END
  END Data_PMOS_NOSF[930]
  PIN BcidMtx[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5231.865 1046.435 5232.145 1047.435 ;
    END
  END BcidMtx[309]
  PIN BcidMtx[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5229.625 1046.435 5229.905 1047.435 ;
    END
  END BcidMtx[307]
  PIN Data_PMOS_NOSF[1074]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5226.825 1046.435 5227.105 1047.435 ;
    END
  END Data_PMOS_NOSF[1074]
  PIN Data_PMOS_NOSF[1086]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5225.145 1046.435 5225.425 1047.435 ;
    END
  END Data_PMOS_NOSF[1086]
  PIN Data_PMOS_NOSF[1087]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5223.465 1046.435 5223.745 1047.435 ;
    END
  END Data_PMOS_NOSF[1087]
  PIN Data_PMOS_NOSF[1071]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5221.785 1046.435 5222.065 1047.435 ;
    END
  END Data_PMOS_NOSF[1071]
  PIN MASKH[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5211.705 1046.435 5211.985 1047.435 ;
    END
  END MASKH[51]
  PIN MASKD[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5206.665 1046.435 5206.945 1047.435 ;
    END
  END MASKD[101]
  PIN MASKV[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5201.905 1046.435 5202.185 1047.435 ;
    END
  END MASKV[101]
  PIN Data_PMOS_NOSF[1062]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5200.225 1046.435 5200.505 1047.435 ;
    END
  END Data_PMOS_NOSF[1062]
  PIN Data_PMOS_NOSF[1063]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5173.065 1046.435 5173.345 1047.435 ;
    END
  END Data_PMOS_NOSF[1063]
  PIN Data_PMOS_NOSF[1057]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5171.385 1046.435 5171.665 1047.435 ;
    END
  END Data_PMOS_NOSF[1057]
  PIN nTOK_PMOS_NOSF[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5168.585 1046.435 5168.865 1047.435 ;
    END
  END nTOK_PMOS_NOSF[50]
  PIN BcidMtx[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5166.345 1046.435 5166.625 1047.435 ;
    END
  END BcidMtx[303]
  PIN BcidMtx[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5164.665 1046.435 5164.945 1047.435 ;
    END
  END BcidMtx[302]
  PIN INJ_IN[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5162.425 1046.435 5162.705 1047.435 ;
    END
  END INJ_IN[100]
  PIN Data_PMOS_NOSF[1059]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5160.185 1046.435 5160.465 1047.435 ;
    END
  END Data_PMOS_NOSF[1059]
  PIN Data_PMOS_NOSF[1054]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5145.625 1046.435 5145.905 1047.435 ;
    END
  END Data_PMOS_NOSF[1054]
  PIN Data_PMOS_NOSF[1051]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5143.945 1046.435 5144.225 1047.435 ;
    END
  END Data_PMOS_NOSF[1051]
  PIN MASKV[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5142.265 1046.435 5142.545 1047.435 ;
    END
  END MASKV[100]
  PIN DIG_MON_PMOS_NOSF[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5140.025 1046.435 5140.305 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[100]
  PIN DIG_MON_SEL[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5137.785 1046.435 5138.065 1047.435 ;
    END
  END DIG_MON_SEL[99]
  PIN DIG_MON_SEL[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18647.785 1046.435 18648.065 1047.435 ;
    END
  END DIG_MON_SEL[437]
  PIN MASKV[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5133.865 1046.435 5134.145 1047.435 ;
    END
  END MASKV[99]
  PIN Data_PMOS_NOSF[1041]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5092.425 1046.435 5092.705 1047.435 ;
    END
  END Data_PMOS_NOSF[1041]
  PIN Data_PMOS_NOSF[1042]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5090.745 1046.435 5091.025 1047.435 ;
    END
  END Data_PMOS_NOSF[1042]
  PIN Data_PMOS_NOSF[1035]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5088.505 1046.435 5088.785 1047.435 ;
    END
  END Data_PMOS_NOSF[1035]
  PIN nTOK_PMOS_NOSF[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5086.265 1046.435 5086.545 1047.435 ;
    END
  END nTOK_PMOS_NOSF[49]
  PIN BcidMtx[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5084.025 1046.435 5084.305 1047.435 ;
    END
  END BcidMtx[297]
  PIN BcidMtx[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5081.785 1046.435 5082.065 1047.435 ;
    END
  END BcidMtx[295]
  PIN Data_PMOS_NOSF[1032]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5070.585 1046.435 5070.865 1047.435 ;
    END
  END Data_PMOS_NOSF[1032]
  PIN Data_PMOS_NOSF[1044]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5068.905 1046.435 5069.185 1047.435 ;
    END
  END Data_PMOS_NOSF[1044]
  PIN Data_PMOS_NOSF[1033]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5067.785 1046.435 5068.065 1047.435 ;
    END
  END Data_PMOS_NOSF[1033]
  PIN Data_PMOS_NOSF[1029]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5065.545 1046.435 5065.825 1047.435 ;
    END
  END Data_PMOS_NOSF[1029]
  PIN MASKH[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5061.905 1046.435 5062.185 1047.435 ;
    END
  END MASKH[49]
  PIN DIG_MON_PMOS_NOSF[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5060.225 1046.435 5060.505 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[98]
  PIN DIG_MON_SEL[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6151.945 1046.435 6152.225 1047.435 ;
    END
  END DIG_MON_SEL[125]
  PIN INJ_ROW[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6148.585 1046.435 6148.865 1047.435 ;
    END
  END INJ_ROW[62]
  PIN Data_PMOS[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6147.465 1046.435 6147.745 1047.435 ;
    END
  END Data_PMOS[144]
  PIN Data_PMOS[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6145.225 1046.435 6145.505 1047.435 ;
    END
  END Data_PMOS[131]
  PIN Data_PMOS[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6143.545 1046.435 6143.825 1047.435 ;
    END
  END Data_PMOS[140]
  PIN Data_PMOS[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6142.425 1046.435 6142.705 1047.435 ;
    END
  END Data_PMOS[132]
  PIN BcidMtx[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6125.065 1046.435 6125.345 1047.435 ;
    END
  END BcidMtx[376]
  PIN Read_PMOS[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6123.385 1046.435 6123.665 1047.435 ;
    END
  END Read_PMOS[6]
  PIN BcidMtx[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6122.265 1046.435 6122.545 1047.435 ;
    END
  END BcidMtx[373]
  PIN Data_PMOS[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6118.905 1046.435 6119.185 1047.435 ;
    END
  END Data_PMOS[128]
  PIN Data_PMOS[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6117.225 1046.435 6117.505 1047.435 ;
    END
  END Data_PMOS[136]
  PIN Data_PMOS[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6116.105 1046.435 6116.385 1047.435 ;
    END
  END Data_PMOS[142]
  PIN Data_PMOS[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6114.985 1046.435 6115.265 1047.435 ;
    END
  END Data_PMOS[127]
  PIN MASKD[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6073.545 1046.435 6073.825 1047.435 ;
    END
  END MASKD[124]
  PIN DIG_MON_SEL[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6070.745 1046.435 6071.025 1047.435 ;
    END
  END DIG_MON_SEL[124]
  PIN DIG_MON_PMOS[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6067.945 1046.435 6068.225 1047.435 ;
    END
  END DIG_MON_PMOS[11]
  PIN Data_PMOS[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6065.145 1046.435 6065.425 1047.435 ;
    END
  END Data_PMOS[113]
  PIN Data_PMOS[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6064.025 1046.435 6064.305 1047.435 ;
    END
  END Data_PMOS[124]
  PIN Data_PMOS[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6062.345 1046.435 6062.625 1047.435 ;
    END
  END Data_PMOS[125]
  PIN INJ_IN[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6051.145 1046.435 6051.425 1047.435 ;
    END
  END INJ_IN[123]
  PIN BcidMtx[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6048.905 1046.435 6049.185 1047.435 ;
    END
  END BcidMtx[371]
  PIN FREEZE_PMOS[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6047.225 1046.435 6047.505 1047.435 ;
    END
  END FREEZE_PMOS[5]
  PIN BcidMtx[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6044.985 1046.435 6045.265 1047.435 ;
    END
  END BcidMtx[366]
  PIN Data_PMOS[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6040.785 1046.435 6041.065 1047.435 ;
    END
  END Data_PMOS[108]
  PIN Data_PMOS[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6039.105 1046.435 6039.385 1047.435 ;
    END
  END Data_PMOS[120]
  PIN Data_PMOS[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6011.385 1046.435 6011.665 1047.435 ;
    END
  END Data_PMOS[116]
  PIN Data_PMOS[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6010.265 1046.435 6010.545 1047.435 ;
    END
  END Data_PMOS[105]
  PIN MASKH[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6008.585 1046.435 6008.865 1047.435 ;
    END
  END MASKH[61]
  PIN DIG_MON_SEL[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6005.225 1046.435 6005.505 1047.435 ;
    END
  END DIG_MON_SEL[122]
  PIN MASKD[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6003.545 1046.435 6003.825 1047.435 ;
    END
  END MASKD[121]
  PIN BcidMtx[1331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18858.905 1046.435 18859.185 1047.435 ;
    END
  END BcidMtx[1331]
  PIN Data_PMOS[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5986.185 1046.435 5986.465 1047.435 ;
    END
  END Data_PMOS[96]
  PIN Data_PMOS[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5985.065 1046.435 5985.345 1047.435 ;
    END
  END Data_PMOS[89]
  PIN Data_PMOS[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5983.385 1046.435 5983.665 1047.435 ;
    END
  END Data_PMOS[98]
  PIN nTOK_PMOS[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5980.025 1046.435 5980.305 1047.435 ;
    END
  END nTOK_PMOS[4]
  PIN BcidMtx[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5978.345 1046.435 5978.625 1047.435 ;
    END
  END BcidMtx[364]
  PIN Read_PMOS[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5976.665 1046.435 5976.945 1047.435 ;
    END
  END Read_PMOS[4]
  PIN INJ_IN[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5973.865 1046.435 5974.145 1047.435 ;
    END
  END INJ_IN[120]
  PIN Data_PMOS[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5933.545 1046.435 5933.825 1047.435 ;
    END
  END Data_PMOS[86]
  PIN Data_PMOS[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5931.865 1046.435 5932.145 1047.435 ;
    END
  END Data_PMOS[94]
  PIN Data_PMOS[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5929.625 1046.435 5929.905 1047.435 ;
    END
  END Data_PMOS[85]
  PIN Data_PMOS[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5928.505 1046.435 5928.785 1047.435 ;
    END
  END Data_PMOS[101]
  PIN MASKD[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5926.825 1046.435 5927.105 1047.435 ;
    END
  END MASKD[120]
  PIN DIG_MON_SEL[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5923.465 1046.435 5923.745 1047.435 ;
    END
  END DIG_MON_SEL[119]
  PIN DIG_MON_PMOS[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5921.225 1046.435 5921.505 1047.435 ;
    END
  END DIG_MON_PMOS[7]
  PIN Data_PMOS[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5910.585 1046.435 5910.865 1047.435 ;
    END
  END Data_PMOS[81]
  PIN Data_PMOS[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5908.345 1046.435 5908.625 1047.435 ;
    END
  END Data_PMOS[68]
  PIN Data_PMOS[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5907.225 1046.435 5907.505 1047.435 ;
    END
  END Data_PMOS[83]
  PIN Data_PMOS[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5905.545 1046.435 5905.825 1047.435 ;
    END
  END Data_PMOS[69]
  PIN BcidMtx[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5899.665 1046.435 5899.945 1047.435 ;
    END
  END BcidMtx[358]
  PIN Read_PMOS[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5872.505 1046.435 5872.785 1047.435 ;
    END
  END Read_PMOS[3]
  PIN BcidMtx[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5870.825 1046.435 5871.105 1047.435 ;
    END
  END BcidMtx[354]
  PIN Data_PMOS[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5867.465 1046.435 5867.745 1047.435 ;
    END
  END Data_PMOS[72]
  PIN Data_PMOS[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5865.785 1046.435 5866.065 1047.435 ;
    END
  END Data_PMOS[67]
  PIN Data_PMOS[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5864.665 1046.435 5864.945 1047.435 ;
    END
  END Data_PMOS[74]
  PIN Data_PMOS[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5862.985 1046.435 5863.265 1047.435 ;
    END
  END Data_PMOS[80]
  PIN DIG_MON_PMOS[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5860.185 1046.435 5860.465 1047.435 ;
    END
  END DIG_MON_PMOS[6]
  PIN DIG_MON_SEL[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5845.065 1046.435 5845.345 1047.435 ;
    END
  END DIG_MON_SEL[117]
  PIN INJ_ROW[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5841.705 1046.435 5841.985 1047.435 ;
    END
  END INJ_ROW[58]
  PIN Data_PMOS[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5840.025 1046.435 5840.305 1047.435 ;
    END
  END Data_PMOS[50]
  PIN Data_PMOS[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5838.345 1046.435 5838.625 1047.435 ;
    END
  END Data_PMOS[47]
  PIN Data_PMOS[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5836.665 1046.435 5836.945 1047.435 ;
    END
  END Data_PMOS[56]
  PIN INJ_IN[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5834.425 1046.435 5834.705 1047.435 ;
    END
  END INJ_IN[117]
  PIN BcidMtx[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5792.425 1046.435 5792.705 1047.435 ;
    END
  END BcidMtx[352]
  PIN BcidMtx[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3549.065 1046.435 3549.345 1047.435 ;
    END
  END BcidMtx[180]
  PIN Data_PMOS_NOSF[633]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3546.825 1046.435 3547.105 1047.435 ;
    END
  END Data_PMOS_NOSF[633]
  PIN Data_PMOS_NOSF[639]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3545.705 1046.435 3545.985 1047.435 ;
    END
  END Data_PMOS_NOSF[639]
  PIN Data_PMOS_NOSF[631]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3542.345 1046.435 3542.625 1047.435 ;
    END
  END Data_PMOS_NOSF[631]
  PIN Data_PMOS_NOSF[647]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3541.225 1046.435 3541.505 1047.435 ;
    END
  END Data_PMOS_NOSF[647]
  PIN MASKD[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3531.145 1046.435 3531.425 1047.435 ;
    END
  END MASKD[60]
  PIN MASKD[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3526.665 1046.435 3526.945 1047.435 ;
    END
  END MASKD[59]
  PIN INJ_ROW[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3522.465 1046.435 3522.745 1047.435 ;
    END
  END INJ_ROW[29]
  PIN Data_PMOS_NOSF[617]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3520.785 1046.435 3521.065 1047.435 ;
    END
  END Data_PMOS_NOSF[617]
  PIN Data_PMOS_NOSF[622]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3493.065 1046.435 3493.345 1047.435 ;
    END
  END Data_PMOS_NOSF[622]
  PIN Data_PMOS_NOSF[623]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3491.945 1046.435 3492.225 1047.435 ;
    END
  END Data_PMOS_NOSF[623]
  PIN INJ_IN[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3489.705 1046.435 3489.985 1047.435 ;
    END
  END INJ_IN[59]
  PIN BcidMtx[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3486.905 1046.435 3487.185 1047.435 ;
    END
  END BcidMtx[178]
  PIN FREEZE_PMOS_NOSF[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3485.785 1046.435 3486.065 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[29]
  PIN BcidMtx[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3484.105 1046.435 3484.385 1047.435 ;
    END
  END BcidMtx[175]
  PIN Data_PMOS_NOSF[611]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3480.745 1046.435 3481.025 1047.435 ;
    END
  END Data_PMOS_NOSF[611]
  PIN Data_PMOS_NOSF[624]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3466.745 1046.435 3467.025 1047.435 ;
    END
  END Data_PMOS_NOSF[624]
  PIN Data_PMOS_NOSF[625]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3465.065 1046.435 3465.345 1047.435 ;
    END
  END Data_PMOS_NOSF[625]
  PIN Data_PMOS_NOSF[609]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3463.385 1046.435 3463.665 1047.435 ;
    END
  END Data_PMOS_NOSF[609]
  PIN MASKV[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3462.265 1046.435 3462.545 1047.435 ;
    END
  END MASKV[58]
  PIN MASKD[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3461.145 1046.435 3461.425 1047.435 ;
    END
  END MASKD[58]
  PIN MASKD[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3456.665 1046.435 3456.945 1047.435 ;
    END
  END MASKD[57]
  PIN INJ_ROW[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3454.425 1046.435 3454.705 1047.435 ;
    END
  END INJ_ROW[28]
  PIN Data_PMOS_NOSF[606]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3413.545 1046.435 3413.825 1047.435 ;
    END
  END Data_PMOS_NOSF[606]
  PIN Data_PMOS_NOSF[601]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3410.745 1046.435 3411.025 1047.435 ;
    END
  END Data_PMOS_NOSF[601]
  PIN Data_PMOS_NOSF[602]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3409.625 1046.435 3409.905 1047.435 ;
    END
  END Data_PMOS_NOSF[602]
  PIN Data_PMOS_NOSF[594]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3408.505 1046.435 3408.785 1047.435 ;
    END
  END Data_PMOS_NOSF[594]
  PIN BcidMtx[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3404.585 1046.435 3404.865 1047.435 ;
    END
  END BcidMtx[172]
  PIN INJ_ROW[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18881.305 1046.435 18881.585 1047.435 ;
    END
  END INJ_ROW[221]
  PIN Read_PMOS_NOSF[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3402.905 1046.435 3403.185 1047.435 ;
    END
  END Read_PMOS_NOSF[28]
  PIN Data_PMOS_NOSF[591]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3390.585 1046.435 3390.865 1047.435 ;
    END
  END Data_PMOS_NOSF[591]
  PIN Data_PMOS_NOSF[597]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3389.465 1046.435 3389.745 1047.435 ;
    END
  END Data_PMOS_NOSF[597]
  PIN Data_PMOS_NOSF[598]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3388.345 1046.435 3388.625 1047.435 ;
    END
  END Data_PMOS_NOSF[598]
  PIN Data_PMOS_NOSF[588]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3385.545 1046.435 3385.825 1047.435 ;
    END
  END Data_PMOS_NOSF[588]
  PIN MASKV[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3382.465 1046.435 3382.745 1047.435 ;
    END
  END MASKV[56]
  PIN MASKD[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3381.345 1046.435 3381.625 1047.435 ;
    END
  END MASKD[56]
  PIN DIG_MON_SEL[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4471.945 1046.435 4472.225 1047.435 ;
    END
  END DIG_MON_SEL[83]
  PIN DIG_MON_PMOS_NOSF[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4469.705 1046.435 4469.985 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[83]
  PIN MASKV[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4468.025 1046.435 4468.305 1047.435 ;
    END
  END MASKV[83]
  PIN Data_PMOS_NOSF[866]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4465.225 1046.435 4465.505 1047.435 ;
    END
  END Data_PMOS_NOSF[866]
  PIN Data_PMOS_NOSF[881]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4464.105 1046.435 4464.385 1047.435 ;
    END
  END Data_PMOS_NOSF[881]
  PIN Data_PMOS_NOSF[868]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4462.985 1046.435 4463.265 1047.435 ;
    END
  END Data_PMOS_NOSF[868]
  PIN BcidMtx[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4445.065 1046.435 4445.345 1047.435 ;
    END
  END BcidMtx[250]
  PIN FREEZE_PMOS_NOSF[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4443.945 1046.435 4444.225 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[41]
  PIN Read_PMOS_NOSF[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4443.385 1046.435 4443.665 1047.435 ;
    END
  END Read_PMOS_NOSF[41]
  PIN Data_PMOS_NOSF[864]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4439.465 1046.435 4439.745 1047.435 ;
    END
  END Data_PMOS_NOSF[864]
  PIN Data_PMOS_NOSF[870]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4438.345 1046.435 4438.625 1047.435 ;
    END
  END Data_PMOS_NOSF[870]
  PIN Data_PMOS_NOSF[871]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4437.225 1046.435 4437.505 1047.435 ;
    END
  END Data_PMOS_NOSF[871]
  PIN Data_PMOS_NOSF[861]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4434.425 1046.435 4434.705 1047.435 ;
    END
  END Data_PMOS_NOSF[861]
  PIN MASKV[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4394.665 1046.435 4394.945 1047.435 ;
    END
  END MASKV[82]
  PIN MASKD[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4393.545 1046.435 4393.825 1047.435 ;
    END
  END MASKD[82]
  PIN MASKD[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4389.065 1046.435 4389.345 1047.435 ;
    END
  END MASKD[81]
  PIN INJ_ROW[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4386.825 1046.435 4387.105 1047.435 ;
    END
  END INJ_ROW[40]
  PIN Data_PMOS_NOSF[858]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4385.705 1046.435 4385.985 1047.435 ;
    END
  END Data_PMOS_NOSF[858]
  PIN Data_PMOS_NOSF[853]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4382.905 1046.435 4383.185 1047.435 ;
    END
  END Data_PMOS_NOSF[853]
  PIN Data_PMOS_NOSF[854]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4381.785 1046.435 4382.065 1047.435 ;
    END
  END Data_PMOS_NOSF[854]
  PIN Data_PMOS_NOSF[846]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4372.265 1046.435 4372.545 1047.435 ;
    END
  END Data_PMOS_NOSF[846]
  PIN BcidMtx[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4367.785 1046.435 4368.065 1047.435 ;
    END
  END BcidMtx[243]
  PIN Read_PMOS_NOSF[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4366.665 1046.435 4366.945 1047.435 ;
    END
  END Read_PMOS_NOSF[40]
  PIN BcidMtx[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4365.545 1046.435 4365.825 1047.435 ;
    END
  END BcidMtx[241]
  PIN Data_PMOS_NOSF[849]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4359.665 1046.435 4359.945 1047.435 ;
    END
  END Data_PMOS_NOSF[849]
  PIN Data_PMOS_NOSF[850]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4358.545 1046.435 4358.825 1047.435 ;
    END
  END Data_PMOS_NOSF[850]
  PIN Data_PMOS_NOSF[856]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4331.945 1046.435 4332.225 1047.435 ;
    END
  END Data_PMOS_NOSF[856]
  PIN MASKV[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4329.145 1046.435 4329.425 1047.435 ;
    END
  END MASKV[80]
  PIN MASKD[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4328.025 1046.435 4328.305 1047.435 ;
    END
  END MASKD[80]
  PIN MASKD[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4323.545 1046.435 4323.825 1047.435 ;
    END
  END MASKD[79]
  PIN MASKV[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4320.745 1046.435 4321.025 1047.435 ;
    END
  END MASKV[79]
  PIN Data_PMOS_NOSF[831]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4306.185 1046.435 4306.465 1047.435 ;
    END
  END Data_PMOS_NOSF[831]
  PIN Data_PMOS_NOSF[832]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4304.505 1046.435 4304.785 1047.435 ;
    END
  END Data_PMOS_NOSF[832]
  PIN Data_PMOS_NOSF[826]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4302.825 1046.435 4303.105 1047.435 ;
    END
  END Data_PMOS_NOSF[826]
  PIN INJ_IN[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4301.145 1046.435 4301.425 1047.435 ;
    END
  END INJ_IN[79]
  PIN BcidMtx[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4298.905 1046.435 4299.185 1047.435 ;
    END
  END BcidMtx[239]
  PIN Data_HV[1131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18880.185 1046.435 18880.465 1047.435 ;
    END
  END Data_HV[1131]
  PIN BcidMtx[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4295.545 1046.435 4295.825 1047.435 ;
    END
  END BcidMtx[235]
  PIN INJ_IN[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4293.865 1046.435 4294.145 1047.435 ;
    END
  END INJ_IN[78]
  PIN Data_PMOS_NOSF[829]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4251.865 1046.435 4252.145 1047.435 ;
    END
  END Data_PMOS_NOSF[829]
  PIN Data_PMOS_NOSF[835]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4250.745 1046.435 4251.025 1047.435 ;
    END
  END Data_PMOS_NOSF[835]
  PIN Data_PMOS_NOSF[820]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4249.625 1046.435 4249.905 1047.435 ;
    END
  END Data_PMOS_NOSF[820]
  PIN MASKD[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4246.825 1046.435 4247.105 1047.435 ;
    END
  END MASKD[78]
  PIN DIG_MON_SEL[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4243.465 1046.435 4243.745 1047.435 ;
    END
  END DIG_MON_SEL[77]
  PIN MASKV[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4231.145 1046.435 4231.425 1047.435 ;
    END
  END MASKV[77]
  PIN Data_PMOS_NOSF[806]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4230.025 1046.435 4230.305 1047.435 ;
    END
  END Data_PMOS_NOSF[806]
  PIN Data_PMOS_NOSF[803]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4228.345 1046.435 4228.625 1047.435 ;
    END
  END Data_PMOS_NOSF[803]
  PIN Data_PMOS_NOSF[805]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4226.105 1046.435 4226.385 1047.435 ;
    END
  END Data_PMOS_NOSF[805]
  PIN INJ_IN[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4222.465 1046.435 4222.745 1047.435 ;
    END
  END INJ_IN[77]
  PIN BcidMtx[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4219.665 1046.435 4219.945 1047.435 ;
    END
  END BcidMtx[232]
  PIN BcidMtx[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4191.385 1046.435 4191.665 1047.435 ;
    END
  END BcidMtx[229]
  PIN INJ_IN[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4189.705 1046.435 4189.985 1047.435 ;
    END
  END INJ_IN[76]
  PIN Data_PMOS_NOSF[807]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4187.465 1046.435 4187.745 1047.435 ;
    END
  END Data_PMOS_NOSF[807]
  PIN Data_PMOS_NOSF[814]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4185.225 1046.435 4185.505 1047.435 ;
    END
  END Data_PMOS_NOSF[814]
  PIN Data_PMOS_NOSF[799]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4184.105 1046.435 4184.385 1047.435 ;
    END
  END Data_PMOS_NOSF[799]
  PIN MASKV[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4182.425 1046.435 4182.705 1047.435 ;
    END
  END MASKV[76]
  PIN DIG_MON_SEL[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4165.625 1046.435 4165.905 1047.435 ;
    END
  END DIG_MON_SEL[76]
  PIN DIG_MON_PMOS_NOSF[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4162.825 1046.435 4163.105 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[75]
  PIN Data_PMOS_NOSF[789]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4159.465 1046.435 4159.745 1047.435 ;
    END
  END Data_PMOS_NOSF[789]
  PIN Data_PMOS_NOSF[796]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4158.905 1046.435 4159.185 1047.435 ;
    END
  END Data_PMOS_NOSF[796]
  PIN Data_PMOS_NOSF[797]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4157.225 1046.435 4157.505 1047.435 ;
    END
  END Data_PMOS_NOSF[797]
  PIN nTOK_PMOS_NOSF[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4114.105 1046.435 4114.385 1047.435 ;
    END
  END nTOK_PMOS_NOSF[37]
  PIN BcidMtx[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4112.985 1046.435 4113.265 1047.435 ;
    END
  END BcidMtx[227]
  PIN INJ_IN[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2427.945 1046.435 2428.225 1047.435 ;
    END
  END INJ_IN[32]
  PIN Data_PMOS_NOSF[338]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2426.265 1046.435 2426.545 1047.435 ;
    END
  END Data_PMOS_NOSF[338]
  PIN Data_PMOS_NOSF[346]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2424.585 1046.435 2424.865 1047.435 ;
    END
  END Data_PMOS_NOSF[346]
  PIN Data_PMOS_NOSF[352]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2423.465 1046.435 2423.745 1047.435 ;
    END
  END Data_PMOS_NOSF[352]
  PIN Data_PMOS_NOSF[336]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2421.785 1046.435 2422.065 1047.435 ;
    END
  END Data_PMOS_NOSF[336]
  PIN MASKD[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2411.145 1046.435 2411.425 1047.435 ;
    END
  END MASKD[32]
  PIN DIG_MON_SEL[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2407.785 1046.435 2408.065 1047.435 ;
    END
  END DIG_MON_SEL[31]
  PIN INJ_ROW[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2402.465 1046.435 2402.745 1047.435 ;
    END
  END INJ_ROW[15]
  PIN Data_PMOS_NOSF[327]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2400.225 1046.435 2400.505 1047.435 ;
    END
  END Data_PMOS_NOSF[327]
  PIN Data_PMOS_NOSF[320]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2399.105 1046.435 2399.385 1047.435 ;
    END
  END Data_PMOS_NOSF[320]
  PIN Data_PMOS_NOSF[322]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2371.385 1046.435 2371.665 1047.435 ;
    END
  END Data_PMOS_NOSF[322]
  PIN INJ_IN[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2369.705 1046.435 2369.985 1047.435 ;
    END
  END INJ_IN[31]
  PIN BcidMtx[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2367.465 1046.435 2367.745 1047.435 ;
    END
  END BcidMtx[95]
  PIN Read_PMOS_NOSF[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2365.225 1046.435 2365.505 1047.435 ;
    END
  END Read_PMOS_NOSF[15]
  PIN BcidMtx[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2363.545 1046.435 2363.825 1047.435 ;
    END
  END BcidMtx[90]
  PIN Data_PMOS_NOSF[317]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2360.745 1046.435 2361.025 1047.435 ;
    END
  END Data_PMOS_NOSF[317]
  PIN Data_PMOS_NOSF[330]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2346.745 1046.435 2347.025 1047.435 ;
    END
  END Data_PMOS_NOSF[330]
  PIN Data_PMOS_NOSF[331]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2345.065 1046.435 2345.345 1047.435 ;
    END
  END Data_PMOS_NOSF[331]
  PIN Data_PMOS_NOSF[315]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2343.385 1046.435 2343.665 1047.435 ;
    END
  END Data_PMOS_NOSF[315]
  PIN MASKH[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2341.705 1046.435 2341.985 1047.435 ;
    END
  END MASKH[15]
  PIN DIG_MON_SEL[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2337.785 1046.435 2338.065 1047.435 ;
    END
  END DIG_MON_SEL[29]
  PIN Data_PMOS_NOSF[312]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2293.545 1046.435 2293.825 1047.435 ;
    END
  END Data_PMOS_NOSF[312]
  PIN Data_PMOS_NOSF[313]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2291.865 1046.435 2292.145 1047.435 ;
    END
  END Data_PMOS_NOSF[313]
  PIN Data_PMOS_NOSF[307]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2290.745 1046.435 2291.025 1047.435 ;
    END
  END Data_PMOS_NOSF[307]
  PIN Data_PMOS_NOSF[300]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2288.505 1046.435 2288.785 1047.435 ;
    END
  END Data_PMOS_NOSF[300]
  PIN BcidMtx[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2285.145 1046.435 2285.425 1047.435 ;
    END
  END BcidMtx[89]
  PIN Read_PMOS_NOSF[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2282.905 1046.435 2283.185 1047.435 ;
    END
  END Read_PMOS_NOSF[14]
  PIN BcidMtx[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2281.785 1046.435 2282.065 1047.435 ;
    END
  END BcidMtx[85]
  PIN Data_PMOS_NOSF[297]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2270.585 1046.435 2270.865 1047.435 ;
    END
  END Data_PMOS_NOSF[297]
  PIN Data_PMOS_NOSF[303]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2269.465 1046.435 2269.745 1047.435 ;
    END
  END Data_PMOS_NOSF[303]
  PIN Data_PMOS_NOSF[298]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2267.785 1046.435 2268.065 1047.435 ;
    END
  END Data_PMOS_NOSF[298]
  PIN Data_PMOS_NOSF[295]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2266.105 1046.435 2266.385 1047.435 ;
    END
  END Data_PMOS_NOSF[295]
  PIN Data_PMOS_NOSF[311]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2264.985 1046.435 2265.265 1047.435 ;
    END
  END Data_PMOS_NOSF[311]
  PIN DIG_MON_PMOS_NOSF[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2260.225 1046.435 2260.505 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[28]
  PIN FREEZE_PMOS_NOSF[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2513.065 1046.435 2513.345 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[17]
  PIN INJ_ROW[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3348.585 1046.435 3348.865 1047.435 ;
    END
  END INJ_ROW[27]
  PIN Data_PMOS_NOSF[575]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3346.905 1046.435 3347.185 1047.435 ;
    END
  END Data_PMOS_NOSF[575]
  PIN Data_PMOS_NOSF[586]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3345.785 1046.435 3346.065 1047.435 ;
    END
  END Data_PMOS_NOSF[586]
  PIN Data_PMOS_NOSF[587]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3344.105 1046.435 3344.385 1047.435 ;
    END
  END Data_PMOS_NOSF[587]
  PIN INJ_IN[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3341.305 1046.435 3341.585 1047.435 ;
    END
  END INJ_IN[55]
  PIN BcidMtx[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3325.065 1046.435 3325.345 1047.435 ;
    END
  END BcidMtx[166]
  PIN FREEZE_PMOS_NOSF[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3323.945 1046.435 3324.225 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[27]
  PIN BcidMtx[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3321.705 1046.435 3321.985 1047.435 ;
    END
  END BcidMtx[162]
  PIN MASKV[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18652.265 1046.435 18652.545 1047.435 ;
    END
  END MASKV[438]
  PIN Data_PMOS_NOSF[576]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3318.345 1046.435 3318.625 1047.435 ;
    END
  END Data_PMOS_NOSF[576]
  PIN Data_PMOS_NOSF[583]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3316.105 1046.435 3316.385 1047.435 ;
    END
  END Data_PMOS_NOSF[583]
  PIN Data_PMOS_NOSF[568]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3314.985 1046.435 3315.265 1047.435 ;
    END
  END Data_PMOS_NOSF[568]
  PIN Data_PMOS_NOSF[584]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3313.865 1046.435 3314.145 1047.435 ;
    END
  END Data_PMOS_NOSF[584]
  PIN DIG_MON_PMOS_NOSF[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3272.425 1046.435 3272.705 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[54]
  PIN DIG_MON_SEL[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3270.185 1046.435 3270.465 1047.435 ;
    END
  END DIG_MON_SEL[53]
  PIN DIG_MON_PMOS_NOSF[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3267.945 1046.435 3268.225 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[53]
  PIN Data_PMOS_NOSF[554]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3265.145 1046.435 3265.425 1047.435 ;
    END
  END Data_PMOS_NOSF[554]
  PIN Data_PMOS_NOSF[551]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3263.465 1046.435 3263.745 1047.435 ;
    END
  END Data_PMOS_NOSF[551]
  PIN Data_PMOS_NOSF[566]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3262.345 1046.435 3262.625 1047.435 ;
    END
  END Data_PMOS_NOSF[566]
  PIN INJ_IN[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3251.145 1046.435 3251.425 1047.435 ;
    END
  END INJ_IN[53]
  PIN BcidMtx[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3248.345 1046.435 3248.625 1047.435 ;
    END
  END BcidMtx[160]
  PIN FREEZE_PMOS_NOSF[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3247.225 1046.435 3247.505 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[26]
  PIN BcidMtx[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3245.545 1046.435 3245.825 1047.435 ;
    END
  END BcidMtx[157]
  PIN Data_PMOS_NOSF[549]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3240.785 1046.435 3241.065 1047.435 ;
    END
  END Data_PMOS_NOSF[549]
  PIN Data_PMOS_NOSF[556]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3238.545 1046.435 3238.825 1047.435 ;
    END
  END Data_PMOS_NOSF[556]
  PIN Data_PMOS_NOSF[557]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3211.385 1046.435 3211.665 1047.435 ;
    END
  END Data_PMOS_NOSF[557]
  PIN Data_PMOS_NOSF[563]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3209.705 1046.435 3209.985 1047.435 ;
    END
  END Data_PMOS_NOSF[563]
  PIN MASKH[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3208.585 1046.435 3208.865 1047.435 ;
    END
  END MASKH[26]
  PIN DIG_MON_SEL[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3205.225 1046.435 3205.505 1047.435 ;
    END
  END DIG_MON_SEL[52]
  PIN DIG_MON_PMOS_NOSF[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3202.425 1046.435 3202.705 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[51]
  PIN Data_PMOS_NOSF[543]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3200.185 1046.435 3200.465 1047.435 ;
    END
  END Data_PMOS_NOSF[543]
  PIN Data_PMOS_NOSF[544]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3185.625 1046.435 3185.905 1047.435 ;
    END
  END Data_PMOS_NOSF[544]
  PIN Data_PMOS_NOSF[545]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3183.945 1046.435 3184.225 1047.435 ;
    END
  END Data_PMOS_NOSF[545]
  PIN Data_PMOS_NOSF[531]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3182.265 1046.435 3182.545 1047.435 ;
    END
  END Data_PMOS_NOSF[531]
  PIN BcidMtx[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3178.905 1046.435 3179.185 1047.435 ;
    END
  END BcidMtx[155]
  PIN FREEZE_PMOS_NOSF[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3177.225 1046.435 3177.505 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[25]
  PIN BcidMtx[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3175.545 1046.435 3175.825 1047.435 ;
    END
  END BcidMtx[151]
  PIN Data_PMOS_NOSF[528]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3134.105 1046.435 3134.385 1047.435 ;
    END
  END Data_PMOS_NOSF[528]
  PIN Data_PMOS_NOSF[540]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3132.425 1046.435 3132.705 1047.435 ;
    END
  END Data_PMOS_NOSF[540]
  PIN Data_PMOS_NOSF[541]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3130.745 1046.435 3131.025 1047.435 ;
    END
  END Data_PMOS_NOSF[541]
  PIN Data_PMOS_NOSF[526]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3129.625 1046.435 3129.905 1047.435 ;
    END
  END Data_PMOS_NOSF[526]
  PIN MASKV[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3127.945 1046.435 3128.225 1047.435 ;
    END
  END MASKV[50]
  PIN DIG_MON_PMOS_NOSF[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3125.705 1046.435 3125.985 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[50]
  PIN DIG_MON_SEL[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3123.465 1046.435 3123.745 1047.435 ;
    END
  END DIG_MON_SEL[49]
  PIN INJ_ROW[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3111.705 1046.435 3111.985 1047.435 ;
    END
  END INJ_ROW[24]
  PIN Data_PMOS_NOSF[512]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3110.025 1046.435 3110.305 1047.435 ;
    END
  END Data_PMOS_NOSF[512]
  PIN Data_PMOS_NOSF[509]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3108.345 1046.435 3108.625 1047.435 ;
    END
  END Data_PMOS_NOSF[509]
  PIN Data_PMOS_NOSF[518]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3106.665 1046.435 3106.945 1047.435 ;
    END
  END Data_PMOS_NOSF[518]
  PIN INJ_IN[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3102.465 1046.435 3102.745 1047.435 ;
    END
  END INJ_IN[49]
  PIN BcidMtx[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3099.665 1046.435 3099.945 1047.435 ;
    END
  END BcidMtx[148]
  PIN BcidMtx[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3071.945 1046.435 3072.225 1047.435 ;
    END
  END BcidMtx[146]
  PIN INJ_IN[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3069.705 1046.435 3069.985 1047.435 ;
    END
  END INJ_IN[48]
  PIN Data_PMOS_NOSF[513]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3067.465 1046.435 3067.745 1047.435 ;
    END
  END Data_PMOS_NOSF[513]
  PIN Data_PMOS_NOSF[508]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3065.785 1046.435 3066.065 1047.435 ;
    END
  END Data_PMOS_NOSF[508]
  PIN Data_PMOS_NOSF[505]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3064.105 1046.435 3064.385 1047.435 ;
    END
  END Data_PMOS_NOSF[505]
  PIN MASKV[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3062.425 1046.435 3062.705 1047.435 ;
    END
  END MASKV[48]
  PIN DIG_MON_PMOS_NOSF[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3060.185 1046.435 3060.465 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[48]
  PIN DIG_MON_SEL[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3045.065 1046.435 3045.345 1047.435 ;
    END
  END DIG_MON_SEL[47]
  PIN INJ_ROW[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3041.705 1046.435 3041.985 1047.435 ;
    END
  END INJ_ROW[23]
  PIN Data_PMOS_NOSF[491]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3040.025 1046.435 3040.305 1047.435 ;
    END
  END Data_PMOS_NOSF[491]
  PIN Data_PMOS_NOSF[488]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3038.345 1046.435 3038.625 1047.435 ;
    END
  END Data_PMOS_NOSF[488]
  PIN Data_PMOS_NOSF[497]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3036.665 1046.435 3036.945 1047.435 ;
    END
  END Data_PMOS_NOSF[497]
  PIN INJ_IN[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3034.425 1046.435 3034.705 1047.435 ;
    END
  END INJ_IN[47]
  PIN BcidMtx[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2992.425 1046.435 2992.705 1047.435 ;
    END
  END BcidMtx[142]
  PIN Read_PMOS_NOSF[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2990.745 1046.435 2991.025 1047.435 ;
    END
  END Read_PMOS_NOSF[23]
  PIN BcidMtx[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2989.065 1046.435 2989.345 1047.435 ;
    END
  END BcidMtx[138]
  PIN Data_PMOS_NOSF[485]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2986.265 1046.435 2986.545 1047.435 ;
    END
  END Data_PMOS_NOSF[485]
  PIN Data_PMOS_NOSF[493]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2984.585 1046.435 2984.865 1047.435 ;
    END
  END Data_PMOS_NOSF[493]
  PIN Data_PMOS_NOSF[494]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2982.905 1046.435 2983.185 1047.435 ;
    END
  END Data_PMOS_NOSF[494]
  PIN Data_PMOS_NOSF[500]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2981.225 1046.435 2981.505 1047.435 ;
    END
  END Data_PMOS_NOSF[500]
  PIN DIG_MON_PMOS_NOSF[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2970.025 1046.435 2970.305 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[46]
  PIN DIG_MON_SEL[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2968.345 1046.435 2968.625 1047.435 ;
    END
  END DIG_MON_SEL[46]
  PIN DIG_MON_PMOS_NOSF[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2965.545 1046.435 2965.825 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[45]
  PIN Data_PMOS_NOSF[470]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2960.785 1046.435 2961.065 1047.435 ;
    END
  END Data_PMOS_NOSF[470]
  PIN Data_PMOS_NOSF[481]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2959.665 1046.435 2959.945 1047.435 ;
    END
  END Data_PMOS_NOSF[481]
  PIN Data_PMOS_NOSF[482]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2932.505 1046.435 2932.785 1047.435 ;
    END
  END Data_PMOS_NOSF[482]
  PIN INJ_IN[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2929.705 1046.435 2929.985 1047.435 ;
    END
  END INJ_IN[45]
  PIN BcidMtx[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2927.465 1046.435 2927.745 1047.435 ;
    END
  END BcidMtx[137]
  PIN FREEZE_PMOS_NOSF[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2925.785 1046.435 2926.065 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[22]
  PIN BcidMtx[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2924.665 1046.435 2924.945 1047.435 ;
    END
  END BcidMtx[134]
  PIN BcidMtx[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2923.545 1046.435 2923.825 1047.435 ;
    END
  END BcidMtx[132]
  PIN Data_PMOS_NOSF[464]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2920.745 1046.435 2921.025 1047.435 ;
    END
  END Data_PMOS_NOSF[464]
  PIN Data_PMOS_NOSF[466]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2905.625 1046.435 2905.905 1047.435 ;
    END
  END Data_PMOS_NOSF[466]
  PIN Data_PMOS_NOSF[473]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2904.505 1046.435 2904.785 1047.435 ;
    END
  END Data_PMOS_NOSF[473]
  PIN Data_PMOS_NOSF[479]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2902.825 1046.435 2903.105 1047.435 ;
    END
  END Data_PMOS_NOSF[479]
  PIN MASKD[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2901.145 1046.435 2901.425 1047.435 ;
    END
  END MASKD[44]
  PIN DIG_MON_SEL[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2898.345 1046.435 2898.625 1047.435 ;
    END
  END DIG_MON_SEL[44]
  PIN DIG_MON_PMOS_NOSF[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2895.545 1046.435 2895.825 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[43]
  PIN Data_PMOS_NOSF[449]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2852.985 1046.435 2853.265 1047.435 ;
    END
  END Data_PMOS_NOSF[449]
  PIN Data_PMOS_NOSF[460]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2851.865 1046.435 2852.145 1047.435 ;
    END
  END Data_PMOS_NOSF[460]
  PIN Data_PMOS_NOSF[461]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2850.185 1046.435 2850.465 1047.435 ;
    END
  END Data_PMOS_NOSF[461]
  PIN Data_PMOS_NOSF[447]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2848.505 1046.435 2848.785 1047.435 ;
    END
  END Data_PMOS_NOSF[447]
  PIN BcidMtx[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2845.145 1046.435 2845.425 1047.435 ;
    END
  END BcidMtx[131]
  PIN FREEZE_PMOS_NOSF[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2843.465 1046.435 2843.745 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[21]
  PIN MASKH[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18651.705 1046.435 18651.985 1047.435 ;
    END
  END MASKH[219]
  PIN INJ_IN[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2831.705 1046.435 2831.985 1047.435 ;
    END
  END INJ_IN[42]
  PIN Data_PMOS_NOSF[450]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2829.465 1046.435 2829.745 1047.435 ;
    END
  END Data_PMOS_NOSF[450]
  PIN Data_PMOS_NOSF[445]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2827.785 1046.435 2828.065 1047.435 ;
    END
  END Data_PMOS_NOSF[445]
  PIN Data_PMOS_NOSF[442]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2826.105 1046.435 2826.385 1047.435 ;
    END
  END Data_PMOS_NOSF[442]
  PIN MASKV[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2822.465 1046.435 2822.745 1047.435 ;
    END
  END MASKV[42]
  PIN FREEZE_PMOS_NOSF[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3073.065 1046.435 3073.345 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[24]
  PIN DIG_MON_PMOS_NOSF[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3909.705 1046.435 3909.985 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[69]
  PIN Data_PMOS_NOSF[722]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3906.905 1046.435 3907.185 1047.435 ;
    END
  END Data_PMOS_NOSF[722]
  PIN Data_PMOS_NOSF[733]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3905.785 1046.435 3906.065 1047.435 ;
    END
  END Data_PMOS_NOSF[733]
  PIN Data_PMOS_NOSF[734]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3904.105 1046.435 3904.385 1047.435 ;
    END
  END Data_PMOS_NOSF[734]
  PIN INJ_IN[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3901.305 1046.435 3901.585 1047.435 ;
    END
  END INJ_IN[69]
  PIN BcidMtx[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3885.625 1046.435 3885.905 1047.435 ;
    END
  END BcidMtx[209]
  PIN FREEZE_PMOS_NOSF[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3883.945 1046.435 3884.225 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[34]
  PIN BcidMtx[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3882.265 1046.435 3882.545 1047.435 ;
    END
  END BcidMtx[205]
  PIN INJ_IN[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3880.585 1046.435 3880.865 1047.435 ;
    END
  END INJ_IN[68]
  PIN Data_PMOS_NOSF[723]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3878.345 1046.435 3878.625 1047.435 ;
    END
  END Data_PMOS_NOSF[723]
  PIN Data_PMOS_NOSF[730]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3876.105 1046.435 3876.385 1047.435 ;
    END
  END Data_PMOS_NOSF[730]
  PIN Data_PMOS_NOSF[715]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3874.985 1046.435 3875.265 1047.435 ;
    END
  END Data_PMOS_NOSF[715]
  PIN MASKV[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3834.665 1046.435 3834.945 1047.435 ;
    END
  END MASKV[68]
  PIN MASKD[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3829.065 1046.435 3829.345 1047.435 ;
    END
  END MASKD[67]
  PIN INJ_ROW[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3826.825 1046.435 3827.105 1047.435 ;
    END
  END INJ_ROW[33]
  PIN Data_PMOS_NOSF[701]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3825.145 1046.435 3825.425 1047.435 ;
    END
  END Data_PMOS_NOSF[701]
  PIN Data_PMOS_NOSF[698]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3823.465 1046.435 3823.745 1047.435 ;
    END
  END Data_PMOS_NOSF[698]
  PIN Data_PMOS_NOSF[707]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3821.785 1046.435 3822.065 1047.435 ;
    END
  END Data_PMOS_NOSF[707]
  PIN INJ_IN[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3811.145 1046.435 3811.425 1047.435 ;
    END
  END INJ_IN[67]
  PIN BcidMtx[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3808.345 1046.435 3808.625 1047.435 ;
    END
  END BcidMtx[202]
  PIN Read_PMOS_NOSF[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3806.665 1046.435 3806.945 1047.435 ;
    END
  END Read_PMOS_NOSF[33]
  PIN BcidMtx[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3804.985 1046.435 3805.265 1047.435 ;
    END
  END BcidMtx[198]
  PIN INJ_IN[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3801.905 1046.435 3802.185 1047.435 ;
    END
  END INJ_IN[66]
  PIN Data_PMOS_NOSF[702]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3799.665 1046.435 3799.945 1047.435 ;
    END
  END Data_PMOS_NOSF[702]
  PIN Data_PMOS_NOSF[697]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3772.505 1046.435 3772.785 1047.435 ;
    END
  END Data_PMOS_NOSF[697]
  PIN Data_PMOS_NOSF[694]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3770.825 1046.435 3771.105 1047.435 ;
    END
  END Data_PMOS_NOSF[694]
  PIN MASKV[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3769.145 1046.435 3769.425 1047.435 ;
    END
  END MASKV[66]
  PIN DIG_MON_PMOS_NOSF[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3766.905 1046.435 3767.185 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[66]
  PIN DIG_MON_SEL[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3764.665 1046.435 3764.945 1047.435 ;
    END
  END DIG_MON_SEL[65]
  PIN INJ_ROW[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3761.305 1046.435 3761.585 1047.435 ;
    END
  END INJ_ROW[32]
  PIN Data_PMOS_NOSF[684]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3746.185 1046.435 3746.465 1047.435 ;
    END
  END Data_PMOS_NOSF[684]
  PIN Data_PMOS_NOSF[685]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3744.505 1046.435 3744.785 1047.435 ;
    END
  END Data_PMOS_NOSF[685]
  PIN Data_PMOS_NOSF[686]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3743.385 1046.435 3743.665 1047.435 ;
    END
  END Data_PMOS_NOSF[686]
  PIN INJ_IN[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3741.145 1046.435 3741.425 1047.435 ;
    END
  END INJ_IN[65]
  PIN BcidMtx[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3738.345 1046.435 3738.625 1047.435 ;
    END
  END BcidMtx[196]
  PIN Read_PMOS_NOSF[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3736.665 1046.435 3736.945 1047.435 ;
    END
  END Read_PMOS_NOSF[32]
  PIN BcidMtx[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3734.985 1046.435 3735.265 1047.435 ;
    END
  END BcidMtx[192]
  PIN Data_PMOS_NOSF[674]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3693.545 1046.435 3693.825 1047.435 ;
    END
  END Data_PMOS_NOSF[674]
  PIN Data_PMOS_NOSF[682]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3691.865 1046.435 3692.145 1047.435 ;
    END
  END Data_PMOS_NOSF[682]
  PIN Data_PMOS_NOSF[683]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3690.185 1046.435 3690.465 1047.435 ;
    END
  END Data_PMOS_NOSF[683]
  PIN Data_PMOS_NOSF[689]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3688.505 1046.435 3688.785 1047.435 ;
    END
  END Data_PMOS_NOSF[689]
  PIN MASKD[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3686.825 1046.435 3687.105 1047.435 ;
    END
  END MASKD[64]
  PIN DIG_MON_SEL[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3684.025 1046.435 3684.305 1047.435 ;
    END
  END DIG_MON_SEL[64]
  PIN DIG_MON_PMOS_NOSF[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3681.225 1046.435 3681.505 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[63]
  PIN Data_PMOS_NOSF[669]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3670.585 1046.435 3670.865 1047.435 ;
    END
  END Data_PMOS_NOSF[669]
  PIN Data_PMOS_NOSF[670]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3668.905 1046.435 3669.185 1047.435 ;
    END
  END Data_PMOS_NOSF[670]
  PIN Data_PMOS_NOSF[664]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3667.785 1046.435 3668.065 1047.435 ;
    END
  END Data_PMOS_NOSF[664]
  PIN Data_PMOS_NOSF[658]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3666.105 1046.435 3666.385 1047.435 ;
    END
  END Data_PMOS_NOSF[658]
  PIN nTOK_PMOS_NOSF[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3661.345 1046.435 3661.625 1047.435 ;
    END
  END nTOK_PMOS_NOSF[31]
  PIN BcidMtx[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3659.105 1046.435 3659.385 1047.435 ;
    END
  END BcidMtx[189]
  PIN BcidMtx[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3631.385 1046.435 3631.665 1047.435 ;
    END
  END BcidMtx[187]
  PIN Data_PMOS_NOSF[654]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3628.585 1046.435 3628.865 1047.435 ;
    END
  END Data_PMOS_NOSF[654]
  PIN Data_PMOS_NOSF[666]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3626.905 1046.435 3627.185 1047.435 ;
    END
  END Data_PMOS_NOSF[666]
  PIN Data_PMOS_NOSF[667]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3625.225 1046.435 3625.505 1047.435 ;
    END
  END Data_PMOS_NOSF[667]
  PIN Data_PMOS_NOSF[651]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3623.545 1046.435 3623.825 1047.435 ;
    END
  END Data_PMOS_NOSF[651]
  PIN DIG_MON_PMOS_NOSF[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3620.185 1046.435 3620.465 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[62]
  PIN DIG_MON_SEL[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3605.625 1046.435 3605.905 1047.435 ;
    END
  END DIG_MON_SEL[62]
  PIN MASKD[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3603.945 1046.435 3604.225 1047.435 ;
    END
  END MASKD[61]
  PIN Data_PMOS_NOSF[638]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3600.025 1046.435 3600.305 1047.435 ;
    END
  END Data_PMOS_NOSF[638]
  PIN Data_PMOS_NOSF[649]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3598.905 1046.435 3599.185 1047.435 ;
    END
  END Data_PMOS_NOSF[649]
  PIN Data_PMOS_NOSF[643]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3597.785 1046.435 3598.065 1047.435 ;
    END
  END Data_PMOS_NOSF[643]
  PIN INJ_IN[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3594.425 1046.435 3594.705 1047.435 ;
    END
  END INJ_IN[61]
  PIN BcidMtx[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3552.985 1046.435 3553.265 1047.435 ;
    END
  END BcidMtx[185]
  PIN BcidMtx[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3551.865 1046.435 3552.145 1047.435 ;
    END
  END BcidMtx[183]
  PIN nRST[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18951.305 1046.435 18951.585 1047.435 ;
    END
  END nRST[223]
  PIN Data_HV[1037]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18532.985 1046.435 18533.265 1047.435 ;
    END
  END Data_HV[1037]
  PIN Data_HV[1041]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18532.425 1046.435 18532.705 1047.435 ;
    END
  END Data_HV[1041]
  PIN Data_HV[1048]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18531.865 1046.435 18532.145 1047.435 ;
    END
  END Data_HV[1048]
  PIN Data_HV[1034]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18531.305 1046.435 18531.585 1047.435 ;
    END
  END Data_HV[1034]
  PIN Data_HV[1042]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18530.745 1046.435 18531.025 1047.435 ;
    END
  END Data_HV[1042]
  PIN Data_HV[1049]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18530.185 1046.435 18530.465 1047.435 ;
    END
  END Data_HV[1049]
  PIN Data_HV[1137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18920.785 1046.435 18921.065 1047.435 ;
    END
  END Data_HV[1137]
  PIN Data_HV[1136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18920.225 1046.435 18920.505 1047.435 ;
    END
  END Data_HV[1136]
  PIN INJ_IN[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18527.385 1046.435 18527.665 1047.435 ;
    END
  END INJ_IN[435]
  PIN MASKD[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1670.825 1046.435 1671.105 1047.435 ;
    END
  END MASKD[13]
  PIN INJ_ROW[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1668.585 1046.435 1668.865 1047.435 ;
    END
  END INJ_ROW[6]
  PIN Data_PMOS_NOSF[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1666.905 1046.435 1667.185 1047.435 ;
    END
  END Data_PMOS_NOSF[134]
  PIN Data_PMOS_NOSF[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1664.665 1046.435 1664.945 1047.435 ;
    END
  END Data_PMOS_NOSF[139]
  PIN Data_PMOS_NOSF[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1663.545 1046.435 1663.825 1047.435 ;
    END
  END Data_PMOS_NOSF[140]
  PIN INJ_IN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1661.305 1046.435 1661.585 1047.435 ;
    END
  END INJ_IN[13]
  PIN BcidMtx[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1644.505 1046.435 1644.785 1047.435 ;
    END
  END BcidMtx[39]
  PIN Read_PMOS_NOSF[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1643.385 1046.435 1643.665 1047.435 ;
    END
  END Read_PMOS_NOSF[6]
  PIN BcidMtx[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1641.705 1046.435 1641.985 1047.435 ;
    END
  END BcidMtx[36]
  PIN Data_PMOS_NOSF[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1638.345 1046.435 1638.625 1047.435 ;
    END
  END Data_PMOS_NOSF[135]
  PIN Data_PMOS_NOSF[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1637.225 1046.435 1637.505 1047.435 ;
    END
  END Data_PMOS_NOSF[136]
  PIN Data_PMOS_NOSF[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1635.545 1046.435 1635.825 1047.435 ;
    END
  END Data_PMOS_NOSF[137]
  PIN MASKV[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1594.665 1046.435 1594.945 1047.435 ;
    END
  END MASKV[12]
  PIN MASKD[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1593.545 1046.435 1593.825 1047.435 ;
    END
  END MASKD[12]
  PIN DIG_MON_PMOS_NOSF[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1587.945 1046.435 1588.225 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[11]
  PIN MASKV[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1586.265 1046.435 1586.545 1047.435 ;
    END
  END MASKV[11]
  PIN Data_PMOS_NOSF[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1584.585 1046.435 1584.865 1047.435 ;
    END
  END Data_PMOS_NOSF[117]
  PIN Data_PMOS_NOSF[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1582.345 1046.435 1582.625 1047.435 ;
    END
  END Data_PMOS_NOSF[125]
  PIN Data_PMOS_NOSF[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1581.225 1046.435 1581.505 1047.435 ;
    END
  END Data_PMOS_NOSF[112]
  PIN nTOK_PMOS_NOSF[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1570.025 1046.435 1570.305 1047.435 ;
    END
  END nTOK_PMOS_NOSF[5]
  PIN FREEZE_PMOS_NOSF[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1567.225 1046.435 1567.505 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[5]
  PIN BcidMtx[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1566.105 1046.435 1566.385 1047.435 ;
    END
  END BcidMtx[32]
  PIN INJ_IN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1561.905 1046.435 1562.185 1047.435 ;
    END
  END INJ_IN[10]
  PIN Data_PMOS_NOSF[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1559.105 1046.435 1559.385 1047.435 ;
    END
  END Data_PMOS_NOSF[120]
  PIN Data_PMOS_NOSF[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1532.505 1046.435 1532.785 1047.435 ;
    END
  END Data_PMOS_NOSF[109]
  PIN Data_PMOS_NOSF[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1530.825 1046.435 1531.105 1047.435 ;
    END
  END Data_PMOS_NOSF[106]
  PIN MASKH[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1528.585 1046.435 1528.865 1047.435 ;
    END
  END MASKH[5]
  PIN DIG_MON_PMOS_NOSF[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1526.905 1046.435 1527.185 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[10]
  PIN DIG_MON_SEL[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1525.225 1046.435 1525.505 1047.435 ;
    END
  END DIG_MON_SEL[10]
  PIN INJ_ROW[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1521.305 1046.435 1521.585 1047.435 ;
    END
  END INJ_ROW[4]
  PIN Data_PMOS_NOSF[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1520.185 1046.435 1520.465 1047.435 ;
    END
  END Data_PMOS_NOSF[102]
  PIN Data_PMOS_NOSF[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1505.625 1046.435 1505.905 1047.435 ;
    END
  END Data_PMOS_NOSF[103]
  PIN Data_PMOS_NOSF[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1503.385 1046.435 1503.665 1047.435 ;
    END
  END Data_PMOS_NOSF[98]
  PIN Data_PMOS_NOSF[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1502.265 1046.435 1502.545 1047.435 ;
    END
  END Data_PMOS_NOSF[90]
  PIN BcidMtx[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1498.905 1046.435 1499.185 1047.435 ;
    END
  END BcidMtx[29]
  PIN Read_PMOS_NOSF[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1496.665 1046.435 1496.945 1047.435 ;
    END
  END Read_PMOS_NOSF[4]
  PIN BcidMtx[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1495.545 1046.435 1495.825 1047.435 ;
    END
  END BcidMtx[25]
  PIN Data_PMOS_NOSF[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1454.105 1046.435 1454.385 1047.435 ;
    END
  END Data_PMOS_NOSF[87]
  PIN Data_PMOS_NOSF[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1451.865 1046.435 1452.145 1047.435 ;
    END
  END Data_PMOS_NOSF[94]
  PIN Data_PMOS_NOSF[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1450.745 1046.435 1451.025 1047.435 ;
    END
  END Data_PMOS_NOSF[100]
  PIN Data_PMOS_NOSF[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1448.505 1046.435 1448.785 1047.435 ;
    END
  END Data_PMOS_NOSF[101]
  PIN MASKD[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1446.825 1046.435 1447.105 1047.435 ;
    END
  END MASKD[8]
  PIN DIG_MON_PMOS_NOSF[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1445.705 1046.435 1445.985 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[8]
  PIN DIG_MON_SEL[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1443.465 1046.435 1443.745 1047.435 ;
    END
  END DIG_MON_SEL[7]
  PIN MASKV[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1431.145 1046.435 1431.425 1047.435 ;
    END
  END MASKV[7]
  PIN Data_PMOS_NOSF[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1430.025 1046.435 1430.305 1047.435 ;
    END
  END Data_PMOS_NOSF[71]
  PIN Data_PMOS_NOSF[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1428.345 1046.435 1428.625 1047.435 ;
    END
  END Data_PMOS_NOSF[68]
  PIN Data_PMOS_NOSF[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1426.105 1046.435 1426.385 1047.435 ;
    END
  END Data_PMOS_NOSF[70]
  PIN INJ_IN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1422.465 1046.435 1422.745 1047.435 ;
    END
  END INJ_IN[7]
  PIN BcidMtx[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1420.225 1046.435 1420.505 1047.435 ;
    END
  END BcidMtx[23]
  PIN BcidMtx[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1391.945 1046.435 1392.225 1047.435 ;
    END
  END BcidMtx[20]
  PIN BcidMtx[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1390.825 1046.435 1391.105 1047.435 ;
    END
  END BcidMtx[18]
  PIN Data_PMOS_NOSF[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1388.025 1046.435 1388.305 1047.435 ;
    END
  END Data_PMOS_NOSF[65]
  PIN Data_PMOS_NOSF[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1386.345 1046.435 1386.625 1047.435 ;
    END
  END Data_PMOS_NOSF[73]
  PIN Data_PMOS_NOSF[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1384.665 1046.435 1384.945 1047.435 ;
    END
  END Data_PMOS_NOSF[74]
  PIN Data_PMOS_NOSF[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1382.985 1046.435 1383.265 1047.435 ;
    END
  END Data_PMOS_NOSF[80]
  PIN MASKD[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1381.305 1046.435 1381.585 1047.435 ;
    END
  END MASKD[6]
  PIN MASKD[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1363.945 1046.435 1364.225 1047.435 ;
    END
  END MASKD[5]
  PIN MASKV[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1361.145 1046.435 1361.425 1047.435 ;
    END
  END MASKV[5]
  PIN Data_PMOS_NOSF[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1359.465 1046.435 1359.745 1047.435 ;
    END
  END Data_PMOS_NOSF[54]
  PIN Data_PMOS_NOSF[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1357.785 1046.435 1358.065 1047.435 ;
    END
  END Data_PMOS_NOSF[55]
  PIN Data_PMOS_NOSF[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1356.105 1046.435 1356.385 1047.435 ;
    END
  END Data_PMOS_NOSF[49]
  PIN nTOK_PMOS_NOSF[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1314.105 1046.435 1314.385 1047.435 ;
    END
  END nTOK_PMOS_NOSF[2]
  PIN BcidMtx[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1311.865 1046.435 1312.145 1047.435 ;
    END
  END BcidMtx[15]
  PIN Read_PMOS_NOSF[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1310.745 1046.435 1311.025 1047.435 ;
    END
  END Read_PMOS_NOSF[2]
  PIN INJ_IN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1307.945 1046.435 1308.225 1047.435 ;
    END
  END INJ_IN[4]
  PIN Read_PMOS_NOSF[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1870.745 1046.435 1871.025 1047.435 ;
    END
  END Read_PMOS_NOSF[9]
  PIN Data_PMOS_NOSF[192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1866.825 1046.435 1867.105 1047.435 ;
    END
  END Data_PMOS_NOSF[192]
  PIN Data_PMOS_NOSF[204]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1865.145 1046.435 1865.425 1047.435 ;
    END
  END Data_PMOS_NOSF[204]
  PIN Data_PMOS_NOSF[199]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1864.585 1046.435 1864.865 1047.435 ;
    END
  END Data_PMOS_NOSF[199]
  PIN Data_PMOS_NOSF[200]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1862.905 1046.435 1863.185 1047.435 ;
    END
  END Data_PMOS_NOSF[200]
  PIN MASKV[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1852.265 1046.435 1852.545 1047.435 ;
    END
  END MASKV[18]
  PIN MASKD[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1851.145 1046.435 1851.425 1047.435 ;
    END
  END MASKD[18]
  PIN DIG_MON_SEL[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1848.345 1046.435 1848.625 1047.435 ;
    END
  END DIG_MON_SEL[18]
  PIN MASKV[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1841.905 1046.435 1842.185 1047.435 ;
    END
  END MASKV[17]
  PIN Data_PMOS_NOSF[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1841.345 1046.435 1841.625 1047.435 ;
    END
  END Data_PMOS_NOSF[186]
  PIN Data_PMOS_NOSF[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1839.665 1046.435 1839.945 1047.435 ;
    END
  END Data_PMOS_NOSF[187]
  PIN Data_PMOS_NOSF[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1812.505 1046.435 1812.785 1047.435 ;
    END
  END Data_PMOS_NOSF[188]
  PIN Data_PMOS_NOSF[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1810.825 1046.435 1811.105 1047.435 ;
    END
  END Data_PMOS_NOSF[174]
  PIN BcidMtx[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1807.465 1046.435 1807.745 1047.435 ;
    END
  END BcidMtx[53]
  PIN FREEZE_PMOS_NOSF[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1805.785 1046.435 1806.065 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[8]
  PIN BcidMtx[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1804.665 1046.435 1804.945 1047.435 ;
    END
  END BcidMtx[50]
  PIN BcidMtx[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1803.545 1046.435 1803.825 1047.435 ;
    END
  END BcidMtx[48]
  PIN Data_PMOS_NOSF[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1800.185 1046.435 1800.465 1047.435 ;
    END
  END Data_PMOS_NOSF[177]
  PIN Data_PMOS_NOSF[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1785.065 1046.435 1785.345 1047.435 ;
    END
  END Data_PMOS_NOSF[184]
  PIN Data_PMOS_NOSF[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1783.945 1046.435 1784.225 1047.435 ;
    END
  END Data_PMOS_NOSF[169]
  PIN MASKV[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1782.265 1046.435 1782.545 1047.435 ;
    END
  END MASKV[16]
  PIN DIG_MON_PMOS_NOSF[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1780.025 1046.435 1780.305 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[16]
  PIN MASKV[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1773.865 1046.435 1774.145 1047.435 ;
    END
  END MASKV[15]
  PIN Data_PMOS_NOSF[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1732.425 1046.435 1732.705 1047.435 ;
    END
  END Data_PMOS_NOSF[159]
  PIN Data_PMOS_NOSF[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1731.865 1046.435 1732.145 1047.435 ;
    END
  END Data_PMOS_NOSF[166]
  PIN Data_PMOS_NOSF[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1729.065 1046.435 1729.345 1047.435 ;
    END
  END Data_PMOS_NOSF[154]
  PIN nTOK_PMOS_NOSF[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1726.265 1046.435 1726.545 1047.435 ;
    END
  END nTOK_PMOS_NOSF[7]
  PIN BcidMtx[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1724.025 1046.435 1724.305 1047.435 ;
    END
  END BcidMtx[45]
  PIN BcidMtx[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1722.345 1046.435 1722.625 1047.435 ;
    END
  END BcidMtx[44]
  PIN INJ_IN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1711.705 1046.435 1711.985 1047.435 ;
    END
  END INJ_IN[14]
  PIN Data_PMOS_NOSF[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1709.465 1046.435 1709.745 1047.435 ;
    END
  END Data_PMOS_NOSF[156]
  PIN Data_PMOS_NOSF[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1707.785 1046.435 1708.065 1047.435 ;
    END
  END Data_PMOS_NOSF[151]
  PIN Data_PMOS_NOSF[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1705.545 1046.435 1705.825 1047.435 ;
    END
  END Data_PMOS_NOSF[147]
  PIN Data_PMOS_NOSF[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1706.105 1046.435 1706.385 1047.435 ;
    END
  END Data_PMOS_NOSF[148]
  PIN MASKD[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1701.345 1046.435 1701.625 1047.435 ;
    END
  END MASKD[14]
  PIN DIG_MON_SEL[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1698.545 1046.435 1698.825 1047.435 ;
    END
  END DIG_MON_SEL[14]
  PIN MASKD[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2790.825 1046.435 2791.105 1047.435 ;
    END
  END MASKD[41]
  PIN MASKV[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2788.025 1046.435 2788.305 1047.435 ;
    END
  END MASKV[41]
  PIN Data_PMOS_NOSF[432]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2786.345 1046.435 2786.625 1047.435 ;
    END
  END Data_PMOS_NOSF[432]
  PIN Data_PMOS_NOSF[433]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2784.665 1046.435 2784.945 1047.435 ;
    END
  END Data_PMOS_NOSF[433]
  PIN Data_PMOS_NOSF[427]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2782.985 1046.435 2783.265 1047.435 ;
    END
  END Data_PMOS_NOSF[427]
  PIN nTOK_PMOS_NOSF[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2780.185 1046.435 2780.465 1047.435 ;
    END
  END nTOK_PMOS_NOSF[20]
  PIN BcidMtx[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2764.505 1046.435 2764.785 1047.435 ;
    END
  END BcidMtx[123]
  PIN BcidMtx[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2762.825 1046.435 2763.105 1047.435 ;
    END
  END BcidMtx[122]
  PIN INJ_IN[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2760.585 1046.435 2760.865 1047.435 ;
    END
  END INJ_IN[40]
  PIN Data_PMOS_NOSF[423]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2759.465 1046.435 2759.745 1047.435 ;
    END
  END Data_PMOS_NOSF[423]
  PIN Data_PMOS_NOSF[424]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2756.665 1046.435 2756.945 1047.435 ;
    END
  END Data_PMOS_NOSF[424]
  PIN Data_PMOS_NOSF[431]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2755.545 1046.435 2755.825 1047.435 ;
    END
  END Data_PMOS_NOSF[431]
  PIN Data_PMOS_NOSF[421]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2754.985 1046.435 2755.265 1047.435 ;
    END
  END Data_PMOS_NOSF[421]
  PIN MASKD[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2713.545 1046.435 2713.825 1047.435 ;
    END
  END MASKD[40]
  PIN DIG_MON_SEL[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2710.745 1046.435 2711.025 1047.435 ;
    END
  END DIG_MON_SEL[40]
  PIN DIG_MON_PMOS_NOSF[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2707.945 1046.435 2708.225 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[39]
  PIN Data_PMOS_NOSF[417]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2705.705 1046.435 2705.985 1047.435 ;
    END
  END Data_PMOS_NOSF[417]
  PIN Data_PMOS_NOSF[404]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2703.465 1046.435 2703.745 1047.435 ;
    END
  END Data_PMOS_NOSF[404]
  PIN Data_PMOS_NOSF[412]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2702.905 1046.435 2703.185 1047.435 ;
    END
  END Data_PMOS_NOSF[412]
  PIN Data_PMOS_NOSF[405]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2692.265 1046.435 2692.545 1047.435 ;
    END
  END Data_PMOS_NOSF[405]
  PIN BcidMtx[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2688.905 1046.435 2689.185 1047.435 ;
    END
  END BcidMtx[119]
  PIN FREEZE_PMOS_NOSF[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2687.225 1046.435 2687.505 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[19]
  PIN BcidMtx[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2685.545 1046.435 2685.825 1047.435 ;
    END
  END BcidMtx[115]
  PIN Data_PMOS_NOSF[402]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2680.785 1046.435 2681.065 1047.435 ;
    END
  END Data_PMOS_NOSF[402]
  PIN Data_PMOS_NOSF[408]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2679.665 1046.435 2679.945 1047.435 ;
    END
  END Data_PMOS_NOSF[408]
  PIN Data_PMOS_NOSF[403]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2652.505 1046.435 2652.785 1047.435 ;
    END
  END Data_PMOS_NOSF[403]
  PIN Data_PMOS_NOSF[400]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2650.825 1046.435 2651.105 1047.435 ;
    END
  END Data_PMOS_NOSF[400]
  PIN Data_PMOS_NOSF[416]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2649.705 1046.435 2649.985 1047.435 ;
    END
  END Data_PMOS_NOSF[416]
  PIN MASKD[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2648.025 1046.435 2648.305 1047.435 ;
    END
  END MASKD[38]
  PIN DIG_MON_SEL[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2645.225 1046.435 2645.505 1047.435 ;
    END
  END DIG_MON_SEL[38]
  PIN DIG_MON_SEL[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2644.665 1046.435 2644.945 1047.435 ;
    END
  END DIG_MON_SEL[37]
  PIN Data_PMOS_NOSF[396]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2640.185 1046.435 2640.465 1047.435 ;
    END
  END Data_PMOS_NOSF[396]
  PIN Data_PMOS_NOSF[397]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2625.625 1046.435 2625.905 1047.435 ;
    END
  END Data_PMOS_NOSF[397]
  PIN Data_PMOS_NOSF[391]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2624.505 1046.435 2624.785 1047.435 ;
    END
  END Data_PMOS_NOSF[391]
  PIN INJ_IN[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2621.145 1046.435 2621.425 1047.435 ;
    END
  END INJ_IN[37]
  PIN BcidMtx[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2618.905 1046.435 2619.185 1047.435 ;
    END
  END BcidMtx[113]
  PIN BcidMtx[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2617.785 1046.435 2618.065 1047.435 ;
    END
  END BcidMtx[111]
  PIN BcidMtx[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2614.985 1046.435 2615.265 1047.435 ;
    END
  END BcidMtx[108]
  PIN Data_PMOS_NOSF[380]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2573.545 1046.435 2573.825 1047.435 ;
    END
  END Data_PMOS_NOSF[380]
  PIN Data_PMOS_NOSF[388]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2571.865 1046.435 2572.145 1047.435 ;
    END
  END Data_PMOS_NOSF[388]
  PIN Data_PMOS_NOSF[389]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2570.185 1046.435 2570.465 1047.435 ;
    END
  END Data_PMOS_NOSF[389]
  PIN Data_PMOS_NOSF[395]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2568.505 1046.435 2568.785 1047.435 ;
    END
  END Data_PMOS_NOSF[395]
  PIN MASKD[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2566.825 1046.435 2567.105 1047.435 ;
    END
  END MASKD[36]
  PIN DIG_MON_SEL[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2564.025 1046.435 2564.305 1047.435 ;
    END
  END DIG_MON_SEL[36]
  PIN DIG_MON_PMOS_NOSF[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2561.225 1046.435 2561.505 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[35]
  PIN MASKV[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2551.145 1046.435 2551.425 1047.435 ;
    END
  END MASKV[35]
  PIN Data_PMOS_NOSF[376]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2548.905 1046.435 2549.185 1047.435 ;
    END
  END Data_PMOS_NOSF[376]
  PIN Data_PMOS_NOSF[377]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2547.225 1046.435 2547.505 1047.435 ;
    END
  END Data_PMOS_NOSF[377]
  PIN INJ_IN[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2542.465 1046.435 2542.745 1047.435 ;
    END
  END INJ_IN[35]
  PIN BcidMtx[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2539.665 1046.435 2539.945 1047.435 ;
    END
  END BcidMtx[106]
  PIN Read_PMOS_NOSF[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2512.505 1046.435 2512.785 1047.435 ;
    END
  END Read_PMOS_NOSF[17]
  PIN INJ_IN[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2509.705 1046.435 2509.985 1047.435 ;
    END
  END INJ_IN[34]
  PIN Data_PMOS_NOSF[366]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2507.465 1046.435 2507.745 1047.435 ;
    END
  END Data_PMOS_NOSF[366]
  PIN Data_PMOS_NOSF[367]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2506.345 1046.435 2506.625 1047.435 ;
    END
  END Data_PMOS_NOSF[367]
  PIN Data_PMOS_NOSF[368]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2504.665 1046.435 2504.945 1047.435 ;
    END
  END Data_PMOS_NOSF[368]
  PIN MASKV[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2502.425 1046.435 2502.705 1047.435 ;
    END
  END MASKV[34]
  PIN DIG_MON_PMOS_NOSF[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2500.185 1046.435 2500.465 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[34]
  PIN INJ_ROW[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2481.705 1046.435 2481.985 1047.435 ;
    END
  END INJ_ROW[16]
  PIN Data_PMOS_NOSF[344]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2480.025 1046.435 2480.305 1047.435 ;
    END
  END Data_PMOS_NOSF[344]
  PIN Data_PMOS_NOSF[356]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2477.225 1046.435 2477.505 1047.435 ;
    END
  END Data_PMOS_NOSF[356]
  PIN Data_PMOS_NOSF[343]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2476.105 1046.435 2476.385 1047.435 ;
    END
  END Data_PMOS_NOSF[343]
  PIN nTOK_PMOS_NOSF[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2434.105 1046.435 2434.385 1047.435 ;
    END
  END nTOK_PMOS_NOSF[16]
  PIN BcidMtx[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2431.865 1046.435 2432.145 1047.435 ;
    END
  END BcidMtx[99]
  PIN BcidMtx[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2430.185 1046.435 2430.465 1047.435 ;
    END
  END BcidMtx[98]
  PIN Data_PMOS_NOSF[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1305.705 1046.435 1305.985 1047.435 ;
    END
  END Data_PMOS_NOSF[51]
  PIN Data_PMOS_NOSF[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1304.025 1046.435 1304.305 1047.435 ;
    END
  END Data_PMOS_NOSF[46]
  PIN Data_PMOS_NOSF[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1302.345 1046.435 1302.625 1047.435 ;
    END
  END Data_PMOS_NOSF[43]
  PIN MASKV[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1292.265 1046.435 1292.545 1047.435 ;
    END
  END MASKV[4]
  PIN Data_HV[1145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18891.385 1046.435 18891.665 1047.435 ;
    END
  END Data_HV[1145]
  PIN DIG_MON_SEL[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1288.345 1046.435 1288.625 1047.435 ;
    END
  END DIG_MON_SEL[4]
  PIN DIG_MON_PMOS_NOSF[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1285.545 1046.435 1285.825 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[3]
  PIN Data_PMOS_NOSF[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1281.345 1046.435 1281.625 1047.435 ;
    END
  END Data_PMOS_NOSF[39]
  PIN Data_PMOS_NOSF[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1279.665 1046.435 1279.945 1047.435 ;
    END
  END Data_PMOS_NOSF[40]
  PIN Data_PMOS_NOSF[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1252.505 1046.435 1252.785 1047.435 ;
    END
  END Data_PMOS_NOSF[41]
  PIN Data_PMOS_NOSF[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1250.825 1046.435 1251.105 1047.435 ;
    END
  END Data_PMOS_NOSF[27]
  PIN INJ_IN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1249.705 1046.435 1249.985 1047.435 ;
    END
  END INJ_IN[3]
  PIN BcidMtx[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1246.905 1046.435 1247.185 1047.435 ;
    END
  END BcidMtx[10]
  PIN BcidMtx[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1244.105 1046.435 1244.385 1047.435 ;
    END
  END BcidMtx[7]
  PIN INJ_IN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1242.425 1046.435 1242.705 1047.435 ;
    END
  END INJ_IN[2]
  PIN Data_PMOS_NOSF[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1240.185 1046.435 1240.465 1047.435 ;
    END
  END Data_PMOS_NOSF[30]
  PIN Data_PMOS_NOSF[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1225.065 1046.435 1225.345 1047.435 ;
    END
  END Data_PMOS_NOSF[37]
  PIN Data_PMOS_NOSF[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1223.945 1046.435 1224.225 1047.435 ;
    END
  END Data_PMOS_NOSF[22]
  PIN MASKV[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1222.265 1046.435 1222.545 1047.435 ;
    END
  END MASKV[2]
  PIN DIG_MON_PMOS_NOSF[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1220.025 1046.435 1220.305 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[2]
  PIN DIG_MON_SEL[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1218.345 1046.435 1218.625 1047.435 ;
    END
  END DIG_MON_SEL[2]
  PIN DIG_MON_PMOS_NOSF[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1215.545 1046.435 1215.825 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[1]
  PIN Data_PMOS_NOSF[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1172.985 1046.435 1173.265 1047.435 ;
    END
  END Data_PMOS_NOSF[8]
  PIN Data_PMOS_NOSF[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1171.865 1046.435 1172.145 1047.435 ;
    END
  END Data_PMOS_NOSF[19]
  PIN Data_PMOS_NOSF[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1170.185 1046.435 1170.465 1047.435 ;
    END
  END Data_PMOS_NOSF[20]
  PIN INJ_IN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1167.385 1046.435 1167.665 1047.435 ;
    END
  END INJ_IN[1]
  PIN BcidMtx[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1165.145 1046.435 1165.425 1047.435 ;
    END
  END BcidMtx[5]
  PIN FREEZE_PMOS_NOSF[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1163.465 1046.435 1163.745 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[0]
  PIN BcidMtx[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1161.225 1046.435 1161.505 1047.435 ;
    END
  END BcidMtx[0]
  PIN Data_PMOS_NOSF[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1150.585 1046.435 1150.865 1047.435 ;
    END
  END Data_PMOS_NOSF[3]
  PIN Data_PMOS_NOSF[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1148.905 1046.435 1149.185 1047.435 ;
    END
  END Data_PMOS_NOSF[15]
  PIN Data_PMOS_NOSF[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1146.665 1046.435 1146.945 1047.435 ;
    END
  END Data_PMOS_NOSF[11]
  PIN Data_PMOS_NOSF[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1145.545 1046.435 1145.825 1047.435 ;
    END
  END Data_PMOS_NOSF[0]
  PIN MASKD[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1141.345 1046.435 1141.625 1047.435 ;
    END
  END MASKD[0]
  PIN Data_HV[1050]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18583.385 1046.435 18583.665 1047.435 ;
    END
  END Data_HV[1050]
  PIN DIG_MON_SEL[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1138.545 1046.435 1138.825 1047.435 ;
    END
  END DIG_MON_SEL[0]
  PIN DIG_MON_SEL[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2231.945 1046.435 2232.225 1047.435 ;
    END
  END DIG_MON_SEL[27]
  PIN MASKV[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2228.025 1046.435 2228.305 1047.435 ;
    END
  END MASKV[27]
  PIN Data_PMOS_NOSF[281]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2226.905 1046.435 2227.185 1047.435 ;
    END
  END Data_PMOS_NOSF[281]
  PIN Data_PMOS_NOSF[278]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2225.225 1046.435 2225.505 1047.435 ;
    END
  END Data_PMOS_NOSF[278]
  PIN Data_PMOS_NOSF[280]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2222.985 1046.435 2223.265 1047.435 ;
    END
  END Data_PMOS_NOSF[280]
  PIN INJ_IN[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2221.305 1046.435 2221.585 1047.435 ;
    END
  END INJ_IN[27]
  PIN BcidMtx[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2205.065 1046.435 2205.345 1047.435 ;
    END
  END BcidMtx[82]
  PIN BcidMtx[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2202.825 1046.435 2203.105 1047.435 ;
    END
  END BcidMtx[80]
  PIN BcidMtx[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2201.705 1046.435 2201.985 1047.435 ;
    END
  END BcidMtx[78]
  PIN Data_PMOS_NOSF[275]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2198.905 1046.435 2199.185 1047.435 ;
    END
  END Data_PMOS_NOSF[275]
  PIN Data_PMOS_NOSF[277]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2196.665 1046.435 2196.945 1047.435 ;
    END
  END Data_PMOS_NOSF[277]
  PIN Data_PMOS_NOSF[284]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2195.545 1046.435 2195.825 1047.435 ;
    END
  END Data_PMOS_NOSF[284]
  PIN Data_PMOS_NOSF[290]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2193.865 1046.435 2194.145 1047.435 ;
    END
  END Data_PMOS_NOSF[290]
  PIN MASKV[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18582.265 1046.435 18582.545 1047.435 ;
    END
  END MASKV[436]
  PIN MASKD[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18581.145 1046.435 18581.425 1047.435 ;
    END
  END MASKD[436]
  PIN Data_PMOS_NOSF[270]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2145.705 1046.435 2145.985 1047.435 ;
    END
  END Data_PMOS_NOSF[270]
  PIN Data_PMOS_NOSF[264]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2144.585 1046.435 2144.865 1047.435 ;
    END
  END Data_PMOS_NOSF[264]
  PIN Data_PMOS_NOSF[271]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2144.025 1046.435 2144.305 1047.435 ;
    END
  END Data_PMOS_NOSF[271]
  PIN Data_PMOS_NOSF[258]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2132.265 1046.435 2132.545 1047.435 ;
    END
  END Data_PMOS_NOSF[258]
  PIN INJ_IN[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2131.145 1046.435 2131.425 1047.435 ;
    END
  END INJ_IN[25]
  PIN BcidMtx[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2128.345 1046.435 2128.625 1047.435 ;
    END
  END BcidMtx[76]
  PIN BcidMtx[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2125.545 1046.435 2125.825 1047.435 ;
    END
  END BcidMtx[73]
  PIN BcidMtx[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2124.985 1046.435 2125.265 1047.435 ;
    END
  END BcidMtx[72]
  PIN Data_PMOS_NOSF[255]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2120.785 1046.435 2121.065 1047.435 ;
    END
  END Data_PMOS_NOSF[255]
  PIN Data_PMOS_NOSF[262]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2118.545 1046.435 2118.825 1047.435 ;
    END
  END Data_PMOS_NOSF[262]
  PIN Data_PMOS_NOSF[263]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2091.385 1046.435 2091.665 1047.435 ;
    END
  END Data_PMOS_NOSF[263]
  PIN Data_PMOS_NOSF[252]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2090.265 1046.435 2090.545 1047.435 ;
    END
  END Data_PMOS_NOSF[252]
  PIN MASKD[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2088.025 1046.435 2088.305 1047.435 ;
    END
  END MASKD[24]
  PIN MASKD[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2083.545 1046.435 2083.825 1047.435 ;
    END
  END MASKD[23]
  PIN Data_PMOS_NOSF[249]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2080.185 1046.435 2080.465 1047.435 ;
    END
  END Data_PMOS_NOSF[249]
  PIN Data_PMOS_NOSF[243]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2066.185 1046.435 2066.465 1047.435 ;
    END
  END Data_PMOS_NOSF[243]
  PIN Data_PMOS_NOSF[244]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2064.505 1046.435 2064.785 1047.435 ;
    END
  END Data_PMOS_NOSF[244]
  PIN Data_PMOS_NOSF[237]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2062.265 1046.435 2062.545 1047.435 ;
    END
  END Data_PMOS_NOSF[237]
  PIN nTOK_PMOS_NOSF[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2060.025 1046.435 2060.305 1047.435 ;
    END
  END nTOK_PMOS_NOSF[11]
  PIN BcidMtx[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2057.785 1046.435 2058.065 1047.435 ;
    END
  END BcidMtx[69]
  PIN BcidMtx[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2054.985 1046.435 2055.265 1047.435 ;
    END
  END BcidMtx[66]
  PIN Data_PMOS_NOSF[234]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2014.105 1046.435 2014.385 1047.435 ;
    END
  END Data_PMOS_NOSF[234]
  PIN Data_PMOS_NOSF[246]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2012.425 1046.435 2012.705 1047.435 ;
    END
  END Data_PMOS_NOSF[246]
  PIN Data_PMOS_NOSF[242]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2010.185 1046.435 2010.465 1047.435 ;
    END
  END Data_PMOS_NOSF[242]
  PIN Data_PMOS_NOSF[231]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2009.065 1046.435 2009.345 1047.435 ;
    END
  END Data_PMOS_NOSF[231]
  PIN MASKH[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2007.385 1046.435 2007.665 1047.435 ;
    END
  END MASKH[11]
  PIN DIG_MON_HV[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18580.025 1046.435 18580.305 1047.435 ;
    END
  END DIG_MON_HV[100]
  PIN DIG_MON_SEL[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2003.465 1046.435 2003.745 1047.435 ;
    END
  END DIG_MON_SEL[21]
  PIN INJ_ROW[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1991.705 1046.435 1991.985 1047.435 ;
    END
  END INJ_ROW[10]
  PIN Data_PMOS_NOSF[222]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1989.465 1046.435 1989.745 1047.435 ;
    END
  END Data_PMOS_NOSF[222]
  PIN Data_PMOS_NOSF[215]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1988.345 1046.435 1988.625 1047.435 ;
    END
  END Data_PMOS_NOSF[215]
  PIN Data_PMOS_NOSF[224]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1986.665 1046.435 1986.945 1047.435 ;
    END
  END Data_PMOS_NOSF[224]
  PIN nTOK_PMOS_NOSF[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1981.345 1046.435 1981.625 1047.435 ;
    END
  END nTOK_PMOS_NOSF[10]
  PIN BcidMtx[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1979.665 1046.435 1979.945 1047.435 ;
    END
  END BcidMtx[64]
  PIN BcidMtx[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1951.945 1046.435 1952.225 1047.435 ;
    END
  END BcidMtx[62]
  PIN DIG_MON_SEL[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1777.785 1046.435 1778.065 1047.435 ;
    END
  END DIG_MON_SEL[15]
  PIN Data_PMOS_NOSF[212]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1948.025 1046.435 1948.305 1047.435 ;
    END
  END Data_PMOS_NOSF[212]
  PIN Data_PMOS_NOSF[219]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1947.465 1046.435 1947.745 1047.435 ;
    END
  END Data_PMOS_NOSF[219]
  PIN Data_PMOS_NOSF[221]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1944.665 1046.435 1944.945 1047.435 ;
    END
  END Data_PMOS_NOSF[221]
  PIN Data_PMOS_NOSF[210]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1943.545 1046.435 1943.825 1047.435 ;
    END
  END Data_PMOS_NOSF[210]
  PIN MASKH[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1941.865 1046.435 1942.145 1047.435 ;
    END
  END MASKH[10]
  PIN DIG_MON_PMOS_NOSF[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1922.825 1046.435 1923.105 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[19]
  PIN Data_PMOS_NOSF[207]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1920.585 1046.435 1920.865 1047.435 ;
    END
  END Data_PMOS_NOSF[207]
  PIN Data_PMOS_NOSF[208]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1918.905 1046.435 1919.185 1047.435 ;
    END
  END Data_PMOS_NOSF[208]
  PIN Data_PMOS_NOSF[209]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1917.225 1046.435 1917.505 1047.435 ;
    END
  END Data_PMOS_NOSF[209]
  PIN Data_PMOS_NOSF[195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1915.545 1046.435 1915.825 1047.435 ;
    END
  END Data_PMOS_NOSF[195]
  PIN BcidMtx[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1872.985 1046.435 1873.265 1047.435 ;
    END
  END BcidMtx[59]
  PIN FREEZE_PMOS_NOSF[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1871.305 1046.435 1871.585 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[9]
  PIN BcidMtx[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4672.985 1046.435 4673.265 1047.435 ;
    END
  END BcidMtx[269]
  PIN BcidMtx[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4670.185 1046.435 4670.465 1047.435 ;
    END
  END BcidMtx[266]
  PIN BcidMtx[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4669.625 1046.435 4669.905 1047.435 ;
    END
  END BcidMtx[265]
  PIN Data_PMOS_NOSF[927]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4666.825 1046.435 4667.105 1047.435 ;
    END
  END Data_PMOS_NOSF[927]
  PIN Data_PMOS_NOSF[928]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4664.025 1046.435 4664.305 1047.435 ;
    END
  END Data_PMOS_NOSF[928]
  PIN Data_PMOS_NOSF[940]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4663.465 1046.435 4663.745 1047.435 ;
    END
  END Data_PMOS_NOSF[940]
  PIN Data_PMOS_NOSF[924]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4661.785 1046.435 4662.065 1047.435 ;
    END
  END Data_PMOS_NOSF[924]
  PIN DIG_MON_PMOS_NOSF[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4650.025 1046.435 4650.305 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[88]
  PIN MASKD[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4646.665 1046.435 4646.945 1047.435 ;
    END
  END MASKD[87]
  PIN Data_PMOS_NOSF[911]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4640.785 1046.435 4641.065 1047.435 ;
    END
  END Data_PMOS_NOSF[911]
  PIN Data_PMOS_NOSF[915]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4640.225 1046.435 4640.505 1047.435 ;
    END
  END Data_PMOS_NOSF[915]
  PIN Data_PMOS_NOSF[916]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4613.065 1046.435 4613.345 1047.435 ;
    END
  END Data_PMOS_NOSF[916]
  PIN INJ_IN[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4609.705 1046.435 4609.985 1047.435 ;
    END
  END INJ_IN[87]
  PIN nTOK_PMOS_NOSF[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4608.585 1046.435 4608.865 1047.435 ;
    END
  END nTOK_PMOS_NOSF[43]
  PIN BcidMtx[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4606.345 1046.435 4606.625 1047.435 ;
    END
  END BcidMtx[261]
  PIN BcidMtx[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4603.545 1046.435 4603.825 1047.435 ;
    END
  END BcidMtx[258]
  PIN INJ_IN[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4602.425 1046.435 4602.705 1047.435 ;
    END
  END INJ_IN[86]
  PIN Data_PMOS_NOSF[912]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4600.185 1046.435 4600.465 1047.435 ;
    END
  END Data_PMOS_NOSF[912]
  PIN Data_PMOS_NOSF[914]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4584.505 1046.435 4584.785 1047.435 ;
    END
  END Data_PMOS_NOSF[914]
  PIN Data_PMOS_NOSF[904]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4583.945 1046.435 4584.225 1047.435 ;
    END
  END Data_PMOS_NOSF[904]
  PIN MASKV[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4582.265 1046.435 4582.545 1047.435 ;
    END
  END MASKV[86]
  PIN DIG_MON_SEL[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4578.345 1046.435 4578.625 1047.435 ;
    END
  END DIG_MON_SEL[86]
  PIN DIG_MON_SEL[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4577.785 1046.435 4578.065 1047.435 ;
    END
  END DIG_MON_SEL[85]
  PIN INJ_ROW[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4574.425 1046.435 4574.705 1047.435 ;
    END
  END INJ_ROW[42]
  PIN Data_PMOS_NOSF[894]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4532.425 1046.435 4532.705 1047.435 ;
    END
  END Data_PMOS_NOSF[894]
  PIN Data_PMOS_NOSF[901]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4531.865 1046.435 4532.145 1047.435 ;
    END
  END Data_PMOS_NOSF[901]
  PIN Data_PMOS_NOSF[895]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4530.745 1046.435 4531.025 1047.435 ;
    END
  END Data_PMOS_NOSF[895]
  PIN INJ_IN[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4527.385 1046.435 4527.665 1047.435 ;
    END
  END INJ_IN[85]
  PIN nTOK_PMOS_NOSF[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4526.265 1046.435 4526.545 1047.435 ;
    END
  END nTOK_PMOS_NOSF[42]
  PIN BcidMtx[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4521.785 1046.435 4522.065 1047.435 ;
    END
  END BcidMtx[253]
  PIN BcidMtx[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4521.225 1046.435 4521.505 1047.435 ;
    END
  END BcidMtx[252]
  PIN Data_PMOS_NOSF[884]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4510.025 1046.435 4510.305 1047.435 ;
    END
  END Data_PMOS_NOSF[884]
  PIN Data_PMOS_NOSF[898]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4507.225 1046.435 4507.505 1047.435 ;
    END
  END Data_PMOS_NOSF[898]
  PIN Data_PMOS_NOSF[893]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4506.665 1046.435 4506.945 1047.435 ;
    END
  END Data_PMOS_NOSF[893]
  PIN Data_PMOS_NOSF[899]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4504.985 1046.435 4505.265 1047.435 ;
    END
  END Data_PMOS_NOSF[899]
  PIN DIG_MON_SEL[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4498.545 1046.435 4498.825 1047.435 ;
    END
  END DIG_MON_SEL[84]
  PIN MASKD[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5590.825 1046.435 5591.105 1047.435 ;
    END
  END MASKD[111]
  PIN Data_PMOS_NOSF[1163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5586.905 1046.435 5587.185 1047.435 ;
    END
  END Data_PMOS_NOSF[1163]
  PIN Data_PMOS_NOSF[1167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5586.345 1046.435 5586.625 1047.435 ;
    END
  END Data_PMOS_NOSF[1167]
  PIN Data_HV[1119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18862.265 1046.435 18862.545 1047.435 ;
    END
  END Data_HV[1119]
  PIN Data_PMOS_NOSF[1161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5582.425 1046.435 5582.705 1047.435 ;
    END
  END Data_PMOS_NOSF[1161]
  PIN INJ_IN[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5581.305 1046.435 5581.585 1047.435 ;
    END
  END INJ_IN[111]
  PIN BcidMtx[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5565.065 1046.435 5565.345 1047.435 ;
    END
  END BcidMtx[334]
  PIN BcidMtx[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5562.265 1046.435 5562.545 1047.435 ;
    END
  END BcidMtx[331]
  PIN BcidMtx[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5561.705 1046.435 5561.985 1047.435 ;
    END
  END BcidMtx[330]
  PIN Data_PMOS_NOSF[1157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5558.905 1046.435 5559.185 1047.435 ;
    END
  END Data_PMOS_NOSF[1157]
  PIN Data_PMOS_NOSF[1171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5556.105 1046.435 5556.385 1047.435 ;
    END
  END Data_PMOS_NOSF[1171]
  PIN Data_PMOS_NOSF[1166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5555.545 1046.435 5555.825 1047.435 ;
    END
  END Data_PMOS_NOSF[1166]
  PIN Data_PMOS_NOSF[1172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5553.865 1046.435 5554.145 1047.435 ;
    END
  END Data_PMOS_NOSF[1172]
  PIN DIG_MON_SEL[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5510.745 1046.435 5511.025 1047.435 ;
    END
  END DIG_MON_SEL[110]
  PIN DIG_MON_PMOS_NOSF[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5507.945 1046.435 5508.225 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[109]
  PIN Data_PMOS_NOSF[1146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5504.585 1046.435 5504.865 1047.435 ;
    END
  END Data_PMOS_NOSF[1146]
  PIN Data_PMOS_NOSF[1153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5504.025 1046.435 5504.305 1047.435 ;
    END
  END Data_PMOS_NOSF[1153]
  PIN Data_PMOS_NOSF[1154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5502.345 1046.435 5502.625 1047.435 ;
    END
  END Data_PMOS_NOSF[1154]
  PIN nTOK_PMOS_NOSF[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5490.025 1046.435 5490.305 1047.435 ;
    END
  END nTOK_PMOS_NOSF[54]
  PIN BcidMtx[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5488.905 1046.435 5489.185 1047.435 ;
    END
  END BcidMtx[329]
  PIN FREEZE_PMOS_NOSF[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5487.225 1046.435 5487.505 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[54]
  PIN INJ_IN[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5481.905 1046.435 5482.185 1047.435 ;
    END
  END INJ_IN[108]
  PIN Data_PMOS_NOSF[1137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5480.785 1046.435 5481.065 1047.435 ;
    END
  END Data_PMOS_NOSF[1137]
  PIN Data_PMOS_NOSF[1149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5479.105 1046.435 5479.385 1047.435 ;
    END
  END Data_PMOS_NOSF[1149]
  PIN Data_PMOS_NOSF[1135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5450.825 1046.435 5451.105 1047.435 ;
    END
  END Data_PMOS_NOSF[1135]
  PIN Data_PMOS_NOSF[1134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5450.265 1046.435 5450.545 1047.435 ;
    END
  END Data_PMOS_NOSF[1134]
  PIN MASKH[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5448.585 1046.435 5448.865 1047.435 ;
    END
  END MASKH[54]
  PIN DIG_MON_SEL[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5444.665 1046.435 5444.945 1047.435 ;
    END
  END DIG_MON_SEL[107]
  PIN MASKD[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5443.545 1046.435 5443.825 1047.435 ;
    END
  END MASKD[107]
  PIN MASKV[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5440.745 1046.435 5441.025 1047.435 ;
    END
  END MASKV[107]
  PIN Data_PMOS_NOSF[1118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5425.065 1046.435 5425.345 1047.435 ;
    END
  END Data_PMOS_NOSF[1118]
  PIN Data_PMOS_NOSF[1126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5424.505 1046.435 5424.785 1047.435 ;
    END
  END Data_PMOS_NOSF[1126]
  PIN Data_PMOS_NOSF[1133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5423.945 1046.435 5424.225 1047.435 ;
    END
  END Data_PMOS_NOSF[1133]
  PIN nTOK_PMOS_NOSF[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5420.025 1046.435 5420.305 1047.435 ;
    END
  END nTOK_PMOS_NOSF[53]
  PIN BcidMtx[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5418.905 1046.435 5419.185 1047.435 ;
    END
  END BcidMtx[323]
  PIN FREEZE_PMOS_NOSF[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5417.225 1046.435 5417.505 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[53]
  PIN INJ_IN[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5413.865 1046.435 5414.145 1047.435 ;
    END
  END INJ_IN[106]
  PIN Data_PMOS_NOSF[1116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5374.105 1046.435 5374.385 1047.435 ;
    END
  END Data_PMOS_NOSF[1116]
  PIN Data_PMOS_NOSF[1128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5372.425 1046.435 5372.705 1047.435 ;
    END
  END Data_PMOS_NOSF[1128]
  PIN Data_PMOS_NOSF[1114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5369.625 1046.435 5369.905 1047.435 ;
    END
  END Data_PMOS_NOSF[1114]
  PIN Data_PMOS_NOSF[1113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5369.065 1046.435 5369.345 1047.435 ;
    END
  END Data_PMOS_NOSF[1113]
  PIN MASKH[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5367.385 1046.435 5367.665 1047.435 ;
    END
  END MASKH[53]
  PIN DIG_MON_SEL[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5363.465 1046.435 5363.745 1047.435 ;
    END
  END DIG_MON_SEL[105]
  PIN MASKD[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5362.345 1046.435 5362.625 1047.435 ;
    END
  END MASKD[105]
  PIN MASKV[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5351.145 1046.435 5351.425 1047.435 ;
    END
  END MASKV[105]
  PIN Data_PMOS_NOSF[1097]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5348.345 1046.435 5348.625 1047.435 ;
    END
  END Data_PMOS_NOSF[1097]
  PIN Data_PMOS_NOSF[1105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5347.785 1046.435 5348.065 1047.435 ;
    END
  END Data_PMOS_NOSF[1105]
  PIN Data_PMOS_NOSF[1099]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5346.105 1046.435 5346.385 1047.435 ;
    END
  END Data_PMOS_NOSF[1099]
  PIN BcidMtx[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5339.665 1046.435 5339.945 1047.435 ;
    END
  END BcidMtx[316]
  PIN BcidMtx[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5339.105 1046.435 5339.385 1047.435 ;
    END
  END BcidMtx[315]
  PIN BcidMtx[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5311.385 1046.435 5311.665 1047.435 ;
    END
  END BcidMtx[313]
  PIN Data_PMOS_NOSF[1101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5307.465 1046.435 5307.745 1047.435 ;
    END
  END Data_PMOS_NOSF[1101]
  PIN Data_PMOS_NOSF[1107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5306.905 1046.435 5307.185 1047.435 ;
    END
  END Data_PMOS_NOSF[1107]
  PIN Data_PMOS_NOSF[1108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5305.225 1046.435 5305.505 1047.435 ;
    END
  END Data_PMOS_NOSF[1108]
  PIN MASKV[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5302.425 1046.435 5302.705 1047.435 ;
    END
  END MASKV[104]
  PIN MASKH[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5301.865 1046.435 5302.145 1047.435 ;
    END
  END MASKH[52]
  PIN INJ_ROW[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5281.705 1046.435 5281.985 1047.435 ;
    END
  END INJ_ROW[51]
  PIN MASKV[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5281.145 1046.435 5281.425 1047.435 ;
    END
  END MASKV[103]
  PIN Data_PMOS_NOSF[1083]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5279.465 1046.435 5279.745 1047.435 ;
    END
  END Data_PMOS_NOSF[1083]
  PIN Data_PMOS_NOSF[1085]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5276.665 1046.435 5276.945 1047.435 ;
    END
  END Data_PMOS_NOSF[1085]
  PIN Data_PMOS_NOSF[1078]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5276.105 1046.435 5276.385 1047.435 ;
    END
  END Data_PMOS_NOSF[1078]
  PIN nTOK_PMOS_NOSF[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5234.105 1046.435 5234.385 1047.435 ;
    END
  END nTOK_PMOS_NOSF[51]
  PIN Read_PMOS[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5790.745 1046.435 5791.025 1047.435 ;
    END
  END Read_PMOS[2]
  PIN BcidMtx[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5789.065 1046.435 5789.345 1047.435 ;
    END
  END BcidMtx[348]
  PIN Data_PMOS[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5786.265 1046.435 5786.545 1047.435 ;
    END
  END Data_PMOS[44]
  PIN Data_PMOS[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5784.025 1046.435 5784.305 1047.435 ;
    END
  END Data_PMOS[46]
  PIN Data_PMOS[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5782.345 1046.435 5782.625 1047.435 ;
    END
  END Data_PMOS[43]
  PIN MASKV[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5772.265 1046.435 5772.545 1047.435 ;
    END
  END MASKV[116]
  PIN DIG_MON_PMOS[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5770.025 1046.435 5770.305 1047.435 ;
    END
  END DIG_MON_PMOS[4]
  PIN DIG_MON_SEL[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5767.785 1046.435 5768.065 1047.435 ;
    END
  END DIG_MON_SEL[115]
  PIN DIG_MON_PMOS[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5765.545 1046.435 5765.825 1047.435 ;
    END
  END DIG_MON_PMOS[3]
  PIN Data_PMOS[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5760.785 1046.435 5761.065 1047.435 ;
    END
  END Data_PMOS[29]
  PIN Data_PMOS[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5759.105 1046.435 5759.385 1047.435 ;
    END
  END Data_PMOS[26]
  PIN Data_PMOS[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5731.945 1046.435 5732.225 1047.435 ;
    END
  END Data_PMOS[35]
  PIN Data_PMOS[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5730.825 1046.435 5731.105 1047.435 ;
    END
  END Data_PMOS[27]
  PIN BcidMtx[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5726.345 1046.435 5726.625 1047.435 ;
    END
  END BcidMtx[345]
  PIN BcidMtx[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5723.545 1046.435 5723.825 1047.435 ;
    END
  END BcidMtx[342]
  PIN Data_PMOS[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5720.745 1046.435 5721.025 1047.435 ;
    END
  END Data_PMOS[23]
  PIN Data_PMOS[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5720.185 1046.435 5720.465 1047.435 ;
    END
  END Data_PMOS[30]
  PIN Data_PMOS[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5705.625 1046.435 5705.905 1047.435 ;
    END
  END Data_PMOS[25]
  PIN Data_PMOS[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5702.825 1046.435 5703.105 1047.435 ;
    END
  END Data_PMOS[38]
  PIN BcidMtx[1330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18858.345 1046.435 18858.625 1047.435 ;
    END
  END BcidMtx[1330]
  PIN MASKD[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5701.145 1046.435 5701.425 1047.435 ;
    END
  END MASKD[114]
  PIN DIG_MON_SEL[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5697.785 1046.435 5698.065 1047.435 ;
    END
  END DIG_MON_SEL[113]
  PIN INJ_ROW[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5694.425 1046.435 5694.705 1047.435 ;
    END
  END INJ_ROW[56]
  PIN MASKV[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5693.865 1046.435 5694.145 1047.435 ;
    END
  END MASKV[113]
  PIN Data_PMOS[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5651.305 1046.435 5651.585 1047.435 ;
    END
  END Data_PMOS[5]
  PIN Data_PMOS[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5649.625 1046.435 5649.905 1047.435 ;
    END
  END Data_PMOS[14]
  PIN Data_PMOS[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5648.505 1046.435 5648.785 1047.435 ;
    END
  END Data_PMOS[6]
  PIN BcidMtx[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5644.585 1046.435 5644.865 1047.435 ;
    END
  END BcidMtx[340]
  PIN Read_PMOS[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5642.905 1046.435 5643.185 1047.435 ;
    END
  END Read_PMOS[0]
  PIN BcidMtx[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5641.785 1046.435 5642.065 1047.435 ;
    END
  END BcidMtx[337]
  PIN Data_PMOS[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5629.465 1046.435 5629.745 1047.435 ;
    END
  END Data_PMOS[9]
  PIN Data_PMOS[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5628.345 1046.435 5628.625 1047.435 ;
    END
  END Data_PMOS[10]
  PIN Data_PMOS[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5627.225 1046.435 5627.505 1047.435 ;
    END
  END Data_PMOS[16]
  PIN Data_PMOS[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5624.985 1046.435 5625.265 1047.435 ;
    END
  END Data_PMOS[17]
  PIN MASKH[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5621.905 1046.435 5622.185 1047.435 ;
    END
  END MASKH[56]
  PIN DIG_MON_PMOS[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5620.225 1046.435 5620.505 1047.435 ;
    END
  END DIG_MON_PMOS[0]
  PIN DIG_MON_SEL[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6711.945 1046.435 6712.225 1047.435 ;
    END
  END DIG_MON_SEL[139]
  PIN DIG_MON_PMOS[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6709.705 1046.435 6709.985 1047.435 ;
    END
  END DIG_MON_PMOS[27]
  PIN Data_PMOS[291]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6707.465 1046.435 6707.745 1047.435 ;
    END
  END Data_PMOS[291]
  PIN Data_PMOS[278]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6705.225 1046.435 6705.505 1047.435 ;
    END
  END Data_PMOS[278]
  PIN Data_PMOS[286]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6704.665 1046.435 6704.945 1047.435 ;
    END
  END Data_PMOS[286]
  PIN Data_PMOS[280]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6702.985 1046.435 6703.265 1047.435 ;
    END
  END Data_PMOS[280]
  PIN nTOK_PMOS[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6700.185 1046.435 6700.465 1047.435 ;
    END
  END nTOK_PMOS[13]
  PIN BcidMtx[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6684.505 1046.435 6684.785 1047.435 ;
    END
  END BcidMtx[417]
  PIN BcidMtx[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6682.825 1046.435 6683.105 1047.435 ;
    END
  END BcidMtx[416]
  PIN INJ_IN[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6680.585 1046.435 6680.865 1047.435 ;
    END
  END INJ_IN[138]
  PIN Data_PMOS[282]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6678.345 1046.435 6678.625 1047.435 ;
    END
  END Data_PMOS[282]
  PIN Data_PMOS[277]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6676.665 1046.435 6676.945 1047.435 ;
    END
  END Data_PMOS[277]
  PIN Data_PMOS[273]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6674.425 1046.435 6674.705 1047.435 ;
    END
  END Data_PMOS[273]
  PIN MASKV[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6634.665 1046.435 6634.945 1047.435 ;
    END
  END MASKV[138]
  PIN MASKD[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6633.545 1046.435 6633.825 1047.435 ;
    END
  END MASKD[138]
  PIN DIG_MON_SEL[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6630.745 1046.435 6631.025 1047.435 ;
    END
  END DIG_MON_SEL[138]
  PIN DIG_MON_PMOS[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6627.945 1046.435 6628.225 1047.435 ;
    END
  END DIG_MON_PMOS[25]
  PIN Data_PMOS[270]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6625.705 1046.435 6625.985 1047.435 ;
    END
  END Data_PMOS[270]
  PIN Data_PMOS[271]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6624.025 1046.435 6624.305 1047.435 ;
    END
  END Data_PMOS[271]
  PIN Data_PMOS[272]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6622.345 1046.435 6622.625 1047.435 ;
    END
  END Data_PMOS[272]
  PIN Data_PMOS[258]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6612.265 1046.435 6612.545 1047.435 ;
    END
  END Data_PMOS[258]
  PIN BcidMtx[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6608.905 1046.435 6609.185 1047.435 ;
    END
  END BcidMtx[413]
  PIN FREEZE_PMOS[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6607.225 1046.435 6607.505 1047.435 ;
    END
  END FREEZE_PMOS[12]
  PIN BcidMtx[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6605.545 1046.435 6605.825 1047.435 ;
    END
  END BcidMtx[409]
  PIN Data_PMOS[254]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6600.225 1046.435 6600.505 1047.435 ;
    END
  END Data_PMOS[254]
  PIN Data_PMOS[267]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6599.105 1046.435 6599.385 1047.435 ;
    END
  END Data_PMOS[267]
  PIN Data_PMOS[268]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6571.945 1046.435 6572.225 1047.435 ;
    END
  END Data_PMOS[268]
  PIN Data_PMOS[269]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6569.705 1046.435 6569.985 1047.435 ;
    END
  END Data_PMOS[269]
  PIN MASKH[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6568.585 1046.435 6568.865 1047.435 ;
    END
  END MASKH[68]
  PIN DIG_MON_SEL[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6564.665 1046.435 6564.945 1047.435 ;
    END
  END DIG_MON_SEL[135]
  PIN INJ_ROW[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6561.305 1046.435 6561.585 1047.435 ;
    END
  END INJ_ROW[67]
  PIN Data_PMOS[239]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6559.625 1046.435 6559.905 1047.435 ;
    END
  END Data_PMOS[239]
  PIN Data_PMOS[236]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6545.065 1046.435 6545.345 1047.435 ;
    END
  END Data_PMOS[236]
  PIN Data_PMOS[245]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6543.385 1046.435 6543.665 1047.435 ;
    END
  END Data_PMOS[245]
  PIN INJ_IN[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6541.145 1046.435 6541.425 1047.435 ;
    END
  END INJ_IN[135]
  PIN BcidMtx[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6537.785 1046.435 6538.065 1047.435 ;
    END
  END BcidMtx[405]
  PIN Read_PMOS[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6536.665 1046.435 6536.945 1047.435 ;
    END
  END Read_PMOS[11]
  PIN BcidMtx[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6534.985 1046.435 6535.265 1047.435 ;
    END
  END BcidMtx[402]
  PIN Data_PMOS[233]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6493.545 1046.435 6493.825 1047.435 ;
    END
  END Data_PMOS[233]
  PIN Data_PMOS[241]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6491.865 1046.435 6492.145 1047.435 ;
    END
  END Data_PMOS[241]
  PIN Data_PMOS[242]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6490.185 1046.435 6490.465 1047.435 ;
    END
  END Data_PMOS[242]
  PIN Data_PMOS[248]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6488.505 1046.435 6488.785 1047.435 ;
    END
  END Data_PMOS[248]
  PIN MASKD[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6486.825 1046.435 6487.105 1047.435 ;
    END
  END MASKD[134]
  PIN DIG_MON_SEL[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6484.025 1046.435 6484.305 1047.435 ;
    END
  END DIG_MON_SEL[134]
  PIN INJ_ROW[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6471.705 1046.435 6471.985 1047.435 ;
    END
  END INJ_ROW[66]
  PIN Data_PMOS[228]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6470.585 1046.435 6470.865 1047.435 ;
    END
  END Data_PMOS[228]
  PIN Data_PMOS[229]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6468.905 1046.435 6469.185 1047.435 ;
    END
  END Data_PMOS[229]
  PIN Data_PMOS[224]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6466.665 1046.435 6466.945 1047.435 ;
    END
  END Data_PMOS[224]
  PIN Data_PMOS[216]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6465.545 1046.435 6465.825 1047.435 ;
    END
  END Data_PMOS[216]
  PIN BcidMtx[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6460.225 1046.435 6460.505 1047.435 ;
    END
  END BcidMtx[401]
  PIN BcidMtx[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6431.945 1046.435 6432.225 1047.435 ;
    END
  END BcidMtx[398]
  PIN BcidMtx[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6430.825 1046.435 6431.105 1047.435 ;
    END
  END BcidMtx[396]
  PIN Data_PMOS[212]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6428.025 1046.435 6428.305 1047.435 ;
    END
  END Data_PMOS[212]
  PIN Data_PMOS[220]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6426.345 1046.435 6426.625 1047.435 ;
    END
  END Data_PMOS[220]
  PIN Data_PMOS[221]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6424.665 1046.435 6424.945 1047.435 ;
    END
  END Data_PMOS[221]
  PIN Data_PMOS[227]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6422.985 1046.435 6423.265 1047.435 ;
    END
  END Data_PMOS[227]
  PIN MASKD[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6421.305 1046.435 6421.585 1047.435 ;
    END
  END MASKD[132]
  PIN DIG_MON_SEL[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6405.625 1046.435 6405.905 1047.435 ;
    END
  END DIG_MON_SEL[132]
  PIN DIG_MON_PMOS[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6402.825 1046.435 6403.105 1047.435 ;
    END
  END DIG_MON_PMOS[19]
  PIN Data_PMOS[197]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6400.025 1046.435 6400.305 1047.435 ;
    END
  END Data_PMOS[197]
  PIN Data_PMOS[208]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6398.905 1046.435 6399.185 1047.435 ;
    END
  END Data_PMOS[208]
  PIN Data_PMOS[209]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6397.225 1046.435 6397.505 1047.435 ;
    END
  END Data_PMOS[209]
  PIN Data_PMOS[195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6395.545 1046.435 6395.825 1047.435 ;
    END
  END Data_PMOS[195]
  PIN BcidMtx[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6352.985 1046.435 6353.265 1047.435 ;
    END
  END BcidMtx[395]
  PIN FREEZE_PMOS[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6351.305 1046.435 6351.585 1047.435 ;
    END
  END FREEZE_PMOS[9]
  PIN Data_PMOS[1077]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9755.545 1046.435 9755.825 1047.435 ;
    END
  END Data_PMOS[1077]
  PIN BcidMtx[647]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9712.985 1046.435 9713.265 1047.435 ;
    END
  END BcidMtx[647]
  PIN FREEZE_PMOS[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9711.305 1046.435 9711.585 1047.435 ;
    END
  END FREEZE_PMOS[51]
  PIN BcidMtx[643]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9709.625 1046.435 9709.905 1047.435 ;
    END
  END BcidMtx[643]
  PIN Data_PMOS[1074]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9706.825 1046.435 9707.105 1047.435 ;
    END
  END Data_PMOS[1074]
  PIN Data_PMOS[1086]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9705.145 1046.435 9705.425 1047.435 ;
    END
  END Data_PMOS[1086]
  PIN Data_PMOS[1087]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9703.465 1046.435 9703.745 1047.435 ;
    END
  END Data_PMOS[1087]
  PIN Data_PMOS[1071]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9701.785 1046.435 9702.065 1047.435 ;
    END
  END Data_PMOS[1071]
  PIN MASKH[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9691.705 1046.435 9691.985 1047.435 ;
    END
  END MASKH[107]
  PIN DIG_MON_SEL[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9687.785 1046.435 9688.065 1047.435 ;
    END
  END DIG_MON_SEL[213]
  PIN MASKV[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9681.905 1046.435 9682.185 1047.435 ;
    END
  END MASKV[213]
  PIN Data_PMOS[1062]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9680.225 1046.435 9680.505 1047.435 ;
    END
  END Data_PMOS[1062]
  PIN Data_PMOS[1063]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9653.065 1046.435 9653.345 1047.435 ;
    END
  END Data_PMOS[1063]
  PIN Data_PMOS[1057]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9651.385 1046.435 9651.665 1047.435 ;
    END
  END Data_PMOS[1057]
  PIN BcidMtx[640]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9646.905 1046.435 9647.185 1047.435 ;
    END
  END BcidMtx[640]
  PIN FREEZE_PMOS[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9645.785 1046.435 9646.065 1047.435 ;
    END
  END FREEZE_PMOS[50]
  PIN BcidMtx[638]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9644.665 1046.435 9644.945 1047.435 ;
    END
  END BcidMtx[638]
  PIN Data_PMOS[1052]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9640.745 1046.435 9641.025 1047.435 ;
    END
  END Data_PMOS[1052]
  PIN Data_PMOS[1065]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9626.745 1046.435 9627.025 1047.435 ;
    END
  END Data_PMOS[1065]
  PIN Data_PMOS[1054]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9625.625 1046.435 9625.905 1047.435 ;
    END
  END Data_PMOS[1054]
  PIN Data_PMOS[1067]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9622.825 1046.435 9623.105 1047.435 ;
    END
  END Data_PMOS[1067]
  PIN MASKH[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9621.705 1046.435 9621.985 1047.435 ;
    END
  END MASKH[106]
  PIN MASKV[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18791.145 1046.435 18791.425 1047.435 ;
    END
  END MASKV[441]
  PIN MASKD[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9616.665 1046.435 9616.945 1047.435 ;
    END
  END MASKD[211]
  PIN DIG_MON_PMOS[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9615.545 1046.435 9615.825 1047.435 ;
    END
  END DIG_MON_PMOS[99]
  PIN MASKV[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9613.865 1046.435 9614.145 1047.435 ;
    END
  END MASKV[211]
  PIN Data_PMOS[1042]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9570.745 1046.435 9571.025 1047.435 ;
    END
  END Data_PMOS[1042]
  PIN Data_PMOS[1043]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9569.625 1046.435 9569.905 1047.435 ;
    END
  END Data_PMOS[1043]
  PIN INJ_IN[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9567.385 1046.435 9567.665 1047.435 ;
    END
  END INJ_IN[211]
  PIN BcidMtx[633]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9564.025 1046.435 9564.305 1047.435 ;
    END
  END BcidMtx[633]
  PIN Read_PMOS[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9562.905 1046.435 9563.185 1047.435 ;
    END
  END Read_PMOS[49]
  PIN BcidMtx[630]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9561.225 1046.435 9561.505 1047.435 ;
    END
  END BcidMtx[630]
  PIN Data_PMOS[1038]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9549.465 1046.435 9549.745 1047.435 ;
    END
  END Data_PMOS[1038]
  PIN Data_PMOS[1039]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9548.345 1046.435 9548.625 1047.435 ;
    END
  END Data_PMOS[1039]
  PIN Data_PMOS[1040]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9546.665 1046.435 9546.945 1047.435 ;
    END
  END Data_PMOS[1040]
  PIN MASKV[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9542.465 1046.435 9542.745 1047.435 ;
    END
  END MASKV[210]
  PIN MASKD[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9541.345 1046.435 9541.625 1047.435 ;
    END
  END MASKD[210]
  PIN MASKD[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10630.825 1046.435 10631.105 1047.435 ;
    END
  END MASKD[237]
  PIN INJ_ROW[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10628.585 1046.435 10628.865 1047.435 ;
    END
  END INJ_ROW[118]
  PIN Data_COMP[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10626.905 1046.435 10627.185 1047.435 ;
    END
  END Data_COMP[134]
  PIN Data_COMP[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10625.225 1046.435 10625.505 1047.435 ;
    END
  END Data_COMP[131]
  PIN Data_COMP[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10624.105 1046.435 10624.385 1047.435 ;
    END
  END Data_COMP[146]
  PIN Data_COMP[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10622.985 1046.435 10623.265 1047.435 ;
    END
  END Data_COMP[133]
  PIN BcidMtx[712]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10605.065 1046.435 10605.345 1047.435 ;
    END
  END BcidMtx[712]
  PIN FREEZE_COMP[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10603.945 1046.435 10604.225 1047.435 ;
    END
  END FREEZE_COMP[6]
  PIN BcidMtx[710]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10602.825 1046.435 10603.105 1047.435 ;
    END
  END BcidMtx[710]
  PIN Data_COMP[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10598.905 1046.435 10599.185 1047.435 ;
    END
  END Data_COMP[128]
  PIN Data_COMP[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10597.785 1046.435 10598.065 1047.435 ;
    END
  END Data_COMP[141]
  PIN Data_COMP[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10596.665 1046.435 10596.945 1047.435 ;
    END
  END Data_COMP[130]
  PIN Data_COMP[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10593.865 1046.435 10594.145 1047.435 ;
    END
  END Data_COMP[143]
  PIN MASKH[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10554.105 1046.435 10554.385 1047.435 ;
    END
  END MASKH[118]
  PIN DIG_MON_COMP[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10552.425 1046.435 10552.705 1047.435 ;
    END
  END DIG_MON_COMP[12]
  PIN MASKD[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10549.065 1046.435 10549.345 1047.435 ;
    END
  END MASKD[235]
  PIN INJ_ROW[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10546.825 1046.435 10547.105 1047.435 ;
    END
  END INJ_ROW[117]
  PIN Data_COMP[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10545.705 1046.435 10545.985 1047.435 ;
    END
  END Data_COMP[123]
  PIN Data_COMP[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10542.905 1046.435 10543.185 1047.435 ;
    END
  END Data_COMP[118]
  PIN Data_COMP[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10541.785 1046.435 10542.065 1047.435 ;
    END
  END Data_COMP[119]
  PIN Data_COMP[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10532.265 1046.435 10532.545 1047.435 ;
    END
  END Data_COMP[111]
  PIN BcidMtx[705]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10527.785 1046.435 10528.065 1047.435 ;
    END
  END BcidMtx[705]
  PIN Read_COMP[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10526.665 1046.435 10526.945 1047.435 ;
    END
  END Read_COMP[5]
  PIN BcidMtx[703]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10525.545 1046.435 10525.825 1047.435 ;
    END
  END BcidMtx[703]
  PIN Data_COMP[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10519.665 1046.435 10519.945 1047.435 ;
    END
  END Data_COMP[114]
  PIN Data_COMP[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10518.545 1046.435 10518.825 1047.435 ;
    END
  END Data_COMP[115]
  PIN Data_COMP[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10491.945 1046.435 10492.225 1047.435 ;
    END
  END Data_COMP[121]
  PIN MASKV[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10489.145 1046.435 10489.425 1047.435 ;
    END
  END MASKV[234]
  PIN MASKD[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10488.025 1046.435 10488.305 1047.435 ;
    END
  END MASKD[234]
  PIN MASKD[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10483.545 1046.435 10483.825 1047.435 ;
    END
  END MASKD[233]
  PIN MASKV[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10480.745 1046.435 10481.025 1047.435 ;
    END
  END MASKV[233]
  PIN Data_COMP[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10479.625 1046.435 10479.905 1047.435 ;
    END
  END Data_COMP[92]
  PIN Data_COMP[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10464.505 1046.435 10464.785 1047.435 ;
    END
  END Data_COMP[97]
  PIN Data_COMP[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10462.825 1046.435 10463.105 1047.435 ;
    END
  END Data_COMP[91]
  PIN INJ_IN[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10461.145 1046.435 10461.425 1047.435 ;
    END
  END INJ_IN[233]
  PIN BcidMtx[701]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10458.905 1046.435 10459.185 1047.435 ;
    END
  END BcidMtx[701]
  PIN BcidMtx[698]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10456.105 1046.435 10456.385 1047.435 ;
    END
  END BcidMtx[698]
  PIN BcidMtx[696]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10454.985 1046.435 10455.265 1047.435 ;
    END
  END BcidMtx[696]
  PIN Data_COMP[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10414.105 1046.435 10414.385 1047.435 ;
    END
  END Data_COMP[87]
  PIN Data_COMP[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10411.305 1046.435 10411.585 1047.435 ;
    END
  END Data_COMP[88]
  PIN Data_COMP[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10410.185 1046.435 10410.465 1047.435 ;
    END
  END Data_COMP[95]
  PIN Data_COMP[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10409.065 1046.435 10409.345 1047.435 ;
    END
  END Data_COMP[84]
  PIN DIG_MON_COMP[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10405.705 1046.435 10405.985 1047.435 ;
    END
  END DIG_MON_COMP[8]
  PIN DIG_MON_SEL[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10404.025 1046.435 10404.305 1047.435 ;
    END
  END DIG_MON_SEL[232]
  PIN MASKD[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10402.345 1046.435 10402.625 1047.435 ;
    END
  END MASKD[231]
  PIN Data_COMP[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10390.025 1046.435 10390.305 1047.435 ;
    END
  END Data_COMP[71]
  PIN Data_COMP[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10388.905 1046.435 10389.185 1047.435 ;
    END
  END Data_COMP[82]
  PIN Data_COMP[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10387.785 1046.435 10388.065 1047.435 ;
    END
  END Data_COMP[76]
  PIN INJ_IN[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10382.465 1046.435 10382.745 1047.435 ;
    END
  END INJ_IN[231]
  PIN BcidMtx[695]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10380.225 1046.435 10380.505 1047.435 ;
    END
  END BcidMtx[695]
  PIN BcidMtx[693]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10379.105 1046.435 10379.385 1047.435 ;
    END
  END BcidMtx[693]
  PIN INJ_IN[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10349.705 1046.435 10349.985 1047.435 ;
    END
  END INJ_IN[230]
  PIN Data_COMP[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10348.025 1046.435 10348.305 1047.435 ;
    END
  END Data_COMP[65]
  PIN Data_COMP[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10346.905 1046.435 10347.185 1047.435 ;
    END
  END Data_COMP[78]
  PIN Data_COMP[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10344.665 1046.435 10344.945 1047.435 ;
    END
  END Data_COMP[74]
  PIN Data_COMP[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10343.545 1046.435 10343.825 1047.435 ;
    END
  END Data_COMP[63]
  PIN MASKV[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10342.425 1046.435 10342.705 1047.435 ;
    END
  END MASKV[230]
  PIN DIG_MON_SEL[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10325.625 1046.435 10325.905 1047.435 ;
    END
  END DIG_MON_SEL[230]
  PIN MASKD[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10323.945 1046.435 10324.225 1047.435 ;
    END
  END MASKD[229]
  PIN INJ_ROW[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10321.705 1046.435 10321.985 1047.435 ;
    END
  END INJ_ROW[114]
  PIN Data_COMP[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10318.905 1046.435 10319.185 1047.435 ;
    END
  END Data_COMP[61]
  PIN Data_COMP[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10317.785 1046.435 10318.065 1047.435 ;
    END
  END Data_COMP[55]
  PIN INJ_IN[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9194.425 1046.435 9194.705 1047.435 ;
    END
  END INJ_IN[201]
  PIN BcidMtx[604]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9152.425 1046.435 9152.705 1047.435 ;
    END
  END BcidMtx[604]
  PIN Read_PMOS[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9150.745 1046.435 9151.025 1047.435 ;
    END
  END Read_PMOS[44]
  PIN BcidMtx[600]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9149.065 1046.435 9149.345 1047.435 ;
    END
  END BcidMtx[600]
  PIN Data_PMOS[926]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9146.265 1046.435 9146.545 1047.435 ;
    END
  END Data_PMOS[926]
  PIN Data_PMOS[934]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9144.585 1046.435 9144.865 1047.435 ;
    END
  END Data_PMOS[934]
  PIN Data_PMOS[935]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9142.905 1046.435 9143.185 1047.435 ;
    END
  END Data_PMOS[935]
  PIN Data_PMOS[941]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9141.225 1046.435 9141.505 1047.435 ;
    END
  END Data_PMOS[941]
  PIN MASKD[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9131.145 1046.435 9131.425 1047.435 ;
    END
  END MASKD[200]
  PIN DIG_MON_SEL[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9128.345 1046.435 9128.625 1047.435 ;
    END
  END DIG_MON_SEL[200]
  PIN DIG_MON_SEL[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18803.465 1046.435 18803.745 1047.435 ;
    END
  END DIG_MON_SEL[441]
  PIN MASKD[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18802.345 1046.435 18802.625 1047.435 ;
    END
  END MASKD[441]
  PIN Data_PMOS[911]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9120.785 1046.435 9121.065 1047.435 ;
    END
  END Data_PMOS[911]
  PIN Data_PMOS[908]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9119.105 1046.435 9119.385 1047.435 ;
    END
  END Data_PMOS[908]
  PIN Data_PMOS[917]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9091.945 1046.435 9092.225 1047.435 ;
    END
  END Data_PMOS[917]
  PIN INJ_IN[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9089.705 1046.435 9089.985 1047.435 ;
    END
  END INJ_IN[199]
  PIN BcidMtx[598]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9086.905 1046.435 9087.185 1047.435 ;
    END
  END BcidMtx[598]
  PIN Read_PMOS[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9085.225 1046.435 9085.505 1047.435 ;
    END
  END Read_PMOS[43]
  PIN BcidMtx[594]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9083.545 1046.435 9083.825 1047.435 ;
    END
  END BcidMtx[594]
  PIN Data_PMOS[905]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9080.745 1046.435 9081.025 1047.435 ;
    END
  END Data_PMOS[905]
  PIN Data_PMOS[913]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9066.185 1046.435 9066.465 1047.435 ;
    END
  END Data_PMOS[913]
  PIN Data_PMOS[914]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9064.505 1046.435 9064.785 1047.435 ;
    END
  END Data_PMOS[914]
  PIN Data_PMOS[920]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9062.825 1046.435 9063.105 1047.435 ;
    END
  END Data_PMOS[920]
  PIN MASKD[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9061.145 1046.435 9061.425 1047.435 ;
    END
  END MASKD[198]
  PIN DIG_MON_SEL[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9058.345 1046.435 9058.625 1047.435 ;
    END
  END DIG_MON_SEL[198]
  PIN DIG_MON_PMOS[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9055.545 1046.435 9055.825 1047.435 ;
    END
  END DIG_MON_PMOS[85]
  PIN Data_PMOS[900]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9013.545 1046.435 9013.825 1047.435 ;
    END
  END Data_PMOS[900]
  PIN Data_PMOS[901]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9011.865 1046.435 9012.145 1047.435 ;
    END
  END Data_PMOS[901]
  PIN Data_PMOS[902]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9010.185 1046.435 9010.465 1047.435 ;
    END
  END Data_PMOS[902]
  PIN INJ_IN[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9007.385 1046.435 9007.665 1047.435 ;
    END
  END INJ_IN[197]
  PIN BcidMtx[593]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9005.145 1046.435 9005.425 1047.435 ;
    END
  END BcidMtx[593]
  PIN FREEZE_PMOS[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9003.465 1046.435 9003.745 1047.435 ;
    END
  END FREEZE_PMOS[42]
  PIN BcidMtx[588]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9001.225 1046.435 9001.505 1047.435 ;
    END
  END BcidMtx[588]
  PIN Data_PMOS[885]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8990.585 1046.435 8990.865 1047.435 ;
    END
  END Data_PMOS[885]
  PIN Data_PMOS[897]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8988.905 1046.435 8989.185 1047.435 ;
    END
  END Data_PMOS[897]
  PIN Data_PMOS[893]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8986.665 1046.435 8986.945 1047.435 ;
    END
  END Data_PMOS[893]
  PIN Data_PMOS[882]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8985.545 1046.435 8985.825 1047.435 ;
    END
  END Data_PMOS[882]
  PIN MASKH[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8981.905 1046.435 8982.185 1047.435 ;
    END
  END MASKH[98]
  PIN DIG_MON_SEL[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8978.545 1046.435 8978.825 1047.435 ;
    END
  END DIG_MON_SEL[196]
  PIN DIG_MON_SEL[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10071.945 1046.435 10072.225 1047.435 ;
    END
  END DIG_MON_SEL[223]
  PIN DIG_MON_PMOS[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10069.705 1046.435 10069.985 1047.435 ;
    END
  END DIG_MON_PMOS[111]
  PIN Data_PMOS[1163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10066.905 1046.435 10067.185 1047.435 ;
    END
  END Data_PMOS[1163]
  PIN Data_PMOS[1174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10065.785 1046.435 10066.065 1047.435 ;
    END
  END Data_PMOS[1174]
  PIN Data_PMOS[1175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10064.105 1046.435 10064.385 1047.435 ;
    END
  END Data_PMOS[1175]
  PIN Data_PMOS[1161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10062.425 1046.435 10062.705 1047.435 ;
    END
  END Data_PMOS[1161]
  PIN BcidMtx[671]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10045.625 1046.435 10045.905 1047.435 ;
    END
  END BcidMtx[671]
  PIN FREEZE_PMOS[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10043.945 1046.435 10044.225 1047.435 ;
    END
  END FREEZE_PMOS[55]
  PIN BcidMtx[666]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10041.705 1046.435 10041.985 1047.435 ;
    END
  END BcidMtx[666]
  PIN Data_PMOS[1158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10039.465 1046.435 10039.745 1047.435 ;
    END
  END Data_PMOS[1158]
  PIN Data_PMOS[1170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10037.785 1046.435 10038.065 1047.435 ;
    END
  END Data_PMOS[1170]
  PIN Data_PMOS[1171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10036.105 1046.435 10036.385 1047.435 ;
    END
  END Data_PMOS[1171]
  PIN Data_PMOS[1155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10034.425 1046.435 10034.705 1047.435 ;
    END
  END Data_PMOS[1155]
  PIN MASKH[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9994.105 1046.435 9994.385 1047.435 ;
    END
  END MASKH[111]
  PIN MASKD[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9989.065 1046.435 9989.345 1047.435 ;
    END
  END MASKD[221]
  PIN MASKV[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9986.265 1046.435 9986.545 1047.435 ;
    END
  END MASKV[221]
  PIN Data_PMOS[1142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9985.145 1046.435 9985.425 1047.435 ;
    END
  END Data_PMOS[1142]
  PIN Data_PMOS[1139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9983.465 1046.435 9983.745 1047.435 ;
    END
  END Data_PMOS[1139]
  PIN Data_PMOS[1148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9981.785 1046.435 9982.065 1047.435 ;
    END
  END Data_PMOS[1148]
  PIN nTOK_PMOS[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9970.025 1046.435 9970.305 1047.435 ;
    END
  END nTOK_PMOS[54]
  PIN BcidMtx[664]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9968.345 1046.435 9968.625 1047.435 ;
    END
  END BcidMtx[664]
  PIN Read_PMOS[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9966.665 1046.435 9966.945 1047.435 ;
    END
  END Read_PMOS[54]
  PIN INJ_IN[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9961.905 1046.435 9962.185 1047.435 ;
    END
  END INJ_IN[220]
  PIN Data_PMOS[1136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9960.225 1046.435 9960.505 1047.435 ;
    END
  END Data_PMOS[1136]
  PIN Data_PMOS[1144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9958.545 1046.435 9958.825 1047.435 ;
    END
  END Data_PMOS[1144]
  PIN Data_PMOS[1135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9930.825 1046.435 9931.105 1047.435 ;
    END
  END Data_PMOS[1135]
  PIN Data_PMOS[1151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9929.705 1046.435 9929.985 1047.435 ;
    END
  END Data_PMOS[1151]
  PIN MASKD[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9928.025 1046.435 9928.305 1047.435 ;
    END
  END MASKD[220]
  PIN DIG_MON_SEL[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9924.665 1046.435 9924.945 1047.435 ;
    END
  END DIG_MON_SEL[219]
  PIN DIG_MON_PMOS[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9922.425 1046.435 9922.705 1047.435 ;
    END
  END DIG_MON_PMOS[107]
  PIN Data_PMOS[1131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9920.185 1046.435 9920.465 1047.435 ;
    END
  END Data_PMOS[1131]
  PIN Data_PMOS[1126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9904.505 1046.435 9904.785 1047.435 ;
    END
  END Data_PMOS[1126]
  PIN Data_PMOS[1133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9903.945 1046.435 9904.225 1047.435 ;
    END
  END Data_PMOS[1133]
  PIN Data_PMOS[1119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9902.265 1046.435 9902.545 1047.435 ;
    END
  END Data_PMOS[1119]
  PIN BcidMtx[658]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9898.345 1046.435 9898.625 1047.435 ;
    END
  END BcidMtx[658]
  PIN Read_PMOS[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9896.665 1046.435 9896.945 1047.435 ;
    END
  END Read_PMOS[53]
  PIN BcidMtx[655]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9895.545 1046.435 9895.825 1047.435 ;
    END
  END BcidMtx[655]
  PIN Data_PMOS[1116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9854.105 1046.435 9854.385 1047.435 ;
    END
  END Data_PMOS[1116]
  PIN Data_PMOS[1128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9852.425 1046.435 9852.705 1047.435 ;
    END
  END Data_PMOS[1128]
  PIN Data_PMOS[1129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9850.745 1046.435 9851.025 1047.435 ;
    END
  END Data_PMOS[1129]
  PIN Data_PMOS[1113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9849.065 1046.435 9849.345 1047.435 ;
    END
  END Data_PMOS[1113]
  PIN MASKH[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9847.385 1046.435 9847.665 1047.435 ;
    END
  END MASKH[109]
  PIN MASKD[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9842.345 1046.435 9842.625 1047.435 ;
    END
  END MASKD[217]
  PIN MASKV[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9831.145 1046.435 9831.425 1047.435 ;
    END
  END MASKV[217]
  PIN Data_PMOS[1104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9829.465 1046.435 9829.745 1047.435 ;
    END
  END Data_PMOS[1104]
  PIN Data_PMOS[1112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9827.225 1046.435 9827.505 1047.435 ;
    END
  END Data_PMOS[1112]
  PIN Data_PMOS[1099]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9826.105 1046.435 9826.385 1047.435 ;
    END
  END Data_PMOS[1099]
  PIN nTOK_PMOS[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9821.345 1046.435 9821.625 1047.435 ;
    END
  END nTOK_PMOS[52]
  PIN BcidMtx[651]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9819.105 1046.435 9819.385 1047.435 ;
    END
  END BcidMtx[651]
  PIN BcidMtx[649]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9791.385 1046.435 9791.665 1047.435 ;
    END
  END BcidMtx[649]
  PIN Data_PMOS[1095]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9788.585 1046.435 9788.865 1047.435 ;
    END
  END Data_PMOS[1095]
  PIN Data_PMOS[1107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9786.905 1046.435 9787.185 1047.435 ;
    END
  END Data_PMOS[1107]
  PIN Data_PMOS[1108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9785.225 1046.435 9785.505 1047.435 ;
    END
  END Data_PMOS[1108]
  PIN Data_PMOS[1092]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9783.545 1046.435 9783.825 1047.435 ;
    END
  END Data_PMOS[1092]
  PIN MASKH[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9781.865 1046.435 9782.145 1047.435 ;
    END
  END MASKH[108]
  PIN MASKD[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9781.305 1046.435 9781.585 1047.435 ;
    END
  END MASKD[216]
  PIN DIG_MON_SEL[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9765.625 1046.435 9765.905 1047.435 ;
    END
  END DIG_MON_SEL[216]
  PIN DIG_MON_PMOS[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9762.825 1046.435 9763.105 1047.435 ;
    END
  END DIG_MON_PMOS[103]
  PIN Data_PMOS[1089]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9760.585 1046.435 9760.865 1047.435 ;
    END
  END Data_PMOS[1089]
  PIN Data_PMOS[1090]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9758.905 1046.435 9759.185 1047.435 ;
    END
  END Data_PMOS[1090]
  PIN Data_PMOS[1091]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9757.225 1046.435 9757.505 1047.435 ;
    END
  END Data_PMOS[1091]
  PIN nTOK_PMOS[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8034.105 1046.435 8034.385 1047.435 ;
    END
  END nTOK_PMOS[30]
  PIN FREEZE_PMOS[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8031.305 1046.435 8031.585 1047.435 ;
    END
  END FREEZE_PMOS[30]
  PIN BcidMtx[518]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8030.185 1046.435 8030.465 1047.435 ;
    END
  END BcidMtx[518]
  PIN INJ_IN[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8027.945 1046.435 8028.225 1047.435 ;
    END
  END INJ_IN[172]
  PIN Data_PMOS[645]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8025.145 1046.435 8025.425 1047.435 ;
    END
  END Data_PMOS[645]
  PIN Data_PMOS[634]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8024.025 1046.435 8024.305 1047.435 ;
    END
  END Data_PMOS[634]
  PIN Data_PMOS[631]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8022.345 1046.435 8022.625 1047.435 ;
    END
  END Data_PMOS[631]
  PIN MASKH[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8011.705 1046.435 8011.985 1047.435 ;
    END
  END MASKH[86]
  PIN DIG_MON_PMOS[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8010.025 1046.435 8010.305 1047.435 ;
    END
  END DIG_MON_PMOS[60]
  PIN DIG_MON_SEL[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8007.785 1046.435 8008.065 1047.435 ;
    END
  END DIG_MON_SEL[171]
  PIN INJ_ROW[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8002.465 1046.435 8002.745 1047.435 ;
    END
  END INJ_ROW[85]
  PIN Data_PMOS[627]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8001.345 1046.435 8001.625 1047.435 ;
    END
  END Data_PMOS[627]
  PIN Data_PMOS[621]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8000.225 1046.435 8000.505 1047.435 ;
    END
  END Data_PMOS[621]
  PIN Data_PMOS[623]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7971.945 1046.435 7972.225 1047.435 ;
    END
  END Data_PMOS[623]
  PIN Data_PMOS[615]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7970.825 1046.435 7971.105 1047.435 ;
    END
  END Data_PMOS[615]
  PIN nTOK_PMOS[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7968.585 1046.435 7968.865 1047.435 ;
    END
  END nTOK_PMOS[29]
  PIN BcidMtx[514]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7966.905 1046.435 7967.185 1047.435 ;
    END
  END BcidMtx[514]
  PIN BcidMtx[512]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7964.665 1046.435 7964.945 1047.435 ;
    END
  END BcidMtx[512]
  PIN INJ_IN[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7962.425 1046.435 7962.705 1047.435 ;
    END
  END INJ_IN[170]
  PIN Data_PMOS[618]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7960.185 1046.435 7960.465 1047.435 ;
    END
  END Data_PMOS[618]
  PIN Data_PMOS[613]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7945.625 1046.435 7945.905 1047.435 ;
    END
  END Data_PMOS[613]
  PIN Data_PMOS[610]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7943.945 1046.435 7944.225 1047.435 ;
    END
  END Data_PMOS[610]
  PIN MASKV[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7942.265 1046.435 7942.545 1047.435 ;
    END
  END MASKV[170]
  PIN DIG_MON_PMOS[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7940.025 1046.435 7940.305 1047.435 ;
    END
  END DIG_MON_PMOS[58]
  PIN INJ_ROW[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7934.425 1046.435 7934.705 1047.435 ;
    END
  END INJ_ROW[84]
  PIN Data_PMOS[596]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7892.985 1046.435 7893.265 1047.435 ;
    END
  END Data_PMOS[596]
  PIN Data_PMOS[600]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7892.425 1046.435 7892.705 1047.435 ;
    END
  END Data_PMOS[600]
  PIN Data_PMOS[601]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7890.745 1046.435 7891.025 1047.435 ;
    END
  END Data_PMOS[601]
  PIN INJ_IN[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7887.385 1046.435 7887.665 1047.435 ;
    END
  END INJ_IN[169]
  PIN nTOK_PMOS[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7886.265 1046.435 7886.545 1047.435 ;
    END
  END nTOK_PMOS[28]
  PIN BcidMtx[508]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7884.585 1046.435 7884.865 1047.435 ;
    END
  END BcidMtx[508]
  PIN BcidMtx[505]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7881.785 1046.435 7882.065 1047.435 ;
    END
  END BcidMtx[505]
  PIN BcidMtx[504]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7881.225 1046.435 7881.505 1047.435 ;
    END
  END BcidMtx[504]
  PIN Data_PMOS[590]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7870.025 1046.435 7870.305 1047.435 ;
    END
  END Data_PMOS[590]
  PIN Data_PMOS[598]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7868.345 1046.435 7868.625 1047.435 ;
    END
  END Data_PMOS[598]
  PIN Data_PMOS[599]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7866.665 1046.435 7866.945 1047.435 ;
    END
  END Data_PMOS[599]
  PIN Data_PMOS[605]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7864.985 1046.435 7865.265 1047.435 ;
    END
  END Data_PMOS[605]
  PIN MASKD[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7861.345 1046.435 7861.625 1047.435 ;
    END
  END MASKD[168]
  PIN DIG_MON_SEL[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7858.545 1046.435 7858.825 1047.435 ;
    END
  END DIG_MON_SEL[168]
  PIN FREEZE_PMOS[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8113.065 1046.435 8113.345 1047.435 ;
    END
  END FREEZE_PMOS[31]
  PIN MASKV[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8948.025 1046.435 8948.305 1047.435 ;
    END
  END MASKV[195]
  PIN Data_PMOS[873]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8946.345 1046.435 8946.625 1047.435 ;
    END
  END Data_PMOS[873]
  PIN Data_PMOS[874]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8944.665 1046.435 8944.945 1047.435 ;
    END
  END Data_PMOS[874]
  PIN Data_PMOS[868]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8942.985 1046.435 8943.265 1047.435 ;
    END
  END Data_PMOS[868]
  PIN nTOK_PMOS[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8940.185 1046.435 8940.465 1047.435 ;
    END
  END nTOK_PMOS[41]
  PIN BcidMtx[587]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8925.625 1046.435 8925.905 1047.435 ;
    END
  END BcidMtx[587]
  PIN BcidMtx[584]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8922.825 1046.435 8923.105 1047.435 ;
    END
  END BcidMtx[584]
  PIN INJ_IN[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8920.585 1046.435 8920.865 1047.435 ;
    END
  END INJ_IN[194]
  PIN Data_PMOS[864]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8919.465 1046.435 8919.745 1047.435 ;
    END
  END Data_PMOS[864]
  PIN Data_PMOS[865]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8916.665 1046.435 8916.945 1047.435 ;
    END
  END Data_PMOS[865]
  PIN Data_PMOS[862]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8914.985 1046.435 8915.265 1047.435 ;
    END
  END Data_PMOS[862]
  PIN MASKV[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8874.665 1046.435 8874.945 1047.435 ;
    END
  END MASKV[194]
  PIN DIG_MON_PMOS[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8872.425 1046.435 8872.705 1047.435 ;
    END
  END DIG_MON_PMOS[82]
  PIN DIG_MON_SEL[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8870.185 1046.435 8870.465 1047.435 ;
    END
  END DIG_MON_SEL[193]
  PIN INJ_ROW[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8866.825 1046.435 8867.105 1047.435 ;
    END
  END INJ_ROW[96]
  PIN Data_PMOS[848]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8865.145 1046.435 8865.425 1047.435 ;
    END
  END Data_PMOS[848]
  PIN Data_PMOS[845]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8863.465 1046.435 8863.745 1047.435 ;
    END
  END Data_PMOS[845]
  PIN Data_PMOS[853]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8862.905 1046.435 8863.185 1047.435 ;
    END
  END Data_PMOS[853]
  PIN INJ_IN[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8851.145 1046.435 8851.425 1047.435 ;
    END
  END INJ_IN[193]
  PIN BcidMtx[581]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8848.905 1046.435 8849.185 1047.435 ;
    END
  END BcidMtx[581]
  PIN FREEZE_PMOS[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8847.225 1046.435 8847.505 1047.435 ;
    END
  END FREEZE_PMOS[40]
  PIN BcidMtx[577]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8845.545 1046.435 8845.825 1047.435 ;
    END
  END BcidMtx[577]
  PIN Data_PMOS[843]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8840.785 1046.435 8841.065 1047.435 ;
    END
  END Data_PMOS[843]
  PIN Data_PMOS[855]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8839.105 1046.435 8839.385 1047.435 ;
    END
  END Data_PMOS[855]
  PIN Data_PMOS[856]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8811.945 1046.435 8812.225 1047.435 ;
    END
  END Data_PMOS[856]
  PIN Data_PMOS[840]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8810.265 1046.435 8810.545 1047.435 ;
    END
  END Data_PMOS[840]
  PIN MASKH[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8808.585 1046.435 8808.865 1047.435 ;
    END
  END MASKH[96]
  PIN MASKD[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8803.545 1046.435 8803.825 1047.435 ;
    END
  END MASKD[191]
  PIN DIG_MON_PMOS[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8802.425 1046.435 8802.705 1047.435 ;
    END
  END DIG_MON_PMOS[79]
  PIN Data_PMOS[831]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8786.185 1046.435 8786.465 1047.435 ;
    END
  END Data_PMOS[831]
  PIN Data_PMOS[832]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8784.505 1046.435 8784.785 1047.435 ;
    END
  END Data_PMOS[832]
  PIN Data_PMOS[839]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8783.945 1046.435 8784.225 1047.435 ;
    END
  END Data_PMOS[839]
  PIN nTOK_PMOS[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8780.025 1046.435 8780.305 1047.435 ;
    END
  END nTOK_PMOS[39]
  PIN BcidMtx[573]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8777.785 1046.435 8778.065 1047.435 ;
    END
  END BcidMtx[573]
  PIN BcidMtx[572]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8776.105 1046.435 8776.385 1047.435 ;
    END
  END BcidMtx[572]
  PIN INJ_IN[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8773.865 1046.435 8774.145 1047.435 ;
    END
  END INJ_IN[190]
  PIN Data_PMOS[828]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8732.985 1046.435 8733.265 1047.435 ;
    END
  END Data_PMOS[828]
  PIN Data_PMOS[823]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8731.305 1046.435 8731.585 1047.435 ;
    END
  END Data_PMOS[823]
  PIN Data_PMOS[820]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8729.625 1046.435 8729.905 1047.435 ;
    END
  END Data_PMOS[820]
  PIN MASKV[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8727.945 1046.435 8728.225 1047.435 ;
    END
  END MASKV[190]
  PIN DIG_MON_PMOS[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8725.705 1046.435 8725.985 1047.435 ;
    END
  END DIG_MON_PMOS[78]
  PIN DIG_MON_SEL[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8723.465 1046.435 8723.745 1047.435 ;
    END
  END DIG_MON_SEL[189]
  PIN INJ_ROW[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8711.705 1046.435 8711.985 1047.435 ;
    END
  END INJ_ROW[94]
  PIN Data_PMOS[806]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8710.025 1046.435 8710.305 1047.435 ;
    END
  END Data_PMOS[806]
  PIN Data_PMOS[803]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8708.345 1046.435 8708.625 1047.435 ;
    END
  END Data_PMOS[803]
  PIN Data_PMOS[812]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8706.665 1046.435 8706.945 1047.435 ;
    END
  END Data_PMOS[812]
  PIN INJ_IN[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8702.465 1046.435 8702.745 1047.435 ;
    END
  END INJ_IN[189]
  PIN BcidMtx[568]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8699.665 1046.435 8699.945 1047.435 ;
    END
  END BcidMtx[568]
  PIN BcidMtx[566]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8671.945 1046.435 8672.225 1047.435 ;
    END
  END BcidMtx[566]
  PIN BcidMtx[565]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8671.385 1046.435 8671.665 1047.435 ;
    END
  END BcidMtx[565]
  PIN Data_PMOS[807]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8667.465 1046.435 8667.745 1047.435 ;
    END
  END Data_PMOS[807]
  PIN Data_PMOS[802]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8665.785 1046.435 8666.065 1047.435 ;
    END
  END Data_PMOS[802]
  PIN Data_PMOS[809]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8664.665 1046.435 8664.945 1047.435 ;
    END
  END Data_PMOS[809]
  PIN MASKH[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8661.865 1046.435 8662.145 1047.435 ;
    END
  END MASKH[94]
  PIN DIG_MON_PMOS[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8660.185 1046.435 8660.465 1047.435 ;
    END
  END DIG_MON_PMOS[76]
  PIN DIG_MON_SEL[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8645.625 1046.435 8645.905 1047.435 ;
    END
  END DIG_MON_SEL[188]
  PIN MASKV[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8641.145 1046.435 8641.425 1047.435 ;
    END
  END MASKV[187]
  PIN Data_PMOS[795]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8640.585 1046.435 8640.865 1047.435 ;
    END
  END Data_PMOS[795]
  PIN Data_PMOS[796]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8638.905 1046.435 8639.185 1047.435 ;
    END
  END Data_PMOS[796]
  PIN Data_PMOS[797]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8637.225 1046.435 8637.505 1047.435 ;
    END
  END Data_PMOS[797]
  PIN Data_PMOS[783]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8635.545 1046.435 8635.825 1047.435 ;
    END
  END Data_PMOS[783]
  PIN BcidMtx[563]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8592.985 1046.435 8593.265 1047.435 ;
    END
  END BcidMtx[563]
  PIN FREEZE_PMOS[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8591.305 1046.435 8591.585 1047.435 ;
    END
  END FREEZE_PMOS[37]
  PIN BcidMtx[559]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8589.625 1046.435 8589.905 1047.435 ;
    END
  END BcidMtx[559]
  PIN INJ_IN[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8587.945 1046.435 8588.225 1047.435 ;
    END
  END INJ_IN[186]
  PIN Data_PMOS[787]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8584.585 1046.435 8584.865 1047.435 ;
    END
  END Data_PMOS[787]
  PIN Data_PMOS[793]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8583.465 1046.435 8583.745 1047.435 ;
    END
  END Data_PMOS[793]
  PIN Data_PMOS[794]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8581.225 1046.435 8581.505 1047.435 ;
    END
  END Data_PMOS[794]
  PIN MASKD[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8571.145 1046.435 8571.425 1047.435 ;
    END
  END MASKD[186]
  PIN DIG_MON_SEL[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8568.345 1046.435 8568.625 1047.435 ;
    END
  END DIG_MON_SEL[186]
  PIN INJ_ROW[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8562.465 1046.435 8562.745 1047.435 ;
    END
  END INJ_ROW[92]
  PIN Data_PMOS[764]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8560.785 1046.435 8561.065 1047.435 ;
    END
  END Data_PMOS[764]
  PIN Data_PMOS[775]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8559.665 1046.435 8559.945 1047.435 ;
    END
  END Data_PMOS[775]
  PIN Data_PMOS[769]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8533.065 1046.435 8533.345 1047.435 ;
    END
  END Data_PMOS[769]
  PIN Data_PMOS[762]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8530.825 1046.435 8531.105 1047.435 ;
    END
  END Data_PMOS[762]
  PIN nTOK_PMOS[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8528.585 1046.435 8528.865 1047.435 ;
    END
  END nTOK_PMOS[36]
  PIN BcidMtx[556]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8526.905 1046.435 8527.185 1047.435 ;
    END
  END BcidMtx[556]
  PIN BcidMtx[553]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8524.105 1046.435 8524.385 1047.435 ;
    END
  END BcidMtx[553]
  PIN Data_PMOS[759]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8521.305 1046.435 8521.585 1047.435 ;
    END
  END Data_PMOS[759]
  PIN Data_PMOS[771]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8506.745 1046.435 8507.025 1047.435 ;
    END
  END Data_PMOS[771]
  PIN Data_PMOS[772]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8505.065 1046.435 8505.345 1047.435 ;
    END
  END Data_PMOS[772]
  PIN Data_PMOS[756]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8503.385 1046.435 8503.665 1047.435 ;
    END
  END Data_PMOS[756]
  PIN MASKD[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8501.145 1046.435 8501.425 1047.435 ;
    END
  END MASKD[184]
  PIN MASKD[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8496.665 1046.435 8496.945 1047.435 ;
    END
  END MASKD[183]
  PIN INJ_ROW[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8494.425 1046.435 8494.705 1047.435 ;
    END
  END INJ_ROW[91]
  PIN Data_PMOS[747]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8452.425 1046.435 8452.705 1047.435 ;
    END
  END Data_PMOS[747]
  PIN Data_PMOS[748]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8450.745 1046.435 8451.025 1047.435 ;
    END
  END Data_PMOS[748]
  PIN Data_PMOS[749]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8449.625 1046.435 8449.905 1047.435 ;
    END
  END Data_PMOS[749]
  PIN Data_PMOS[741]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8448.505 1046.435 8448.785 1047.435 ;
    END
  END Data_PMOS[741]
  PIN BcidMtx[551]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8445.145 1046.435 8445.425 1047.435 ;
    END
  END BcidMtx[551]
  PIN BcidMtx[549]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8444.025 1046.435 8444.305 1047.435 ;
    END
  END BcidMtx[549]
  PIN BcidMtx[547]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8441.785 1046.435 8442.065 1047.435 ;
    END
  END BcidMtx[547]
  PIN Data_PMOS[738]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8430.585 1046.435 8430.865 1047.435 ;
    END
  END Data_PMOS[738]
  PIN Data_PMOS[744]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8429.465 1046.435 8429.745 1047.435 ;
    END
  END Data_PMOS[744]
  PIN Data_PMOS[751]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8427.225 1046.435 8427.505 1047.435 ;
    END
  END Data_PMOS[751]
  PIN Data_PMOS[735]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8425.545 1046.435 8425.825 1047.435 ;
    END
  END Data_PMOS[735]
  PIN MASKV[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8422.465 1046.435 8422.745 1047.435 ;
    END
  END MASKV[182]
  PIN DIG_MON_PMOS[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8420.225 1046.435 8420.505 1047.435 ;
    END
  END DIG_MON_PMOS[70]
  PIN FREEZE_PMOS[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8673.065 1046.435 8673.345 1047.435 ;
    END
  END FREEZE_PMOS[38]
  PIN MASKV[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9508.025 1046.435 9508.305 1047.435 ;
    END
  END MASKV[209]
  PIN Data_PMOS[1016]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9506.905 1046.435 9507.185 1047.435 ;
    END
  END Data_PMOS[1016]
  PIN Data_PMOS[1013]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9505.225 1046.435 9505.505 1047.435 ;
    END
  END Data_PMOS[1013]
  PIN Data_PMOS[1022]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9503.545 1046.435 9503.825 1047.435 ;
    END
  END Data_PMOS[1022]
  PIN INJ_IN[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9501.305 1046.435 9501.585 1047.435 ;
    END
  END INJ_IN[209]
  PIN BcidMtx[628]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9485.065 1046.435 9485.345 1047.435 ;
    END
  END BcidMtx[628]
  PIN FREEZE_PMOS[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9483.945 1046.435 9484.225 1047.435 ;
    END
  END FREEZE_PMOS[48]
  PIN BcidMtx[624]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9481.705 1046.435 9481.985 1047.435 ;
    END
  END BcidMtx[624]
  PIN Data_PMOS[1010]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9478.905 1046.435 9479.185 1047.435 ;
    END
  END Data_PMOS[1010]
  PIN Data_PMOS[1023]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9477.785 1046.435 9478.065 1047.435 ;
    END
  END Data_PMOS[1023]
  PIN Data_PMOS[1019]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9475.545 1046.435 9475.825 1047.435 ;
    END
  END Data_PMOS[1019]
  PIN Data_PMOS[1025]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9473.865 1046.435 9474.145 1047.435 ;
    END
  END Data_PMOS[1025]
  PIN DIG_MON_PMOS[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9432.425 1046.435 9432.705 1047.435 ;
    END
  END DIG_MON_PMOS[96]
  PIN DIG_MON_SEL[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9430.745 1046.435 9431.025 1047.435 ;
    END
  END DIG_MON_SEL[208]
  PIN DIG_MON_PMOS[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9427.945 1046.435 9428.225 1047.435 ;
    END
  END DIG_MON_PMOS[95]
  PIN MASKV[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9426.265 1046.435 9426.545 1047.435 ;
    END
  END MASKV[207]
  PIN Data_PMOS[1006]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9424.025 1046.435 9424.305 1047.435 ;
    END
  END Data_PMOS[1006]
  PIN Data_PMOS[1007]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9422.345 1046.435 9422.625 1047.435 ;
    END
  END Data_PMOS[1007]
  PIN Data_PMOS[1001]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9421.785 1046.435 9422.065 1047.435 ;
    END
  END Data_PMOS[1001]
  PIN nTOK_PMOS[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9410.025 1046.435 9410.305 1047.435 ;
    END
  END nTOK_PMOS[47]
  PIN BcidMtx[621]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9407.785 1046.435 9408.065 1047.435 ;
    END
  END BcidMtx[621]
  PIN BcidMtx[620]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9406.105 1046.435 9406.385 1047.435 ;
    END
  END BcidMtx[620]
  PIN INJ_IN[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9401.905 1046.435 9402.185 1047.435 ;
    END
  END INJ_IN[206]
  PIN Data_PMOS[996]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9399.665 1046.435 9399.945 1047.435 ;
    END
  END Data_PMOS[996]
  PIN Data_PMOS[997]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9398.545 1046.435 9398.825 1047.435 ;
    END
  END Data_PMOS[997]
  PIN Data_PMOS[998]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9371.385 1046.435 9371.665 1047.435 ;
    END
  END Data_PMOS[998]
  PIN Data_PMOS[1004]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9369.705 1046.435 9369.985 1047.435 ;
    END
  END Data_PMOS[1004]
  PIN MASKD[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9368.025 1046.435 9368.305 1047.435 ;
    END
  END MASKD[206]
  PIN DIG_MON_SEL[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9365.225 1046.435 9365.505 1047.435 ;
    END
  END DIG_MON_SEL[206]
  PIN DIG_MON_PMOS[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9362.425 1046.435 9362.705 1047.435 ;
    END
  END DIG_MON_PMOS[93]
  PIN Data_PMOS[984]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9360.185 1046.435 9360.465 1047.435 ;
    END
  END Data_PMOS[984]
  PIN Data_PMOS[985]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9345.625 1046.435 9345.905 1047.435 ;
    END
  END Data_PMOS[985]
  PIN Data_PMOS[986]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9343.945 1046.435 9344.225 1047.435 ;
    END
  END Data_PMOS[986]
  PIN Data_PMOS[972]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9342.265 1046.435 9342.545 1047.435 ;
    END
  END Data_PMOS[972]
  PIN BcidMtx[617]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9338.905 1046.435 9339.185 1047.435 ;
    END
  END BcidMtx[617]
  PIN FREEZE_PMOS[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9337.225 1046.435 9337.505 1047.435 ;
    END
  END FREEZE_PMOS[46]
  PIN BcidMtx[613]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9335.545 1046.435 9335.825 1047.435 ;
    END
  END BcidMtx[613]
  PIN Data_PMOS[969]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9294.105 1046.435 9294.385 1047.435 ;
    END
  END Data_PMOS[969]
  PIN Data_PMOS[981]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9292.425 1046.435 9292.705 1047.435 ;
    END
  END Data_PMOS[981]
  PIN Data_PMOS[982]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9290.745 1046.435 9291.025 1047.435 ;
    END
  END Data_PMOS[982]
  PIN Data_PMOS[966]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9289.065 1046.435 9289.345 1047.435 ;
    END
  END Data_PMOS[966]
  PIN MASKH[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9287.385 1046.435 9287.665 1047.435 ;
    END
  END MASKH[102]
  PIN MASKD[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9282.345 1046.435 9282.625 1047.435 ;
    END
  END MASKD[203]
  PIN MASKV[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9271.145 1046.435 9271.425 1047.435 ;
    END
  END MASKV[203]
  PIN Data_PMOS[957]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9269.465 1046.435 9269.745 1047.435 ;
    END
  END Data_PMOS[957]
  PIN Data_PMOS[958]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9267.785 1046.435 9268.065 1047.435 ;
    END
  END Data_PMOS[958]
  PIN Data_PMOS[952]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9266.105 1046.435 9266.385 1047.435 ;
    END
  END Data_PMOS[952]
  PIN nTOK_PMOS[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9261.345 1046.435 9261.625 1047.435 ;
    END
  END nTOK_PMOS[45]
  PIN BcidMtx[609]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9259.105 1046.435 9259.385 1047.435 ;
    END
  END BcidMtx[609]
  PIN BcidMtx[607]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9231.385 1046.435 9231.665 1047.435 ;
    END
  END BcidMtx[607]
  PIN Data_PMOS[948]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9228.585 1046.435 9228.865 1047.435 ;
    END
  END Data_PMOS[948]
  PIN Data_PMOS[960]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9226.905 1046.435 9227.185 1047.435 ;
    END
  END Data_PMOS[960]
  PIN Data_PMOS[961]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9225.225 1046.435 9225.505 1047.435 ;
    END
  END Data_PMOS[961]
  PIN Data_PMOS[945]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9223.545 1046.435 9223.825 1047.435 ;
    END
  END Data_PMOS[945]
  PIN MASKH[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9221.865 1046.435 9222.145 1047.435 ;
    END
  END MASKH[101]
  PIN DIG_MON_HV[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18805.705 1046.435 18805.985 1047.435 ;
    END
  END DIG_MON_HV[106]
  PIN INJ_ROW[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9201.705 1046.435 9201.985 1047.435 ;
    END
  END INJ_ROW[100]
  PIN Data_PMOS[932]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9200.025 1046.435 9200.305 1047.435 ;
    END
  END Data_PMOS[932]
  PIN Data_PMOS[929]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9198.345 1046.435 9198.625 1047.435 ;
    END
  END Data_PMOS[929]
  PIN Data_PMOS[938]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9196.665 1046.435 9196.945 1047.435 ;
    END
  END Data_PMOS[938]
  PIN BcidMtx[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6349.625 1046.435 6349.905 1047.435 ;
    END
  END BcidMtx[391]
  PIN Data_PMOS[192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6346.825 1046.435 6347.105 1047.435 ;
    END
  END Data_PMOS[192]
  PIN Data_PMOS[204]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6345.145 1046.435 6345.425 1047.435 ;
    END
  END Data_PMOS[204]
  PIN Data_PMOS[200]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6342.905 1046.435 6343.185 1047.435 ;
    END
  END Data_PMOS[200]
  PIN Data_PMOS[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6341.785 1046.435 6342.065 1047.435 ;
    END
  END Data_PMOS[189]
  PIN MASKH[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6331.705 1046.435 6331.985 1047.435 ;
    END
  END MASKH[65]
  PIN DIG_MON_SEL[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6328.345 1046.435 6328.625 1047.435 ;
    END
  END DIG_MON_SEL[130]
  PIN MASKD[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6326.665 1046.435 6326.945 1047.435 ;
    END
  END MASKD[129]
  PIN MASKV[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6321.905 1046.435 6322.185 1047.435 ;
    END
  END MASKV[129]
  PIN Data_PMOS[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6320.225 1046.435 6320.505 1047.435 ;
    END
  END Data_PMOS[180]
  PIN Data_PMOS[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6293.065 1046.435 6293.345 1047.435 ;
    END
  END Data_PMOS[181]
  PIN Data_PMOS[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6291.385 1046.435 6291.665 1047.435 ;
    END
  END Data_PMOS[175]
  PIN nTOK_PMOS[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6288.585 1046.435 6288.865 1047.435 ;
    END
  END nTOK_PMOS[8]
  PIN BcidMtx[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6286.345 1046.435 6286.625 1047.435 ;
    END
  END BcidMtx[387]
  PIN BcidMtx[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6284.665 1046.435 6284.945 1047.435 ;
    END
  END BcidMtx[386]
  PIN Data_PMOS[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6281.305 1046.435 6281.585 1047.435 ;
    END
  END Data_PMOS[171]
  PIN Data_PMOS[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6280.185 1046.435 6280.465 1047.435 ;
    END
  END Data_PMOS[177]
  PIN BcidMtx[1327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18855.545 1046.435 18855.825 1047.435 ;
    END
  END BcidMtx[1327]
  PIN Data_PMOS[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6263.945 1046.435 6264.225 1047.435 ;
    END
  END Data_PMOS[169]
  PIN Data_PMOS[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6262.825 1046.435 6263.105 1047.435 ;
    END
  END Data_PMOS[185]
  PIN MASKD[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6261.145 1046.435 6261.425 1047.435 ;
    END
  END MASKD[128]
  PIN DIG_MON_SEL[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6257.785 1046.435 6258.065 1047.435 ;
    END
  END DIG_MON_SEL[127]
  PIN DIG_MON_PMOS[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6255.545 1046.435 6255.825 1047.435 ;
    END
  END DIG_MON_PMOS[15]
  PIN Data_PMOS[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6213.545 1046.435 6213.825 1047.435 ;
    END
  END Data_PMOS[165]
  PIN Data_PMOS[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6211.305 1046.435 6211.585 1047.435 ;
    END
  END Data_PMOS[152]
  PIN Data_PMOS[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6210.185 1046.435 6210.465 1047.435 ;
    END
  END Data_PMOS[167]
  PIN Data_PMOS[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6208.505 1046.435 6208.785 1047.435 ;
    END
  END Data_PMOS[153]
  PIN BcidMtx[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6204.585 1046.435 6204.865 1047.435 ;
    END
  END BcidMtx[382]
  PIN FREEZE_PMOS[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6203.465 1046.435 6203.745 1047.435 ;
    END
  END FREEZE_PMOS[7]
  PIN BcidMtx[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6201.785 1046.435 6202.065 1047.435 ;
    END
  END BcidMtx[379]
  PIN Data_PMOS[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6190.585 1046.435 6190.865 1047.435 ;
    END
  END Data_PMOS[150]
  PIN Data_PMOS[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6188.905 1046.435 6189.185 1047.435 ;
    END
  END Data_PMOS[162]
  PIN Data_PMOS[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6187.225 1046.435 6187.505 1047.435 ;
    END
  END Data_PMOS[163]
  PIN Data_PMOS[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6185.545 1046.435 6185.825 1047.435 ;
    END
  END Data_PMOS[147]
  PIN Data_HV[1065]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18586.745 1046.435 18587.025 1047.435 ;
    END
  END Data_HV[1065]
  PIN MASKD[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6181.345 1046.435 6181.625 1047.435 ;
    END
  END MASKD[126]
  PIN FREEZE_PMOS[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6433.065 1046.435 6433.345 1047.435 ;
    END
  END FREEZE_PMOS[10]
  PIN MASKD[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7270.825 1046.435 7271.105 1047.435 ;
    END
  END MASKD[153]
  PIN MASKV[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7268.025 1046.435 7268.305 1047.435 ;
    END
  END MASKV[153]
  PIN Data_PMOS[439]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7265.785 1046.435 7266.065 1047.435 ;
    END
  END Data_PMOS[439]
  PIN Data_PMOS[433]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7264.665 1046.435 7264.945 1047.435 ;
    END
  END Data_PMOS[433]
  PIN Data_PMOS[427]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7262.985 1046.435 7263.265 1047.435 ;
    END
  END Data_PMOS[427]
  PIN nTOK_PMOS[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7260.185 1046.435 7260.465 1047.435 ;
    END
  END nTOK_PMOS[20]
  PIN BcidMtx[459]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7244.505 1046.435 7244.785 1047.435 ;
    END
  END BcidMtx[459]
  PIN BcidMtx[458]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7242.825 1046.435 7243.105 1047.435 ;
    END
  END BcidMtx[458]
  PIN Data_PMOS[423]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7239.465 1046.435 7239.745 1047.435 ;
    END
  END Data_PMOS[423]
  PIN Data_PMOS[429]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7238.345 1046.435 7238.625 1047.435 ;
    END
  END Data_PMOS[429]
  PIN Data_PMOS[424]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7236.665 1046.435 7236.945 1047.435 ;
    END
  END Data_PMOS[424]
  PIN Data_PMOS[420]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7234.425 1046.435 7234.705 1047.435 ;
    END
  END Data_PMOS[420]
  PIN MASKV[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7194.665 1046.435 7194.945 1047.435 ;
    END
  END MASKV[152]
  PIN DIG_MON_PMOS[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7192.425 1046.435 7192.705 1047.435 ;
    END
  END DIG_MON_PMOS[40]
  PIN DIG_MON_SEL[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7190.185 1046.435 7190.465 1047.435 ;
    END
  END DIG_MON_SEL[151]
  PIN INJ_ROW[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7186.825 1046.435 7187.105 1047.435 ;
    END
  END INJ_ROW[75]
  PIN Data_PMOS[407]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7185.145 1046.435 7185.425 1047.435 ;
    END
  END Data_PMOS[407]
  PIN Data_PMOS[412]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7182.905 1046.435 7183.185 1047.435 ;
    END
  END Data_PMOS[412]
  PIN Data_PMOS[413]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7181.785 1046.435 7182.065 1047.435 ;
    END
  END Data_PMOS[413]
  PIN INJ_IN[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7171.145 1046.435 7171.425 1047.435 ;
    END
  END INJ_IN[151]
  PIN BcidMtx[453]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7167.785 1046.435 7168.065 1047.435 ;
    END
  END BcidMtx[453]
  PIN Read_PMOS[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7166.665 1046.435 7166.945 1047.435 ;
    END
  END Read_PMOS[19]
  PIN BcidMtx[450]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7164.985 1046.435 7165.265 1047.435 ;
    END
  END BcidMtx[450]
  PIN Data_PMOS[408]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7159.665 1046.435 7159.945 1047.435 ;
    END
  END Data_PMOS[408]
  PIN Data_PMOS[409]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7158.545 1046.435 7158.825 1047.435 ;
    END
  END Data_PMOS[409]
  PIN Data_PMOS[399]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7130.265 1046.435 7130.545 1047.435 ;
    END
  END Data_PMOS[399]
  PIN Data_HV[1116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18814.105 1046.435 18814.385 1047.435 ;
    END
  END Data_HV[1116]
  PIN MASKH[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7128.585 1046.435 7128.865 1047.435 ;
    END
  END MASKH[75]
  PIN DIG_MON_PMOS[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7122.425 1046.435 7122.705 1047.435 ;
    END
  END DIG_MON_PMOS[37]
  PIN MASKV[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7120.745 1046.435 7121.025 1047.435 ;
    END
  END MASKV[149]
  PIN Data_PMOS[390]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7106.185 1046.435 7106.465 1047.435 ;
    END
  END Data_PMOS[390]
  PIN Data_PMOS[398]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7103.945 1046.435 7104.225 1047.435 ;
    END
  END Data_PMOS[398]
  PIN Data_PMOS[385]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7102.825 1046.435 7103.105 1047.435 ;
    END
  END Data_PMOS[385]
  PIN nTOK_PMOS[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7100.025 1046.435 7100.305 1047.435 ;
    END
  END nTOK_PMOS[18]
  PIN FREEZE_PMOS[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7097.225 1046.435 7097.505 1047.435 ;
    END
  END FREEZE_PMOS[18]
  PIN BcidMtx[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7096.105 1046.435 7096.385 1047.435 ;
    END
  END BcidMtx[446]
  PIN INJ_IN[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7093.865 1046.435 7094.145 1047.435 ;
    END
  END INJ_IN[148]
  PIN Data_PMOS[387]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7052.985 1046.435 7053.265 1047.435 ;
    END
  END Data_PMOS[387]
  PIN Data_PMOS[382]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7051.305 1046.435 7051.585 1047.435 ;
    END
  END Data_PMOS[382]
  PIN Data_PMOS[379]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7049.625 1046.435 7049.905 1047.435 ;
    END
  END Data_PMOS[379]
  PIN MASKH[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7047.385 1046.435 7047.665 1047.435 ;
    END
  END MASKH[74]
  PIN DIG_MON_PMOS[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7045.705 1046.435 7045.985 1047.435 ;
    END
  END DIG_MON_PMOS[36]
  PIN DIG_MON_SEL[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7043.465 1046.435 7043.745 1047.435 ;
    END
  END DIG_MON_SEL[147]
  PIN MASKV[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7031.145 1046.435 7031.425 1047.435 ;
    END
  END MASKV[147]
  PIN Data_PMOS[365]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7030.025 1046.435 7030.305 1047.435 ;
    END
  END Data_PMOS[365]
  PIN Data_PMOS[362]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7028.345 1046.435 7028.625 1047.435 ;
    END
  END Data_PMOS[362]
  PIN Data_PMOS[371]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7026.665 1046.435 7026.945 1047.435 ;
    END
  END Data_PMOS[371]
  PIN INJ_IN[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7022.465 1046.435 7022.745 1047.435 ;
    END
  END INJ_IN[147]
  PIN BcidMtx[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7019.665 1046.435 7019.945 1047.435 ;
    END
  END BcidMtx[442]
  PIN BcidMtx[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6991.385 1046.435 6991.665 1047.435 ;
    END
  END BcidMtx[439]
  PIN INJ_IN[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6989.705 1046.435 6989.985 1047.435 ;
    END
  END INJ_IN[146]
  PIN Data_PMOS[366]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6987.465 1046.435 6987.745 1047.435 ;
    END
  END Data_PMOS[366]
  PIN Data_PMOS[373]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6985.225 1046.435 6985.505 1047.435 ;
    END
  END Data_PMOS[373]
  PIN Data_PMOS[358]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6984.105 1046.435 6984.385 1047.435 ;
    END
  END Data_PMOS[358]
  PIN MASKV[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6982.425 1046.435 6982.705 1047.435 ;
    END
  END MASKV[146]
  PIN DIG_MON_SEL[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6965.065 1046.435 6965.345 1047.435 ;
    END
  END DIG_MON_SEL[145]
  PIN INJ_ROW[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6961.705 1046.435 6961.985 1047.435 ;
    END
  END INJ_ROW[72]
  PIN Data_PMOS[348]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6959.465 1046.435 6959.745 1047.435 ;
    END
  END Data_PMOS[348]
  PIN Data_PMOS[341]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6958.345 1046.435 6958.625 1047.435 ;
    END
  END Data_PMOS[341]
  PIN Data_PMOS[350]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6956.665 1046.435 6956.945 1047.435 ;
    END
  END Data_PMOS[350]
  PIN nTOK_PMOS[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6914.105 1046.435 6914.385 1047.435 ;
    END
  END nTOK_PMOS[16]
  PIN BcidMtx[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6912.425 1046.435 6912.705 1047.435 ;
    END
  END BcidMtx[436]
  PIN Read_PMOS[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6910.745 1046.435 6911.025 1047.435 ;
    END
  END Read_PMOS[16]
  PIN Read_PMOS[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7470.745 1046.435 7471.025 1047.435 ;
    END
  END Read_PMOS[23]
  PIN BcidMtx[475]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7469.625 1046.435 7469.905 1047.435 ;
    END
  END BcidMtx[475]
  PIN Data_PMOS[486]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7466.825 1046.435 7467.105 1047.435 ;
    END
  END Data_PMOS[486]
  PIN Data_PMOS[493]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7464.585 1046.435 7464.865 1047.435 ;
    END
  END Data_PMOS[493]
  PIN Data_PMOS[499]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7463.465 1046.435 7463.745 1047.435 ;
    END
  END Data_PMOS[499]
  PIN Data_PMOS[483]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7461.785 1046.435 7462.065 1047.435 ;
    END
  END Data_PMOS[483]
  PIN MASKD[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7451.145 1046.435 7451.425 1047.435 ;
    END
  END MASKD[158]
  PIN MASKD[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7446.665 1046.435 7446.945 1047.435 ;
    END
  END MASKD[157]
  PIN MASKV[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7441.905 1046.435 7442.185 1047.435 ;
    END
  END MASKV[157]
  PIN Data_PMOS[474]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7440.225 1046.435 7440.505 1047.435 ;
    END
  END Data_PMOS[474]
  PIN Data_PMOS[475]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7413.065 1046.435 7413.345 1047.435 ;
    END
  END Data_PMOS[475]
  PIN Data_PMOS[469]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7411.385 1046.435 7411.665 1047.435 ;
    END
  END Data_PMOS[469]
  PIN nTOK_PMOS[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7408.585 1046.435 7408.865 1047.435 ;
    END
  END nTOK_PMOS[22]
  PIN BcidMtx[472]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7406.905 1046.435 7407.185 1047.435 ;
    END
  END BcidMtx[472]
  PIN Read_PMOS[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7405.225 1046.435 7405.505 1047.435 ;
    END
  END Read_PMOS[22]
  PIN BcidMtx[470]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7404.665 1046.435 7404.945 1047.435 ;
    END
  END BcidMtx[470]
  PIN INJ_IN[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7402.425 1046.435 7402.705 1047.435 ;
    END
  END INJ_IN[156]
  PIN Data_PMOS[471]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7400.185 1046.435 7400.465 1047.435 ;
    END
  END Data_PMOS[471]
  PIN Data_PMOS[466]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7385.625 1046.435 7385.905 1047.435 ;
    END
  END Data_PMOS[466]
  PIN Data_PMOS[463]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7383.945 1046.435 7384.225 1047.435 ;
    END
  END Data_PMOS[463]
  PIN Data_PMOS[479]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7382.825 1046.435 7383.105 1047.435 ;
    END
  END Data_PMOS[479]
  PIN MASKD[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7381.145 1046.435 7381.425 1047.435 ;
    END
  END MASKD[156]
  PIN DIG_MON_SEL[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7378.345 1046.435 7378.625 1047.435 ;
    END
  END DIG_MON_SEL[156]
  PIN DIG_MON_PMOS[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7375.545 1046.435 7375.825 1047.435 ;
    END
  END DIG_MON_PMOS[43]
  PIN Data_PMOS[459]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7333.545 1046.435 7333.825 1047.435 ;
    END
  END Data_PMOS[459]
  PIN Data_PMOS[460]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7331.865 1046.435 7332.145 1047.435 ;
    END
  END Data_PMOS[460]
  PIN Data_PMOS[461]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7330.185 1046.435 7330.465 1047.435 ;
    END
  END Data_PMOS[461]
  PIN Data_PMOS[447]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7328.505 1046.435 7328.785 1047.435 ;
    END
  END Data_PMOS[447]
  PIN BcidMtx[467]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7325.145 1046.435 7325.425 1047.435 ;
    END
  END BcidMtx[467]
  PIN BcidMtx[465]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7324.025 1046.435 7324.305 1047.435 ;
    END
  END BcidMtx[465]
  PIN BcidMtx[464]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7322.345 1046.435 7322.625 1047.435 ;
    END
  END BcidMtx[464]
  PIN Data_HV[1113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18809.065 1046.435 18809.345 1047.435 ;
    END
  END Data_HV[1113]
  PIN Data_PMOS[443]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7310.025 1046.435 7310.305 1047.435 ;
    END
  END Data_PMOS[443]
  PIN Data_PMOS[450]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7309.465 1046.435 7309.745 1047.435 ;
    END
  END Data_PMOS[450]
  PIN Data_PMOS[445]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7307.785 1046.435 7308.065 1047.435 ;
    END
  END Data_PMOS[445]
  PIN Data_PMOS[442]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7306.105 1046.435 7306.385 1047.435 ;
    END
  END Data_PMOS[442]
  PIN MASKV[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7302.465 1046.435 7302.745 1047.435 ;
    END
  END MASKV[154]
  PIN MASKD[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7301.345 1046.435 7301.625 1047.435 ;
    END
  END MASKD[154]
  PIN DIG_MON_SEL[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7298.545 1046.435 7298.825 1047.435 ;
    END
  END DIG_MON_SEL[154]
  PIN DIG_MON_PMOS[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8389.705 1046.435 8389.985 1047.435 ;
    END
  END DIG_MON_PMOS[69]
  PIN MASKV[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8388.025 1046.435 8388.305 1047.435 ;
    END
  END MASKV[181]
  PIN Data_PMOS[726]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8386.345 1046.435 8386.625 1047.435 ;
    END
  END Data_PMOS[726]
  PIN Data_PMOS[734]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8384.105 1046.435 8384.385 1047.435 ;
    END
  END Data_PMOS[734]
  PIN Data_PMOS[721]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8382.985 1046.435 8383.265 1047.435 ;
    END
  END Data_PMOS[721]
  PIN nTOK_PMOS[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8380.185 1046.435 8380.465 1047.435 ;
    END
  END nTOK_PMOS[34]
  PIN FREEZE_PMOS[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8363.945 1046.435 8364.225 1047.435 ;
    END
  END FREEZE_PMOS[34]
  PIN BcidMtx[542]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8362.825 1046.435 8363.105 1047.435 ;
    END
  END BcidMtx[542]
  PIN INJ_IN[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8360.585 1046.435 8360.865 1047.435 ;
    END
  END INJ_IN[180]
  PIN Data_PMOS[729]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8357.785 1046.435 8358.065 1047.435 ;
    END
  END Data_PMOS[729]
  PIN Data_PMOS[718]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8356.665 1046.435 8356.945 1047.435 ;
    END
  END Data_PMOS[718]
  PIN Data_PMOS[715]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8354.985 1046.435 8355.265 1047.435 ;
    END
  END Data_PMOS[715]
  PIN MASKH[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8314.105 1046.435 8314.385 1047.435 ;
    END
  END MASKH[90]
  PIN DIG_MON_PMOS[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8312.425 1046.435 8312.705 1047.435 ;
    END
  END DIG_MON_PMOS[68]
  PIN DIG_MON_SEL[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8310.185 1046.435 8310.465 1047.435 ;
    END
  END DIG_MON_SEL[179]
  PIN MASKV[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8306.265 1046.435 8306.545 1047.435 ;
    END
  END MASKV[179]
  PIN Data_PMOS[701]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8305.145 1046.435 8305.425 1047.435 ;
    END
  END Data_PMOS[701]
  PIN Data_PMOS[698]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8303.465 1046.435 8303.745 1047.435 ;
    END
  END Data_PMOS[698]
  PIN Data_PMOS[700]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8301.225 1046.435 8301.505 1047.435 ;
    END
  END Data_PMOS[700]
  PIN INJ_IN[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8291.145 1046.435 8291.425 1047.435 ;
    END
  END INJ_IN[179]
  PIN BcidMtx[538]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8288.345 1046.435 8288.625 1047.435 ;
    END
  END BcidMtx[538]
  PIN BcidMtx[536]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8286.105 1046.435 8286.385 1047.435 ;
    END
  END BcidMtx[536]
  PIN Data_HV[1130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18808.505 1046.435 18808.785 1047.435 ;
    END
  END Data_HV[1130]
  PIN Data_PMOS[696]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8280.785 1046.435 8281.065 1047.435 ;
    END
  END Data_PMOS[696]
  PIN Data_PMOS[703]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8278.545 1046.435 8278.825 1047.435 ;
    END
  END Data_PMOS[703]
  PIN Data_PMOS[709]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8251.945 1046.435 8252.225 1047.435 ;
    END
  END Data_PMOS[709]
  PIN Data_PMOS[693]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8250.265 1046.435 8250.545 1047.435 ;
    END
  END Data_PMOS[693]
  PIN MASKD[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8248.025 1046.435 8248.305 1047.435 ;
    END
  END MASKD[178]
  PIN MASKD[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8243.545 1046.435 8243.825 1047.435 ;
    END
  END MASKD[177]
  PIN Data_PMOS[690]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8240.185 1046.435 8240.465 1047.435 ;
    END
  END Data_PMOS[690]
  PIN Data_PMOS[684]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8226.185 1046.435 8226.465 1047.435 ;
    END
  END Data_PMOS[684]
  PIN Data_PMOS[685]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8224.505 1046.435 8224.785 1047.435 ;
    END
  END Data_PMOS[685]
  PIN Data_PMOS[678]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8222.265 1046.435 8222.545 1047.435 ;
    END
  END Data_PMOS[678]
  PIN nTOK_PMOS[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8220.025 1046.435 8220.305 1047.435 ;
    END
  END nTOK_PMOS[32]
  PIN BcidMtx[531]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8217.785 1046.435 8218.065 1047.435 ;
    END
  END BcidMtx[531]
  PIN BcidMtx[528]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8214.985 1046.435 8215.265 1047.435 ;
    END
  END BcidMtx[528]
  PIN Data_PMOS[675]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8174.105 1046.435 8174.385 1047.435 ;
    END
  END Data_PMOS[675]
  PIN Data_PMOS[687]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8172.425 1046.435 8172.705 1047.435 ;
    END
  END Data_PMOS[687]
  PIN Data_PMOS[683]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8170.185 1046.435 8170.465 1047.435 ;
    END
  END Data_PMOS[683]
  PIN Data_PMOS[672]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8169.065 1046.435 8169.345 1047.435 ;
    END
  END Data_PMOS[672]
  PIN MASKH[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8167.385 1046.435 8167.665 1047.435 ;
    END
  END MASKH[88]
  PIN DIG_MON_SEL[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8164.025 1046.435 8164.305 1047.435 ;
    END
  END DIG_MON_SEL[176]
  PIN MASKD[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8162.345 1046.435 8162.625 1047.435 ;
    END
  END MASKD[175]
  PIN MASKV[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8151.145 1046.435 8151.425 1047.435 ;
    END
  END MASKV[175]
  PIN Data_PMOS[670]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8148.905 1046.435 8149.185 1047.435 ;
    END
  END Data_PMOS[670]
  PIN Data_PMOS[664]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8147.785 1046.435 8148.065 1047.435 ;
    END
  END Data_PMOS[664]
  PIN Data_PMOS[658]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8146.105 1046.435 8146.385 1047.435 ;
    END
  END Data_PMOS[658]
  PIN BcidMtx[527]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8140.225 1046.435 8140.505 1047.435 ;
    END
  END BcidMtx[527]
  PIN BcidMtx[525]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8139.105 1046.435 8139.385 1047.435 ;
    END
  END BcidMtx[525]
  PIN BcidMtx[523]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8111.385 1046.435 8111.665 1047.435 ;
    END
  END BcidMtx[523]
  PIN Data_PMOS[653]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8108.025 1046.435 8108.305 1047.435 ;
    END
  END Data_PMOS[653]
  PIN Data_PMOS[666]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8106.905 1046.435 8107.185 1047.435 ;
    END
  END Data_PMOS[666]
  PIN Data_PMOS[667]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8105.225 1046.435 8105.505 1047.435 ;
    END
  END Data_PMOS[667]
  PIN Data_PMOS[668]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8102.985 1046.435 8103.265 1047.435 ;
    END
  END Data_PMOS[668]
  PIN MASKH[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8101.865 1046.435 8102.145 1047.435 ;
    END
  END MASKH[87]
  PIN DIG_MON_PMOS[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8082.825 1046.435 8083.105 1047.435 ;
    END
  END DIG_MON_PMOS[61]
  PIN MASKV[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8081.145 1046.435 8081.425 1047.435 ;
    END
  END MASKV[173]
  PIN Data_PMOS[642]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8079.465 1046.435 8079.745 1047.435 ;
    END
  END Data_PMOS[642]
  PIN Data_PMOS[650]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8077.225 1046.435 8077.505 1047.435 ;
    END
  END Data_PMOS[650]
  PIN Data_PMOS[637]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8076.105 1046.435 8076.385 1047.435 ;
    END
  END Data_PMOS[637]
  PIN BcidMtx[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6909.065 1046.435 6909.345 1047.435 ;
    END
  END BcidMtx[432]
  PIN Data_PMOS[339]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6906.825 1046.435 6907.105 1047.435 ;
    END
  END Data_PMOS[339]
  PIN Data_PMOS[351]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6905.145 1046.435 6905.425 1047.435 ;
    END
  END Data_PMOS[351]
  PIN Data_PMOS[347]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6902.905 1046.435 6903.185 1047.435 ;
    END
  END Data_PMOS[347]
  PIN Data_PMOS[336]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6901.785 1046.435 6902.065 1047.435 ;
    END
  END Data_PMOS[336]
  PIN MASKH[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6891.705 1046.435 6891.985 1047.435 ;
    END
  END MASKH[72]
  PIN DIG_MON_SEL[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6888.345 1046.435 6888.625 1047.435 ;
    END
  END DIG_MON_SEL[144]
  PIN MASKD[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6886.665 1046.435 6886.945 1047.435 ;
    END
  END MASKD[143]
  PIN INJ_ROW[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6882.465 1046.435 6882.745 1047.435 ;
    END
  END INJ_ROW[71]
  PIN Data_PMOS[327]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6880.225 1046.435 6880.505 1047.435 ;
    END
  END Data_PMOS[327]
  PIN Data_PMOS[328]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6853.065 1046.435 6853.345 1047.435 ;
    END
  END Data_PMOS[328]
  PIN Data_PMOS[322]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6851.385 1046.435 6851.665 1047.435 ;
    END
  END Data_PMOS[322]
  PIN nTOK_PMOS[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6848.585 1046.435 6848.865 1047.435 ;
    END
  END nTOK_PMOS[15]
  PIN BcidMtx[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6846.905 1046.435 6847.185 1047.435 ;
    END
  END BcidMtx[430]
  PIN Read_PMOS[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6845.225 1046.435 6845.505 1047.435 ;
    END
  END Read_PMOS[15]
  PIN INJ_IN[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6842.425 1046.435 6842.705 1047.435 ;
    END
  END INJ_IN[142]
  PIN Data_PMOS[317]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6840.745 1046.435 6841.025 1047.435 ;
    END
  END Data_PMOS[317]
  PIN Data_PMOS[325]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6826.185 1046.435 6826.465 1047.435 ;
    END
  END Data_PMOS[325]
  PIN Data_PMOS[316]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6823.945 1046.435 6824.225 1047.435 ;
    END
  END Data_PMOS[316]
  PIN Data_PMOS[332]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6822.825 1046.435 6823.105 1047.435 ;
    END
  END Data_PMOS[332]
  PIN MASKD[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6821.145 1046.435 6821.425 1047.435 ;
    END
  END MASKD[142]
  PIN DIG_MON_SEL[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6817.785 1046.435 6818.065 1047.435 ;
    END
  END DIG_MON_SEL[141]
  PIN DIG_MON_PMOS[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6815.545 1046.435 6815.825 1047.435 ;
    END
  END DIG_MON_PMOS[29]
  PIN Data_PMOS[312]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6773.545 1046.435 6773.825 1047.435 ;
    END
  END Data_PMOS[312]
  PIN Data_PMOS[299]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6771.305 1046.435 6771.585 1047.435 ;
    END
  END Data_PMOS[299]
  PIN Data_PMOS[314]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6770.185 1046.435 6770.465 1047.435 ;
    END
  END Data_PMOS[314]
  PIN Data_PMOS[300]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6768.505 1046.435 6768.785 1047.435 ;
    END
  END Data_PMOS[300]
  PIN BcidMtx[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6764.585 1046.435 6764.865 1047.435 ;
    END
  END BcidMtx[424]
  PIN FREEZE_PMOS[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6763.465 1046.435 6763.745 1047.435 ;
    END
  END FREEZE_PMOS[14]
  PIN BcidMtx[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6761.785 1046.435 6762.065 1047.435 ;
    END
  END BcidMtx[421]
  PIN Data_PMOS[297]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6750.585 1046.435 6750.865 1047.435 ;
    END
  END Data_PMOS[297]
  PIN Data_PMOS[303]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6749.465 1046.435 6749.745 1047.435 ;
    END
  END Data_PMOS[303]
  PIN Data_HV[1128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18812.425 1046.435 18812.705 1047.435 ;
    END
  END Data_HV[1128]
  PIN Data_PMOS[295]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6746.105 1046.435 6746.385 1047.435 ;
    END
  END Data_PMOS[295]
  PIN Data_PMOS[311]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6744.985 1046.435 6745.265 1047.435 ;
    END
  END Data_PMOS[311]
  PIN MASKD[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6741.345 1046.435 6741.625 1047.435 ;
    END
  END MASKD[140]
  PIN FREEZE_PMOS[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6993.065 1046.435 6993.345 1047.435 ;
    END
  END FREEZE_PMOS[17]
  PIN MASKD[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7830.825 1046.435 7831.105 1047.435 ;
    END
  END MASKD[167]
  PIN MASKV[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7828.025 1046.435 7828.305 1047.435 ;
    END
  END MASKV[167]
  PIN Data_PMOS[586]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7825.785 1046.435 7826.065 1047.435 ;
    END
  END Data_PMOS[586]
  PIN Data_PMOS[580]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7824.665 1046.435 7824.945 1047.435 ;
    END
  END Data_PMOS[580]
  PIN Data_PMOS[574]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7822.985 1046.435 7823.265 1047.435 ;
    END
  END Data_PMOS[574]
  PIN BcidMtx[503]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7805.625 1046.435 7805.905 1047.435 ;
    END
  END BcidMtx[503]
  PIN BcidMtx[501]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7804.505 1046.435 7804.785 1047.435 ;
    END
  END BcidMtx[501]
  PIN BcidMtx[500]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7802.825 1046.435 7803.105 1047.435 ;
    END
  END BcidMtx[500]
  PIN Data_HV[1123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18811.865 1046.435 18812.145 1047.435 ;
    END
  END Data_HV[1123]
  PIN Data_PMOS[569]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7798.905 1046.435 7799.185 1047.435 ;
    END
  END Data_PMOS[569]
  PIN Data_PMOS[577]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7797.225 1046.435 7797.505 1047.435 ;
    END
  END Data_PMOS[577]
  PIN Data_PMOS[568]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7794.985 1046.435 7795.265 1047.435 ;
    END
  END Data_PMOS[568]
  PIN Data_PMOS[584]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7793.865 1046.435 7794.145 1047.435 ;
    END
  END Data_PMOS[584]
  PIN MASKD[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7753.545 1046.435 7753.825 1047.435 ;
    END
  END MASKD[166]
  PIN DIG_MON_SEL[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7750.185 1046.435 7750.465 1047.435 ;
    END
  END DIG_MON_SEL[165]
  PIN DIG_MON_PMOS[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7747.945 1046.435 7748.225 1047.435 ;
    END
  END DIG_MON_PMOS[53]
  PIN Data_PMOS[564]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7745.705 1046.435 7745.985 1047.435 ;
    END
  END Data_PMOS[564]
  PIN Data_PMOS[551]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7743.465 1046.435 7743.745 1047.435 ;
    END
  END Data_PMOS[551]
  PIN Data_PMOS[566]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7742.345 1046.435 7742.625 1047.435 ;
    END
  END Data_PMOS[566]
  PIN Data_PMOS[552]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7732.265 1046.435 7732.545 1047.435 ;
    END
  END Data_PMOS[552]
  PIN BcidMtx[496]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7728.345 1046.435 7728.625 1047.435 ;
    END
  END BcidMtx[496]
  PIN FREEZE_PMOS[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7727.225 1046.435 7727.505 1047.435 ;
    END
  END FREEZE_PMOS[26]
  PIN BcidMtx[493]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7725.545 1046.435 7725.825 1047.435 ;
    END
  END BcidMtx[493]
  PIN Data_PMOS[548]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7720.225 1046.435 7720.505 1047.435 ;
    END
  END Data_PMOS[548]
  PIN Data_PMOS[561]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7719.105 1046.435 7719.385 1047.435 ;
    END
  END Data_PMOS[561]
  PIN Data_PMOS[550]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7692.505 1046.435 7692.785 1047.435 ;
    END
  END Data_PMOS[550]
  PIN Data_PMOS[546]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7690.265 1046.435 7690.545 1047.435 ;
    END
  END Data_PMOS[546]
  PIN MASKV[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7689.145 1046.435 7689.425 1047.435 ;
    END
  END MASKV[164]
  PIN DIG_MON_PMOS[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7686.905 1046.435 7687.185 1047.435 ;
    END
  END DIG_MON_PMOS[52]
  PIN MASKD[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7683.545 1046.435 7683.825 1047.435 ;
    END
  END MASKD[163]
  PIN INJ_ROW[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7681.305 1046.435 7681.585 1047.435 ;
    END
  END INJ_ROW[81]
  PIN Data_PMOS[533]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7679.625 1046.435 7679.905 1047.435 ;
    END
  END Data_PMOS[533]
  PIN Data_PMOS[538]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7664.505 1046.435 7664.785 1047.435 ;
    END
  END Data_PMOS[538]
  PIN Data_PMOS[539]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7663.385 1046.435 7663.665 1047.435 ;
    END
  END Data_PMOS[539]
  PIN INJ_IN[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7661.145 1046.435 7661.425 1047.435 ;
    END
  END INJ_IN[163]
  PIN BcidMtx[489]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7657.785 1046.435 7658.065 1047.435 ;
    END
  END BcidMtx[489]
  PIN Read_PMOS[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7656.665 1046.435 7656.945 1047.435 ;
    END
  END Read_PMOS[25]
  PIN BcidMtx[486]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7654.985 1046.435 7655.265 1047.435 ;
    END
  END BcidMtx[486]
  PIN Data_PMOS[534]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7612.985 1046.435 7613.265 1047.435 ;
    END
  END Data_PMOS[534]
  PIN Data_PMOS[535]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7611.865 1046.435 7612.145 1047.435 ;
    END
  END Data_PMOS[535]
  PIN Data_PMOS[536]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7610.185 1046.435 7610.465 1047.435 ;
    END
  END Data_PMOS[536]
  PIN MASKV[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7607.945 1046.435 7608.225 1047.435 ;
    END
  END MASKV[162]
  PIN MASKD[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7606.825 1046.435 7607.105 1047.435 ;
    END
  END MASKD[162]
  PIN DIG_MON_SEL[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7604.025 1046.435 7604.305 1047.435 ;
    END
  END DIG_MON_SEL[162]
  PIN INJ_ROW[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7591.705 1046.435 7591.985 1047.435 ;
    END
  END INJ_ROW[80]
  PIN Data_PMOS[522]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7590.585 1046.435 7590.865 1047.435 ;
    END
  END Data_PMOS[522]
  PIN Data_PMOS[523]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7588.905 1046.435 7589.185 1047.435 ;
    END
  END Data_PMOS[523]
  PIN Data_PMOS[518]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7586.665 1046.435 7586.945 1047.435 ;
    END
  END Data_PMOS[518]
  PIN Data_PMOS[510]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7585.545 1046.435 7585.825 1047.435 ;
    END
  END Data_PMOS[510]
  PIN BcidMtx[485]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7580.225 1046.435 7580.505 1047.435 ;
    END
  END BcidMtx[485]
  PIN BcidMtx[482]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7551.945 1046.435 7552.225 1047.435 ;
    END
  END BcidMtx[482]
  PIN BcidMtx[480]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7550.825 1046.435 7551.105 1047.435 ;
    END
  END BcidMtx[480]
  PIN Data_PMOS[506]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7548.025 1046.435 7548.305 1047.435 ;
    END
  END Data_PMOS[506]
  PIN Data_PMOS[508]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7545.785 1046.435 7546.065 1047.435 ;
    END
  END Data_PMOS[508]
  PIN Data_PMOS[515]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7544.665 1046.435 7544.945 1047.435 ;
    END
  END Data_PMOS[515]
  PIN Data_PMOS[521]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7542.985 1046.435 7543.265 1047.435 ;
    END
  END Data_PMOS[521]
  PIN DIG_MON_PMOS[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7540.185 1046.435 7540.465 1047.435 ;
    END
  END DIG_MON_PMOS[48]
  PIN DIG_MON_SEL[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7525.625 1046.435 7525.905 1047.435 ;
    END
  END DIG_MON_SEL[160]
  PIN DIG_MON_PMOS[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7522.825 1046.435 7523.105 1047.435 ;
    END
  END DIG_MON_PMOS[47]
  PIN Data_PMOS[491]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7520.025 1046.435 7520.305 1047.435 ;
    END
  END Data_PMOS[491]
  PIN Data_PMOS[502]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7518.905 1046.435 7519.185 1047.435 ;
    END
  END Data_PMOS[502]
  PIN Data_PMOS[503]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7517.225 1046.435 7517.505 1047.435 ;
    END
  END Data_PMOS[503]
  PIN INJ_IN[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7514.425 1046.435 7514.705 1047.435 ;
    END
  END INJ_IN[159]
  PIN Data_HV[1115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18813.545 1046.435 18813.825 1047.435 ;
    END
  END Data_HV[1115]
  PIN BcidMtx[479]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7472.985 1046.435 7473.265 1047.435 ;
    END
  END BcidMtx[479]
  PIN Data_COMP[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10316.665 1046.435 10316.945 1047.435 ;
    END
  END Data_COMP[56]
  PIN BcidMtx[689]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10272.985 1046.435 10273.265 1047.435 ;
    END
  END BcidMtx[689]
  PIN BcidMtx[687]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10271.865 1046.435 10272.145 1047.435 ;
    END
  END BcidMtx[687]
  PIN Read_COMP[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10270.745 1046.435 10271.025 1047.435 ;
    END
  END Read_COMP[2]
  PIN INJ_IN[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10267.945 1046.435 10268.225 1047.435 ;
    END
  END INJ_IN[228]
  PIN Data_COMP[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10266.265 1046.435 10266.545 1047.435 ;
    END
  END Data_COMP[44]
  PIN Data_COMP[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10264.585 1046.435 10264.865 1047.435 ;
    END
  END Data_COMP[52]
  PIN Data_COMP[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10262.905 1046.435 10263.185 1047.435 ;
    END
  END Data_COMP[53]
  PIN Data_COMP[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10261.785 1046.435 10262.065 1047.435 ;
    END
  END Data_COMP[42]
  PIN MASKV[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10252.265 1046.435 10252.545 1047.435 ;
    END
  END MASKV[228]
  PIN DIG_MON_SEL[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10247.785 1046.435 10248.065 1047.435 ;
    END
  END DIG_MON_SEL[227]
  PIN INJ_ROW[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10242.465 1046.435 10242.745 1047.435 ;
    END
  END INJ_ROW[113]
  PIN Data_COMP[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10240.225 1046.435 10240.505 1047.435 ;
    END
  END Data_COMP[33]
  PIN Data_COMP[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10239.105 1046.435 10239.385 1047.435 ;
    END
  END Data_COMP[26]
  PIN Data_COMP[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10211.945 1046.435 10212.225 1047.435 ;
    END
  END Data_COMP[35]
  PIN nTOK_COMP[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10208.585 1046.435 10208.865 1047.435 ;
    END
  END nTOK_COMP[1]
  PIN BcidMtx[683]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10207.465 1046.435 10207.745 1047.435 ;
    END
  END BcidMtx[683]
  PIN FREEZE_COMP[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10205.785 1046.435 10206.065 1047.435 ;
    END
  END FREEZE_COMP[1]
  PIN INJ_IN[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10202.425 1046.435 10202.705 1047.435 ;
    END
  END INJ_IN[226]
  PIN Data_COMP[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10201.305 1046.435 10201.585 1047.435 ;
    END
  END Data_COMP[24]
  PIN Data_COMP[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10186.745 1046.435 10187.025 1047.435 ;
    END
  END Data_COMP[36]
  PIN Data_COMP[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10184.505 1046.435 10184.785 1047.435 ;
    END
  END Data_COMP[32]
  PIN Data_COMP[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10183.945 1046.435 10184.225 1047.435 ;
    END
  END Data_COMP[22]
  PIN MASKV[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10182.265 1046.435 10182.545 1047.435 ;
    END
  END MASKV[226]
  PIN DIG_MON_SEL[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10178.345 1046.435 10178.625 1047.435 ;
    END
  END DIG_MON_SEL[226]
  PIN DIG_MON_COMP[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10175.545 1046.435 10175.825 1047.435 ;
    END
  END DIG_MON_COMP[1]
  PIN Data_COMP[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10132.425 1046.435 10132.705 1047.435 ;
    END
  END Data_COMP[12]
  PIN Data_COMP[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10131.865 1046.435 10132.145 1047.435 ;
    END
  END Data_COMP[19]
  PIN Data_COMP[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10130.185 1046.435 10130.465 1047.435 ;
    END
  END Data_COMP[20]
  PIN nTOK_COMP[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10126.265 1046.435 10126.545 1047.435 ;
    END
  END nTOK_COMP[0]
  PIN BcidMtx[676]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10124.585 1046.435 10124.865 1047.435 ;
    END
  END BcidMtx[676]
  PIN Read_COMP[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10122.905 1046.435 10123.185 1047.435 ;
    END
  END Read_COMP[0]
  PIN INJ_IN[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10111.705 1046.435 10111.985 1047.435 ;
    END
  END INJ_IN[224]
  PIN Data_COMP[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10110.025 1046.435 10110.305 1047.435 ;
    END
  END Data_COMP[2]
  PIN Data_COMP[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10108.345 1046.435 10108.625 1047.435 ;
    END
  END Data_COMP[10]
  PIN Data_COMP[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10106.105 1046.435 10106.385 1047.435 ;
    END
  END Data_COMP[1]
  PIN Data_COMP[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10104.985 1046.435 10105.265 1047.435 ;
    END
  END Data_COMP[17]
  PIN MASKD[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10101.345 1046.435 10101.625 1047.435 ;
    END
  END MASKD[224]
  PIN FREEZE_COMP[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10353.065 1046.435 10353.345 1047.435 ;
    END
  END FREEZE_COMP[3]
  PIN MASKD[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11190.825 1046.435 11191.105 1047.435 ;
    END
  END MASKD[251]
  PIN MASKV[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11188.025 1046.435 11188.305 1047.435 ;
    END
  END MASKV[251]
  PIN Data_COMP[292]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11185.785 1046.435 11186.065 1047.435 ;
    END
  END Data_COMP[292]
  PIN Data_COMP[286]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11184.665 1046.435 11184.945 1047.435 ;
    END
  END Data_COMP[286]
  PIN Data_COMP[280]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11182.985 1046.435 11183.265 1047.435 ;
    END
  END Data_COMP[280]
  PIN BcidMtx[755]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11165.625 1046.435 11165.905 1047.435 ;
    END
  END BcidMtx[755]
  PIN BcidMtx[753]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11164.505 1046.435 11164.785 1047.435 ;
    END
  END BcidMtx[753]
  PIN BcidMtx[752]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11162.825 1046.435 11163.105 1047.435 ;
    END
  END BcidMtx[752]
  PIN Data_COMP[276]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11159.465 1046.435 11159.745 1047.435 ;
    END
  END Data_COMP[276]
  PIN Data_COMP[282]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11158.345 1046.435 11158.625 1047.435 ;
    END
  END Data_COMP[282]
  PIN Data_COMP[277]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11156.665 1046.435 11156.945 1047.435 ;
    END
  END Data_COMP[277]
  PIN Data_COMP[273]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11154.425 1046.435 11154.705 1047.435 ;
    END
  END Data_COMP[273]
  PIN MASKV[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11114.665 1046.435 11114.945 1047.435 ;
    END
  END MASKV[250]
  PIN MASKH[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11114.105 1046.435 11114.385 1047.435 ;
    END
  END MASKH[125]
  PIN DIG_MON_SEL[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11110.185 1046.435 11110.465 1047.435 ;
    END
  END DIG_MON_SEL[249]
  PIN MASKD[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11109.065 1046.435 11109.345 1047.435 ;
    END
  END MASKD[249]
  PIN INJ_ROW[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11106.825 1046.435 11107.105 1047.435 ;
    END
  END INJ_ROW[124]
  PIN Data_COMP[271]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11104.025 1046.435 11104.305 1047.435 ;
    END
  END Data_COMP[271]
  PIN Data_COMP[265]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11102.905 1046.435 11103.185 1047.435 ;
    END
  END Data_COMP[265]
  PIN Data_COMP[259]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11101.225 1046.435 11101.505 1047.435 ;
    END
  END Data_COMP[259]
  PIN BcidMtx[748]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11088.345 1046.435 11088.625 1047.435 ;
    END
  END BcidMtx[748]
  PIN BcidMtx[747]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11087.785 1046.435 11088.065 1047.435 ;
    END
  END BcidMtx[747]
  PIN BcidMtx[746]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11086.105 1046.435 11086.385 1047.435 ;
    END
  END BcidMtx[746]
  PIN Data_COMP[254]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11080.225 1046.435 11080.505 1047.435 ;
    END
  END Data_COMP[254]
  PIN Data_COMP[261]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11079.665 1046.435 11079.945 1047.435 ;
    END
  END Data_COMP[261]
  PIN Data_COMP[256]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11052.505 1046.435 11052.785 1047.435 ;
    END
  END Data_COMP[256]
  PIN Data_COMP[269]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11049.705 1046.435 11049.985 1047.435 ;
    END
  END Data_COMP[269]
  PIN MASKV[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11049.145 1046.435 11049.425 1047.435 ;
    END
  END MASKV[248]
  PIN DIG_MON_COMP[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11046.905 1046.435 11047.185 1047.435 ;
    END
  END DIG_MON_COMP[24]
  PIN DIG_MON_COMP[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11042.425 1046.435 11042.705 1047.435 ;
    END
  END DIG_MON_COMP[23]
  PIN INJ_ROW[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11041.305 1046.435 11041.585 1047.435 ;
    END
  END INJ_ROW[123]
  PIN Data_COMP[239]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11039.625 1046.435 11039.905 1047.435 ;
    END
  END Data_COMP[239]
  PIN Data_COMP[251]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11023.945 1046.435 11024.225 1047.435 ;
    END
  END Data_COMP[251]
  PIN Data_COMP[245]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11023.385 1046.435 11023.665 1047.435 ;
    END
  END Data_COMP[245]
  PIN INJ_IN[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11021.145 1046.435 11021.425 1047.435 ;
    END
  END INJ_IN[247]
  PIN FREEZE_COMP[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11017.225 1046.435 11017.505 1047.435 ;
    END
  END FREEZE_COMP[11]
  PIN Read_COMP[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11016.665 1046.435 11016.945 1047.435 ;
    END
  END Read_COMP[11]
  PIN BcidMtx[738]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11014.985 1046.435 11015.265 1047.435 ;
    END
  END BcidMtx[738]
  PIN Data_COMP[246]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10972.425 1046.435 10972.705 1047.435 ;
    END
  END Data_COMP[246]
  PIN Data_COMP[241]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10971.865 1046.435 10972.145 1047.435 ;
    END
  END Data_COMP[241]
  PIN Data_COMP[242]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10970.185 1046.435 10970.465 1047.435 ;
    END
  END Data_COMP[242]
  PIN MASKH[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10967.385 1046.435 10967.665 1047.435 ;
    END
  END MASKH[123]
  PIN DIG_MON_COMP[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10965.705 1046.435 10965.985 1047.435 ;
    END
  END DIG_MON_COMP[22]
  PIN DIG_MON_SEL[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10964.025 1046.435 10964.305 1047.435 ;
    END
  END DIG_MON_SEL[246]
  PIN MASKV[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10951.145 1046.435 10951.425 1047.435 ;
    END
  END MASKV[245]
  PIN Data_COMP[228]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10950.585 1046.435 10950.865 1047.435 ;
    END
  END Data_COMP[228]
  PIN Data_COMP[229]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10948.905 1046.435 10949.185 1047.435 ;
    END
  END Data_COMP[229]
  PIN Data_COMP[217]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10946.105 1046.435 10946.385 1047.435 ;
    END
  END Data_COMP[217]
  PIN Data_COMP[216]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10945.545 1046.435 10945.825 1047.435 ;
    END
  END Data_COMP[216]
  PIN BcidMtx[737]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10940.225 1046.435 10940.505 1047.435 ;
    END
  END BcidMtx[737]
  PIN BcidMtx[733]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10911.385 1046.435 10911.665 1047.435 ;
    END
  END BcidMtx[733]
  PIN BcidMtx[732]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10910.825 1046.435 10911.105 1047.435 ;
    END
  END BcidMtx[732]
  PIN INJ_IN[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10909.705 1046.435 10909.985 1047.435 ;
    END
  END INJ_IN[244]
  PIN Data_COMP[220]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10906.345 1046.435 10906.625 1047.435 ;
    END
  END Data_COMP[220]
  PIN Data_COMP[214]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10905.785 1046.435 10906.065 1047.435 ;
    END
  END Data_COMP[214]
  PIN Data_COMP[211]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10904.105 1046.435 10904.385 1047.435 ;
    END
  END Data_COMP[211]
  PIN MASKD[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10901.305 1046.435 10901.585 1047.435 ;
    END
  END MASKD[244]
  PIN DIG_MON_COMP[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10900.185 1046.435 10900.465 1047.435 ;
    END
  END DIG_MON_COMP[20]
  PIN DIG_MON_SEL[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10885.065 1046.435 10885.345 1047.435 ;
    END
  END DIG_MON_SEL[243]
  PIN Data_COMP[207]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10880.585 1046.435 10880.865 1047.435 ;
    END
  END Data_COMP[207]
  PIN Data_COMP[197]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10880.025 1046.435 10880.305 1047.435 ;
    END
  END Data_COMP[197]
  PIN nRST[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17379.105 1046.435 17379.385 1047.435 ;
    END
  END nRST[203]
  PIN nRST[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14579.105 1046.435 14579.385 1047.435 ;
    END
  END nRST[168]
  PIN nRST[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14019.105 1046.435 14019.385 1047.435 ;
    END
  END nRST[161]
  PIN nRST[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18499.105 1046.435 18499.385 1047.435 ;
    END
  END nRST[217]
  PIN nRST[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17939.105 1046.435 17939.385 1047.435 ;
    END
  END nRST[210]
  PIN nRST[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4578.905 1046.435 4579.185 1047.435 ;
    END
  END nRST[43]
  PIN nRST[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4018.905 1046.435 4019.185 1047.435 ;
    END
  END nRST[36]
  PIN nRST[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3458.905 1046.435 3459.185 1047.435 ;
    END
  END nRST[29]
  PIN nRST[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2898.905 1046.435 2899.185 1047.435 ;
    END
  END nRST[22]
  PIN nRST[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2338.905 1046.435 2339.185 1047.435 ;
    END
  END nRST[15]
  PIN nRST[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1778.905 1046.435 1779.185 1047.435 ;
    END
  END nRST[8]
  PIN nRST[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1218.905 1046.435 1219.185 1047.435 ;
    END
  END nRST[1]
  PIN nRST[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7125.785 1046.435 7126.065 1047.435 ;
    END
  END nRST[75]
  PIN nRST[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7685.785 1046.435 7686.065 1047.435 ;
    END
  END nRST[82]
  PIN nRST[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8245.785 1046.435 8246.065 1047.435 ;
    END
  END nRST[89]
  PIN nRST[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8805.785 1046.435 8806.065 1047.435 ;
    END
  END nRST[96]
  PIN nRST[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5698.905 1046.435 5699.185 1047.435 ;
    END
  END nRST[57]
  PIN nRST[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5138.905 1046.435 5139.185 1047.435 ;
    END
  END nRST[50]
  PIN nRST[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9365.785 1046.435 9366.065 1047.435 ;
    END
  END nRST[103]
  PIN nRST[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9925.785 1046.435 9926.065 1047.435 ;
    END
  END nRST[110]
  PIN nRST[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10485.785 1046.435 10486.065 1047.435 ;
    END
  END nRST[117]
  PIN nRST[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11045.785 1046.435 11046.065 1047.435 ;
    END
  END nRST[124]
  PIN nRST[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16819.105 1046.435 16819.385 1047.435 ;
    END
  END nRST[196]
  PIN nRST[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16259.105 1046.435 16259.385 1047.435 ;
    END
  END nRST[189]
  PIN nRST[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15699.105 1046.435 15699.385 1047.435 ;
    END
  END nRST[182]
  PIN nRST[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15139.105 1046.435 15139.385 1047.435 ;
    END
  END nRST[175]
  PIN nRST[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13459.105 1046.435 13459.385 1047.435 ;
    END
  END nRST[154]
  PIN nRST[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12899.105 1046.435 12899.385 1047.435 ;
    END
  END nRST[147]
  PIN nRST[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12339.105 1046.435 12339.385 1047.435 ;
    END
  END nRST[140]
  PIN nRST[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11779.105 1046.435 11779.385 1047.435 ;
    END
  END nRST[133]
  PIN nRST[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11219.105 1046.435 11219.385 1047.435 ;
    END
  END nRST[126]
  PIN nRST[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2819.105 1046.435 2819.385 1047.435 ;
    END
  END nRST[21]
  PIN nRST[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2259.105 1046.435 2259.385 1047.435 ;
    END
  END nRST[14]
  PIN nRST[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1139.105 1046.435 1139.385 1047.435 ;
    END
  END nRST[0]
  PIN nRST[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10326.185 1046.435 10326.465 1047.435 ;
    END
  END nRST[115]
  PIN nRST[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10886.185 1046.435 10886.465 1047.435 ;
    END
  END nRST[122]
  PIN nRST[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11446.185 1046.435 11446.465 1047.435 ;
    END
  END nRST[129]
  PIN nRST[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4499.105 1046.435 4499.385 1047.435 ;
    END
  END nRST[42]
  PIN nRST[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3939.105 1046.435 3939.385 1047.435 ;
    END
  END nRST[35]
  PIN nRST[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3379.105 1046.435 3379.385 1047.435 ;
    END
  END nRST[28]
  PIN nRST[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6739.105 1046.435 6739.385 1047.435 ;
    END
  END nRST[70]
  PIN nRST[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6179.105 1046.435 6179.385 1047.435 ;
    END
  END nRST[63]
  PIN nRST[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5619.105 1046.435 5619.385 1047.435 ;
    END
  END nRST[56]
  PIN nRST[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5059.105 1046.435 5059.385 1047.435 ;
    END
  END nRST[49]
  PIN nRST[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10659.105 1046.435 10659.385 1047.435 ;
    END
  END nRST[119]
  PIN nRST[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10099.105 1046.435 10099.385 1047.435 ;
    END
  END nRST[112]
  PIN nRST[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9539.105 1046.435 9539.385 1047.435 ;
    END
  END nRST[105]
  PIN nRST[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7299.105 1046.435 7299.385 1047.435 ;
    END
  END nRST[77]
  PIN nRST[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8979.105 1046.435 8979.385 1047.435 ;
    END
  END nRST[98]
  PIN nRST[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8419.105 1046.435 8419.385 1047.435 ;
    END
  END nRST[91]
  PIN nRST[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7859.105 1046.435 7859.385 1047.435 ;
    END
  END nRST[84]
  PIN nRST[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1699.105 1046.435 1699.385 1047.435 ;
    END
  END nRST[7]
  PIN nRST[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12006.185 1046.435 12006.465 1047.435 ;
    END
  END nRST[136]
  PIN nRST[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12566.185 1046.435 12566.465 1047.435 ;
    END
  END nRST[143]
  PIN nRST[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13126.185 1046.435 13126.465 1047.435 ;
    END
  END nRST[150]
  PIN nRST[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13686.185 1046.435 13686.465 1047.435 ;
    END
  END nRST[157]
  PIN nRST[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4244.585 1046.435 4244.865 1047.435 ;
    END
  END nRST[39]
  PIN nRST[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5924.585 1046.435 5924.865 1047.435 ;
    END
  END nRST[60]
  PIN nRST[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6484.585 1046.435 6484.865 1047.435 ;
    END
  END nRST[67]
  PIN nRST[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7044.585 1046.435 7044.865 1047.435 ;
    END
  END nRST[74]
  PIN nRST[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2564.585 1046.435 2564.865 1047.435 ;
    END
  END nRST[18]
  PIN nRST[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3124.585 1046.435 3124.865 1047.435 ;
    END
  END nRST[25]
  PIN nRST[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3684.585 1046.435 3684.865 1047.435 ;
    END
  END nRST[32]
  PIN nRST[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18726.185 1046.435 18726.465 1047.435 ;
    END
  END nRST[220]
  PIN nRST[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1444.585 1046.435 1444.865 1047.435 ;
    END
  END nRST[4]
  PIN nRST[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2004.585 1046.435 2004.865 1047.435 ;
    END
  END nRST[11]
  PIN nRST[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14246.185 1046.435 14246.465 1047.435 ;
    END
  END nRST[164]
  PIN nRST[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14806.185 1046.435 14806.465 1047.435 ;
    END
  END nRST[171]
  PIN nRST[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15366.185 1046.435 15366.465 1047.435 ;
    END
  END nRST[178]
  PIN nRST[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17046.185 1046.435 17046.465 1047.435 ;
    END
  END nRST[199]
  PIN nRST[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17606.185 1046.435 17606.465 1047.435 ;
    END
  END nRST[206]
  PIN nRST[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18166.185 1046.435 18166.465 1047.435 ;
    END
  END nRST[213]
  PIN nRST[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15926.185 1046.435 15926.465 1047.435 ;
    END
  END nRST[185]
  PIN nRST[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16486.185 1046.435 16486.465 1047.435 ;
    END
  END nRST[192]
  PIN nRST[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4804.585 1046.435 4804.865 1047.435 ;
    END
  END nRST[46]
  PIN nRST[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5364.585 1046.435 5364.865 1047.435 ;
    END
  END nRST[53]
  PIN nRST[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7604.585 1046.435 7604.865 1047.435 ;
    END
  END nRST[81]
  PIN nRST[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16004.585 1046.435 16004.865 1047.435 ;
    END
  END nRST[186]
  PIN nRST[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16564.585 1046.435 16564.865 1047.435 ;
    END
  END nRST[193]
  PIN nRST[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12084.585 1046.435 12084.865 1047.435 ;
    END
  END nRST[137]
  PIN nRST[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12644.585 1046.435 12644.865 1047.435 ;
    END
  END nRST[144]
  PIN nRST[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13204.585 1046.435 13204.865 1047.435 ;
    END
  END nRST[151]
  PIN nRST[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13764.585 1046.435 13764.865 1047.435 ;
    END
  END nRST[158]
  PIN nRST[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14324.585 1046.435 14324.865 1047.435 ;
    END
  END nRST[165]
  PIN nRST[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14884.585 1046.435 14884.865 1047.435 ;
    END
  END nRST[172]
  PIN nRST[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15444.585 1046.435 15444.865 1047.435 ;
    END
  END nRST[179]
  PIN nRST[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8164.585 1046.435 8164.865 1047.435 ;
    END
  END nRST[88]
  PIN nRST[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8724.585 1046.435 8724.865 1047.435 ;
    END
  END nRST[95]
  PIN nRST[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9284.585 1046.435 9284.865 1047.435 ;
    END
  END nRST[102]
  PIN nRST[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10404.585 1046.435 10404.865 1047.435 ;
    END
  END nRST[116]
  PIN nRST[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10964.585 1046.435 10964.865 1047.435 ;
    END
  END nRST[123]
  PIN nRST[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11524.585 1046.435 11524.865 1047.435 ;
    END
  END nRST[130]
  PIN nRST[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9844.585 1046.435 9844.865 1047.435 ;
    END
  END nRST[109]
  PIN nRST[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17124.585 1046.435 17124.865 1047.435 ;
    END
  END nRST[200]
  PIN nRST[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17684.585 1046.435 17684.865 1047.435 ;
    END
  END nRST[207]
  PIN nRST[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18244.585 1046.435 18244.865 1047.435 ;
    END
  END nRST[214]
  PIN nRST[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18804.585 1046.435 18804.865 1047.435 ;
    END
  END nRST[221]
  PIN nRST[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1525.785 1046.435 1526.065 1047.435 ;
    END
  END nRST[5]
  PIN nRST[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2085.785 1046.435 2086.065 1047.435 ;
    END
  END nRST[12]
  PIN nRST[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2645.785 1046.435 2646.065 1047.435 ;
    END
  END nRST[19]
  PIN nRST[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7938.905 1046.435 7939.185 1047.435 ;
    END
  END nRST[85]
  PIN nRST[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7378.905 1046.435 7379.185 1047.435 ;
    END
  END nRST[78]
  PIN nRST[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6818.905 1046.435 6819.185 1047.435 ;
    END
  END nRST[71]
  PIN nRST[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6258.905 1046.435 6259.185 1047.435 ;
    END
  END nRST[64]
  PIN nRST[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3205.785 1046.435 3206.065 1047.435 ;
    END
  END nRST[26]
  PIN nRST[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3765.785 1046.435 3766.065 1047.435 ;
    END
  END nRST[33]
  PIN nRST[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5445.785 1046.435 5446.065 1047.435 ;
    END
  END nRST[54]
  PIN nRST[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6005.785 1046.435 6006.065 1047.435 ;
    END
  END nRST[61]
  PIN nRST[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6565.785 1046.435 6566.065 1047.435 ;
    END
  END nRST[68]
  PIN nRST[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4325.785 1046.435 4326.065 1047.435 ;
    END
  END nRST[40]
  PIN nRST[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4885.785 1046.435 4886.065 1047.435 ;
    END
  END nRST[47]
  PIN SET_VCASN[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13427.955 1046.435 13428.235 1047.435 ;
    END
  END SET_VCASN[87]
  PIN SET_VCASN[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13567.955 1046.435 13568.235 1047.435 ;
    END
  END SET_VCASN[88]
  PIN SET_VCASN[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13707.955 1046.435 13708.235 1047.435 ;
    END
  END SET_VCASN[89]
  PIN SET_VCASN[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13847.955 1046.435 13848.235 1047.435 ;
    END
  END SET_VCASN[90]
  PIN SET_VCASN[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13987.955 1046.435 13988.235 1047.435 ;
    END
  END SET_VCASN[91]
  PIN SET_VCASN[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14127.955 1046.435 14128.235 1047.435 ;
    END
  END SET_VCASN[92]
  PIN SET_VCASN[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14267.955 1046.435 14268.235 1047.435 ;
    END
  END SET_VCASN[93]
  PIN SET_VCASN[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14407.955 1046.435 14408.235 1047.435 ;
    END
  END SET_VCASN[94]
  PIN SET_VCASN[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14547.955 1046.435 14548.235 1047.435 ;
    END
  END SET_VCASN[95]
  PIN SET_VCASN[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14687.955 1046.435 14688.235 1047.435 ;
    END
  END SET_VCASN[96]
  PIN SET_VCASN[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14827.955 1046.435 14828.235 1047.435 ;
    END
  END SET_VCASN[97]
  PIN SET_VCASN[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14967.955 1046.435 14968.235 1047.435 ;
    END
  END SET_VCASN[98]
  PIN SET_VCASN[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15107.955 1046.435 15108.235 1047.435 ;
    END
  END SET_VCASN[99]
  PIN SET_VCASN[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15247.955 1046.435 15248.235 1047.435 ;
    END
  END SET_VCASN[100]
  PIN SET_VCASN[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15387.955 1046.435 15388.235 1047.435 ;
    END
  END SET_VCASN[101]
  PIN SET_VCASN[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15527.955 1046.435 15528.235 1047.435 ;
    END
  END SET_VCASN[102]
  PIN SET_VCASN[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15667.955 1046.435 15668.235 1047.435 ;
    END
  END SET_VCASN[103]
  PIN SET_VCASN[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15807.955 1046.435 15808.235 1047.435 ;
    END
  END SET_VCASN[104]
  PIN SET_VCASN[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15947.955 1046.435 15948.235 1047.435 ;
    END
  END SET_VCASN[105]
  PIN SET_VCASN[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16087.955 1046.435 16088.235 1047.435 ;
    END
  END SET_VCASN[106]
  PIN SET_VCASN[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16227.955 1046.435 16228.235 1047.435 ;
    END
  END SET_VCASN[107]
  PIN SET_VCASN[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16367.955 1046.435 16368.235 1047.435 ;
    END
  END SET_VCASN[108]
  PIN SET_VCASN[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16507.955 1046.435 16508.235 1047.435 ;
    END
  END SET_VCASN[109]
  PIN SET_VCASN[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16647.955 1046.435 16648.235 1047.435 ;
    END
  END SET_VCASN[110]
  PIN SET_VCASN[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16787.955 1046.435 16788.235 1047.435 ;
    END
  END SET_VCASN[111]
  PIN SET_VCASN[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16927.955 1046.435 16928.235 1047.435 ;
    END
  END SET_VCASN[112]
  PIN SET_VCASN[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17067.955 1046.435 17068.235 1047.435 ;
    END
  END SET_VCASN[113]
  PIN SET_VCASN[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17207.955 1046.435 17208.235 1047.435 ;
    END
  END SET_VCASN[114]
  PIN SET_VCASN[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17347.955 1046.435 17348.235 1047.435 ;
    END
  END SET_VCASN[115]
  PIN SET_VCASN[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17487.955 1046.435 17488.235 1047.435 ;
    END
  END SET_VCASN[116]
  PIN SET_VCASN[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17627.955 1046.435 17628.235 1047.435 ;
    END
  END SET_VCASN[117]
  PIN SET_VCASN[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17767.955 1046.435 17768.235 1047.435 ;
    END
  END SET_VCASN[118]
  PIN SET_VCASN[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17907.955 1046.435 17908.235 1047.435 ;
    END
  END SET_VCASN[119]
  PIN SET_VCASN[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18047.955 1046.435 18048.235 1047.435 ;
    END
  END SET_VCASN[120]
  PIN SET_VCASN[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18187.955 1046.435 18188.235 1047.435 ;
    END
  END SET_VCASN[121]
  PIN SET_VCASN[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18327.955 1046.435 18328.235 1047.435 ;
    END
  END SET_VCASN[122]
  PIN SET_VCASN[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18467.955 1046.435 18468.235 1047.435 ;
    END
  END SET_VCASN[123]
  PIN SET_VCASN[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18607.955 1046.435 18608.235 1047.435 ;
    END
  END SET_VCASN[124]
  PIN SET_VCASN[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18747.955 1046.435 18748.235 1047.435 ;
    END
  END SET_VCASN[125]
  PIN SET_VCASN[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18887.955 1046.435 18888.235 1047.435 ;
    END
  END SET_VCASN[126]
  PIN SET_VCASN[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19027.955 1046.435 19028.235 1047.435 ;
    END
  END SET_VCASN[127]
  PIN SET_VRESET_P[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6560.675 1046.435 6560.955 1047.435 ;
    END
  END SET_VRESET_P[38]
  PIN SET_VRESET_P[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6700.675 1046.435 6700.955 1047.435 ;
    END
  END SET_VRESET_P[39]
  PIN SET_VRESET_P[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6840.675 1046.435 6840.955 1047.435 ;
    END
  END SET_VRESET_P[40]
  PIN SET_VRESET_P[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6980.675 1046.435 6980.955 1047.435 ;
    END
  END SET_VRESET_P[41]
  PIN SET_VRESET_P[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7120.675 1046.435 7120.955 1047.435 ;
    END
  END SET_VRESET_P[42]
  PIN SET_VRESET_P[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7260.675 1046.435 7260.955 1047.435 ;
    END
  END SET_VRESET_P[43]
  PIN SET_VRESET_P[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7400.675 1046.435 7400.955 1047.435 ;
    END
  END SET_VRESET_P[44]
  PIN SET_VRESET_P[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7540.675 1046.435 7540.955 1047.435 ;
    END
  END SET_VRESET_P[45]
  PIN SET_VRESET_P[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7680.675 1046.435 7680.955 1047.435 ;
    END
  END SET_VRESET_P[46]
  PIN SET_VRESET_P[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7820.675 1046.435 7820.955 1047.435 ;
    END
  END SET_VRESET_P[47]
  PIN SET_VRESET_P[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7960.675 1046.435 7960.955 1047.435 ;
    END
  END SET_VRESET_P[48]
  PIN SET_VRESET_P[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8100.675 1046.435 8100.955 1047.435 ;
    END
  END SET_VRESET_P[49]
  PIN SET_VRESET_P[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8240.675 1046.435 8240.955 1047.435 ;
    END
  END SET_VRESET_P[50]
  PIN SET_VRESET_P[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8380.675 1046.435 8380.955 1047.435 ;
    END
  END SET_VRESET_P[51]
  PIN SET_VRESET_P[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8520.675 1046.435 8520.955 1047.435 ;
    END
  END SET_VRESET_P[52]
  PIN SET_VRESET_P[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8660.675 1046.435 8660.955 1047.435 ;
    END
  END SET_VRESET_P[53]
  PIN SET_VRESET_P[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8800.675 1046.435 8800.955 1047.435 ;
    END
  END SET_VRESET_P[54]
  PIN SET_VRESET_P[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8940.675 1046.435 8940.955 1047.435 ;
    END
  END SET_VRESET_P[55]
  PIN SET_VRESET_P[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9080.675 1046.435 9080.955 1047.435 ;
    END
  END SET_VRESET_P[56]
  PIN SET_VRESET_P[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9220.675 1046.435 9220.955 1047.435 ;
    END
  END SET_VRESET_P[57]
  PIN SET_VRESET_P[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9360.675 1046.435 9360.955 1047.435 ;
    END
  END SET_VRESET_P[58]
  PIN SET_VRESET_P[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9500.675 1046.435 9500.955 1047.435 ;
    END
  END SET_VRESET_P[59]
  PIN SET_VRESET_P[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9640.675 1046.435 9640.955 1047.435 ;
    END
  END SET_VRESET_P[60]
  PIN SET_VRESET_P[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9780.675 1046.435 9780.955 1047.435 ;
    END
  END SET_VRESET_P[61]
  PIN SET_VRESET_P[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9920.675 1046.435 9920.955 1047.435 ;
    END
  END SET_VRESET_P[62]
  PIN SET_VRESET_P[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10060.675 1046.435 10060.955 1047.435 ;
    END
  END SET_VRESET_P[63]
  PIN SET_VRESET_P[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10200.675 1046.435 10200.955 1047.435 ;
    END
  END SET_VRESET_P[64]
  PIN SET_VRESET_P[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10340.675 1046.435 10340.955 1047.435 ;
    END
  END SET_VRESET_P[65]
  PIN SET_VRESET_P[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10480.675 1046.435 10480.955 1047.435 ;
    END
  END SET_VRESET_P[66]
  PIN SET_VRESET_P[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10620.675 1046.435 10620.955 1047.435 ;
    END
  END SET_VRESET_P[67]
  PIN SET_VRESET_P[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10760.675 1046.435 10760.955 1047.435 ;
    END
  END SET_VRESET_P[68]
  PIN SET_VRESET_P[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10900.675 1046.435 10900.955 1047.435 ;
    END
  END SET_VRESET_P[69]
  PIN SET_VRESET_P[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11040.675 1046.435 11040.955 1047.435 ;
    END
  END SET_VRESET_P[70]
  PIN SET_VRESET_P[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11180.675 1046.435 11180.955 1047.435 ;
    END
  END SET_VRESET_P[71]
  PIN SET_VRESET_P[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11320.675 1046.435 11320.955 1047.435 ;
    END
  END SET_VRESET_P[72]
  PIN SET_VRESET_P[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11460.675 1046.435 11460.955 1047.435 ;
    END
  END SET_VRESET_P[73]
  PIN SET_VRESET_P[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11600.675 1046.435 11600.955 1047.435 ;
    END
  END SET_VRESET_P[74]
  PIN SET_VRESET_P[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11740.675 1046.435 11740.955 1047.435 ;
    END
  END SET_VRESET_P[75]
  PIN SET_VRESET_P[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11880.675 1046.435 11880.955 1047.435 ;
    END
  END SET_VRESET_P[76]
  PIN SET_VRESET_P[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12020.675 1046.435 12020.955 1047.435 ;
    END
  END SET_VRESET_P[77]
  PIN SET_VRESET_P[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12160.675 1046.435 12160.955 1047.435 ;
    END
  END SET_VRESET_P[78]
  PIN SET_VRESET_P[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12300.675 1046.435 12300.955 1047.435 ;
    END
  END SET_VRESET_P[79]
  PIN SET_VRESET_P[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12440.675 1046.435 12440.955 1047.435 ;
    END
  END SET_VRESET_P[80]
  PIN SET_VRESET_P[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12580.675 1046.435 12580.955 1047.435 ;
    END
  END SET_VRESET_P[81]
  PIN SET_VRESET_P[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12720.675 1046.435 12720.955 1047.435 ;
    END
  END SET_VRESET_P[82]
  PIN SET_VRESET_P[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12860.675 1046.435 12860.955 1047.435 ;
    END
  END SET_VRESET_P[83]
  PIN SET_VRESET_P[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13000.675 1046.435 13000.955 1047.435 ;
    END
  END SET_VRESET_P[84]
  PIN SET_VRESET_P[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13140.675 1046.435 13140.955 1047.435 ;
    END
  END SET_VRESET_P[85]
  PIN SET_VRESET_P[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13280.675 1046.435 13280.955 1047.435 ;
    END
  END SET_VRESET_P[86]
  PIN SET_VRESET_P[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13420.675 1046.435 13420.955 1047.435 ;
    END
  END SET_VRESET_P[87]
  PIN SET_VRESET_P[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13560.675 1046.435 13560.955 1047.435 ;
    END
  END SET_VRESET_P[88]
  PIN SET_VRESET_P[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13700.675 1046.435 13700.955 1047.435 ;
    END
  END SET_VRESET_P[89]
  PIN SET_VRESET_P[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13840.675 1046.435 13840.955 1047.435 ;
    END
  END SET_VRESET_P[90]
  PIN SET_VRESET_P[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13980.675 1046.435 13980.955 1047.435 ;
    END
  END SET_VRESET_P[91]
  PIN SET_VRESET_P[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14120.675 1046.435 14120.955 1047.435 ;
    END
  END SET_VRESET_P[92]
  PIN SET_VRESET_P[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14260.675 1046.435 14260.955 1047.435 ;
    END
  END SET_VRESET_P[93]
  PIN SET_VRESET_P[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14400.675 1046.435 14400.955 1047.435 ;
    END
  END SET_VRESET_P[94]
  PIN SET_VRESET_P[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14540.675 1046.435 14540.955 1047.435 ;
    END
  END SET_VRESET_P[95]
  PIN SET_VRESET_P[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14680.675 1046.435 14680.955 1047.435 ;
    END
  END SET_VRESET_P[96]
  PIN SET_VRESET_P[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14820.675 1046.435 14820.955 1047.435 ;
    END
  END SET_VRESET_P[97]
  PIN SET_VRESET_P[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14960.675 1046.435 14960.955 1047.435 ;
    END
  END SET_VRESET_P[98]
  PIN SET_VH[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8097.035 1046.435 8097.315 1047.435 ;
    END
  END SET_VH[49]
  PIN SET_VH[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8237.035 1046.435 8237.315 1047.435 ;
    END
  END SET_VH[50]
  PIN SET_VH[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8377.035 1046.435 8377.315 1047.435 ;
    END
  END SET_VH[51]
  PIN SET_VH[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8517.035 1046.435 8517.315 1047.435 ;
    END
  END SET_VH[52]
  PIN SET_VH[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8657.035 1046.435 8657.315 1047.435 ;
    END
  END SET_VH[53]
  PIN SET_VH[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8797.035 1046.435 8797.315 1047.435 ;
    END
  END SET_VH[54]
  PIN SET_VH[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8937.035 1046.435 8937.315 1047.435 ;
    END
  END SET_VH[55]
  PIN SET_VH[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9077.035 1046.435 9077.315 1047.435 ;
    END
  END SET_VH[56]
  PIN SET_VH[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9217.035 1046.435 9217.315 1047.435 ;
    END
  END SET_VH[57]
  PIN SET_VH[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9357.035 1046.435 9357.315 1047.435 ;
    END
  END SET_VH[58]
  PIN SET_VH[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9497.035 1046.435 9497.315 1047.435 ;
    END
  END SET_VH[59]
  PIN SET_VH[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9637.035 1046.435 9637.315 1047.435 ;
    END
  END SET_VH[60]
  PIN SET_VH[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9777.035 1046.435 9777.315 1047.435 ;
    END
  END SET_VH[61]
  PIN SET_VH[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9917.035 1046.435 9917.315 1047.435 ;
    END
  END SET_VH[62]
  PIN SET_VH[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10057.035 1046.435 10057.315 1047.435 ;
    END
  END SET_VH[63]
  PIN SET_VH[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10197.035 1046.435 10197.315 1047.435 ;
    END
  END SET_VH[64]
  PIN SET_VH[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10337.035 1046.435 10337.315 1047.435 ;
    END
  END SET_VH[65]
  PIN SET_VH[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10477.035 1046.435 10477.315 1047.435 ;
    END
  END SET_VH[66]
  PIN SET_VH[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10617.035 1046.435 10617.315 1047.435 ;
    END
  END SET_VH[67]
  PIN SET_VH[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10757.035 1046.435 10757.315 1047.435 ;
    END
  END SET_VH[68]
  PIN SET_VH[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10897.035 1046.435 10897.315 1047.435 ;
    END
  END SET_VH[69]
  PIN SET_VH[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11037.035 1046.435 11037.315 1047.435 ;
    END
  END SET_VH[70]
  PIN SET_VH[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11177.035 1046.435 11177.315 1047.435 ;
    END
  END SET_VH[71]
  PIN SET_VH[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11317.035 1046.435 11317.315 1047.435 ;
    END
  END SET_VH[72]
  PIN SET_VH[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11457.035 1046.435 11457.315 1047.435 ;
    END
  END SET_VH[73]
  PIN SET_VH[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11597.035 1046.435 11597.315 1047.435 ;
    END
  END SET_VH[74]
  PIN SET_VH[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11737.035 1046.435 11737.315 1047.435 ;
    END
  END SET_VH[75]
  PIN SET_VH[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11877.035 1046.435 11877.315 1047.435 ;
    END
  END SET_VH[76]
  PIN SET_VH[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12017.035 1046.435 12017.315 1047.435 ;
    END
  END SET_VH[77]
  PIN SET_VH[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12157.035 1046.435 12157.315 1047.435 ;
    END
  END SET_VH[78]
  PIN SET_VH[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12297.035 1046.435 12297.315 1047.435 ;
    END
  END SET_VH[79]
  PIN SET_VH[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12437.035 1046.435 12437.315 1047.435 ;
    END
  END SET_VH[80]
  PIN SET_VH[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12577.035 1046.435 12577.315 1047.435 ;
    END
  END SET_VH[81]
  PIN SET_VH[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12717.035 1046.435 12717.315 1047.435 ;
    END
  END SET_VH[82]
  PIN SET_VH[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12857.035 1046.435 12857.315 1047.435 ;
    END
  END SET_VH[83]
  PIN SET_VH[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12997.035 1046.435 12997.315 1047.435 ;
    END
  END SET_VH[84]
  PIN SET_VH[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13137.035 1046.435 13137.315 1047.435 ;
    END
  END SET_VH[85]
  PIN SET_VH[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13277.035 1046.435 13277.315 1047.435 ;
    END
  END SET_VH[86]
  PIN SET_VH[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13417.035 1046.435 13417.315 1047.435 ;
    END
  END SET_VH[87]
  PIN SET_VH[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13557.035 1046.435 13557.315 1047.435 ;
    END
  END SET_VH[88]
  PIN SET_VH[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13697.035 1046.435 13697.315 1047.435 ;
    END
  END SET_VH[89]
  PIN SET_VH[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13837.035 1046.435 13837.315 1047.435 ;
    END
  END SET_VH[90]
  PIN SET_VH[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13977.035 1046.435 13977.315 1047.435 ;
    END
  END SET_VH[91]
  PIN SET_VH[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14117.035 1046.435 14117.315 1047.435 ;
    END
  END SET_VH[92]
  PIN SET_VH[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14257.035 1046.435 14257.315 1047.435 ;
    END
  END SET_VH[93]
  PIN SET_VH[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14397.035 1046.435 14397.315 1047.435 ;
    END
  END SET_VH[94]
  PIN SET_VH[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14537.035 1046.435 14537.315 1047.435 ;
    END
  END SET_VH[95]
  PIN SET_VH[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14677.035 1046.435 14677.315 1047.435 ;
    END
  END SET_VH[96]
  PIN SET_VH[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14817.035 1046.435 14817.315 1047.435 ;
    END
  END SET_VH[97]
  PIN SET_VH[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14957.035 1046.435 14957.315 1047.435 ;
    END
  END SET_VH[98]
  PIN SET_VH[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15097.035 1046.435 15097.315 1047.435 ;
    END
  END SET_VH[99]
  PIN SET_VH[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15237.035 1046.435 15237.315 1047.435 ;
    END
  END SET_VH[100]
  PIN SET_VH[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15377.035 1046.435 15377.315 1047.435 ;
    END
  END SET_VH[101]
  PIN SET_VH[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15517.035 1046.435 15517.315 1047.435 ;
    END
  END SET_VH[102]
  PIN SET_VH[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15657.035 1046.435 15657.315 1047.435 ;
    END
  END SET_VH[103]
  PIN SET_VH[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15797.035 1046.435 15797.315 1047.435 ;
    END
  END SET_VH[104]
  PIN SET_VH[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15937.035 1046.435 15937.315 1047.435 ;
    END
  END SET_VH[105]
  PIN SET_VH[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16077.035 1046.435 16077.315 1047.435 ;
    END
  END SET_VH[106]
  PIN SET_VH[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16217.035 1046.435 16217.315 1047.435 ;
    END
  END SET_VH[107]
  PIN SET_VH[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16357.035 1046.435 16357.315 1047.435 ;
    END
  END SET_VH[108]
  PIN SET_VH[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16497.035 1046.435 16497.315 1047.435 ;
    END
  END SET_VH[109]
  PIN SET_VH[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16637.035 1046.435 16637.315 1047.435 ;
    END
  END SET_VH[110]
  PIN SET_VH[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16777.035 1046.435 16777.315 1047.435 ;
    END
  END SET_VH[111]
  PIN SET_VH[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16917.035 1046.435 16917.315 1047.435 ;
    END
  END SET_VH[112]
  PIN SET_VH[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17057.035 1046.435 17057.315 1047.435 ;
    END
  END SET_VH[113]
  PIN SET_VH[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17197.035 1046.435 17197.315 1047.435 ;
    END
  END SET_VH[114]
  PIN SET_VH[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17337.035 1046.435 17337.315 1047.435 ;
    END
  END SET_VH[115]
  PIN SET_VH[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17477.035 1046.435 17477.315 1047.435 ;
    END
  END SET_VH[116]
  PIN SET_VH[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17617.035 1046.435 17617.315 1047.435 ;
    END
  END SET_VH[117]
  PIN SET_VH[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17757.035 1046.435 17757.315 1047.435 ;
    END
  END SET_VH[118]
  PIN SET_VH[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17897.035 1046.435 17897.315 1047.435 ;
    END
  END SET_VH[119]
  PIN SET_VH[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18037.035 1046.435 18037.315 1047.435 ;
    END
  END SET_VH[120]
  PIN SET_VH[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18177.035 1046.435 18177.315 1047.435 ;
    END
  END SET_VH[121]
  PIN SET_VH[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18317.035 1046.435 18317.315 1047.435 ;
    END
  END SET_VH[122]
  PIN SET_VH[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18457.035 1046.435 18457.315 1047.435 ;
    END
  END SET_VH[123]
  PIN SET_VH[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18597.035 1046.435 18597.315 1047.435 ;
    END
  END SET_VH[124]
  PIN SET_VH[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18737.035 1046.435 18737.315 1047.435 ;
    END
  END SET_VH[125]
  PIN SET_VH[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18877.035 1046.435 18877.315 1047.435 ;
    END
  END SET_VH[126]
  PIN SET_VH[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19017.035 1046.435 19017.315 1047.435 ;
    END
  END SET_VH[127]
  PIN SET_VRESET_P[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1240.675 1046.435 1240.955 1047.435 ;
    END
  END SET_VRESET_P[0]
  PIN SET_VRESET_P[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1380.675 1046.435 1380.955 1047.435 ;
    END
  END SET_VRESET_P[1]
  PIN SET_VRESET_P[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1520.675 1046.435 1520.955 1047.435 ;
    END
  END SET_VRESET_P[2]
  PIN SET_VRESET_P[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1660.675 1046.435 1660.955 1047.435 ;
    END
  END SET_VRESET_P[3]
  PIN SET_VRESET_P[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1800.675 1046.435 1800.955 1047.435 ;
    END
  END SET_VRESET_P[4]
  PIN SET_VRESET_P[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1940.675 1046.435 1940.955 1047.435 ;
    END
  END SET_VRESET_P[5]
  PIN SET_VRESET_P[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2080.675 1046.435 2080.955 1047.435 ;
    END
  END SET_VRESET_P[6]
  PIN SET_VRESET_P[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2220.675 1046.435 2220.955 1047.435 ;
    END
  END SET_VRESET_P[7]
  PIN SET_VRESET_P[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2360.675 1046.435 2360.955 1047.435 ;
    END
  END SET_VRESET_P[8]
  PIN SET_VRESET_P[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2500.675 1046.435 2500.955 1047.435 ;
    END
  END SET_VRESET_P[9]
  PIN SET_VRESET_P[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2640.675 1046.435 2640.955 1047.435 ;
    END
  END SET_VRESET_P[10]
  PIN SET_VRESET_P[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2780.675 1046.435 2780.955 1047.435 ;
    END
  END SET_VRESET_P[11]
  PIN SET_VRESET_P[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2920.675 1046.435 2920.955 1047.435 ;
    END
  END SET_VRESET_P[12]
  PIN SET_VRESET_P[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3060.675 1046.435 3060.955 1047.435 ;
    END
  END SET_VRESET_P[13]
  PIN SET_VRESET_P[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3200.675 1046.435 3200.955 1047.435 ;
    END
  END SET_VRESET_P[14]
  PIN SET_VRESET_P[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3340.675 1046.435 3340.955 1047.435 ;
    END
  END SET_VRESET_P[15]
  PIN SET_VRESET_P[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3480.675 1046.435 3480.955 1047.435 ;
    END
  END SET_VRESET_P[16]
  PIN SET_VRESET_P[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3620.675 1046.435 3620.955 1047.435 ;
    END
  END SET_VRESET_P[17]
  PIN SET_VRESET_P[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3760.675 1046.435 3760.955 1047.435 ;
    END
  END SET_VRESET_P[18]
  PIN SET_VRESET_P[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3900.675 1046.435 3900.955 1047.435 ;
    END
  END SET_VRESET_P[19]
  PIN SET_VRESET_P[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4040.675 1046.435 4040.955 1047.435 ;
    END
  END SET_VRESET_P[20]
  PIN SET_VRESET_P[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4180.675 1046.435 4180.955 1047.435 ;
    END
  END SET_VRESET_P[21]
  PIN SET_VRESET_P[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4320.675 1046.435 4320.955 1047.435 ;
    END
  END SET_VRESET_P[22]
  PIN SET_VRESET_P[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4460.675 1046.435 4460.955 1047.435 ;
    END
  END SET_VRESET_P[23]
  PIN SET_VRESET_P[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4600.675 1046.435 4600.955 1047.435 ;
    END
  END SET_VRESET_P[24]
  PIN SET_VRESET_P[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4740.675 1046.435 4740.955 1047.435 ;
    END
  END SET_VRESET_P[25]
  PIN SET_VRESET_P[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4880.675 1046.435 4880.955 1047.435 ;
    END
  END SET_VRESET_P[26]
  PIN SET_VRESET_P[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5020.675 1046.435 5020.955 1047.435 ;
    END
  END SET_VRESET_P[27]
  PIN SET_VRESET_P[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5160.675 1046.435 5160.955 1047.435 ;
    END
  END SET_VRESET_P[28]
  PIN SET_VRESET_P[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5300.675 1046.435 5300.955 1047.435 ;
    END
  END SET_VRESET_P[29]
  PIN SET_VRESET_P[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5440.675 1046.435 5440.955 1047.435 ;
    END
  END SET_VRESET_P[30]
  PIN SET_VRESET_P[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5580.675 1046.435 5580.955 1047.435 ;
    END
  END SET_VRESET_P[31]
  PIN SET_VRESET_P[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5720.675 1046.435 5720.955 1047.435 ;
    END
  END SET_VRESET_P[32]
  PIN SET_VRESET_P[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5860.675 1046.435 5860.955 1047.435 ;
    END
  END SET_VRESET_P[33]
  PIN SET_VRESET_P[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6000.675 1046.435 6000.955 1047.435 ;
    END
  END SET_VRESET_P[34]
  PIN SET_VRESET_P[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6140.675 1046.435 6140.955 1047.435 ;
    END
  END SET_VRESET_P[35]
  PIN SET_VRESET_P[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6280.675 1046.435 6280.955 1047.435 ;
    END
  END SET_VRESET_P[36]
  PIN SET_VRESET_P[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6420.675 1046.435 6420.955 1047.435 ;
    END
  END SET_VRESET_P[37]
  PIN SET_VCASN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1247.955 1046.435 1248.235 1047.435 ;
    END
  END SET_VCASN[0]
  PIN SET_VCASN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1387.955 1046.435 1388.235 1047.435 ;
    END
  END SET_VCASN[1]
  PIN SET_VCASN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1527.955 1046.435 1528.235 1047.435 ;
    END
  END SET_VCASN[2]
  PIN SET_VCASN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1667.955 1046.435 1668.235 1047.435 ;
    END
  END SET_VCASN[3]
  PIN SET_VCASN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1807.955 1046.435 1808.235 1047.435 ;
    END
  END SET_VCASN[4]
  PIN SET_VCASN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1947.955 1046.435 1948.235 1047.435 ;
    END
  END SET_VCASN[5]
  PIN SET_VCASN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2087.955 1046.435 2088.235 1047.435 ;
    END
  END SET_VCASN[6]
  PIN SET_VCASN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2227.955 1046.435 2228.235 1047.435 ;
    END
  END SET_VCASN[7]
  PIN SET_VCASN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2367.955 1046.435 2368.235 1047.435 ;
    END
  END SET_VCASN[8]
  PIN SET_VCASN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2507.955 1046.435 2508.235 1047.435 ;
    END
  END SET_VCASN[9]
  PIN SET_VCASN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2647.955 1046.435 2648.235 1047.435 ;
    END
  END SET_VCASN[10]
  PIN SET_VCASN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2787.955 1046.435 2788.235 1047.435 ;
    END
  END SET_VCASN[11]
  PIN SET_VCASN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2927.955 1046.435 2928.235 1047.435 ;
    END
  END SET_VCASN[12]
  PIN SET_VCASN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3067.955 1046.435 3068.235 1047.435 ;
    END
  END SET_VCASN[13]
  PIN SET_VCASN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3207.955 1046.435 3208.235 1047.435 ;
    END
  END SET_VCASN[14]
  PIN SET_VCASN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3347.955 1046.435 3348.235 1047.435 ;
    END
  END SET_VCASN[15]
  PIN SET_VCASN[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3487.955 1046.435 3488.235 1047.435 ;
    END
  END SET_VCASN[16]
  PIN SET_VCASN[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3627.955 1046.435 3628.235 1047.435 ;
    END
  END SET_VCASN[17]
  PIN SET_VCASN[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3767.955 1046.435 3768.235 1047.435 ;
    END
  END SET_VCASN[18]
  PIN SET_VCASN[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3907.955 1046.435 3908.235 1047.435 ;
    END
  END SET_VCASN[19]
  PIN SET_VCASN[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4047.955 1046.435 4048.235 1047.435 ;
    END
  END SET_VCASN[20]
  PIN SET_VCASN[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4187.955 1046.435 4188.235 1047.435 ;
    END
  END SET_VCASN[21]
  PIN SET_VCASN[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4327.955 1046.435 4328.235 1047.435 ;
    END
  END SET_VCASN[22]
  PIN SET_VCASN[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4467.955 1046.435 4468.235 1047.435 ;
    END
  END SET_VCASN[23]
  PIN SET_VCASN[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4607.955 1046.435 4608.235 1047.435 ;
    END
  END SET_VCASN[24]
  PIN SET_VCASN[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4747.955 1046.435 4748.235 1047.435 ;
    END
  END SET_VCASN[25]
  PIN SET_VCASN[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4887.955 1046.435 4888.235 1047.435 ;
    END
  END SET_VCASN[26]
  PIN SET_VCASN[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5027.955 1046.435 5028.235 1047.435 ;
    END
  END SET_VCASN[27]
  PIN SET_VCASN[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5167.955 1046.435 5168.235 1047.435 ;
    END
  END SET_VCASN[28]
  PIN SET_VCASN[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5307.955 1046.435 5308.235 1047.435 ;
    END
  END SET_VCASN[29]
  PIN SET_VCASN[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5447.955 1046.435 5448.235 1047.435 ;
    END
  END SET_VCASN[30]
  PIN SET_VCASN[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5587.955 1046.435 5588.235 1047.435 ;
    END
  END SET_VCASN[31]
  PIN SET_VCASN[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5727.955 1046.435 5728.235 1047.435 ;
    END
  END SET_VCASN[32]
  PIN SET_VCASN[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5867.955 1046.435 5868.235 1047.435 ;
    END
  END SET_VCASN[33]
  PIN SET_VCASN[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6007.955 1046.435 6008.235 1047.435 ;
    END
  END SET_VCASN[34]
  PIN SET_VCASN[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6147.955 1046.435 6148.235 1047.435 ;
    END
  END SET_VCASN[35]
  PIN SET_VCASN[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6287.955 1046.435 6288.235 1047.435 ;
    END
  END SET_VCASN[36]
  PIN SET_VCASN[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6427.955 1046.435 6428.235 1047.435 ;
    END
  END SET_VCASN[37]
  PIN SET_VCASN[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6567.955 1046.435 6568.235 1047.435 ;
    END
  END SET_VCASN[38]
  PIN SET_VCASN[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6707.955 1046.435 6708.235 1047.435 ;
    END
  END SET_VCASN[39]
  PIN SET_VCASN[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6847.955 1046.435 6848.235 1047.435 ;
    END
  END SET_VCASN[40]
  PIN SET_VCASN[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6987.955 1046.435 6988.235 1047.435 ;
    END
  END SET_VCASN[41]
  PIN SET_VCASN[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7127.955 1046.435 7128.235 1047.435 ;
    END
  END SET_VCASN[42]
  PIN SET_VCASN[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7267.955 1046.435 7268.235 1047.435 ;
    END
  END SET_VCASN[43]
  PIN SET_VCASN[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7407.955 1046.435 7408.235 1047.435 ;
    END
  END SET_VCASN[44]
  PIN SET_VCASN[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7547.955 1046.435 7548.235 1047.435 ;
    END
  END SET_VCASN[45]
  PIN SET_VCASN[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7687.955 1046.435 7688.235 1047.435 ;
    END
  END SET_VCASN[46]
  PIN SET_VCASN[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7827.955 1046.435 7828.235 1047.435 ;
    END
  END SET_VCASN[47]
  PIN SET_VCASN[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7967.955 1046.435 7968.235 1047.435 ;
    END
  END SET_VCASN[48]
  PIN SET_VCASN[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8107.955 1046.435 8108.235 1047.435 ;
    END
  END SET_VCASN[49]
  PIN SET_VCASN[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8247.955 1046.435 8248.235 1047.435 ;
    END
  END SET_VCASN[50]
  PIN SET_VCASN[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8387.955 1046.435 8388.235 1047.435 ;
    END
  END SET_VCASN[51]
  PIN SET_VCASN[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8527.955 1046.435 8528.235 1047.435 ;
    END
  END SET_VCASN[52]
  PIN SET_VCASN[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8667.955 1046.435 8668.235 1047.435 ;
    END
  END SET_VCASN[53]
  PIN SET_VCASN[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8807.955 1046.435 8808.235 1047.435 ;
    END
  END SET_VCASN[54]
  PIN SET_VCASN[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8947.955 1046.435 8948.235 1047.435 ;
    END
  END SET_VCASN[55]
  PIN SET_VCASN[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9087.955 1046.435 9088.235 1047.435 ;
    END
  END SET_VCASN[56]
  PIN SET_VCASN[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9227.955 1046.435 9228.235 1047.435 ;
    END
  END SET_VCASN[57]
  PIN SET_VCASN[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9367.955 1046.435 9368.235 1047.435 ;
    END
  END SET_VCASN[58]
  PIN SET_VCASN[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9507.955 1046.435 9508.235 1047.435 ;
    END
  END SET_VCASN[59]
  PIN SET_VCASN[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9647.955 1046.435 9648.235 1047.435 ;
    END
  END SET_VCASN[60]
  PIN SET_VCASN[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9787.955 1046.435 9788.235 1047.435 ;
    END
  END SET_VCASN[61]
  PIN SET_VCASN[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9927.955 1046.435 9928.235 1047.435 ;
    END
  END SET_VCASN[62]
  PIN SET_VCASN[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10067.955 1046.435 10068.235 1047.435 ;
    END
  END SET_VCASN[63]
  PIN SET_VCASN[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10207.955 1046.435 10208.235 1047.435 ;
    END
  END SET_VCASN[64]
  PIN SET_VCASN[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10347.955 1046.435 10348.235 1047.435 ;
    END
  END SET_VCASN[65]
  PIN SET_VCASN[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10487.955 1046.435 10488.235 1047.435 ;
    END
  END SET_VCASN[66]
  PIN SET_VCASN[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10627.955 1046.435 10628.235 1047.435 ;
    END
  END SET_VCASN[67]
  PIN SET_VCASN[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10767.955 1046.435 10768.235 1047.435 ;
    END
  END SET_VCASN[68]
  PIN SET_VCASN[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10907.955 1046.435 10908.235 1047.435 ;
    END
  END SET_VCASN[69]
  PIN SET_VCASN[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11047.955 1046.435 11048.235 1047.435 ;
    END
  END SET_VCASN[70]
  PIN SET_VCASN[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11187.955 1046.435 11188.235 1047.435 ;
    END
  END SET_VCASN[71]
  PIN SET_VCASN[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11327.955 1046.435 11328.235 1047.435 ;
    END
  END SET_VCASN[72]
  PIN SET_VCASN[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11467.955 1046.435 11468.235 1047.435 ;
    END
  END SET_VCASN[73]
  PIN SET_VCASN[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11607.955 1046.435 11608.235 1047.435 ;
    END
  END SET_VCASN[74]
  PIN SET_VCASN[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11747.955 1046.435 11748.235 1047.435 ;
    END
  END SET_VCASN[75]
  PIN SET_VCASN[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11887.955 1046.435 11888.235 1047.435 ;
    END
  END SET_VCASN[76]
  PIN SET_VCASN[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12027.955 1046.435 12028.235 1047.435 ;
    END
  END SET_VCASN[77]
  PIN SET_VCASN[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12167.955 1046.435 12168.235 1047.435 ;
    END
  END SET_VCASN[78]
  PIN SET_VCASN[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12307.955 1046.435 12308.235 1047.435 ;
    END
  END SET_VCASN[79]
  PIN SET_VCASN[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12447.955 1046.435 12448.235 1047.435 ;
    END
  END SET_VCASN[80]
  PIN SET_VCASN[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12587.955 1046.435 12588.235 1047.435 ;
    END
  END SET_VCASN[81]
  PIN SET_VCASN[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12727.955 1046.435 12728.235 1047.435 ;
    END
  END SET_VCASN[82]
  PIN SET_VCASN[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12867.955 1046.435 12868.235 1047.435 ;
    END
  END SET_VCASN[83]
  PIN SET_VCASN[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13007.955 1046.435 13008.235 1047.435 ;
    END
  END SET_VCASN[84]
  PIN SET_VCASN[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13147.955 1046.435 13148.235 1047.435 ;
    END
  END SET_VCASN[85]
  PIN SET_VCASN[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13287.955 1046.435 13288.235 1047.435 ;
    END
  END SET_VCASN[86]
  PIN SET_ICASN[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18950.675 1046.435 18950.955 1047.435 ;
    END
  END SET_ICASN[127]
  PIN SET_VRESET_D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1229.755 1046.435 1230.035 1047.435 ;
    END
  END SET_VRESET_D[0]
  PIN SET_VRESET_D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1369.755 1046.435 1370.035 1047.435 ;
    END
  END SET_VRESET_D[1]
  PIN SET_VRESET_D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1509.755 1046.435 1510.035 1047.435 ;
    END
  END SET_VRESET_D[2]
  PIN SET_VRESET_D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1649.755 1046.435 1650.035 1047.435 ;
    END
  END SET_VRESET_D[3]
  PIN SET_VRESET_D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1789.755 1046.435 1790.035 1047.435 ;
    END
  END SET_VRESET_D[4]
  PIN SET_VRESET_D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1929.755 1046.435 1930.035 1047.435 ;
    END
  END SET_VRESET_D[5]
  PIN SET_VRESET_D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2069.755 1046.435 2070.035 1047.435 ;
    END
  END SET_VRESET_D[6]
  PIN SET_VRESET_D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2209.755 1046.435 2210.035 1047.435 ;
    END
  END SET_VRESET_D[7]
  PIN SET_VRESET_D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2349.755 1046.435 2350.035 1047.435 ;
    END
  END SET_VRESET_D[8]
  PIN SET_VRESET_D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2489.755 1046.435 2490.035 1047.435 ;
    END
  END SET_VRESET_D[9]
  PIN SET_VRESET_D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2629.755 1046.435 2630.035 1047.435 ;
    END
  END SET_VRESET_D[10]
  PIN SET_VRESET_D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2769.755 1046.435 2770.035 1047.435 ;
    END
  END SET_VRESET_D[11]
  PIN SET_VRESET_D[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2909.755 1046.435 2910.035 1047.435 ;
    END
  END SET_VRESET_D[12]
  PIN SET_VRESET_D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3049.755 1046.435 3050.035 1047.435 ;
    END
  END SET_VRESET_D[13]
  PIN SET_VRESET_D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3189.755 1046.435 3190.035 1047.435 ;
    END
  END SET_VRESET_D[14]
  PIN SET_VRESET_D[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3329.755 1046.435 3330.035 1047.435 ;
    END
  END SET_VRESET_D[15]
  PIN SET_VRESET_D[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3469.755 1046.435 3470.035 1047.435 ;
    END
  END SET_VRESET_D[16]
  PIN SET_VRESET_D[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3609.755 1046.435 3610.035 1047.435 ;
    END
  END SET_VRESET_D[17]
  PIN SET_VRESET_D[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3749.755 1046.435 3750.035 1047.435 ;
    END
  END SET_VRESET_D[18]
  PIN SET_VRESET_D[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3889.755 1046.435 3890.035 1047.435 ;
    END
  END SET_VRESET_D[19]
  PIN SET_VRESET_D[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4029.755 1046.435 4030.035 1047.435 ;
    END
  END SET_VRESET_D[20]
  PIN SET_VRESET_D[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4169.755 1046.435 4170.035 1047.435 ;
    END
  END SET_VRESET_D[21]
  PIN SET_VRESET_D[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4309.755 1046.435 4310.035 1047.435 ;
    END
  END SET_VRESET_D[22]
  PIN SET_VRESET_D[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4449.755 1046.435 4450.035 1047.435 ;
    END
  END SET_VRESET_D[23]
  PIN SET_VRESET_D[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4589.755 1046.435 4590.035 1047.435 ;
    END
  END SET_VRESET_D[24]
  PIN SET_VRESET_D[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4729.755 1046.435 4730.035 1047.435 ;
    END
  END SET_VRESET_D[25]
  PIN SET_VRESET_D[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4869.755 1046.435 4870.035 1047.435 ;
    END
  END SET_VRESET_D[26]
  PIN SET_VRESET_D[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5009.755 1046.435 5010.035 1047.435 ;
    END
  END SET_VRESET_D[27]
  PIN SET_VRESET_D[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5149.755 1046.435 5150.035 1047.435 ;
    END
  END SET_VRESET_D[28]
  PIN SET_VRESET_D[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5289.755 1046.435 5290.035 1047.435 ;
    END
  END SET_VRESET_D[29]
  PIN SET_VRESET_D[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5429.755 1046.435 5430.035 1047.435 ;
    END
  END SET_VRESET_D[30]
  PIN SET_VRESET_D[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5569.755 1046.435 5570.035 1047.435 ;
    END
  END SET_VRESET_D[31]
  PIN SET_VRESET_D[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5709.755 1046.435 5710.035 1047.435 ;
    END
  END SET_VRESET_D[32]
  PIN SET_VRESET_D[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5849.755 1046.435 5850.035 1047.435 ;
    END
  END SET_VRESET_D[33]
  PIN SET_VRESET_D[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5989.755 1046.435 5990.035 1047.435 ;
    END
  END SET_VRESET_D[34]
  PIN SET_VRESET_D[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6129.755 1046.435 6130.035 1047.435 ;
    END
  END SET_VRESET_D[35]
  PIN SET_VRESET_D[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6269.755 1046.435 6270.035 1047.435 ;
    END
  END SET_VRESET_D[36]
  PIN SET_VRESET_D[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6409.755 1046.435 6410.035 1047.435 ;
    END
  END SET_VRESET_D[37]
  PIN SET_VRESET_D[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6549.755 1046.435 6550.035 1047.435 ;
    END
  END SET_VRESET_D[38]
  PIN SET_VRESET_D[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6689.755 1046.435 6690.035 1047.435 ;
    END
  END SET_VRESET_D[39]
  PIN SET_VRESET_D[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6829.755 1046.435 6830.035 1047.435 ;
    END
  END SET_VRESET_D[40]
  PIN SET_VRESET_D[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6969.755 1046.435 6970.035 1047.435 ;
    END
  END SET_VRESET_D[41]
  PIN SET_VRESET_D[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7109.755 1046.435 7110.035 1047.435 ;
    END
  END SET_VRESET_D[42]
  PIN SET_VRESET_D[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7249.755 1046.435 7250.035 1047.435 ;
    END
  END SET_VRESET_D[43]
  PIN SET_VRESET_D[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7389.755 1046.435 7390.035 1047.435 ;
    END
  END SET_VRESET_D[44]
  PIN SET_VRESET_D[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7529.755 1046.435 7530.035 1047.435 ;
    END
  END SET_VRESET_D[45]
  PIN SET_VRESET_D[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7669.755 1046.435 7670.035 1047.435 ;
    END
  END SET_VRESET_D[46]
  PIN SET_VRESET_D[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7809.755 1046.435 7810.035 1047.435 ;
    END
  END SET_VRESET_D[47]
  PIN SET_VRESET_D[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7949.755 1046.435 7950.035 1047.435 ;
    END
  END SET_VRESET_D[48]
  PIN SET_VRESET_D[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8089.755 1046.435 8090.035 1047.435 ;
    END
  END SET_VRESET_D[49]
  PIN SET_VRESET_D[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8229.755 1046.435 8230.035 1047.435 ;
    END
  END SET_VRESET_D[50]
  PIN SET_VRESET_D[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8369.755 1046.435 8370.035 1047.435 ;
    END
  END SET_VRESET_D[51]
  PIN SET_VRESET_D[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8509.755 1046.435 8510.035 1047.435 ;
    END
  END SET_VRESET_D[52]
  PIN SET_VRESET_D[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8649.755 1046.435 8650.035 1047.435 ;
    END
  END SET_VRESET_D[53]
  PIN SET_VRESET_D[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8789.755 1046.435 8790.035 1047.435 ;
    END
  END SET_VRESET_D[54]
  PIN SET_VRESET_D[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8929.755 1046.435 8930.035 1047.435 ;
    END
  END SET_VRESET_D[55]
  PIN SET_VRESET_D[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9069.755 1046.435 9070.035 1047.435 ;
    END
  END SET_VRESET_D[56]
  PIN SET_VRESET_D[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9209.755 1046.435 9210.035 1047.435 ;
    END
  END SET_VRESET_D[57]
  PIN SET_VRESET_D[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9349.755 1046.435 9350.035 1047.435 ;
    END
  END SET_VRESET_D[58]
  PIN SET_VRESET_D[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9489.755 1046.435 9490.035 1047.435 ;
    END
  END SET_VRESET_D[59]
  PIN SET_VRESET_D[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9629.755 1046.435 9630.035 1047.435 ;
    END
  END SET_VRESET_D[60]
  PIN SET_VRESET_D[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9769.755 1046.435 9770.035 1047.435 ;
    END
  END SET_VRESET_D[61]
  PIN SET_VRESET_D[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9909.755 1046.435 9910.035 1047.435 ;
    END
  END SET_VRESET_D[62]
  PIN SET_VRESET_D[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10049.755 1046.435 10050.035 1047.435 ;
    END
  END SET_VRESET_D[63]
  PIN SET_VRESET_D[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10189.755 1046.435 10190.035 1047.435 ;
    END
  END SET_VRESET_D[64]
  PIN SET_VRESET_D[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10329.755 1046.435 10330.035 1047.435 ;
    END
  END SET_VRESET_D[65]
  PIN SET_VRESET_D[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10469.755 1046.435 10470.035 1047.435 ;
    END
  END SET_VRESET_D[66]
  PIN SET_VRESET_D[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10609.755 1046.435 10610.035 1047.435 ;
    END
  END SET_VRESET_D[67]
  PIN SET_VRESET_D[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10749.755 1046.435 10750.035 1047.435 ;
    END
  END SET_VRESET_D[68]
  PIN SET_VRESET_D[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10889.755 1046.435 10890.035 1047.435 ;
    END
  END SET_VRESET_D[69]
  PIN SET_VRESET_D[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11029.755 1046.435 11030.035 1047.435 ;
    END
  END SET_VRESET_D[70]
  PIN SET_VRESET_D[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11169.755 1046.435 11170.035 1047.435 ;
    END
  END SET_VRESET_D[71]
  PIN SET_VRESET_D[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11309.755 1046.435 11310.035 1047.435 ;
    END
  END SET_VRESET_D[72]
  PIN SET_VRESET_D[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11449.755 1046.435 11450.035 1047.435 ;
    END
  END SET_VRESET_D[73]
  PIN SET_VRESET_D[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11589.755 1046.435 11590.035 1047.435 ;
    END
  END SET_VRESET_D[74]
  PIN SET_VRESET_D[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11729.755 1046.435 11730.035 1047.435 ;
    END
  END SET_VRESET_D[75]
  PIN SET_VRESET_D[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11869.755 1046.435 11870.035 1047.435 ;
    END
  END SET_VRESET_D[76]
  PIN SET_VRESET_D[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12009.755 1046.435 12010.035 1047.435 ;
    END
  END SET_VRESET_D[77]
  PIN SET_VRESET_D[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12149.755 1046.435 12150.035 1047.435 ;
    END
  END SET_VRESET_D[78]
  PIN SET_VRESET_D[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12289.755 1046.435 12290.035 1047.435 ;
    END
  END SET_VRESET_D[79]
  PIN SET_VRESET_D[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12429.755 1046.435 12430.035 1047.435 ;
    END
  END SET_VRESET_D[80]
  PIN SET_VRESET_D[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12569.755 1046.435 12570.035 1047.435 ;
    END
  END SET_VRESET_D[81]
  PIN SET_VRESET_D[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12709.755 1046.435 12710.035 1047.435 ;
    END
  END SET_VRESET_D[82]
  PIN SET_VRESET_D[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12849.755 1046.435 12850.035 1047.435 ;
    END
  END SET_VRESET_D[83]
  PIN SET_VRESET_D[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12989.755 1046.435 12990.035 1047.435 ;
    END
  END SET_VRESET_D[84]
  PIN SET_VRESET_D[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13129.755 1046.435 13130.035 1047.435 ;
    END
  END SET_VRESET_D[85]
  PIN SET_VRESET_D[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13269.755 1046.435 13270.035 1047.435 ;
    END
  END SET_VRESET_D[86]
  PIN SET_VRESET_D[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13409.755 1046.435 13410.035 1047.435 ;
    END
  END SET_VRESET_D[87]
  PIN SET_VRESET_D[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13549.755 1046.435 13550.035 1047.435 ;
    END
  END SET_VRESET_D[88]
  PIN SET_VRESET_D[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13689.755 1046.435 13690.035 1047.435 ;
    END
  END SET_VRESET_D[89]
  PIN SET_VRESET_D[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13829.755 1046.435 13830.035 1047.435 ;
    END
  END SET_VRESET_D[90]
  PIN SET_VRESET_D[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13969.755 1046.435 13970.035 1047.435 ;
    END
  END SET_VRESET_D[91]
  PIN SET_VRESET_D[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14109.755 1046.435 14110.035 1047.435 ;
    END
  END SET_VRESET_D[92]
  PIN SET_VRESET_D[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14249.755 1046.435 14250.035 1047.435 ;
    END
  END SET_VRESET_D[93]
  PIN SET_VRESET_D[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14389.755 1046.435 14390.035 1047.435 ;
    END
  END SET_VRESET_D[94]
  PIN SET_VRESET_D[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14529.755 1046.435 14530.035 1047.435 ;
    END
  END SET_VRESET_D[95]
  PIN SET_VRESET_D[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14669.755 1046.435 14670.035 1047.435 ;
    END
  END SET_VRESET_D[96]
  PIN SET_VRESET_D[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14809.755 1046.435 14810.035 1047.435 ;
    END
  END SET_VRESET_D[97]
  PIN SET_VRESET_D[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14949.755 1046.435 14950.035 1047.435 ;
    END
  END SET_VRESET_D[98]
  PIN SET_VRESET_D[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15089.755 1046.435 15090.035 1047.435 ;
    END
  END SET_VRESET_D[99]
  PIN SET_VRESET_D[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15229.755 1046.435 15230.035 1047.435 ;
    END
  END SET_VRESET_D[100]
  PIN SET_VL[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11733.395 1046.435 11733.675 1047.435 ;
    END
  END SET_VL[75]
  PIN SET_VL[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11873.395 1046.435 11873.675 1047.435 ;
    END
  END SET_VL[76]
  PIN SET_VL[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12013.395 1046.435 12013.675 1047.435 ;
    END
  END SET_VL[77]
  PIN SET_VL[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12153.395 1046.435 12153.675 1047.435 ;
    END
  END SET_VL[78]
  PIN SET_VL[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12293.395 1046.435 12293.675 1047.435 ;
    END
  END SET_VL[79]
  PIN SET_VL[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12433.395 1046.435 12433.675 1047.435 ;
    END
  END SET_VL[80]
  PIN SET_VL[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12573.395 1046.435 12573.675 1047.435 ;
    END
  END SET_VL[81]
  PIN SET_VL[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12713.395 1046.435 12713.675 1047.435 ;
    END
  END SET_VL[82]
  PIN SET_VL[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12853.395 1046.435 12853.675 1047.435 ;
    END
  END SET_VL[83]
  PIN SET_VL[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12993.395 1046.435 12993.675 1047.435 ;
    END
  END SET_VL[84]
  PIN SET_VL[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13133.395 1046.435 13133.675 1047.435 ;
    END
  END SET_VL[85]
  PIN SET_VL[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13273.395 1046.435 13273.675 1047.435 ;
    END
  END SET_VL[86]
  PIN SET_VL[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13413.395 1046.435 13413.675 1047.435 ;
    END
  END SET_VL[87]
  PIN SET_VL[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13553.395 1046.435 13553.675 1047.435 ;
    END
  END SET_VL[88]
  PIN SET_VL[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13693.395 1046.435 13693.675 1047.435 ;
    END
  END SET_VL[89]
  PIN SET_VL[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13833.395 1046.435 13833.675 1047.435 ;
    END
  END SET_VL[90]
  PIN SET_VL[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13973.395 1046.435 13973.675 1047.435 ;
    END
  END SET_VL[91]
  PIN SET_VL[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14113.395 1046.435 14113.675 1047.435 ;
    END
  END SET_VL[92]
  PIN SET_VL[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14253.395 1046.435 14253.675 1047.435 ;
    END
  END SET_VL[93]
  PIN SET_VL[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14393.395 1046.435 14393.675 1047.435 ;
    END
  END SET_VL[94]
  PIN SET_VL[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14533.395 1046.435 14533.675 1047.435 ;
    END
  END SET_VL[95]
  PIN SET_VL[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14673.395 1046.435 14673.675 1047.435 ;
    END
  END SET_VL[96]
  PIN SET_VL[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14813.395 1046.435 14813.675 1047.435 ;
    END
  END SET_VL[97]
  PIN SET_VL[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14953.395 1046.435 14953.675 1047.435 ;
    END
  END SET_VL[98]
  PIN SET_VL[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15093.395 1046.435 15093.675 1047.435 ;
    END
  END SET_VL[99]
  PIN SET_VL[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15233.395 1046.435 15233.675 1047.435 ;
    END
  END SET_VL[100]
  PIN SET_VL[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15373.395 1046.435 15373.675 1047.435 ;
    END
  END SET_VL[101]
  PIN SET_VL[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15513.395 1046.435 15513.675 1047.435 ;
    END
  END SET_VL[102]
  PIN SET_VL[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15653.395 1046.435 15653.675 1047.435 ;
    END
  END SET_VL[103]
  PIN SET_VL[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15793.395 1046.435 15793.675 1047.435 ;
    END
  END SET_VL[104]
  PIN SET_VL[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15933.395 1046.435 15933.675 1047.435 ;
    END
  END SET_VL[105]
  PIN SET_VL[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16073.395 1046.435 16073.675 1047.435 ;
    END
  END SET_VL[106]
  PIN SET_VL[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16213.395 1046.435 16213.675 1047.435 ;
    END
  END SET_VL[107]
  PIN SET_VL[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16353.395 1046.435 16353.675 1047.435 ;
    END
  END SET_VL[108]
  PIN SET_VL[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16493.395 1046.435 16493.675 1047.435 ;
    END
  END SET_VL[109]
  PIN SET_VL[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16633.395 1046.435 16633.675 1047.435 ;
    END
  END SET_VL[110]
  PIN SET_VL[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16773.395 1046.435 16773.675 1047.435 ;
    END
  END SET_VL[111]
  PIN SET_VL[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16913.395 1046.435 16913.675 1047.435 ;
    END
  END SET_VL[112]
  PIN SET_VL[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17053.395 1046.435 17053.675 1047.435 ;
    END
  END SET_VL[113]
  PIN SET_VL[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17193.395 1046.435 17193.675 1047.435 ;
    END
  END SET_VL[114]
  PIN SET_VL[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17333.395 1046.435 17333.675 1047.435 ;
    END
  END SET_VL[115]
  PIN SET_VL[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17473.395 1046.435 17473.675 1047.435 ;
    END
  END SET_VL[116]
  PIN SET_VL[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17613.395 1046.435 17613.675 1047.435 ;
    END
  END SET_VL[117]
  PIN SET_VL[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17753.395 1046.435 17753.675 1047.435 ;
    END
  END SET_VL[118]
  PIN SET_VL[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17893.395 1046.435 17893.675 1047.435 ;
    END
  END SET_VL[119]
  PIN SET_VL[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18033.395 1046.435 18033.675 1047.435 ;
    END
  END SET_VL[120]
  PIN SET_VL[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18173.395 1046.435 18173.675 1047.435 ;
    END
  END SET_VL[121]
  PIN SET_VL[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18313.395 1046.435 18313.675 1047.435 ;
    END
  END SET_VL[122]
  PIN SET_VL[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18453.395 1046.435 18453.675 1047.435 ;
    END
  END SET_VL[123]
  PIN SET_VL[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18593.395 1046.435 18593.675 1047.435 ;
    END
  END SET_VL[124]
  PIN SET_VL[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18733.395 1046.435 18733.675 1047.435 ;
    END
  END SET_VL[125]
  PIN SET_VL[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18873.395 1046.435 18873.675 1047.435 ;
    END
  END SET_VL[126]
  PIN SET_VL[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19013.395 1046.435 19013.675 1047.435 ;
    END
  END SET_VL[127]
  PIN SET_VH[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1237.035 1046.435 1237.315 1047.435 ;
    END
  END SET_VH[0]
  PIN SET_VH[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1377.035 1046.435 1377.315 1047.435 ;
    END
  END SET_VH[1]
  PIN SET_VH[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1517.035 1046.435 1517.315 1047.435 ;
    END
  END SET_VH[2]
  PIN SET_VH[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1657.035 1046.435 1657.315 1047.435 ;
    END
  END SET_VH[3]
  PIN SET_VH[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1797.035 1046.435 1797.315 1047.435 ;
    END
  END SET_VH[4]
  PIN SET_VH[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1937.035 1046.435 1937.315 1047.435 ;
    END
  END SET_VH[5]
  PIN SET_VH[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2077.035 1046.435 2077.315 1047.435 ;
    END
  END SET_VH[6]
  PIN SET_VH[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2217.035 1046.435 2217.315 1047.435 ;
    END
  END SET_VH[7]
  PIN SET_VH[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2357.035 1046.435 2357.315 1047.435 ;
    END
  END SET_VH[8]
  PIN SET_VH[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2497.035 1046.435 2497.315 1047.435 ;
    END
  END SET_VH[9]
  PIN SET_VH[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2637.035 1046.435 2637.315 1047.435 ;
    END
  END SET_VH[10]
  PIN SET_VH[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2777.035 1046.435 2777.315 1047.435 ;
    END
  END SET_VH[11]
  PIN SET_VH[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2917.035 1046.435 2917.315 1047.435 ;
    END
  END SET_VH[12]
  PIN SET_VH[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3057.035 1046.435 3057.315 1047.435 ;
    END
  END SET_VH[13]
  PIN SET_VH[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3197.035 1046.435 3197.315 1047.435 ;
    END
  END SET_VH[14]
  PIN SET_VH[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3337.035 1046.435 3337.315 1047.435 ;
    END
  END SET_VH[15]
  PIN SET_VH[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3477.035 1046.435 3477.315 1047.435 ;
    END
  END SET_VH[16]
  PIN SET_VH[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3617.035 1046.435 3617.315 1047.435 ;
    END
  END SET_VH[17]
  PIN SET_VH[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3757.035 1046.435 3757.315 1047.435 ;
    END
  END SET_VH[18]
  PIN SET_VH[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3897.035 1046.435 3897.315 1047.435 ;
    END
  END SET_VH[19]
  PIN SET_VH[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4037.035 1046.435 4037.315 1047.435 ;
    END
  END SET_VH[20]
  PIN SET_VH[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4177.035 1046.435 4177.315 1047.435 ;
    END
  END SET_VH[21]
  PIN SET_VH[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4317.035 1046.435 4317.315 1047.435 ;
    END
  END SET_VH[22]
  PIN SET_VH[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4457.035 1046.435 4457.315 1047.435 ;
    END
  END SET_VH[23]
  PIN SET_VH[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4597.035 1046.435 4597.315 1047.435 ;
    END
  END SET_VH[24]
  PIN SET_VH[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4737.035 1046.435 4737.315 1047.435 ;
    END
  END SET_VH[25]
  PIN SET_VH[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4877.035 1046.435 4877.315 1047.435 ;
    END
  END SET_VH[26]
  PIN SET_VH[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5017.035 1046.435 5017.315 1047.435 ;
    END
  END SET_VH[27]
  PIN SET_VH[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5157.035 1046.435 5157.315 1047.435 ;
    END
  END SET_VH[28]
  PIN SET_VH[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5297.035 1046.435 5297.315 1047.435 ;
    END
  END SET_VH[29]
  PIN SET_VH[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5437.035 1046.435 5437.315 1047.435 ;
    END
  END SET_VH[30]
  PIN SET_VH[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5577.035 1046.435 5577.315 1047.435 ;
    END
  END SET_VH[31]
  PIN SET_VH[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5717.035 1046.435 5717.315 1047.435 ;
    END
  END SET_VH[32]
  PIN SET_VH[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5857.035 1046.435 5857.315 1047.435 ;
    END
  END SET_VH[33]
  PIN SET_VH[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5997.035 1046.435 5997.315 1047.435 ;
    END
  END SET_VH[34]
  PIN SET_VH[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6137.035 1046.435 6137.315 1047.435 ;
    END
  END SET_VH[35]
  PIN SET_VH[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6277.035 1046.435 6277.315 1047.435 ;
    END
  END SET_VH[36]
  PIN SET_VH[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6417.035 1046.435 6417.315 1047.435 ;
    END
  END SET_VH[37]
  PIN SET_VH[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6557.035 1046.435 6557.315 1047.435 ;
    END
  END SET_VH[38]
  PIN SET_VH[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6697.035 1046.435 6697.315 1047.435 ;
    END
  END SET_VH[39]
  PIN SET_VH[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6837.035 1046.435 6837.315 1047.435 ;
    END
  END SET_VH[40]
  PIN SET_VH[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6977.035 1046.435 6977.315 1047.435 ;
    END
  END SET_VH[41]
  PIN SET_VH[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7117.035 1046.435 7117.315 1047.435 ;
    END
  END SET_VH[42]
  PIN SET_VH[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7257.035 1046.435 7257.315 1047.435 ;
    END
  END SET_VH[43]
  PIN SET_VH[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7397.035 1046.435 7397.315 1047.435 ;
    END
  END SET_VH[44]
  PIN SET_VH[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7537.035 1046.435 7537.315 1047.435 ;
    END
  END SET_VH[45]
  PIN SET_VH[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7677.035 1046.435 7677.315 1047.435 ;
    END
  END SET_VH[46]
  PIN SET_VH[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7817.035 1046.435 7817.315 1047.435 ;
    END
  END SET_VH[47]
  PIN SET_VH[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7957.035 1046.435 7957.315 1047.435 ;
    END
  END SET_VH[48]
  PIN SET_VRESET_D[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15369.755 1046.435 15370.035 1047.435 ;
    END
  END SET_VRESET_D[101]
  PIN SET_VRESET_D[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15509.755 1046.435 15510.035 1047.435 ;
    END
  END SET_VRESET_D[102]
  PIN SET_VRESET_D[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15649.755 1046.435 15650.035 1047.435 ;
    END
  END SET_VRESET_D[103]
  PIN SET_VRESET_D[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15789.755 1046.435 15790.035 1047.435 ;
    END
  END SET_VRESET_D[104]
  PIN SET_VRESET_D[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15929.755 1046.435 15930.035 1047.435 ;
    END
  END SET_VRESET_D[105]
  PIN SET_VRESET_D[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16069.755 1046.435 16070.035 1047.435 ;
    END
  END SET_VRESET_D[106]
  PIN SET_VRESET_D[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16209.755 1046.435 16210.035 1047.435 ;
    END
  END SET_VRESET_D[107]
  PIN SET_VRESET_D[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16349.755 1046.435 16350.035 1047.435 ;
    END
  END SET_VRESET_D[108]
  PIN SET_VRESET_D[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16489.755 1046.435 16490.035 1047.435 ;
    END
  END SET_VRESET_D[109]
  PIN SET_VRESET_D[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16629.755 1046.435 16630.035 1047.435 ;
    END
  END SET_VRESET_D[110]
  PIN SET_VRESET_D[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16769.755 1046.435 16770.035 1047.435 ;
    END
  END SET_VRESET_D[111]
  PIN SET_VRESET_D[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16909.755 1046.435 16910.035 1047.435 ;
    END
  END SET_VRESET_D[112]
  PIN SET_VRESET_D[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17049.755 1046.435 17050.035 1047.435 ;
    END
  END SET_VRESET_D[113]
  PIN SET_VRESET_D[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17189.755 1046.435 17190.035 1047.435 ;
    END
  END SET_VRESET_D[114]
  PIN SET_VRESET_D[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17329.755 1046.435 17330.035 1047.435 ;
    END
  END SET_VRESET_D[115]
  PIN SET_VRESET_D[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17469.755 1046.435 17470.035 1047.435 ;
    END
  END SET_VRESET_D[116]
  PIN SET_VRESET_D[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17609.755 1046.435 17610.035 1047.435 ;
    END
  END SET_VRESET_D[117]
  PIN SET_VRESET_D[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17749.755 1046.435 17750.035 1047.435 ;
    END
  END SET_VRESET_D[118]
  PIN SET_VRESET_D[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17889.755 1046.435 17890.035 1047.435 ;
    END
  END SET_VRESET_D[119]
  PIN SET_VRESET_D[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18029.755 1046.435 18030.035 1047.435 ;
    END
  END SET_VRESET_D[120]
  PIN SET_VRESET_D[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18169.755 1046.435 18170.035 1047.435 ;
    END
  END SET_VRESET_D[121]
  PIN SET_VRESET_D[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18309.755 1046.435 18310.035 1047.435 ;
    END
  END SET_VRESET_D[122]
  PIN SET_VRESET_D[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18449.755 1046.435 18450.035 1047.435 ;
    END
  END SET_VRESET_D[123]
  PIN SET_VRESET_D[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18589.755 1046.435 18590.035 1047.435 ;
    END
  END SET_VRESET_D[124]
  PIN SET_VRESET_D[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18729.755 1046.435 18730.035 1047.435 ;
    END
  END SET_VRESET_D[125]
  PIN SET_VRESET_D[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18869.755 1046.435 18870.035 1047.435 ;
    END
  END SET_VRESET_D[126]
  PIN SET_VRESET_D[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19009.755 1046.435 19010.035 1047.435 ;
    END
  END SET_VRESET_D[127]
  PIN SET_VL[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1233.395 1046.435 1233.675 1047.435 ;
    END
  END SET_VL[0]
  PIN SET_VL[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1373.395 1046.435 1373.675 1047.435 ;
    END
  END SET_VL[1]
  PIN SET_VL[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1513.395 1046.435 1513.675 1047.435 ;
    END
  END SET_VL[2]
  PIN SET_VL[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1653.395 1046.435 1653.675 1047.435 ;
    END
  END SET_VL[3]
  PIN SET_VL[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1793.395 1046.435 1793.675 1047.435 ;
    END
  END SET_VL[4]
  PIN SET_VL[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1933.395 1046.435 1933.675 1047.435 ;
    END
  END SET_VL[5]
  PIN SET_VL[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2073.395 1046.435 2073.675 1047.435 ;
    END
  END SET_VL[6]
  PIN SET_VL[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2213.395 1046.435 2213.675 1047.435 ;
    END
  END SET_VL[7]
  PIN SET_VL[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2353.395 1046.435 2353.675 1047.435 ;
    END
  END SET_VL[8]
  PIN SET_VL[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2493.395 1046.435 2493.675 1047.435 ;
    END
  END SET_VL[9]
  PIN SET_VL[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2633.395 1046.435 2633.675 1047.435 ;
    END
  END SET_VL[10]
  PIN SET_VL[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2773.395 1046.435 2773.675 1047.435 ;
    END
  END SET_VL[11]
  PIN SET_VL[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2913.395 1046.435 2913.675 1047.435 ;
    END
  END SET_VL[12]
  PIN SET_VL[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3053.395 1046.435 3053.675 1047.435 ;
    END
  END SET_VL[13]
  PIN SET_VL[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3193.395 1046.435 3193.675 1047.435 ;
    END
  END SET_VL[14]
  PIN SET_VL[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3333.395 1046.435 3333.675 1047.435 ;
    END
  END SET_VL[15]
  PIN SET_VL[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3473.395 1046.435 3473.675 1047.435 ;
    END
  END SET_VL[16]
  PIN SET_VL[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3613.395 1046.435 3613.675 1047.435 ;
    END
  END SET_VL[17]
  PIN SET_VL[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3753.395 1046.435 3753.675 1047.435 ;
    END
  END SET_VL[18]
  PIN SET_VL[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3893.395 1046.435 3893.675 1047.435 ;
    END
  END SET_VL[19]
  PIN SET_VL[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4033.395 1046.435 4033.675 1047.435 ;
    END
  END SET_VL[20]
  PIN SET_VL[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4173.395 1046.435 4173.675 1047.435 ;
    END
  END SET_VL[21]
  PIN SET_VL[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4313.395 1046.435 4313.675 1047.435 ;
    END
  END SET_VL[22]
  PIN SET_VL[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4453.395 1046.435 4453.675 1047.435 ;
    END
  END SET_VL[23]
  PIN SET_VL[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4593.395 1046.435 4593.675 1047.435 ;
    END
  END SET_VL[24]
  PIN SET_VL[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4733.395 1046.435 4733.675 1047.435 ;
    END
  END SET_VL[25]
  PIN SET_VL[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4873.395 1046.435 4873.675 1047.435 ;
    END
  END SET_VL[26]
  PIN SET_VL[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5013.395 1046.435 5013.675 1047.435 ;
    END
  END SET_VL[27]
  PIN SET_VL[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5153.395 1046.435 5153.675 1047.435 ;
    END
  END SET_VL[28]
  PIN SET_VL[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5293.395 1046.435 5293.675 1047.435 ;
    END
  END SET_VL[29]
  PIN SET_VL[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5433.395 1046.435 5433.675 1047.435 ;
    END
  END SET_VL[30]
  PIN SET_VL[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5573.395 1046.435 5573.675 1047.435 ;
    END
  END SET_VL[31]
  PIN SET_VL[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5713.395 1046.435 5713.675 1047.435 ;
    END
  END SET_VL[32]
  PIN SET_VL[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5853.395 1046.435 5853.675 1047.435 ;
    END
  END SET_VL[33]
  PIN SET_VL[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5993.395 1046.435 5993.675 1047.435 ;
    END
  END SET_VL[34]
  PIN SET_VL[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6133.395 1046.435 6133.675 1047.435 ;
    END
  END SET_VL[35]
  PIN SET_VL[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6273.395 1046.435 6273.675 1047.435 ;
    END
  END SET_VL[36]
  PIN SET_VL[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6413.395 1046.435 6413.675 1047.435 ;
    END
  END SET_VL[37]
  PIN SET_VL[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6553.395 1046.435 6553.675 1047.435 ;
    END
  END SET_VL[38]
  PIN SET_VL[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6693.395 1046.435 6693.675 1047.435 ;
    END
  END SET_VL[39]
  PIN SET_VL[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6833.395 1046.435 6833.675 1047.435 ;
    END
  END SET_VL[40]
  PIN SET_VL[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6973.395 1046.435 6973.675 1047.435 ;
    END
  END SET_VL[41]
  PIN SET_VL[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7113.395 1046.435 7113.675 1047.435 ;
    END
  END SET_VL[42]
  PIN SET_VL[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7253.395 1046.435 7253.675 1047.435 ;
    END
  END SET_VL[43]
  PIN SET_VL[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7393.395 1046.435 7393.675 1047.435 ;
    END
  END SET_VL[44]
  PIN SET_VL[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7533.395 1046.435 7533.675 1047.435 ;
    END
  END SET_VL[45]
  PIN SET_VL[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7673.395 1046.435 7673.675 1047.435 ;
    END
  END SET_VL[46]
  PIN SET_VL[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7813.395 1046.435 7813.675 1047.435 ;
    END
  END SET_VL[47]
  PIN SET_VL[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7953.395 1046.435 7953.675 1047.435 ;
    END
  END SET_VL[48]
  PIN SET_VL[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8093.395 1046.435 8093.675 1047.435 ;
    END
  END SET_VL[49]
  PIN SET_VL[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8233.395 1046.435 8233.675 1047.435 ;
    END
  END SET_VL[50]
  PIN SET_VL[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8373.395 1046.435 8373.675 1047.435 ;
    END
  END SET_VL[51]
  PIN SET_VL[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8513.395 1046.435 8513.675 1047.435 ;
    END
  END SET_VL[52]
  PIN SET_VL[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8653.395 1046.435 8653.675 1047.435 ;
    END
  END SET_VL[53]
  PIN SET_VL[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8793.395 1046.435 8793.675 1047.435 ;
    END
  END SET_VL[54]
  PIN SET_VL[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8933.395 1046.435 8933.675 1047.435 ;
    END
  END SET_VL[55]
  PIN SET_VL[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9073.395 1046.435 9073.675 1047.435 ;
    END
  END SET_VL[56]
  PIN SET_VL[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9213.395 1046.435 9213.675 1047.435 ;
    END
  END SET_VL[57]
  PIN SET_VL[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9353.395 1046.435 9353.675 1047.435 ;
    END
  END SET_VL[58]
  PIN SET_VL[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9493.395 1046.435 9493.675 1047.435 ;
    END
  END SET_VL[59]
  PIN SET_VL[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9633.395 1046.435 9633.675 1047.435 ;
    END
  END SET_VL[60]
  PIN SET_VL[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9773.395 1046.435 9773.675 1047.435 ;
    END
  END SET_VL[61]
  PIN SET_VL[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9913.395 1046.435 9913.675 1047.435 ;
    END
  END SET_VL[62]
  PIN SET_VL[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10053.395 1046.435 10053.675 1047.435 ;
    END
  END SET_VL[63]
  PIN SET_VL[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10193.395 1046.435 10193.675 1047.435 ;
    END
  END SET_VL[64]
  PIN SET_VL[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10333.395 1046.435 10333.675 1047.435 ;
    END
  END SET_VL[65]
  PIN SET_VL[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10473.395 1046.435 10473.675 1047.435 ;
    END
  END SET_VL[66]
  PIN SET_VL[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10613.395 1046.435 10613.675 1047.435 ;
    END
  END SET_VL[67]
  PIN SET_VL[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10753.395 1046.435 10753.675 1047.435 ;
    END
  END SET_VL[68]
  PIN SET_VL[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10893.395 1046.435 10893.675 1047.435 ;
    END
  END SET_VL[69]
  PIN SET_VL[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11033.395 1046.435 11033.675 1047.435 ;
    END
  END SET_VL[70]
  PIN SET_VL[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11173.395 1046.435 11173.675 1047.435 ;
    END
  END SET_VL[71]
  PIN SET_VL[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11313.395 1046.435 11313.675 1047.435 ;
    END
  END SET_VL[72]
  PIN SET_VL[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11453.395 1046.435 11453.675 1047.435 ;
    END
  END SET_VL[73]
  PIN SET_VL[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11593.395 1046.435 11593.675 1047.435 ;
    END
  END SET_VL[74]
  PIN SET_VCLIP[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11464.315 1046.435 11464.595 1047.435 ;
    END
  END SET_VCLIP[73]
  PIN SET_VCLIP[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11604.315 1046.435 11604.595 1047.435 ;
    END
  END SET_VCLIP[74]
  PIN SET_VCLIP[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11744.315 1046.435 11744.595 1047.435 ;
    END
  END SET_VCLIP[75]
  PIN SET_VCLIP[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11884.315 1046.435 11884.595 1047.435 ;
    END
  END SET_VCLIP[76]
  PIN SET_VCLIP[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12024.315 1046.435 12024.595 1047.435 ;
    END
  END SET_VCLIP[77]
  PIN SET_VCLIP[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12164.315 1046.435 12164.595 1047.435 ;
    END
  END SET_VCLIP[78]
  PIN SET_VCLIP[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12304.315 1046.435 12304.595 1047.435 ;
    END
  END SET_VCLIP[79]
  PIN SET_VCLIP[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12444.315 1046.435 12444.595 1047.435 ;
    END
  END SET_VCLIP[80]
  PIN SET_VCLIP[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12584.315 1046.435 12584.595 1047.435 ;
    END
  END SET_VCLIP[81]
  PIN SET_VCLIP[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12724.315 1046.435 12724.595 1047.435 ;
    END
  END SET_VCLIP[82]
  PIN SET_VCLIP[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12864.315 1046.435 12864.595 1047.435 ;
    END
  END SET_VCLIP[83]
  PIN SET_VCLIP[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13004.315 1046.435 13004.595 1047.435 ;
    END
  END SET_VCLIP[84]
  PIN SET_VCLIP[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13144.315 1046.435 13144.595 1047.435 ;
    END
  END SET_VCLIP[85]
  PIN SET_VCLIP[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13284.315 1046.435 13284.595 1047.435 ;
    END
  END SET_VCLIP[86]
  PIN SET_VCLIP[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13424.315 1046.435 13424.595 1047.435 ;
    END
  END SET_VCLIP[87]
  PIN SET_VCLIP[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13564.315 1046.435 13564.595 1047.435 ;
    END
  END SET_VCLIP[88]
  PIN SET_VCLIP[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13704.315 1046.435 13704.595 1047.435 ;
    END
  END SET_VCLIP[89]
  PIN SET_VCLIP[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13844.315 1046.435 13844.595 1047.435 ;
    END
  END SET_VCLIP[90]
  PIN SET_VCLIP[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13984.315 1046.435 13984.595 1047.435 ;
    END
  END SET_VCLIP[91]
  PIN SET_VCLIP[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14124.315 1046.435 14124.595 1047.435 ;
    END
  END SET_VCLIP[92]
  PIN SET_VCLIP[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14264.315 1046.435 14264.595 1047.435 ;
    END
  END SET_VCLIP[93]
  PIN SET_VCLIP[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14404.315 1046.435 14404.595 1047.435 ;
    END
  END SET_VCLIP[94]
  PIN SET_VCLIP[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14544.315 1046.435 14544.595 1047.435 ;
    END
  END SET_VCLIP[95]
  PIN SET_VCLIP[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14684.315 1046.435 14684.595 1047.435 ;
    END
  END SET_VCLIP[96]
  PIN SET_VCLIP[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14824.315 1046.435 14824.595 1047.435 ;
    END
  END SET_VCLIP[97]
  PIN SET_VCLIP[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14964.315 1046.435 14964.595 1047.435 ;
    END
  END SET_VCLIP[98]
  PIN SET_VCLIP[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15104.315 1046.435 15104.595 1047.435 ;
    END
  END SET_VCLIP[99]
  PIN SET_VCLIP[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15244.315 1046.435 15244.595 1047.435 ;
    END
  END SET_VCLIP[100]
  PIN SET_VCLIP[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15384.315 1046.435 15384.595 1047.435 ;
    END
  END SET_VCLIP[101]
  PIN SET_VCLIP[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15524.315 1046.435 15524.595 1047.435 ;
    END
  END SET_VCLIP[102]
  PIN SET_VCLIP[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15664.315 1046.435 15664.595 1047.435 ;
    END
  END SET_VCLIP[103]
  PIN SET_VCLIP[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15804.315 1046.435 15804.595 1047.435 ;
    END
  END SET_VCLIP[104]
  PIN SET_VCLIP[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15944.315 1046.435 15944.595 1047.435 ;
    END
  END SET_VCLIP[105]
  PIN SET_VCLIP[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16084.315 1046.435 16084.595 1047.435 ;
    END
  END SET_VCLIP[106]
  PIN SET_VCLIP[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16224.315 1046.435 16224.595 1047.435 ;
    END
  END SET_VCLIP[107]
  PIN SET_VCLIP[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16364.315 1046.435 16364.595 1047.435 ;
    END
  END SET_VCLIP[108]
  PIN SET_VCLIP[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16504.315 1046.435 16504.595 1047.435 ;
    END
  END SET_VCLIP[109]
  PIN SET_VCLIP[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16644.315 1046.435 16644.595 1047.435 ;
    END
  END SET_VCLIP[110]
  PIN SET_VCLIP[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16784.315 1046.435 16784.595 1047.435 ;
    END
  END SET_VCLIP[111]
  PIN SET_VCLIP[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16924.315 1046.435 16924.595 1047.435 ;
    END
  END SET_VCLIP[112]
  PIN SET_VCLIP[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17064.315 1046.435 17064.595 1047.435 ;
    END
  END SET_VCLIP[113]
  PIN SET_VCLIP[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17204.315 1046.435 17204.595 1047.435 ;
    END
  END SET_VCLIP[114]
  PIN SET_VCLIP[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17344.315 1046.435 17344.595 1047.435 ;
    END
  END SET_VCLIP[115]
  PIN SET_VCLIP[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17484.315 1046.435 17484.595 1047.435 ;
    END
  END SET_VCLIP[116]
  PIN SET_VCLIP[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17624.315 1046.435 17624.595 1047.435 ;
    END
  END SET_VCLIP[117]
  PIN SET_VCLIP[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17764.315 1046.435 17764.595 1047.435 ;
    END
  END SET_VCLIP[118]
  PIN SET_VCLIP[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17904.315 1046.435 17904.595 1047.435 ;
    END
  END SET_VCLIP[119]
  PIN SET_VCLIP[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18044.315 1046.435 18044.595 1047.435 ;
    END
  END SET_VCLIP[120]
  PIN SET_VCLIP[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18184.315 1046.435 18184.595 1047.435 ;
    END
  END SET_VCLIP[121]
  PIN SET_VCLIP[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18324.315 1046.435 18324.595 1047.435 ;
    END
  END SET_VCLIP[122]
  PIN SET_VCLIP[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18464.315 1046.435 18464.595 1047.435 ;
    END
  END SET_VCLIP[123]
  PIN SET_VCLIP[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18604.315 1046.435 18604.595 1047.435 ;
    END
  END SET_VCLIP[124]
  PIN SET_VCLIP[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18744.315 1046.435 18744.595 1047.435 ;
    END
  END SET_VCLIP[125]
  PIN SET_VCLIP[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18884.315 1046.435 18884.595 1047.435 ;
    END
  END SET_VCLIP[126]
  PIN SWCNTL_IRESET
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10084.595 1046.435 10085.155 1047.435 ;
    END
  END SWCNTL_IRESET
  PIN SWCNTL_VRESET_D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10087.955 1046.435 10088.515 1047.435 ;
    END
  END SWCNTL_VRESET_D
  PIN SWCNTL_VCLIP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10094.675 1046.435 10095.235 1047.435 ;
    END
  END SWCNTL_VCLIP
  PIN SWCNTL_IREF
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10101.395 1046.435 10101.955 1047.435 ;
    END
  END SWCNTL_IREF
  PIN SWCNTL_DACMONV
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10099.715 1046.435 10100.275 1047.435 ;
    END
  END SWCNTL_DACMONV
  PIN SWCNTL_VRESET_P
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10092.995 1046.435 10093.555 1047.435 ;
    END
  END SWCNTL_VRESET_P
  PIN SWCNTL_IDB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10082.915 1046.435 10083.475 1047.435 ;
    END
  END SWCNTL_IDB
  PIN SET_IBUFP_R[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19151.955 1046.435 19152.235 1047.435 ;
    END
  END SET_IBUFP_R[0]
  PIN SET_IBUFP_R[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19152.515 1046.435 19152.795 1047.435 ;
    END
  END SET_IBUFP_R[1]
  PIN SET_IBUFP_R[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19153.075 1046.435 19153.355 1047.435 ;
    END
  END SET_IBUFP_R[2]
  PIN SET_IBUFP_R[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19153.635 1046.435 19153.915 1047.435 ;
    END
  END SET_IBUFP_R[3]
  PIN SET_IBUFN_R[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19154.195 1046.435 19154.475 1047.435 ;
    END
  END SET_IBUFN_R[0]
  PIN SET_IBUFN_R[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19154.755 1046.435 19155.035 1047.435 ;
    END
  END SET_IBUFN_R[1]
  PIN SET_IBUFN_R[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19155.315 1046.435 19155.595 1047.435 ;
    END
  END SET_IBUFN_R[2]
  PIN SET_IBUFN_R[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19155.875 1046.435 19156.155 1047.435 ;
    END
  END SET_IBUFN_R[3]
  PIN SWCNTL_ICASN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10086.275 1046.435 10086.835 1047.435 ;
    END
  END SWCNTL_ICASN
  PIN SWCNTL_VL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10089.635 1046.435 10090.195 1047.435 ;
    END
  END SWCNTL_VL
  PIN SWCNTL_DACMONI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10098.035 1046.435 10098.595 1047.435 ;
    END
  END SWCNTL_DACMONI
  PIN SWCNTL_IBIAS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10079.555 1046.435 10080.115 1047.435 ;
    END
  END SWCNTL_IBIAS
  PIN SET_IRESET_BIT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10103.075 1046.435 10103.635 1047.29 ;
    END
  END SET_IRESET_BIT
  PIN SWCNTL_VCASN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10096.355 1046.435 10096.915 1047.435 ;
    END
  END SWCNTL_VCASN
  PIN SWCNTL_VH
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10091.315 1046.435 10091.875 1047.435 ;
    END
  END SWCNTL_VH
  PIN SWCNTL_ITHR
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10081.235 1046.435 10081.795 1047.435 ;
    END
  END SWCNTL_ITHR
  PIN nRST[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8646.185 1046.435 8646.465 1047.435 ;
    END
  END nRST[94]
  PIN nRST[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8086.185 1046.435 8086.465 1047.435 ;
    END
  END nRST[87]
  PIN nRST[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7526.185 1046.435 7526.465 1047.435 ;
    END
  END nRST[80]
  PIN nRST[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6966.185 1046.435 6966.465 1047.435 ;
    END
  END nRST[73]
  PIN nRST[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9766.185 1046.435 9766.465 1047.435 ;
    END
  END nRST[108]
  PIN nRST[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9206.185 1046.435 9206.465 1047.435 ;
    END
  END nRST[101]
  PIN nRST[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6406.185 1046.435 6406.465 1047.435 ;
    END
  END nRST[66]
  PIN nRST[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5846.185 1046.435 5846.465 1047.435 ;
    END
  END nRST[59]
  PIN nRST[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5286.185 1046.435 5286.465 1047.435 ;
    END
  END nRST[52]
  PIN nRST[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15848.905 1046.435 15849.185 1047.435 ;
    END
  END nRST[184]
  PIN nRST[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14168.905 1046.435 14169.185 1047.435 ;
    END
  END nRST[163]
  PIN nRST[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1366.185 1046.435 1366.465 1047.435 ;
    END
  END nRST[3]
  PIN nRST[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18648.905 1046.435 18649.185 1047.435 ;
    END
  END nRST[219]
  PIN nRST[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18088.905 1046.435 18089.185 1047.435 ;
    END
  END nRST[212]
  PIN nRST[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17528.905 1046.435 17529.185 1047.435 ;
    END
  END nRST[205]
  PIN nRST[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16968.905 1046.435 16969.185 1047.435 ;
    END
  END nRST[198]
  PIN nRST[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16408.905 1046.435 16409.185 1047.435 ;
    END
  END nRST[191]
  PIN nRST[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4726.185 1046.435 4726.465 1047.435 ;
    END
  END nRST[45]
  PIN nRST[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3606.185 1046.435 3606.465 1047.435 ;
    END
  END nRST[31]
  PIN nRST[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3046.185 1046.435 3046.465 1047.435 ;
    END
  END nRST[24]
  PIN nRST[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2486.185 1046.435 2486.465 1047.435 ;
    END
  END nRST[17]
  PIN nRST[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1926.185 1046.435 1926.465 1047.435 ;
    END
  END nRST[10]
  PIN nRST[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4166.185 1046.435 4166.465 1047.435 ;
    END
  END nRST[38]
  PIN nRST[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15288.905 1046.435 15289.185 1047.435 ;
    END
  END nRST[177]
  PIN nRST[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14728.905 1046.435 14729.185 1047.435 ;
    END
  END nRST[170]
  PIN nRST[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13608.905 1046.435 13609.185 1047.435 ;
    END
  END nRST[156]
  PIN nRST[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13048.905 1046.435 13049.185 1047.435 ;
    END
  END nRST[149]
  PIN nRST[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12488.905 1046.435 12489.185 1047.435 ;
    END
  END nRST[142]
  PIN nRST[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11928.905 1046.435 11929.185 1047.435 ;
    END
  END nRST[135]
  PIN nRST[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11368.905 1046.435 11369.185 1047.435 ;
    END
  END nRST[128]
  PIN nRST[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7448.905 1046.435 7449.185 1047.435 ;
    END
  END nRST[79]
  PIN nRST[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6888.905 1046.435 6889.185 1047.435 ;
    END
  END nRST[72]
  PIN nRST[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6328.905 1046.435 6329.185 1047.435 ;
    END
  END nRST[65]
  PIN nRST[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9688.905 1046.435 9689.185 1047.435 ;
    END
  END nRST[107]
  PIN nRST[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9128.905 1046.435 9129.185 1047.435 ;
    END
  END nRST[100]
  PIN nRST[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8568.905 1046.435 8569.185 1047.435 ;
    END
  END nRST[93]
  PIN nRST[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8008.905 1046.435 8009.185 1047.435 ;
    END
  END nRST[86]
  PIN nRST[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14098.905 1046.435 14099.185 1047.435 ;
    END
  END nRST[162]
  PIN nRST[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13538.905 1046.435 13539.185 1047.435 ;
    END
  END nRST[155]
  PIN nRST[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12978.905 1046.435 12979.185 1047.435 ;
    END
  END nRST[148]
  PIN nRST[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16338.905 1046.435 16339.185 1047.435 ;
    END
  END nRST[190]
  PIN nRST[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15778.905 1046.435 15779.185 1047.435 ;
    END
  END nRST[183]
  PIN nRST[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15218.905 1046.435 15219.185 1047.435 ;
    END
  END nRST[176]
  PIN nRST[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14658.905 1046.435 14659.185 1047.435 ;
    END
  END nRST[169]
  PIN nRST[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18578.905 1046.435 18579.185 1047.435 ;
    END
  END nRST[218]
  PIN nRST[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18018.905 1046.435 18019.185 1047.435 ;
    END
  END nRST[211]
  PIN nRST[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5768.905 1046.435 5769.185 1047.435 ;
    END
  END nRST[58]
  PIN VDDP
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER TOP_M ;
        RECT 746.1 1358.18 748.1 1408.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 1358.18 19453.9 1408.18 ;
    END
    PORT
      LAYER M5 ;
        RECT 1130.48 1046.435 1143.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1176.52 1046.435 1189.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1193.5 1046.435 1206.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1210.48 1046.435 1223.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1256.52 1046.435 1269.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1273.5 1046.435 1286.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1290.48 1046.435 1303.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1336.52 1046.435 1349.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1353.5 1046.435 1366.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1370.48 1046.435 1383.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1416.52 1046.435 1429.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1433.5 1046.435 1446.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1450.48 1046.435 1463.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1496.52 1046.435 1509.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1513.5 1046.435 1526.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1530.48 1046.435 1543.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1576.52 1046.435 1589.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1593.5 1046.435 1606.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1610.48 1046.435 1623.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1656.52 1046.435 1669.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1673.5 1046.435 1686.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1690.48 1046.435 1703.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1736.52 1046.435 1749.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1753.5 1046.435 1766.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1770.48 1046.435 1783.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1816.52 1046.435 1829.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1833.5 1046.435 1846.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1850.48 1046.435 1863.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1896.52 1046.435 1909.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1913.5 1046.435 1926.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1930.48 1046.435 1943.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1976.52 1046.435 1989.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1993.5 1046.435 2006.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2010.48 1046.435 2023.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2056.52 1046.435 2069.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2073.5 1046.435 2086.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2090.48 1046.435 2103.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2136.52 1046.435 2149.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2153.5 1046.435 2166.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2170.48 1046.435 2183.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2216.52 1046.435 2229.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2233.5 1046.435 2246.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2250.48 1046.435 2263.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2296.52 1046.435 2309.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2313.5 1046.435 2326.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2330.48 1046.435 2343.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2376.52 1046.435 2389.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2393.5 1046.435 2406.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2410.48 1046.435 2423.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2456.52 1046.435 2469.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2473.5 1046.435 2486.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2490.48 1046.435 2503.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2536.52 1046.435 2549.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2553.5 1046.435 2566.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2570.48 1046.435 2583.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2616.52 1046.435 2629.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2633.5 1046.435 2646.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2650.48 1046.435 2663.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2696.52 1046.435 2709.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2713.5 1046.435 2726.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2730.48 1046.435 2743.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2776.52 1046.435 2789.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2793.5 1046.435 2806.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2810.48 1046.435 2823.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2856.52 1046.435 2869.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2873.5 1046.435 2886.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2890.48 1046.435 2903.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2936.52 1046.435 2949.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2953.5 1046.435 2966.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2970.48 1046.435 2983.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3016.52 1046.435 3029.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3033.5 1046.435 3046.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3050.48 1046.435 3063.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3096.52 1046.435 3109.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3113.5 1046.435 3126.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3130.48 1046.435 3143.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3176.52 1046.435 3189.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3193.5 1046.435 3206.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3210.48 1046.435 3223.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3256.52 1046.435 3269.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3273.5 1046.435 3286.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3290.48 1046.435 3303.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3336.52 1046.435 3349.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3353.5 1046.435 3366.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3370.48 1046.435 3383.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3416.52 1046.435 3429.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3433.5 1046.435 3446.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3450.48 1046.435 3463.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3496.52 1046.435 3509.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3513.5 1046.435 3526.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3530.48 1046.435 3543.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3576.52 1046.435 3589.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3593.5 1046.435 3606.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3610.48 1046.435 3623.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3656.52 1046.435 3669.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3673.5 1046.435 3686.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3690.48 1046.435 3703.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3736.52 1046.435 3749.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3753.5 1046.435 3766.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3770.48 1046.435 3783.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3816.52 1046.435 3829.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3833.5 1046.435 3846.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3850.48 1046.435 3863.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3896.52 1046.435 3909.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3913.5 1046.435 3926.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3930.48 1046.435 3943.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3976.52 1046.435 3989.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3993.5 1046.435 4006.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4010.48 1046.435 4023.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4056.52 1046.435 4069.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4073.5 1046.435 4086.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4090.48 1046.435 4103.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4136.52 1046.435 4149.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4153.5 1046.435 4166.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4170.48 1046.435 4183.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4216.52 1046.435 4229.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4233.5 1046.435 4246.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4250.48 1046.435 4263.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4296.52 1046.435 4309.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4313.5 1046.435 4326.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4330.48 1046.435 4343.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4376.52 1046.435 4389.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4393.5 1046.435 4406.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4410.48 1046.435 4423.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4456.52 1046.435 4469.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4473.5 1046.435 4486.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4490.48 1046.435 4503.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4536.52 1046.435 4549.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4553.5 1046.435 4566.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4570.48 1046.435 4583.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4616.52 1046.435 4629.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4633.5 1046.435 4646.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4650.48 1046.435 4663.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4696.52 1046.435 4709.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4713.5 1046.435 4726.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4730.48 1046.435 4743.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4776.52 1046.435 4789.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4793.5 1046.435 4806.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4810.48 1046.435 4823.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4856.52 1046.435 4869.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4873.5 1046.435 4886.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4890.48 1046.435 4903.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4936.52 1046.435 4949.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4953.5 1046.435 4966.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4970.48 1046.435 4983.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5016.52 1046.435 5029.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5033.5 1046.435 5046.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5050.48 1046.435 5063.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5096.52 1046.435 5109.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5113.5 1046.435 5126.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5130.48 1046.435 5143.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5176.52 1046.435 5189.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5193.5 1046.435 5206.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5210.48 1046.435 5223.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5256.52 1046.435 5269.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5273.5 1046.435 5286.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5290.48 1046.435 5303.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5336.52 1046.435 5349.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5353.5 1046.435 5366.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5370.48 1046.435 5383.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5416.52 1046.435 5429.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5433.5 1046.435 5446.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5450.48 1046.435 5463.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5496.52 1046.435 5509.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5513.5 1046.435 5526.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5530.48 1046.435 5543.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5576.52 1046.435 5589.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5593.5 1046.435 5606.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5610.48 1046.435 5623.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5656.52 1046.435 5669.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5673.5 1046.435 5686.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5690.48 1046.435 5703.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5736.52 1046.435 5749.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5753.5 1046.435 5766.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5770.48 1046.435 5783.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5816.52 1046.435 5829.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5833.5 1046.435 5846.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5850.48 1046.435 5863.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5896.52 1046.435 5909.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5913.5 1046.435 5926.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5930.48 1046.435 5943.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5976.52 1046.435 5989.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5993.5 1046.435 6006.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6010.48 1046.435 6023.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6056.52 1046.435 6069.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6073.5 1046.435 6086.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6090.48 1046.435 6103.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6136.52 1046.435 6149.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6153.5 1046.435 6166.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6170.48 1046.435 6183.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6216.52 1046.435 6229.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6233.5 1046.435 6246.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6250.48 1046.435 6263.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6296.52 1046.435 6309.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6313.5 1046.435 6326.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6330.48 1046.435 6343.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6376.52 1046.435 6389.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6393.5 1046.435 6406.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6410.48 1046.435 6423.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6456.52 1046.435 6469.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6473.5 1046.435 6486.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6490.48 1046.435 6503.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6536.52 1046.435 6549.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6553.5 1046.435 6566.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6570.48 1046.435 6583.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6616.52 1046.435 6629.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6633.5 1046.435 6646.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6650.48 1046.435 6663.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6696.52 1046.435 6709.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6713.5 1046.435 6726.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6730.48 1046.435 6743.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6776.52 1046.435 6789.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6793.5 1046.435 6806.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6810.48 1046.435 6823.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6856.52 1046.435 6869.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6873.5 1046.435 6886.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6890.48 1046.435 6903.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6936.52 1046.435 6949.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6953.5 1046.435 6966.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6970.48 1046.435 6983.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7016.52 1046.435 7029.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7033.5 1046.435 7046.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7050.48 1046.435 7063.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7096.52 1046.435 7109.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7113.5 1046.435 7126.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7130.48 1046.435 7143.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7176.52 1046.435 7189.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7193.5 1046.435 7206.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7210.48 1046.435 7223.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7256.52 1046.435 7269.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7273.5 1046.435 7286.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7290.48 1046.435 7303.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7336.52 1046.435 7349.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7353.5 1046.435 7366.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7370.48 1046.435 7383.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7416.52 1046.435 7429.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7433.5 1046.435 7446.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7450.48 1046.435 7463.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7496.52 1046.435 7509.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7513.5 1046.435 7526.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7530.48 1046.435 7543.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7576.52 1046.435 7589.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7593.5 1046.435 7606.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7610.48 1046.435 7623.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7656.52 1046.435 7669.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7673.5 1046.435 7686.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7690.48 1046.435 7703.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7736.52 1046.435 7749.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7753.5 1046.435 7766.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7770.48 1046.435 7783.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7816.52 1046.435 7829.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7833.5 1046.435 7846.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7850.48 1046.435 7863.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7896.52 1046.435 7909.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7913.5 1046.435 7926.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7930.48 1046.435 7943.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7976.52 1046.435 7989.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7993.5 1046.435 8006.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8010.48 1046.435 8023.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8056.52 1046.435 8069.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8073.5 1046.435 8086.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8090.48 1046.435 8103.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8136.52 1046.435 8149.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8153.5 1046.435 8166.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8170.48 1046.435 8183.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8216.52 1046.435 8229.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8233.5 1046.435 8246.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8250.48 1046.435 8263.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8296.52 1046.435 8309.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8313.5 1046.435 8326.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8330.48 1046.435 8343.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8376.52 1046.435 8389.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8393.5 1046.435 8406.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8410.48 1046.435 8423.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8456.52 1046.435 8469.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8473.5 1046.435 8486.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8490.48 1046.435 8503.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8536.52 1046.435 8549.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8553.5 1046.435 8566.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8570.48 1046.435 8583.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8616.52 1046.435 8629.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8633.5 1046.435 8646.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8650.48 1046.435 8663.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8696.52 1046.435 8709.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8713.5 1046.435 8726.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8730.48 1046.435 8743.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8776.52 1046.435 8789.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8793.5 1046.435 8806.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8810.48 1046.435 8823.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8856.52 1046.435 8869.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8873.5 1046.435 8886.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8890.48 1046.435 8903.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8936.52 1046.435 8949.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8953.5 1046.435 8966.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8970.48 1046.435 8983.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9016.52 1046.435 9029.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9033.5 1046.435 9046.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9050.48 1046.435 9063.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9096.52 1046.435 9109.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9113.5 1046.435 9126.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9130.48 1046.435 9143.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9176.52 1046.435 9189.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9193.5 1046.435 9206.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9210.48 1046.435 9223.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9256.52 1046.435 9269.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9273.5 1046.435 9286.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9290.48 1046.435 9303.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9336.52 1046.435 9349.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9353.5 1046.435 9366.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9370.48 1046.435 9383.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9416.52 1046.435 9429.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9433.5 1046.435 9446.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9450.48 1046.435 9463.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9496.52 1046.435 9509.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9513.5 1046.435 9526.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9530.48 1046.435 9543.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9576.52 1046.435 9589.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9593.5 1046.435 9606.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9610.48 1046.435 9623.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9656.52 1046.435 9669.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9673.5 1046.435 9686.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9690.48 1046.435 9703.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9736.52 1046.435 9749.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9753.5 1046.435 9766.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9770.48 1046.435 9783.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9816.52 1046.435 9829.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9833.5 1046.435 9846.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9850.48 1046.435 9863.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9896.52 1046.435 9909.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9913.5 1046.435 9926.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9930.48 1046.435 9943.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9976.52 1046.435 9989.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9993.5 1046.435 10006.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10010.48 1046.435 10023.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10056.52 1046.435 10069.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10073.5 1046.435 10086.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10090.48 1046.435 10103.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10136.52 1046.435 10149.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10153.5 1046.435 10166.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10170.48 1046.435 10183.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10216.52 1046.435 10229.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10233.5 1046.435 10246.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10250.48 1046.435 10263.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10296.52 1046.435 10309.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10313.5 1046.435 10326.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10330.48 1046.435 10343.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10376.52 1046.435 10389.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10393.5 1046.435 10406.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10410.48 1046.435 10423.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10456.52 1046.435 10469.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10473.5 1046.435 10486.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10490.48 1046.435 10503.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10536.52 1046.435 10549.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10553.5 1046.435 10566.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10570.48 1046.435 10583.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10616.52 1046.435 10629.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10633.5 1046.435 10646.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10650.48 1046.435 10663.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10696.52 1046.435 10709.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10713.5 1046.435 10726.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10730.48 1046.435 10743.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10776.52 1046.435 10789.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10793.5 1046.435 10806.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10810.48 1046.435 10823.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10856.52 1046.435 10869.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10873.5 1046.435 10886.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10890.48 1046.435 10903.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10936.52 1046.435 10949.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10953.5 1046.435 10966.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10970.48 1046.435 10983.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11016.52 1046.435 11029.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11033.5 1046.435 11046.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11050.48 1046.435 11063.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11096.52 1046.435 11109.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11113.5 1046.435 11126.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11130.48 1046.435 11143.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11176.52 1046.435 11189.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11193.5 1046.435 11206.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11210.48 1046.435 11223.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11256.52 1046.435 11269.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11273.5 1046.435 11286.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11290.48 1046.435 11303.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11336.52 1046.435 11349.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11353.5 1046.435 11366.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11370.48 1046.435 11383.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11416.52 1046.435 11429.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11433.5 1046.435 11446.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11450.48 1046.435 11463.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11496.52 1046.435 11509.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11513.5 1046.435 11526.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11530.48 1046.435 11543.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11576.52 1046.435 11589.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11593.5 1046.435 11606.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11610.48 1046.435 11623.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11656.52 1046.435 11669.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11673.5 1046.435 11686.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11690.48 1046.435 11703.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11736.52 1046.435 11749.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11753.5 1046.435 11766.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11770.48 1046.435 11783.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11816.52 1046.435 11829.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11833.5 1046.435 11846.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11850.48 1046.435 11863.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11896.52 1046.435 11909.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11913.5 1046.435 11926.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11930.48 1046.435 11943.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11976.52 1046.435 11989.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11993.5 1046.435 12006.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12010.48 1046.435 12023.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12056.52 1046.435 12069.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12073.5 1046.435 12086.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12090.48 1046.435 12103.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12136.52 1046.435 12149.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12153.5 1046.435 12166.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12170.48 1046.435 12183.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12216.52 1046.435 12229.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12233.5 1046.435 12246.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12250.48 1046.435 12263.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12296.52 1046.435 12309.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12313.5 1046.435 12326.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12330.48 1046.435 12343.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12376.52 1046.435 12389.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12393.5 1046.435 12406.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12410.48 1046.435 12423.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12456.52 1046.435 12469.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12473.5 1046.435 12486.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12490.48 1046.435 12503.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12536.52 1046.435 12549.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12553.5 1046.435 12566.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12570.48 1046.435 12583.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12616.52 1046.435 12629.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12633.5 1046.435 12646.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12650.48 1046.435 12663.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12696.52 1046.435 12709.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12713.5 1046.435 12726.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12730.48 1046.435 12743.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12776.52 1046.435 12789.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12793.5 1046.435 12806.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12810.48 1046.435 12823.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12856.52 1046.435 12869.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12873.5 1046.435 12886.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12890.48 1046.435 12903.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12936.52 1046.435 12949.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12953.5 1046.435 12966.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12970.48 1046.435 12983.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13016.52 1046.435 13029.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13033.5 1046.435 13046.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13050.48 1046.435 13063.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13096.52 1046.435 13109.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13113.5 1046.435 13126.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13130.48 1046.435 13143.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13176.52 1046.435 13189.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13193.5 1046.435 13206.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13210.48 1046.435 13223.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13256.52 1046.435 13269.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13273.5 1046.435 13286.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13290.48 1046.435 13303.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13336.52 1046.435 13349.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13353.5 1046.435 13366.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13370.48 1046.435 13383.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13416.52 1046.435 13429.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13433.5 1046.435 13446.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13450.48 1046.435 13463.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13496.52 1046.435 13509.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13513.5 1046.435 13526.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13530.48 1046.435 13543.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13576.52 1046.435 13589.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13593.5 1046.435 13606.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13610.48 1046.435 13623.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13656.52 1046.435 13669.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13673.5 1046.435 13686.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13690.48 1046.435 13703.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13736.52 1046.435 13749.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13753.5 1046.435 13766.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13770.48 1046.435 13783.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13816.52 1046.435 13829.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13833.5 1046.435 13846.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13850.48 1046.435 13863.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13896.52 1046.435 13909.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13913.5 1046.435 13926.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13930.48 1046.435 13943.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13976.52 1046.435 13989.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13993.5 1046.435 14006.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14010.48 1046.435 14023.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14056.52 1046.435 14069.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14073.5 1046.435 14086.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14090.48 1046.435 14103.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14136.52 1046.435 14149.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14153.5 1046.435 14166.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14170.48 1046.435 14183.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14216.52 1046.435 14229.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14233.5 1046.435 14246.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14250.48 1046.435 14263.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14296.52 1046.435 14309.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14313.5 1046.435 14326.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14330.48 1046.435 14343.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14376.52 1046.435 14389.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14393.5 1046.435 14406.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14410.48 1046.435 14423.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14456.52 1046.435 14469.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14473.5 1046.435 14486.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14490.48 1046.435 14503.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14536.52 1046.435 14549.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14553.5 1046.435 14566.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14570.48 1046.435 14583.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14616.52 1046.435 14629.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14633.5 1046.435 14646.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14650.48 1046.435 14663.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14696.52 1046.435 14709.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14713.5 1046.435 14726.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14730.48 1046.435 14743.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14776.52 1046.435 14789.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14793.5 1046.435 14806.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14810.48 1046.435 14823.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14856.52 1046.435 14869.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14873.5 1046.435 14886.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14890.48 1046.435 14903.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14936.52 1046.435 14949.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14953.5 1046.435 14966.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14970.48 1046.435 14983.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15016.52 1046.435 15029.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15033.5 1046.435 15046.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15050.48 1046.435 15063.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15096.52 1046.435 15109.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15113.5 1046.435 15126.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15130.48 1046.435 15143.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15176.52 1046.435 15189.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15193.5 1046.435 15206.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15210.48 1046.435 15223.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15256.52 1046.435 15269.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15273.5 1046.435 15286.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15290.48 1046.435 15303.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15336.52 1046.435 15349.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15353.5 1046.435 15366.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15370.48 1046.435 15383.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15416.52 1046.435 15429.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15433.5 1046.435 15446.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15450.48 1046.435 15463.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15496.52 1046.435 15509.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15513.5 1046.435 15526.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15530.48 1046.435 15543.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15576.52 1046.435 15589.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15593.5 1046.435 15606.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15610.48 1046.435 15623.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15656.52 1046.435 15669.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15673.5 1046.435 15686.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15690.48 1046.435 15703.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15736.52 1046.435 15749.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15753.5 1046.435 15766.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15770.48 1046.435 15783.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15816.52 1046.435 15829.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15833.5 1046.435 15846.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15850.48 1046.435 15863.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15896.52 1046.435 15909.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15913.5 1046.435 15926.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15930.48 1046.435 15943.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15976.52 1046.435 15989.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15993.5 1046.435 16006.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16010.48 1046.435 16023.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16056.52 1046.435 16069.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16073.5 1046.435 16086.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16090.48 1046.435 16103.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16136.52 1046.435 16149.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16153.5 1046.435 16166.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16170.48 1046.435 16183.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16216.52 1046.435 16229.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16233.5 1046.435 16246.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16250.48 1046.435 16263.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16296.52 1046.435 16309.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16313.5 1046.435 16326.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16330.48 1046.435 16343.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16376.52 1046.435 16389.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16393.5 1046.435 16406.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16410.48 1046.435 16423.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16456.52 1046.435 16469.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16473.5 1046.435 16486.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16490.48 1046.435 16503.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16536.52 1046.435 16549.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16553.5 1046.435 16566.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16570.48 1046.435 16583.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16616.52 1046.435 16629.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16633.5 1046.435 16646.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16650.48 1046.435 16663.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16696.52 1046.435 16709.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16713.5 1046.435 16726.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16730.48 1046.435 16743.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16776.52 1046.435 16789.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16793.5 1046.435 16806.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16810.48 1046.435 16823.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16856.52 1046.435 16869.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16873.5 1046.435 16886.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16890.48 1046.435 16903.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16936.52 1046.435 16949.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16953.5 1046.435 16966.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16970.48 1046.435 16983.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17016.52 1046.435 17029.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17033.5 1046.435 17046.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17050.48 1046.435 17063.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17096.52 1046.435 17109.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17113.5 1046.435 17126.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17130.48 1046.435 17143.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17176.52 1046.435 17189.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17193.5 1046.435 17206.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17210.48 1046.435 17223.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17256.52 1046.435 17269.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17273.5 1046.435 17286.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17290.48 1046.435 17303.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17336.52 1046.435 17349.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17353.5 1046.435 17366.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17370.48 1046.435 17383.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17416.52 1046.435 17429.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17433.5 1046.435 17446.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17450.48 1046.435 17463.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17496.52 1046.435 17509.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17513.5 1046.435 17526.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17530.48 1046.435 17543.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17576.52 1046.435 17589.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17593.5 1046.435 17606.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17610.48 1046.435 17623.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17656.52 1046.435 17669.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17673.5 1046.435 17686.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17690.48 1046.435 17703.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17736.52 1046.435 17749.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17753.5 1046.435 17766.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17770.48 1046.435 17783.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17816.52 1046.435 17829.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17833.5 1046.435 17846.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17850.48 1046.435 17863.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17896.52 1046.435 17909.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17913.5 1046.435 17926.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17930.48 1046.435 17943.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17976.52 1046.435 17989.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17993.5 1046.435 18006.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18010.48 1046.435 18023.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18056.52 1046.435 18069.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18073.5 1046.435 18086.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18090.48 1046.435 18103.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18136.52 1046.435 18149.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18153.5 1046.435 18166.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18170.48 1046.435 18183.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18216.52 1046.435 18229.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18233.5 1046.435 18246.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18250.48 1046.435 18263.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18296.52 1046.435 18309.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18313.5 1046.435 18326.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18330.48 1046.435 18343.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18376.52 1046.435 18389.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18393.5 1046.435 18406.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18410.48 1046.435 18423.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18456.52 1046.435 18469.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18473.5 1046.435 18486.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18490.48 1046.435 18503.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18536.52 1046.435 18549.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18553.5 1046.435 18566.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18570.48 1046.435 18583.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18616.52 1046.435 18629.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18633.5 1046.435 18646.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18650.48 1046.435 18663.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18696.52 1046.435 18709.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18713.5 1046.435 18726.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18730.48 1046.435 18743.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18776.52 1046.435 18789.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18793.5 1046.435 18806.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18810.48 1046.435 18823.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18856.52 1046.435 18869.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18873.5 1046.435 18886.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18890.48 1046.435 18903.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18936.52 1046.435 18949.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18953.5 1046.435 18966.5 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18970.48 1046.435 18983.48 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 19016.52 1046.435 19029.52 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 19033.5 1046.435 19046.5 1047.435 ;
    END
  END VDDP
  PIN GNDP
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER TOP_M ;
        RECT 746.1 1238.18 748.1 1288.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 1238.18 19453.9 1288.18 ;
    END
    PORT
      LAYER M5 ;
        RECT 1146 1046.435 1174 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1226 1046.435 1254 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1306 1046.435 1334 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1386 1046.435 1414 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1466 1046.435 1494 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1546 1046.435 1574 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1626 1046.435 1654 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1706 1046.435 1734 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1786 1046.435 1814 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1866 1046.435 1894 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 1946 1046.435 1974 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2026 1046.435 2054 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2106 1046.435 2134 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2186 1046.435 2214 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2266 1046.435 2294 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2346 1046.435 2374 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2426 1046.435 2454 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2506 1046.435 2534 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2586 1046.435 2614 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2666 1046.435 2694 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2746 1046.435 2774 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2826 1046.435 2854 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2906 1046.435 2934 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 2986 1046.435 3014 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3066 1046.435 3094 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3146 1046.435 3174 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3226 1046.435 3254 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3306 1046.435 3334 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3386 1046.435 3414 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3466 1046.435 3494 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3546 1046.435 3574 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3626 1046.435 3654 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3706 1046.435 3734 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3786 1046.435 3814 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3866 1046.435 3894 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 3946 1046.435 3974 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4026 1046.435 4054 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4106 1046.435 4134 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4186 1046.435 4214 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4266 1046.435 4294 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4346 1046.435 4374 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4426 1046.435 4454 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4506 1046.435 4534 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4586 1046.435 4614 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4666 1046.435 4694 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4746 1046.435 4774 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4826 1046.435 4854 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4906 1046.435 4934 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 4986 1046.435 5014 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5066 1046.435 5094 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5146 1046.435 5174 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5226 1046.435 5254 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5306 1046.435 5334 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5386 1046.435 5414 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5466 1046.435 5494 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5546 1046.435 5574 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5626 1046.435 5654 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5706 1046.435 5734 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5786 1046.435 5814 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5866 1046.435 5894 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 5946 1046.435 5974 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6026 1046.435 6054 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6106 1046.435 6134 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6186 1046.435 6214 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6266 1046.435 6294 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6346 1046.435 6374 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6426 1046.435 6454 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6506 1046.435 6534 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6586 1046.435 6614 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6666 1046.435 6694 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6746 1046.435 6774 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6826 1046.435 6854 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6906 1046.435 6934 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 6986 1046.435 7014 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7066 1046.435 7094 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7146 1046.435 7174 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7226 1046.435 7254 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7306 1046.435 7334 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7386 1046.435 7414 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7466 1046.435 7494 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7546 1046.435 7574 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7626 1046.435 7654 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7706 1046.435 7734 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7786 1046.435 7814 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7866 1046.435 7894 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 7946 1046.435 7974 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8026 1046.435 8054 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8106 1046.435 8134 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8186 1046.435 8214 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8266 1046.435 8294 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8346 1046.435 8374 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8426 1046.435 8454 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8506 1046.435 8534 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8586 1046.435 8614 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8666 1046.435 8694 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8746 1046.435 8774 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8826 1046.435 8854 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8906 1046.435 8934 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 8986 1046.435 9014 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9066 1046.435 9094 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9146 1046.435 9174 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9226 1046.435 9254 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9306 1046.435 9334 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9386 1046.435 9414 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9466 1046.435 9494 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9546 1046.435 9574 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9626 1046.435 9654 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9706 1046.435 9734 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9786 1046.435 9814 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9866 1046.435 9894 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 9946 1046.435 9974 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10026 1046.435 10054 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10106 1046.435 10134 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10186 1046.435 10214 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10266 1046.435 10294 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10346 1046.435 10374 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10426 1046.435 10454 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10506 1046.435 10534 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10586 1046.435 10614 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10666 1046.435 10694 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10746 1046.435 10774 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10826 1046.435 10854 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10906 1046.435 10934 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 10986 1046.435 11014 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11066 1046.435 11094 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11146 1046.435 11174 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11226 1046.435 11254 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11306 1046.435 11334 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11386 1046.435 11414 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11466 1046.435 11494 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11546 1046.435 11574 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11626 1046.435 11654 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11706 1046.435 11734 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11786 1046.435 11814 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11866 1046.435 11894 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 11946 1046.435 11974 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12026 1046.435 12054 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12106 1046.435 12134 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12186 1046.435 12214 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12266 1046.435 12294 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12346 1046.435 12374 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12426 1046.435 12454 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12506 1046.435 12534 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12586 1046.435 12614 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12666 1046.435 12694 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12746 1046.435 12774 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12826 1046.435 12854 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12906 1046.435 12934 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 12986 1046.435 13014 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13066 1046.435 13094 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13146 1046.435 13174 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13226 1046.435 13254 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13306 1046.435 13334 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13386 1046.435 13414 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13466 1046.435 13494 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13546 1046.435 13574 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13626 1046.435 13654 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13706 1046.435 13734 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13786 1046.435 13814 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13866 1046.435 13894 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 13946 1046.435 13974 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14026 1046.435 14054 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14106 1046.435 14134 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14186 1046.435 14214 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14266 1046.435 14294 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14346 1046.435 14374 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14426 1046.435 14454 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14506 1046.435 14534 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14586 1046.435 14614 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14666 1046.435 14694 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14746 1046.435 14774 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14826 1046.435 14854 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14906 1046.435 14934 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 14986 1046.435 15014 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15066 1046.435 15094 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15146 1046.435 15174 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15226 1046.435 15254 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15306 1046.435 15334 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15386 1046.435 15414 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15466 1046.435 15494 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15546 1046.435 15574 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15626 1046.435 15654 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15706 1046.435 15734 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15786 1046.435 15814 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15866 1046.435 15894 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 15946 1046.435 15974 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16026 1046.435 16054 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16106 1046.435 16134 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16186 1046.435 16214 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16266 1046.435 16294 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16346 1046.435 16374 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16426 1046.435 16454 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16506 1046.435 16534 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16586 1046.435 16614 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16666 1046.435 16694 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16746 1046.435 16774 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16826 1046.435 16854 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16906 1046.435 16934 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 16986 1046.435 17014 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17066 1046.435 17094 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17146 1046.435 17174 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17226 1046.435 17254 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17306 1046.435 17334 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17386 1046.435 17414 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17466 1046.435 17494 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17546 1046.435 17574 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17626 1046.435 17654 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17706 1046.435 17734 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17786 1046.435 17814 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17866 1046.435 17894 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 17946 1046.435 17974 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18026 1046.435 18054 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18106 1046.435 18134 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18186 1046.435 18214 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18266 1046.435 18294 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18346 1046.435 18374 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18426 1046.435 18454 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18506 1046.435 18534 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18586 1046.435 18614 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18666 1046.435 18694 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18746 1046.435 18774 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18826 1046.435 18854 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18906 1046.435 18934 1047.435 ;
    END
    PORT
      LAYER M5 ;
        RECT 18986 1046.435 19014 1047.435 ;
    END
  END GNDP
  PIN SET_IBUFN_L[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1003.845 1046.435 1004.125 1047.435 ;
    END
  END SET_IBUFN_L[3]
  PIN SET_IBUFN_L[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1004.965 1046.435 1005.245 1047.435 ;
    END
  END SET_IBUFN_L[1]
  PIN SET_IBUFN_L[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1004.405 1046.435 1004.685 1047.435 ;
    END
  END SET_IBUFN_L[2]
  PIN SET_IBUFN_L[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1005.525 1046.435 1005.805 1047.435 ;
    END
  END SET_IBUFN_L[0]
  PIN SET_IBUFP_L[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1007.205 1046.435 1007.485 1047.435 ;
    END
  END SET_IBUFP_L[1]
  PIN SET_IBUFP_L[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1007.765 1046.435 1008.045 1047.435 ;
    END
  END SET_IBUFP_L[0]
  PIN SET_IBUFP_L[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1006.645 1046.435 1006.925 1047.435 ;
    END
  END SET_IBUFP_L[2]
  PIN SET_IBUFP_L[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1006.085 1046.435 1006.365 1047.435 ;
    END
  END SET_IBUFP_L[3]
  PIN SET_ITHR[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15578.915 1046.435 15579.195 1047.435 ;
    END
  END SET_ITHR[103]
  PIN SET_ITHR[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15718.915 1046.435 15719.195 1047.435 ;
    END
  END SET_ITHR[104]
  PIN SET_ITHR[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15858.915 1046.435 15859.195 1047.435 ;
    END
  END SET_ITHR[105]
  PIN SET_ITHR[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15998.915 1046.435 15999.195 1047.435 ;
    END
  END SET_ITHR[106]
  PIN SET_ITHR[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16138.915 1046.435 16139.195 1047.435 ;
    END
  END SET_ITHR[107]
  PIN SET_ITHR[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16278.915 1046.435 16279.195 1047.435 ;
    END
  END SET_ITHR[108]
  PIN SET_ITHR[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16418.915 1046.435 16419.195 1047.435 ;
    END
  END SET_ITHR[109]
  PIN SET_ITHR[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16558.915 1046.435 16559.195 1047.435 ;
    END
  END SET_ITHR[110]
  PIN SET_ITHR[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16698.915 1046.435 16699.195 1047.435 ;
    END
  END SET_ITHR[111]
  PIN SET_ITHR[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16838.915 1046.435 16839.195 1047.435 ;
    END
  END SET_ITHR[112]
  PIN SET_ITHR[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16978.915 1046.435 16979.195 1047.435 ;
    END
  END SET_ITHR[113]
  PIN SET_ITHR[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17118.915 1046.435 17119.195 1047.435 ;
    END
  END SET_ITHR[114]
  PIN SET_ITHR[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17258.915 1046.435 17259.195 1047.435 ;
    END
  END SET_ITHR[115]
  PIN SET_ITHR[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17398.915 1046.435 17399.195 1047.435 ;
    END
  END SET_ITHR[116]
  PIN SET_ITHR[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17538.915 1046.435 17539.195 1047.435 ;
    END
  END SET_ITHR[117]
  PIN SET_ITHR[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17678.915 1046.435 17679.195 1047.435 ;
    END
  END SET_ITHR[118]
  PIN SET_ITHR[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17818.915 1046.435 17819.195 1047.435 ;
    END
  END SET_ITHR[119]
  PIN SET_ITHR[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17958.915 1046.435 17959.195 1047.435 ;
    END
  END SET_ITHR[120]
  PIN SET_ITHR[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18098.915 1046.435 18099.195 1047.435 ;
    END
  END SET_ITHR[121]
  PIN SET_ITHR[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18238.915 1046.435 18239.195 1047.435 ;
    END
  END SET_ITHR[122]
  PIN SET_ITHR[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18378.915 1046.435 18379.195 1047.435 ;
    END
  END SET_ITHR[123]
  PIN SET_ITHR[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18518.915 1046.435 18519.195 1047.435 ;
    END
  END SET_ITHR[124]
  PIN SET_ITHR[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18658.915 1046.435 18659.195 1047.435 ;
    END
  END SET_ITHR[125]
  PIN SET_ITHR[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18798.915 1046.435 18799.195 1047.435 ;
    END
  END SET_ITHR[126]
  PIN SET_ITHR[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18938.915 1046.435 18939.195 1047.435 ;
    END
  END SET_ITHR[127]
  PIN SET_IDB[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1162.835 1046.435 1163.115 1047.435 ;
    END
  END SET_IDB[0]
  PIN SET_IDB[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1302.835 1046.435 1303.115 1047.435 ;
    END
  END SET_IDB[1]
  PIN SET_IDB[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1442.835 1046.435 1443.115 1047.435 ;
    END
  END SET_IDB[2]
  PIN SET_IDB[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1582.835 1046.435 1583.115 1047.435 ;
    END
  END SET_IDB[3]
  PIN SET_IDB[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1722.835 1046.435 1723.115 1047.435 ;
    END
  END SET_IDB[4]
  PIN SET_IDB[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1862.835 1046.435 1863.115 1047.435 ;
    END
  END SET_IDB[5]
  PIN SET_IDB[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2002.835 1046.435 2003.115 1047.435 ;
    END
  END SET_IDB[6]
  PIN SET_IDB[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2142.835 1046.435 2143.115 1047.435 ;
    END
  END SET_IDB[7]
  PIN SET_IDB[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2282.835 1046.435 2283.115 1047.435 ;
    END
  END SET_IDB[8]
  PIN SET_IDB[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2422.835 1046.435 2423.115 1047.435 ;
    END
  END SET_IDB[9]
  PIN SET_IDB[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2562.835 1046.435 2563.115 1047.435 ;
    END
  END SET_IDB[10]
  PIN SET_IDB[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2702.835 1046.435 2703.115 1047.435 ;
    END
  END SET_IDB[11]
  PIN SET_IDB[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2842.835 1046.435 2843.115 1047.435 ;
    END
  END SET_IDB[12]
  PIN SET_IDB[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2982.835 1046.435 2983.115 1047.435 ;
    END
  END SET_IDB[13]
  PIN SET_IDB[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3122.835 1046.435 3123.115 1047.435 ;
    END
  END SET_IDB[14]
  PIN SET_IDB[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3262.835 1046.435 3263.115 1047.435 ;
    END
  END SET_IDB[15]
  PIN SET_IDB[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3402.835 1046.435 3403.115 1047.435 ;
    END
  END SET_IDB[16]
  PIN SET_IDB[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3542.835 1046.435 3543.115 1047.435 ;
    END
  END SET_IDB[17]
  PIN SET_IDB[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3682.835 1046.435 3683.115 1047.435 ;
    END
  END SET_IDB[18]
  PIN SET_IDB[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3822.835 1046.435 3823.115 1047.435 ;
    END
  END SET_IDB[19]
  PIN SET_IDB[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3962.835 1046.435 3963.115 1047.435 ;
    END
  END SET_IDB[20]
  PIN SET_IDB[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4102.835 1046.435 4103.115 1047.435 ;
    END
  END SET_IDB[21]
  PIN SET_IDB[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4242.835 1046.435 4243.115 1047.435 ;
    END
  END SET_IDB[22]
  PIN SET_IDB[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4382.835 1046.435 4383.115 1047.435 ;
    END
  END SET_IDB[23]
  PIN SET_IDB[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4522.835 1046.435 4523.115 1047.435 ;
    END
  END SET_IDB[24]
  PIN SET_IDB[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4662.835 1046.435 4663.115 1047.435 ;
    END
  END SET_IDB[25]
  PIN SET_IDB[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4802.835 1046.435 4803.115 1047.435 ;
    END
  END SET_IDB[26]
  PIN SET_IDB[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4942.835 1046.435 4943.115 1047.435 ;
    END
  END SET_IDB[27]
  PIN SET_IDB[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5082.835 1046.435 5083.115 1047.435 ;
    END
  END SET_IDB[28]
  PIN SET_IDB[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5222.835 1046.435 5223.115 1047.435 ;
    END
  END SET_IDB[29]
  PIN SET_IDB[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5362.835 1046.435 5363.115 1047.435 ;
    END
  END SET_IDB[30]
  PIN SET_IDB[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5502.835 1046.435 5503.115 1047.435 ;
    END
  END SET_IDB[31]
  PIN SET_IDB[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5642.835 1046.435 5643.115 1047.435 ;
    END
  END SET_IDB[32]
  PIN SET_IDB[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5782.835 1046.435 5783.115 1047.435 ;
    END
  END SET_IDB[33]
  PIN SET_IDB[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5922.835 1046.435 5923.115 1047.435 ;
    END
  END SET_IDB[34]
  PIN SET_IDB[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6062.835 1046.435 6063.115 1047.435 ;
    END
  END SET_IDB[35]
  PIN SET_IDB[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6202.835 1046.435 6203.115 1047.435 ;
    END
  END SET_IDB[36]
  PIN SET_IDB[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6342.835 1046.435 6343.115 1047.435 ;
    END
  END SET_IDB[37]
  PIN SET_IDB[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6482.835 1046.435 6483.115 1047.435 ;
    END
  END SET_IDB[38]
  PIN SET_IDB[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6622.835 1046.435 6623.115 1047.435 ;
    END
  END SET_IDB[39]
  PIN SET_IDB[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6762.835 1046.435 6763.115 1047.435 ;
    END
  END SET_IDB[40]
  PIN SET_IDB[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6902.835 1046.435 6903.115 1047.435 ;
    END
  END SET_IDB[41]
  PIN SET_IDB[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7042.835 1046.435 7043.115 1047.435 ;
    END
  END SET_IDB[42]
  PIN SET_IDB[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7182.835 1046.435 7183.115 1047.435 ;
    END
  END SET_IDB[43]
  PIN SET_IDB[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7322.835 1046.435 7323.115 1047.435 ;
    END
  END SET_IDB[44]
  PIN SET_IDB[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7462.835 1046.435 7463.115 1047.435 ;
    END
  END SET_IDB[45]
  PIN SET_IDB[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7602.835 1046.435 7603.115 1047.435 ;
    END
  END SET_IDB[46]
  PIN SET_IDB[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7742.835 1046.435 7743.115 1047.435 ;
    END
  END SET_IDB[47]
  PIN SET_IDB[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7882.835 1046.435 7883.115 1047.435 ;
    END
  END SET_IDB[48]
  PIN SET_IDB[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8022.835 1046.435 8023.115 1047.435 ;
    END
  END SET_IDB[49]
  PIN SET_IDB[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8162.835 1046.435 8163.115 1047.435 ;
    END
  END SET_IDB[50]
  PIN SET_IDB[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8302.835 1046.435 8303.115 1047.435 ;
    END
  END SET_IDB[51]
  PIN SET_IDB[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8442.835 1046.435 8443.115 1047.435 ;
    END
  END SET_IDB[52]
  PIN SET_IDB[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8582.835 1046.435 8583.115 1047.435 ;
    END
  END SET_IDB[53]
  PIN SET_IDB[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8722.835 1046.435 8723.115 1047.435 ;
    END
  END SET_IDB[54]
  PIN SET_IDB[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8862.835 1046.435 8863.115 1047.435 ;
    END
  END SET_IDB[55]
  PIN SET_IDB[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9002.835 1046.435 9003.115 1047.435 ;
    END
  END SET_IDB[56]
  PIN SET_IDB[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9142.835 1046.435 9143.115 1047.435 ;
    END
  END SET_IDB[57]
  PIN SET_IDB[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9282.835 1046.435 9283.115 1047.435 ;
    END
  END SET_IDB[58]
  PIN SET_IDB[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9422.835 1046.435 9423.115 1047.435 ;
    END
  END SET_IDB[59]
  PIN SET_IDB[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9562.835 1046.435 9563.115 1047.435 ;
    END
  END SET_IDB[60]
  PIN SET_IDB[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9702.835 1046.435 9703.115 1047.435 ;
    END
  END SET_IDB[61]
  PIN SET_IDB[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9842.835 1046.435 9843.115 1047.435 ;
    END
  END SET_IDB[62]
  PIN SET_IDB[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9982.835 1046.435 9983.115 1047.435 ;
    END
  END SET_IDB[63]
  PIN SET_IDB[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10122.835 1046.435 10123.115 1047.435 ;
    END
  END SET_IDB[64]
  PIN SET_IDB[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10262.835 1046.435 10263.115 1047.435 ;
    END
  END SET_IDB[65]
  PIN SET_IDB[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10402.835 1046.435 10403.115 1047.435 ;
    END
  END SET_IDB[66]
  PIN SET_IDB[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10542.835 1046.435 10543.115 1047.435 ;
    END
  END SET_IDB[67]
  PIN SET_IDB[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10682.835 1046.435 10683.115 1047.435 ;
    END
  END SET_IDB[68]
  PIN SET_IDB[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10822.835 1046.435 10823.115 1047.435 ;
    END
  END SET_IDB[69]
  PIN SET_IDB[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10962.835 1046.435 10963.115 1047.435 ;
    END
  END SET_IDB[70]
  PIN SET_IDB[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11102.835 1046.435 11103.115 1047.435 ;
    END
  END SET_IDB[71]
  PIN SET_IDB[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11242.835 1046.435 11243.115 1047.435 ;
    END
  END SET_IDB[72]
  PIN SET_IDB[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11382.835 1046.435 11383.115 1047.435 ;
    END
  END SET_IDB[73]
  PIN SET_IDB[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11522.835 1046.435 11523.115 1047.435 ;
    END
  END SET_IDB[74]
  PIN SET_IDB[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11662.835 1046.435 11663.115 1047.435 ;
    END
  END SET_IDB[75]
  PIN SET_IDB[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11802.835 1046.435 11803.115 1047.435 ;
    END
  END SET_IDB[76]
  PIN SET_IRESET[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8306.755 1046.435 8307.035 1047.435 ;
    END
  END SET_IRESET[51]
  PIN SET_IRESET[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8446.755 1046.435 8447.035 1047.435 ;
    END
  END SET_IRESET[52]
  PIN SET_IRESET[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8586.755 1046.435 8587.035 1047.435 ;
    END
  END SET_IRESET[53]
  PIN SET_IRESET[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8726.755 1046.435 8727.035 1047.435 ;
    END
  END SET_IRESET[54]
  PIN SET_IRESET[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8866.755 1046.435 8867.035 1047.435 ;
    END
  END SET_IRESET[55]
  PIN SET_IRESET[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9006.755 1046.435 9007.035 1047.435 ;
    END
  END SET_IRESET[56]
  PIN SET_IRESET[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9146.755 1046.435 9147.035 1047.435 ;
    END
  END SET_IRESET[57]
  PIN SET_IRESET[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9286.755 1046.435 9287.035 1047.435 ;
    END
  END SET_IRESET[58]
  PIN SET_IRESET[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9426.755 1046.435 9427.035 1047.435 ;
    END
  END SET_IRESET[59]
  PIN SET_IRESET[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9566.755 1046.435 9567.035 1047.435 ;
    END
  END SET_IRESET[60]
  PIN SET_IRESET[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9706.755 1046.435 9707.035 1047.435 ;
    END
  END SET_IRESET[61]
  PIN SET_IRESET[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9846.755 1046.435 9847.035 1047.435 ;
    END
  END SET_IRESET[62]
  PIN SET_IRESET[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9986.755 1046.435 9987.035 1047.435 ;
    END
  END SET_IRESET[63]
  PIN SET_IRESET[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10126.755 1046.435 10127.035 1047.435 ;
    END
  END SET_IRESET[64]
  PIN SET_IRESET[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10266.755 1046.435 10267.035 1047.435 ;
    END
  END SET_IRESET[65]
  PIN SET_IRESET[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10406.755 1046.435 10407.035 1047.435 ;
    END
  END SET_IRESET[66]
  PIN SET_IRESET[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10546.755 1046.435 10547.035 1047.435 ;
    END
  END SET_IRESET[67]
  PIN SET_IRESET[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10686.755 1046.435 10687.035 1047.435 ;
    END
  END SET_IRESET[68]
  PIN SET_IRESET[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10826.755 1046.435 10827.035 1047.435 ;
    END
  END SET_IRESET[69]
  PIN SET_IRESET[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10966.755 1046.435 10967.035 1047.435 ;
    END
  END SET_IRESET[70]
  PIN SET_IRESET[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11106.755 1046.435 11107.035 1047.435 ;
    END
  END SET_IRESET[71]
  PIN SET_IRESET[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11246.755 1046.435 11247.035 1047.435 ;
    END
  END SET_IRESET[72]
  PIN SET_IRESET[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11386.755 1046.435 11387.035 1047.435 ;
    END
  END SET_IRESET[73]
  PIN SET_IRESET[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11526.755 1046.435 11527.035 1047.435 ;
    END
  END SET_IRESET[74]
  PIN SET_IRESET[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11666.755 1046.435 11667.035 1047.435 ;
    END
  END SET_IRESET[75]
  PIN SET_IRESET[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11806.755 1046.435 11807.035 1047.435 ;
    END
  END SET_IRESET[76]
  PIN SET_IRESET[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11946.755 1046.435 11947.035 1047.435 ;
    END
  END SET_IRESET[77]
  PIN SET_IRESET[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12086.755 1046.435 12087.035 1047.435 ;
    END
  END SET_IRESET[78]
  PIN SET_IRESET[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12226.755 1046.435 12227.035 1047.435 ;
    END
  END SET_IRESET[79]
  PIN SET_IRESET[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12366.755 1046.435 12367.035 1047.435 ;
    END
  END SET_IRESET[80]
  PIN SET_IRESET[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12506.755 1046.435 12507.035 1047.435 ;
    END
  END SET_IRESET[81]
  PIN SET_IRESET[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12646.755 1046.435 12647.035 1047.435 ;
    END
  END SET_IRESET[82]
  PIN SET_IRESET[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12786.755 1046.435 12787.035 1047.435 ;
    END
  END SET_IRESET[83]
  PIN SET_IRESET[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12926.755 1046.435 12927.035 1047.435 ;
    END
  END SET_IRESET[84]
  PIN SET_IRESET[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13066.755 1046.435 13067.035 1047.435 ;
    END
  END SET_IRESET[85]
  PIN SET_IRESET[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13206.755 1046.435 13207.035 1047.435 ;
    END
  END SET_IRESET[86]
  PIN SET_IRESET[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13346.755 1046.435 13347.035 1047.435 ;
    END
  END SET_IRESET[87]
  PIN SET_IRESET[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13486.755 1046.435 13487.035 1047.435 ;
    END
  END SET_IRESET[88]
  PIN SET_IRESET[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13626.755 1046.435 13627.035 1047.435 ;
    END
  END SET_IRESET[89]
  PIN SET_IRESET[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13766.755 1046.435 13767.035 1047.435 ;
    END
  END SET_IRESET[90]
  PIN SET_IRESET[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13906.755 1046.435 13907.035 1047.435 ;
    END
  END SET_IRESET[91]
  PIN SET_IRESET[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14046.755 1046.435 14047.035 1047.435 ;
    END
  END SET_IRESET[92]
  PIN SET_IRESET[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14186.755 1046.435 14187.035 1047.435 ;
    END
  END SET_IRESET[93]
  PIN SET_IRESET[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14326.755 1046.435 14327.035 1047.435 ;
    END
  END SET_IRESET[94]
  PIN SET_IRESET[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14466.755 1046.435 14467.035 1047.435 ;
    END
  END SET_IRESET[95]
  PIN SET_IRESET[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14606.755 1046.435 14607.035 1047.435 ;
    END
  END SET_IRESET[96]
  PIN SET_IRESET[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14746.755 1046.435 14747.035 1047.435 ;
    END
  END SET_IRESET[97]
  PIN SET_IRESET[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14886.755 1046.435 14887.035 1047.435 ;
    END
  END SET_IRESET[98]
  PIN SET_IRESET[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15026.755 1046.435 15027.035 1047.435 ;
    END
  END SET_IRESET[99]
  PIN SET_IRESET[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15166.755 1046.435 15167.035 1047.435 ;
    END
  END SET_IRESET[100]
  PIN SET_IRESET[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15306.755 1046.435 15307.035 1047.435 ;
    END
  END SET_IRESET[101]
  PIN SET_IRESET[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15446.755 1046.435 15447.035 1047.435 ;
    END
  END SET_IRESET[102]
  PIN SET_IRESET[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15586.755 1046.435 15587.035 1047.435 ;
    END
  END SET_IRESET[103]
  PIN SET_IRESET[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15726.755 1046.435 15727.035 1047.435 ;
    END
  END SET_IRESET[104]
  PIN SET_IRESET[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15866.755 1046.435 15867.035 1047.435 ;
    END
  END SET_IRESET[105]
  PIN SET_IRESET[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16006.755 1046.435 16007.035 1047.435 ;
    END
  END SET_IRESET[106]
  PIN SET_IRESET[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16146.755 1046.435 16147.035 1047.435 ;
    END
  END SET_IRESET[107]
  PIN SET_IRESET[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16286.755 1046.435 16287.035 1047.435 ;
    END
  END SET_IRESET[108]
  PIN SET_IRESET[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16426.755 1046.435 16427.035 1047.435 ;
    END
  END SET_IRESET[109]
  PIN SET_IRESET[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16566.755 1046.435 16567.035 1047.435 ;
    END
  END SET_IRESET[110]
  PIN SET_IRESET[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16706.755 1046.435 16707.035 1047.435 ;
    END
  END SET_IRESET[111]
  PIN SET_IRESET[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16846.755 1046.435 16847.035 1047.435 ;
    END
  END SET_IRESET[112]
  PIN SET_IRESET[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16986.755 1046.435 16987.035 1047.435 ;
    END
  END SET_IRESET[113]
  PIN SET_IRESET[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17126.755 1046.435 17127.035 1047.435 ;
    END
  END SET_IRESET[114]
  PIN SET_IRESET[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17266.755 1046.435 17267.035 1047.435 ;
    END
  END SET_IRESET[115]
  PIN SET_IRESET[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17406.755 1046.435 17407.035 1047.435 ;
    END
  END SET_IRESET[116]
  PIN SET_IRESET[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17546.755 1046.435 17547.035 1047.435 ;
    END
  END SET_IRESET[117]
  PIN SET_IRESET[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17686.755 1046.435 17687.035 1047.435 ;
    END
  END SET_IRESET[118]
  PIN SET_IRESET[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17826.755 1046.435 17827.035 1047.435 ;
    END
  END SET_IRESET[119]
  PIN SET_IRESET[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17966.755 1046.435 17967.035 1047.435 ;
    END
  END SET_IRESET[120]
  PIN SET_IRESET[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18106.755 1046.435 18107.035 1047.435 ;
    END
  END SET_IRESET[121]
  PIN SET_IRESET[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18246.755 1046.435 18247.035 1047.435 ;
    END
  END SET_IRESET[122]
  PIN SET_IRESET[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18386.755 1046.435 18387.035 1047.435 ;
    END
  END SET_IRESET[123]
  PIN SET_IRESET[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18526.755 1046.435 18527.035 1047.435 ;
    END
  END SET_IRESET[124]
  PIN SET_IRESET[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18666.755 1046.435 18667.035 1047.435 ;
    END
  END SET_IRESET[125]
  PIN SET_IRESET[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18806.755 1046.435 18807.035 1047.435 ;
    END
  END SET_IRESET[126]
  PIN SET_IRESET[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18946.755 1046.435 18947.035 1047.435 ;
    END
  END SET_IRESET[127]
  PIN SET_ICASN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1170.675 1046.435 1170.955 1047.435 ;
    END
  END SET_ICASN[0]
  PIN SET_ICASN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1310.675 1046.435 1310.955 1047.435 ;
    END
  END SET_ICASN[1]
  PIN SET_ICASN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1450.675 1046.435 1450.955 1047.435 ;
    END
  END SET_ICASN[2]
  PIN SET_ICASN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1590.675 1046.435 1590.955 1047.435 ;
    END
  END SET_ICASN[3]
  PIN SET_ICASN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1730.675 1046.435 1730.955 1047.435 ;
    END
  END SET_ICASN[4]
  PIN SET_ICASN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1870.675 1046.435 1870.955 1047.435 ;
    END
  END SET_ICASN[5]
  PIN SET_ICASN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2010.675 1046.435 2010.955 1047.435 ;
    END
  END SET_ICASN[6]
  PIN SET_ICASN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2150.675 1046.435 2150.955 1047.435 ;
    END
  END SET_ICASN[7]
  PIN SET_ICASN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2290.675 1046.435 2290.955 1047.435 ;
    END
  END SET_ICASN[8]
  PIN SET_ICASN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2430.675 1046.435 2430.955 1047.435 ;
    END
  END SET_ICASN[9]
  PIN SET_ICASN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2570.675 1046.435 2570.955 1047.435 ;
    END
  END SET_ICASN[10]
  PIN SET_ICASN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2710.675 1046.435 2710.955 1047.435 ;
    END
  END SET_ICASN[11]
  PIN SET_ICASN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2850.675 1046.435 2850.955 1047.435 ;
    END
  END SET_ICASN[12]
  PIN SET_ICASN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2990.675 1046.435 2990.955 1047.435 ;
    END
  END SET_ICASN[13]
  PIN SET_ICASN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3130.675 1046.435 3130.955 1047.435 ;
    END
  END SET_ICASN[14]
  PIN SET_ICASN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3270.675 1046.435 3270.955 1047.435 ;
    END
  END SET_ICASN[15]
  PIN SET_ICASN[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3410.675 1046.435 3410.955 1047.435 ;
    END
  END SET_ICASN[16]
  PIN SET_ICASN[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3550.675 1046.435 3550.955 1047.435 ;
    END
  END SET_ICASN[17]
  PIN SET_ICASN[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3690.675 1046.435 3690.955 1047.435 ;
    END
  END SET_ICASN[18]
  PIN SET_ICASN[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3830.675 1046.435 3830.955 1047.435 ;
    END
  END SET_ICASN[19]
  PIN SET_ICASN[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3970.675 1046.435 3970.955 1047.435 ;
    END
  END SET_ICASN[20]
  PIN SET_ICASN[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4110.675 1046.435 4110.955 1047.435 ;
    END
  END SET_ICASN[21]
  PIN SET_ICASN[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4250.675 1046.435 4250.955 1047.435 ;
    END
  END SET_ICASN[22]
  PIN SET_ICASN[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4390.675 1046.435 4390.955 1047.435 ;
    END
  END SET_ICASN[23]
  PIN SET_ICASN[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4530.675 1046.435 4530.955 1047.435 ;
    END
  END SET_ICASN[24]
  PIN SET_ITHR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1438.915 1046.435 1439.195 1047.435 ;
    END
  END SET_ITHR[2]
  PIN SET_ITHR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1578.915 1046.435 1579.195 1047.435 ;
    END
  END SET_ITHR[3]
  PIN SET_ITHR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1718.915 1046.435 1719.195 1047.435 ;
    END
  END SET_ITHR[4]
  PIN SET_ITHR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1858.915 1046.435 1859.195 1047.435 ;
    END
  END SET_ITHR[5]
  PIN SET_ITHR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1998.915 1046.435 1999.195 1047.435 ;
    END
  END SET_ITHR[6]
  PIN SET_ITHR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2138.915 1046.435 2139.195 1047.435 ;
    END
  END SET_ITHR[7]
  PIN SET_ITHR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2278.915 1046.435 2279.195 1047.435 ;
    END
  END SET_ITHR[8]
  PIN SET_ITHR[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2418.915 1046.435 2419.195 1047.435 ;
    END
  END SET_ITHR[9]
  PIN SET_ITHR[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2558.915 1046.435 2559.195 1047.435 ;
    END
  END SET_ITHR[10]
  PIN SET_ITHR[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2698.915 1046.435 2699.195 1047.435 ;
    END
  END SET_ITHR[11]
  PIN SET_ITHR[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2838.915 1046.435 2839.195 1047.435 ;
    END
  END SET_ITHR[12]
  PIN SET_ITHR[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2978.915 1046.435 2979.195 1047.435 ;
    END
  END SET_ITHR[13]
  PIN SET_ITHR[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3118.915 1046.435 3119.195 1047.435 ;
    END
  END SET_ITHR[14]
  PIN SET_ITHR[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3258.915 1046.435 3259.195 1047.435 ;
    END
  END SET_ITHR[15]
  PIN SET_ITHR[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3398.915 1046.435 3399.195 1047.435 ;
    END
  END SET_ITHR[16]
  PIN SET_ITHR[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3538.915 1046.435 3539.195 1047.435 ;
    END
  END SET_ITHR[17]
  PIN SET_ITHR[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3678.915 1046.435 3679.195 1047.435 ;
    END
  END SET_ITHR[18]
  PIN SET_ITHR[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3818.915 1046.435 3819.195 1047.435 ;
    END
  END SET_ITHR[19]
  PIN SET_ITHR[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3958.915 1046.435 3959.195 1047.435 ;
    END
  END SET_ITHR[20]
  PIN SET_ITHR[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4098.915 1046.435 4099.195 1047.435 ;
    END
  END SET_ITHR[21]
  PIN SET_ITHR[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4238.915 1046.435 4239.195 1047.435 ;
    END
  END SET_ITHR[22]
  PIN SET_ITHR[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4378.915 1046.435 4379.195 1047.435 ;
    END
  END SET_ITHR[23]
  PIN SET_ITHR[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4518.915 1046.435 4519.195 1047.435 ;
    END
  END SET_ITHR[24]
  PIN SET_ITHR[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4658.915 1046.435 4659.195 1047.435 ;
    END
  END SET_ITHR[25]
  PIN SET_ITHR[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4798.915 1046.435 4799.195 1047.435 ;
    END
  END SET_ITHR[26]
  PIN SET_ITHR[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4938.915 1046.435 4939.195 1047.435 ;
    END
  END SET_ITHR[27]
  PIN SET_ITHR[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5078.915 1046.435 5079.195 1047.435 ;
    END
  END SET_ITHR[28]
  PIN SET_ITHR[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5218.915 1046.435 5219.195 1047.435 ;
    END
  END SET_ITHR[29]
  PIN SET_ITHR[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5358.915 1046.435 5359.195 1047.435 ;
    END
  END SET_ITHR[30]
  PIN SET_ITHR[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5498.915 1046.435 5499.195 1047.435 ;
    END
  END SET_ITHR[31]
  PIN SET_ITHR[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5638.915 1046.435 5639.195 1047.435 ;
    END
  END SET_ITHR[32]
  PIN SET_VCLIP[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19024.315 1046.435 19024.595 1047.435 ;
    END
  END SET_VCLIP[127]
  PIN SET_ITHR[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5778.915 1046.435 5779.195 1047.435 ;
    END
  END SET_ITHR[33]
  PIN SET_ITHR[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5918.915 1046.435 5919.195 1047.435 ;
    END
  END SET_ITHR[34]
  PIN SET_ITHR[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6058.915 1046.435 6059.195 1047.435 ;
    END
  END SET_ITHR[35]
  PIN SET_ITHR[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6198.915 1046.435 6199.195 1047.435 ;
    END
  END SET_ITHR[36]
  PIN SET_ITHR[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6338.915 1046.435 6339.195 1047.435 ;
    END
  END SET_ITHR[37]
  PIN SET_ITHR[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6478.915 1046.435 6479.195 1047.435 ;
    END
  END SET_ITHR[38]
  PIN SET_ITHR[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6618.915 1046.435 6619.195 1047.435 ;
    END
  END SET_ITHR[39]
  PIN SET_ITHR[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6758.915 1046.435 6759.195 1047.435 ;
    END
  END SET_ITHR[40]
  PIN SET_ITHR[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6898.915 1046.435 6899.195 1047.435 ;
    END
  END SET_ITHR[41]
  PIN SET_ITHR[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7038.915 1046.435 7039.195 1047.435 ;
    END
  END SET_ITHR[42]
  PIN SET_ITHR[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7178.915 1046.435 7179.195 1047.435 ;
    END
  END SET_ITHR[43]
  PIN SET_ITHR[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7318.915 1046.435 7319.195 1047.435 ;
    END
  END SET_ITHR[44]
  PIN SET_ITHR[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7458.915 1046.435 7459.195 1047.435 ;
    END
  END SET_ITHR[45]
  PIN SET_ITHR[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7598.915 1046.435 7599.195 1047.435 ;
    END
  END SET_ITHR[46]
  PIN SET_ITHR[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7738.915 1046.435 7739.195 1047.435 ;
    END
  END SET_ITHR[47]
  PIN SET_ITHR[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7878.915 1046.435 7879.195 1047.435 ;
    END
  END SET_ITHR[48]
  PIN SET_ITHR[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8018.915 1046.435 8019.195 1047.435 ;
    END
  END SET_ITHR[49]
  PIN SET_ITHR[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8158.915 1046.435 8159.195 1047.435 ;
    END
  END SET_ITHR[50]
  PIN SET_ITHR[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8298.915 1046.435 8299.195 1047.435 ;
    END
  END SET_ITHR[51]
  PIN SET_ITHR[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8438.915 1046.435 8439.195 1047.435 ;
    END
  END SET_ITHR[52]
  PIN SET_ITHR[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8578.915 1046.435 8579.195 1047.435 ;
    END
  END SET_ITHR[53]
  PIN SET_ITHR[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8718.915 1046.435 8719.195 1047.435 ;
    END
  END SET_ITHR[54]
  PIN SET_ITHR[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8858.915 1046.435 8859.195 1047.435 ;
    END
  END SET_ITHR[55]
  PIN SET_ITHR[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8998.915 1046.435 8999.195 1047.435 ;
    END
  END SET_ITHR[56]
  PIN SET_ITHR[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9138.915 1046.435 9139.195 1047.435 ;
    END
  END SET_ITHR[57]
  PIN SET_ITHR[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9278.915 1046.435 9279.195 1047.435 ;
    END
  END SET_ITHR[58]
  PIN SET_ITHR[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9418.915 1046.435 9419.195 1047.435 ;
    END
  END SET_ITHR[59]
  PIN SET_ITHR[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9558.915 1046.435 9559.195 1047.435 ;
    END
  END SET_ITHR[60]
  PIN SET_ITHR[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9698.915 1046.435 9699.195 1047.435 ;
    END
  END SET_ITHR[61]
  PIN SET_ITHR[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9838.915 1046.435 9839.195 1047.435 ;
    END
  END SET_ITHR[62]
  PIN SET_ITHR[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9978.915 1046.435 9979.195 1047.435 ;
    END
  END SET_ITHR[63]
  PIN SET_ITHR[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10118.915 1046.435 10119.195 1047.435 ;
    END
  END SET_ITHR[64]
  PIN SET_ITHR[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10258.915 1046.435 10259.195 1047.435 ;
    END
  END SET_ITHR[65]
  PIN SET_ITHR[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10398.915 1046.435 10399.195 1047.435 ;
    END
  END SET_ITHR[66]
  PIN SET_ITHR[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10538.915 1046.435 10539.195 1047.435 ;
    END
  END SET_ITHR[67]
  PIN SET_ITHR[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10678.915 1046.435 10679.195 1047.435 ;
    END
  END SET_ITHR[68]
  PIN SET_ITHR[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10818.915 1046.435 10819.195 1047.435 ;
    END
  END SET_ITHR[69]
  PIN SET_ITHR[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10958.915 1046.435 10959.195 1047.435 ;
    END
  END SET_ITHR[70]
  PIN SET_ITHR[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11098.915 1046.435 11099.195 1047.435 ;
    END
  END SET_ITHR[71]
  PIN SET_ITHR[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11238.915 1046.435 11239.195 1047.435 ;
    END
  END SET_ITHR[72]
  PIN SET_ITHR[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11378.915 1046.435 11379.195 1047.435 ;
    END
  END SET_ITHR[73]
  PIN SET_ITHR[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11518.915 1046.435 11519.195 1047.435 ;
    END
  END SET_ITHR[74]
  PIN SET_ITHR[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11658.915 1046.435 11659.195 1047.435 ;
    END
  END SET_ITHR[75]
  PIN SET_ITHR[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11798.915 1046.435 11799.195 1047.435 ;
    END
  END SET_ITHR[76]
  PIN SET_ITHR[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11938.915 1046.435 11939.195 1047.435 ;
    END
  END SET_ITHR[77]
  PIN SET_ITHR[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12078.915 1046.435 12079.195 1047.435 ;
    END
  END SET_ITHR[78]
  PIN SET_ITHR[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12218.915 1046.435 12219.195 1047.435 ;
    END
  END SET_ITHR[79]
  PIN SET_ITHR[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12358.915 1046.435 12359.195 1047.435 ;
    END
  END SET_ITHR[80]
  PIN SET_ITHR[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12498.915 1046.435 12499.195 1047.435 ;
    END
  END SET_ITHR[81]
  PIN SET_ITHR[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12638.915 1046.435 12639.195 1047.435 ;
    END
  END SET_ITHR[82]
  PIN SET_ITHR[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12778.915 1046.435 12779.195 1047.435 ;
    END
  END SET_ITHR[83]
  PIN SET_ITHR[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12918.915 1046.435 12919.195 1047.435 ;
    END
  END SET_ITHR[84]
  PIN SET_ITHR[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13058.915 1046.435 13059.195 1047.435 ;
    END
  END SET_ITHR[85]
  PIN SET_ITHR[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13198.915 1046.435 13199.195 1047.435 ;
    END
  END SET_ITHR[86]
  PIN SET_ITHR[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13338.915 1046.435 13339.195 1047.435 ;
    END
  END SET_ITHR[87]
  PIN SET_ITHR[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13478.915 1046.435 13479.195 1047.435 ;
    END
  END SET_ITHR[88]
  PIN SET_ITHR[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13618.915 1046.435 13619.195 1047.435 ;
    END
  END SET_ITHR[89]
  PIN SET_ITHR[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13758.915 1046.435 13759.195 1047.435 ;
    END
  END SET_ITHR[90]
  PIN SET_ITHR[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13898.915 1046.435 13899.195 1047.435 ;
    END
  END SET_ITHR[91]
  PIN SET_ITHR[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14038.915 1046.435 14039.195 1047.435 ;
    END
  END SET_ITHR[92]
  PIN SET_ITHR[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14178.915 1046.435 14179.195 1047.435 ;
    END
  END SET_ITHR[93]
  PIN SET_ITHR[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14318.915 1046.435 14319.195 1047.435 ;
    END
  END SET_ITHR[94]
  PIN SET_ITHR[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14458.915 1046.435 14459.195 1047.435 ;
    END
  END SET_ITHR[95]
  PIN SET_ITHR[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14598.915 1046.435 14599.195 1047.435 ;
    END
  END SET_ITHR[96]
  PIN SET_ITHR[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14738.915 1046.435 14739.195 1047.435 ;
    END
  END SET_ITHR[97]
  PIN SET_ITHR[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14878.915 1046.435 14879.195 1047.435 ;
    END
  END SET_ITHR[98]
  PIN SET_ITHR[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15018.915 1046.435 15019.195 1047.435 ;
    END
  END SET_ITHR[99]
  PIN SET_ITHR[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15158.915 1046.435 15159.195 1047.435 ;
    END
  END SET_ITHR[100]
  PIN SET_ITHR[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15298.915 1046.435 15299.195 1047.435 ;
    END
  END SET_ITHR[101]
  PIN SET_ITHR[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15438.915 1046.435 15439.195 1047.435 ;
    END
  END SET_ITHR[102]
  PIN SET_IBIAS[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1154.995 1046.435 1155.275 1047.435 ;
    END
  END SET_IBIAS[0]
  PIN SET_IBIAS[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1294.995 1046.435 1295.275 1047.435 ;
    END
  END SET_IBIAS[1]
  PIN SET_IBIAS[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1434.995 1046.435 1435.275 1047.435 ;
    END
  END SET_IBIAS[2]
  PIN SET_IBIAS[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1574.995 1046.435 1575.275 1047.435 ;
    END
  END SET_IBIAS[3]
  PIN SET_IBIAS[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1714.995 1046.435 1715.275 1047.435 ;
    END
  END SET_IBIAS[4]
  PIN SET_IBIAS[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1854.995 1046.435 1855.275 1047.435 ;
    END
  END SET_IBIAS[5]
  PIN SET_IBIAS[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1994.995 1046.435 1995.275 1047.435 ;
    END
  END SET_IBIAS[6]
  PIN SET_IBIAS[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2134.995 1046.435 2135.275 1047.435 ;
    END
  END SET_IBIAS[7]
  PIN SET_IBIAS[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2274.995 1046.435 2275.275 1047.435 ;
    END
  END SET_IBIAS[8]
  PIN SET_IBIAS[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2414.995 1046.435 2415.275 1047.435 ;
    END
  END SET_IBIAS[9]
  PIN SET_IBIAS[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2554.995 1046.435 2555.275 1047.435 ;
    END
  END SET_IBIAS[10]
  PIN SET_IBIAS[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2694.995 1046.435 2695.275 1047.435 ;
    END
  END SET_IBIAS[11]
  PIN SET_IBIAS[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2834.995 1046.435 2835.275 1047.435 ;
    END
  END SET_IBIAS[12]
  PIN SET_IBIAS[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2974.995 1046.435 2975.275 1047.435 ;
    END
  END SET_IBIAS[13]
  PIN SET_IBIAS[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3114.995 1046.435 3115.275 1047.435 ;
    END
  END SET_IBIAS[14]
  PIN SET_IBIAS[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3254.995 1046.435 3255.275 1047.435 ;
    END
  END SET_IBIAS[15]
  PIN SET_IBIAS[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3394.995 1046.435 3395.275 1047.435 ;
    END
  END SET_IBIAS[16]
  PIN SET_IBIAS[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3534.995 1046.435 3535.275 1047.435 ;
    END
  END SET_IBIAS[17]
  PIN SET_IBIAS[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3674.995 1046.435 3675.275 1047.435 ;
    END
  END SET_IBIAS[18]
  PIN SET_IBIAS[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3814.995 1046.435 3815.275 1047.435 ;
    END
  END SET_IBIAS[19]
  PIN SET_IBIAS[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3954.995 1046.435 3955.275 1047.435 ;
    END
  END SET_IBIAS[20]
  PIN SET_IBIAS[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4094.995 1046.435 4095.275 1047.435 ;
    END
  END SET_IBIAS[21]
  PIN SET_IBIAS[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4234.995 1046.435 4235.275 1047.435 ;
    END
  END SET_IBIAS[22]
  PIN SET_IBIAS[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4374.995 1046.435 4375.275 1047.435 ;
    END
  END SET_IBIAS[23]
  PIN SET_IBIAS[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4514.995 1046.435 4515.275 1047.435 ;
    END
  END SET_IBIAS[24]
  PIN SET_IBIAS[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4654.995 1046.435 4655.275 1047.435 ;
    END
  END SET_IBIAS[25]
  PIN SET_IBIAS[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4794.995 1046.435 4795.275 1047.435 ;
    END
  END SET_IBIAS[26]
  PIN SET_IBIAS[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4934.995 1046.435 4935.275 1047.435 ;
    END
  END SET_IBIAS[27]
  PIN SET_IBIAS[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5074.995 1046.435 5075.275 1047.435 ;
    END
  END SET_IBIAS[28]
  PIN SET_IBIAS[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5214.995 1046.435 5215.275 1047.435 ;
    END
  END SET_IBIAS[29]
  PIN SET_IBIAS[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5354.995 1046.435 5355.275 1047.435 ;
    END
  END SET_IBIAS[30]
  PIN SET_IBIAS[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5494.995 1046.435 5495.275 1047.435 ;
    END
  END SET_IBIAS[31]
  PIN SET_IBIAS[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5634.995 1046.435 5635.275 1047.435 ;
    END
  END SET_IBIAS[32]
  PIN SET_IBIAS[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5774.995 1046.435 5775.275 1047.435 ;
    END
  END SET_IBIAS[33]
  PIN SET_IBIAS[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5914.995 1046.435 5915.275 1047.435 ;
    END
  END SET_IBIAS[34]
  PIN SET_IBIAS[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6054.995 1046.435 6055.275 1047.435 ;
    END
  END SET_IBIAS[35]
  PIN SET_IBIAS[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6194.995 1046.435 6195.275 1047.435 ;
    END
  END SET_IBIAS[36]
  PIN SET_IBIAS[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6334.995 1046.435 6335.275 1047.435 ;
    END
  END SET_IBIAS[37]
  PIN SET_IBIAS[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6474.995 1046.435 6475.275 1047.435 ;
    END
  END SET_IBIAS[38]
  PIN SET_IBIAS[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6614.995 1046.435 6615.275 1047.435 ;
    END
  END SET_IBIAS[39]
  PIN SET_IBIAS[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6754.995 1046.435 6755.275 1047.435 ;
    END
  END SET_IBIAS[40]
  PIN SET_IBIAS[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6894.995 1046.435 6895.275 1047.435 ;
    END
  END SET_IBIAS[41]
  PIN SET_IBIAS[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7034.995 1046.435 7035.275 1047.435 ;
    END
  END SET_IBIAS[42]
  PIN SET_IBIAS[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7174.995 1046.435 7175.275 1047.435 ;
    END
  END SET_IBIAS[43]
  PIN SET_IBIAS[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7314.995 1046.435 7315.275 1047.435 ;
    END
  END SET_IBIAS[44]
  PIN SET_IBIAS[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7454.995 1046.435 7455.275 1047.435 ;
    END
  END SET_IBIAS[45]
  PIN SET_IBIAS[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7594.995 1046.435 7595.275 1047.435 ;
    END
  END SET_IBIAS[46]
  PIN SET_IBIAS[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7734.995 1046.435 7735.275 1047.435 ;
    END
  END SET_IBIAS[47]
  PIN SET_IBIAS[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7874.995 1046.435 7875.275 1047.435 ;
    END
  END SET_IBIAS[48]
  PIN SET_IBIAS[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8014.995 1046.435 8015.275 1047.435 ;
    END
  END SET_IBIAS[49]
  PIN SET_IBIAS[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8154.995 1046.435 8155.275 1047.435 ;
    END
  END SET_IBIAS[50]
  PIN SET_IBIAS[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8294.995 1046.435 8295.275 1047.435 ;
    END
  END SET_IBIAS[51]
  PIN SET_IBIAS[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8434.995 1046.435 8435.275 1047.435 ;
    END
  END SET_IBIAS[52]
  PIN SET_IBIAS[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8574.995 1046.435 8575.275 1047.435 ;
    END
  END SET_IBIAS[53]
  PIN SET_IBIAS[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8714.995 1046.435 8715.275 1047.435 ;
    END
  END SET_IBIAS[54]
  PIN SET_IBIAS[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8854.995 1046.435 8855.275 1047.435 ;
    END
  END SET_IBIAS[55]
  PIN SET_IBIAS[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8994.995 1046.435 8995.275 1047.435 ;
    END
  END SET_IBIAS[56]
  PIN SET_IBIAS[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9134.995 1046.435 9135.275 1047.435 ;
    END
  END SET_IBIAS[57]
  PIN SET_IBIAS[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9274.995 1046.435 9275.275 1047.435 ;
    END
  END SET_IBIAS[58]
  PIN SET_IBIAS[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9414.995 1046.435 9415.275 1047.435 ;
    END
  END SET_IBIAS[59]
  PIN SET_IBIAS[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9554.995 1046.435 9555.275 1047.435 ;
    END
  END SET_IBIAS[60]
  PIN SET_IBIAS[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9694.995 1046.435 9695.275 1047.435 ;
    END
  END SET_IBIAS[61]
  PIN SET_IBIAS[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9834.995 1046.435 9835.275 1047.435 ;
    END
  END SET_IBIAS[62]
  PIN SET_IBIAS[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9974.995 1046.435 9975.275 1047.435 ;
    END
  END SET_IBIAS[63]
  PIN SET_IBIAS[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10114.995 1046.435 10115.275 1047.435 ;
    END
  END SET_IBIAS[64]
  PIN SET_IBIAS[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10254.995 1046.435 10255.275 1047.435 ;
    END
  END SET_IBIAS[65]
  PIN SET_IBIAS[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10394.995 1046.435 10395.275 1047.435 ;
    END
  END SET_IBIAS[66]
  PIN SET_IBIAS[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10534.995 1046.435 10535.275 1047.435 ;
    END
  END SET_IBIAS[67]
  PIN SET_IBIAS[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10674.995 1046.435 10675.275 1047.435 ;
    END
  END SET_IBIAS[68]
  PIN SET_IBIAS[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10814.995 1046.435 10815.275 1047.435 ;
    END
  END SET_IBIAS[69]
  PIN SET_IBIAS[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10954.995 1046.435 10955.275 1047.435 ;
    END
  END SET_IBIAS[70]
  PIN SET_IBIAS[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11094.995 1046.435 11095.275 1047.435 ;
    END
  END SET_IBIAS[71]
  PIN SET_IBIAS[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11234.995 1046.435 11235.275 1047.435 ;
    END
  END SET_IBIAS[72]
  PIN SET_IBIAS[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11374.995 1046.435 11375.275 1047.435 ;
    END
  END SET_IBIAS[73]
  PIN SET_IBIAS[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11514.995 1046.435 11515.275 1047.435 ;
    END
  END SET_IBIAS[74]
  PIN SET_IBIAS[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11654.995 1046.435 11655.275 1047.435 ;
    END
  END SET_IBIAS[75]
  PIN SET_IBIAS[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11794.995 1046.435 11795.275 1047.435 ;
    END
  END SET_IBIAS[76]
  PIN SET_IBIAS[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11934.995 1046.435 11935.275 1047.435 ;
    END
  END SET_IBIAS[77]
  PIN SET_IBIAS[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12074.995 1046.435 12075.275 1047.435 ;
    END
  END SET_IBIAS[78]
  PIN SET_IBIAS[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12214.995 1046.435 12215.275 1047.435 ;
    END
  END SET_IBIAS[79]
  PIN SET_IBIAS[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12354.995 1046.435 12355.275 1047.435 ;
    END
  END SET_IBIAS[80]
  PIN SET_IBIAS[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12494.995 1046.435 12495.275 1047.435 ;
    END
  END SET_IBIAS[81]
  PIN SET_IBIAS[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12634.995 1046.435 12635.275 1047.435 ;
    END
  END SET_IBIAS[82]
  PIN SET_IBIAS[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12774.995 1046.435 12775.275 1047.435 ;
    END
  END SET_IBIAS[83]
  PIN SET_IBIAS[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12914.995 1046.435 12915.275 1047.435 ;
    END
  END SET_IBIAS[84]
  PIN SET_IBIAS[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13054.995 1046.435 13055.275 1047.435 ;
    END
  END SET_IBIAS[85]
  PIN SET_IBIAS[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13194.995 1046.435 13195.275 1047.435 ;
    END
  END SET_IBIAS[86]
  PIN SET_IBIAS[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13334.995 1046.435 13335.275 1047.435 ;
    END
  END SET_IBIAS[87]
  PIN SET_IBIAS[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13474.995 1046.435 13475.275 1047.435 ;
    END
  END SET_IBIAS[88]
  PIN SET_IBIAS[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13614.995 1046.435 13615.275 1047.435 ;
    END
  END SET_IBIAS[89]
  PIN SET_IBIAS[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13754.995 1046.435 13755.275 1047.435 ;
    END
  END SET_IBIAS[90]
  PIN SET_IBIAS[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13894.995 1046.435 13895.275 1047.435 ;
    END
  END SET_IBIAS[91]
  PIN SET_IBIAS[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14034.995 1046.435 14035.275 1047.435 ;
    END
  END SET_IBIAS[92]
  PIN SET_IBIAS[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14174.995 1046.435 14175.275 1047.435 ;
    END
  END SET_IBIAS[93]
  PIN SET_IBIAS[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14314.995 1046.435 14315.275 1047.435 ;
    END
  END SET_IBIAS[94]
  PIN SET_IBIAS[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14454.995 1046.435 14455.275 1047.435 ;
    END
  END SET_IBIAS[95]
  PIN SET_IBIAS[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14594.995 1046.435 14595.275 1047.435 ;
    END
  END SET_IBIAS[96]
  PIN SET_IBIAS[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14734.995 1046.435 14735.275 1047.435 ;
    END
  END SET_IBIAS[97]
  PIN SET_IBIAS[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14874.995 1046.435 14875.275 1047.435 ;
    END
  END SET_IBIAS[98]
  PIN SET_IBIAS[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15014.995 1046.435 15015.275 1047.435 ;
    END
  END SET_IBIAS[99]
  PIN SET_IBIAS[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15154.995 1046.435 15155.275 1047.435 ;
    END
  END SET_IBIAS[100]
  PIN SET_IBIAS[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15294.995 1046.435 15295.275 1047.435 ;
    END
  END SET_IBIAS[101]
  PIN SET_IBIAS[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15434.995 1046.435 15435.275 1047.435 ;
    END
  END SET_IBIAS[102]
  PIN SET_IBIAS[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15574.995 1046.435 15575.275 1047.435 ;
    END
  END SET_IBIAS[103]
  PIN SET_IBIAS[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15714.995 1046.435 15715.275 1047.435 ;
    END
  END SET_IBIAS[104]
  PIN SET_IBIAS[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15854.995 1046.435 15855.275 1047.435 ;
    END
  END SET_IBIAS[105]
  PIN SET_IBIAS[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15994.995 1046.435 15995.275 1047.435 ;
    END
  END SET_IBIAS[106]
  PIN SET_IBIAS[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16134.995 1046.435 16135.275 1047.435 ;
    END
  END SET_IBIAS[107]
  PIN SET_IBIAS[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16274.995 1046.435 16275.275 1047.435 ;
    END
  END SET_IBIAS[108]
  PIN SET_IBIAS[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16414.995 1046.435 16415.275 1047.435 ;
    END
  END SET_IBIAS[109]
  PIN SET_IBIAS[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16554.995 1046.435 16555.275 1047.435 ;
    END
  END SET_IBIAS[110]
  PIN SET_IBIAS[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16694.995 1046.435 16695.275 1047.435 ;
    END
  END SET_IBIAS[111]
  PIN SET_IBIAS[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16834.995 1046.435 16835.275 1047.435 ;
    END
  END SET_IBIAS[112]
  PIN SET_IBIAS[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16974.995 1046.435 16975.275 1047.435 ;
    END
  END SET_IBIAS[113]
  PIN SET_IBIAS[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17114.995 1046.435 17115.275 1047.435 ;
    END
  END SET_IBIAS[114]
  PIN SET_IBIAS[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17254.995 1046.435 17255.275 1047.435 ;
    END
  END SET_IBIAS[115]
  PIN SET_IBIAS[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17394.995 1046.435 17395.275 1047.435 ;
    END
  END SET_IBIAS[116]
  PIN SET_IBIAS[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17534.995 1046.435 17535.275 1047.435 ;
    END
  END SET_IBIAS[117]
  PIN SET_IBIAS[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17674.995 1046.435 17675.275 1047.435 ;
    END
  END SET_IBIAS[118]
  PIN SET_IBIAS[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17814.995 1046.435 17815.275 1047.435 ;
    END
  END SET_IBIAS[119]
  PIN SET_IBIAS[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17954.995 1046.435 17955.275 1047.435 ;
    END
  END SET_IBIAS[120]
  PIN SET_IBIAS[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18094.995 1046.435 18095.275 1047.435 ;
    END
  END SET_IBIAS[121]
  PIN SET_IBIAS[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18234.995 1046.435 18235.275 1047.435 ;
    END
  END SET_IBIAS[122]
  PIN SET_IBIAS[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18374.995 1046.435 18375.275 1047.435 ;
    END
  END SET_IBIAS[123]
  PIN SET_IBIAS[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18514.995 1046.435 18515.275 1047.435 ;
    END
  END SET_IBIAS[124]
  PIN SET_IBIAS[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18654.995 1046.435 18655.275 1047.435 ;
    END
  END SET_IBIAS[125]
  PIN SET_IBIAS[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18794.995 1046.435 18795.275 1047.435 ;
    END
  END SET_IBIAS[126]
  PIN SET_IBIAS[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18934.995 1046.435 18935.275 1047.435 ;
    END
  END SET_IBIAS[127]
  PIN SET_ITHR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1158.915 1046.435 1159.195 1047.435 ;
    END
  END SET_ITHR[0]
  PIN SET_ITHR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1298.915 1046.435 1299.195 1047.435 ;
    END
  END SET_ITHR[1]
  PIN SET_IDB[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11942.835 1046.435 11943.115 1047.435 ;
    END
  END SET_IDB[77]
  PIN SET_IDB[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12082.835 1046.435 12083.115 1047.435 ;
    END
  END SET_IDB[78]
  PIN SET_IDB[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12222.835 1046.435 12223.115 1047.435 ;
    END
  END SET_IDB[79]
  PIN SET_IDB[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12362.835 1046.435 12363.115 1047.435 ;
    END
  END SET_IDB[80]
  PIN SET_IDB[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12502.835 1046.435 12503.115 1047.435 ;
    END
  END SET_IDB[81]
  PIN SET_IDB[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12642.835 1046.435 12643.115 1047.435 ;
    END
  END SET_IDB[82]
  PIN SET_IDB[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12782.835 1046.435 12783.115 1047.435 ;
    END
  END SET_IDB[83]
  PIN SET_IDB[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12922.835 1046.435 12923.115 1047.435 ;
    END
  END SET_IDB[84]
  PIN SET_IDB[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13062.835 1046.435 13063.115 1047.435 ;
    END
  END SET_IDB[85]
  PIN SET_IDB[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13202.835 1046.435 13203.115 1047.435 ;
    END
  END SET_IDB[86]
  PIN SET_IDB[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13342.835 1046.435 13343.115 1047.435 ;
    END
  END SET_IDB[87]
  PIN SET_IDB[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13482.835 1046.435 13483.115 1047.435 ;
    END
  END SET_IDB[88]
  PIN SET_IDB[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13622.835 1046.435 13623.115 1047.435 ;
    END
  END SET_IDB[89]
  PIN SET_IDB[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13762.835 1046.435 13763.115 1047.435 ;
    END
  END SET_IDB[90]
  PIN SET_IDB[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13902.835 1046.435 13903.115 1047.435 ;
    END
  END SET_IDB[91]
  PIN SET_IDB[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14042.835 1046.435 14043.115 1047.435 ;
    END
  END SET_IDB[92]
  PIN SET_IDB[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14182.835 1046.435 14183.115 1047.435 ;
    END
  END SET_IDB[93]
  PIN SET_IDB[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14322.835 1046.435 14323.115 1047.435 ;
    END
  END SET_IDB[94]
  PIN SET_IDB[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14462.835 1046.435 14463.115 1047.435 ;
    END
  END SET_IDB[95]
  PIN SET_IDB[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14602.835 1046.435 14603.115 1047.435 ;
    END
  END SET_IDB[96]
  PIN SET_IDB[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14742.835 1046.435 14743.115 1047.435 ;
    END
  END SET_IDB[97]
  PIN SET_IDB[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14882.835 1046.435 14883.115 1047.435 ;
    END
  END SET_IDB[98]
  PIN SET_IDB[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15022.835 1046.435 15023.115 1047.435 ;
    END
  END SET_IDB[99]
  PIN SET_IDB[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15162.835 1046.435 15163.115 1047.435 ;
    END
  END SET_IDB[100]
  PIN SET_IDB[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15302.835 1046.435 15303.115 1047.435 ;
    END
  END SET_IDB[101]
  PIN SET_IDB[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15442.835 1046.435 15443.115 1047.435 ;
    END
  END SET_IDB[102]
  PIN SET_IDB[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15582.835 1046.435 15583.115 1047.435 ;
    END
  END SET_IDB[103]
  PIN SET_IDB[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15722.835 1046.435 15723.115 1047.435 ;
    END
  END SET_IDB[104]
  PIN SET_IDB[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15862.835 1046.435 15863.115 1047.435 ;
    END
  END SET_IDB[105]
  PIN SET_IDB[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16002.835 1046.435 16003.115 1047.435 ;
    END
  END SET_IDB[106]
  PIN SET_IDB[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16142.835 1046.435 16143.115 1047.435 ;
    END
  END SET_IDB[107]
  PIN SET_IDB[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16282.835 1046.435 16283.115 1047.435 ;
    END
  END SET_IDB[108]
  PIN SET_IDB[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16422.835 1046.435 16423.115 1047.435 ;
    END
  END SET_IDB[109]
  PIN SET_IDB[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16562.835 1046.435 16563.115 1047.435 ;
    END
  END SET_IDB[110]
  PIN SET_IDB[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16702.835 1046.435 16703.115 1047.435 ;
    END
  END SET_IDB[111]
  PIN SET_IDB[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16842.835 1046.435 16843.115 1047.435 ;
    END
  END SET_IDB[112]
  PIN SET_IDB[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16982.835 1046.435 16983.115 1047.435 ;
    END
  END SET_IDB[113]
  PIN SET_IDB[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17122.835 1046.435 17123.115 1047.435 ;
    END
  END SET_IDB[114]
  PIN SET_IDB[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17262.835 1046.435 17263.115 1047.435 ;
    END
  END SET_IDB[115]
  PIN SET_IDB[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17402.835 1046.435 17403.115 1047.435 ;
    END
  END SET_IDB[116]
  PIN SET_IDB[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17542.835 1046.435 17543.115 1047.435 ;
    END
  END SET_IDB[117]
  PIN SET_IDB[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17682.835 1046.435 17683.115 1047.435 ;
    END
  END SET_IDB[118]
  PIN SET_IDB[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17822.835 1046.435 17823.115 1047.435 ;
    END
  END SET_IDB[119]
  PIN SET_IDB[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17962.835 1046.435 17963.115 1047.435 ;
    END
  END SET_IDB[120]
  PIN SET_IDB[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18102.835 1046.435 18103.115 1047.435 ;
    END
  END SET_IDB[121]
  PIN SET_IDB[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18242.835 1046.435 18243.115 1047.435 ;
    END
  END SET_IDB[122]
  PIN SET_IDB[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18382.835 1046.435 18383.115 1047.435 ;
    END
  END SET_IDB[123]
  PIN SET_IDB[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18522.835 1046.435 18523.115 1047.435 ;
    END
  END SET_IDB[124]
  PIN SET_IDB[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18662.835 1046.435 18663.115 1047.435 ;
    END
  END SET_IDB[125]
  PIN SET_IDB[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18802.835 1046.435 18803.115 1047.435 ;
    END
  END SET_IDB[126]
  PIN SET_IDB[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18942.835 1046.435 18943.115 1047.435 ;
    END
  END SET_IDB[127]
  PIN SET_IRESET[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1166.755 1046.435 1167.035 1047.435 ;
    END
  END SET_IRESET[0]
  PIN SET_IRESET[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1306.755 1046.435 1307.035 1047.435 ;
    END
  END SET_IRESET[1]
  PIN SET_IRESET[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1446.755 1046.435 1447.035 1047.435 ;
    END
  END SET_IRESET[2]
  PIN SET_IRESET[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1586.755 1046.435 1587.035 1047.435 ;
    END
  END SET_IRESET[3]
  PIN SET_IRESET[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1726.755 1046.435 1727.035 1047.435 ;
    END
  END SET_IRESET[4]
  PIN SET_IRESET[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1866.755 1046.435 1867.035 1047.435 ;
    END
  END SET_IRESET[5]
  PIN SET_IRESET[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2006.755 1046.435 2007.035 1047.435 ;
    END
  END SET_IRESET[6]
  PIN SET_IRESET[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2146.755 1046.435 2147.035 1047.435 ;
    END
  END SET_IRESET[7]
  PIN SET_IRESET[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2286.755 1046.435 2287.035 1047.435 ;
    END
  END SET_IRESET[8]
  PIN SET_IRESET[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2426.755 1046.435 2427.035 1047.435 ;
    END
  END SET_IRESET[9]
  PIN SET_IRESET[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2566.755 1046.435 2567.035 1047.435 ;
    END
  END SET_IRESET[10]
  PIN SET_IRESET[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2706.755 1046.435 2707.035 1047.435 ;
    END
  END SET_IRESET[11]
  PIN SET_IRESET[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2846.755 1046.435 2847.035 1047.435 ;
    END
  END SET_IRESET[12]
  PIN SET_IRESET[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2986.755 1046.435 2987.035 1047.435 ;
    END
  END SET_IRESET[13]
  PIN SET_IRESET[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3126.755 1046.435 3127.035 1047.435 ;
    END
  END SET_IRESET[14]
  PIN SET_IRESET[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3266.755 1046.435 3267.035 1047.435 ;
    END
  END SET_IRESET[15]
  PIN SET_IRESET[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3406.755 1046.435 3407.035 1047.435 ;
    END
  END SET_IRESET[16]
  PIN SET_IRESET[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3546.755 1046.435 3547.035 1047.435 ;
    END
  END SET_IRESET[17]
  PIN SET_IRESET[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3686.755 1046.435 3687.035 1047.435 ;
    END
  END SET_IRESET[18]
  PIN SET_IRESET[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3826.755 1046.435 3827.035 1047.435 ;
    END
  END SET_IRESET[19]
  PIN SET_IRESET[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3966.755 1046.435 3967.035 1047.435 ;
    END
  END SET_IRESET[20]
  PIN SET_IRESET[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4106.755 1046.435 4107.035 1047.435 ;
    END
  END SET_IRESET[21]
  PIN SET_IRESET[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4246.755 1046.435 4247.035 1047.435 ;
    END
  END SET_IRESET[22]
  PIN SET_IRESET[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4386.755 1046.435 4387.035 1047.435 ;
    END
  END SET_IRESET[23]
  PIN SET_IRESET[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4526.755 1046.435 4527.035 1047.435 ;
    END
  END SET_IRESET[24]
  PIN SET_IRESET[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4666.755 1046.435 4667.035 1047.435 ;
    END
  END SET_IRESET[25]
  PIN SET_IRESET[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4806.755 1046.435 4807.035 1047.435 ;
    END
  END SET_IRESET[26]
  PIN SET_IRESET[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4946.755 1046.435 4947.035 1047.435 ;
    END
  END SET_IRESET[27]
  PIN SET_IRESET[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5086.755 1046.435 5087.035 1047.435 ;
    END
  END SET_IRESET[28]
  PIN SET_IRESET[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5226.755 1046.435 5227.035 1047.435 ;
    END
  END SET_IRESET[29]
  PIN SET_IRESET[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5366.755 1046.435 5367.035 1047.435 ;
    END
  END SET_IRESET[30]
  PIN SET_IRESET[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5506.755 1046.435 5507.035 1047.435 ;
    END
  END SET_IRESET[31]
  PIN SET_IRESET[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5646.755 1046.435 5647.035 1047.435 ;
    END
  END SET_IRESET[32]
  PIN SET_IRESET[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5786.755 1046.435 5787.035 1047.435 ;
    END
  END SET_IRESET[33]
  PIN SET_IRESET[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5926.755 1046.435 5927.035 1047.435 ;
    END
  END SET_IRESET[34]
  PIN SET_IRESET[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6066.755 1046.435 6067.035 1047.435 ;
    END
  END SET_IRESET[35]
  PIN SET_IRESET[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6206.755 1046.435 6207.035 1047.435 ;
    END
  END SET_IRESET[36]
  PIN SET_IRESET[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6346.755 1046.435 6347.035 1047.435 ;
    END
  END SET_IRESET[37]
  PIN SET_IRESET[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6486.755 1046.435 6487.035 1047.435 ;
    END
  END SET_IRESET[38]
  PIN SET_IRESET[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6626.755 1046.435 6627.035 1047.435 ;
    END
  END SET_IRESET[39]
  PIN SET_IRESET[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6766.755 1046.435 6767.035 1047.435 ;
    END
  END SET_IRESET[40]
  PIN SET_IRESET[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6906.755 1046.435 6907.035 1047.435 ;
    END
  END SET_IRESET[41]
  PIN SET_IRESET[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7046.755 1046.435 7047.035 1047.435 ;
    END
  END SET_IRESET[42]
  PIN SET_IRESET[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7186.755 1046.435 7187.035 1047.435 ;
    END
  END SET_IRESET[43]
  PIN SET_IRESET[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7326.755 1046.435 7327.035 1047.435 ;
    END
  END SET_IRESET[44]
  PIN SET_IRESET[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7466.755 1046.435 7467.035 1047.435 ;
    END
  END SET_IRESET[45]
  PIN SET_IRESET[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7606.755 1046.435 7607.035 1047.435 ;
    END
  END SET_IRESET[46]
  PIN SET_IRESET[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7746.755 1046.435 7747.035 1047.435 ;
    END
  END SET_IRESET[47]
  PIN SET_IRESET[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7886.755 1046.435 7887.035 1047.435 ;
    END
  END SET_IRESET[48]
  PIN SET_IRESET[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8026.755 1046.435 8027.035 1047.435 ;
    END
  END SET_IRESET[49]
  PIN SET_IRESET[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8166.755 1046.435 8167.035 1047.435 ;
    END
  END SET_IRESET[50]
  PIN SET_ICASN[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4670.675 1046.435 4670.955 1047.435 ;
    END
  END SET_ICASN[25]
  PIN SET_ICASN[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4810.675 1046.435 4810.955 1047.435 ;
    END
  END SET_ICASN[26]
  PIN SET_ICASN[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4950.675 1046.435 4950.955 1047.435 ;
    END
  END SET_ICASN[27]
  PIN SET_ICASN[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5090.675 1046.435 5090.955 1047.435 ;
    END
  END SET_ICASN[28]
  PIN SET_ICASN[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5230.675 1046.435 5230.955 1047.435 ;
    END
  END SET_ICASN[29]
  PIN SET_ICASN[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5370.675 1046.435 5370.955 1047.435 ;
    END
  END SET_ICASN[30]
  PIN SET_ICASN[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5510.675 1046.435 5510.955 1047.435 ;
    END
  END SET_ICASN[31]
  PIN SET_ICASN[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5650.675 1046.435 5650.955 1047.435 ;
    END
  END SET_ICASN[32]
  PIN SET_ICASN[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5790.675 1046.435 5790.955 1047.435 ;
    END
  END SET_ICASN[33]
  PIN SET_ICASN[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5930.675 1046.435 5930.955 1047.435 ;
    END
  END SET_ICASN[34]
  PIN SET_ICASN[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6070.675 1046.435 6070.955 1047.435 ;
    END
  END SET_ICASN[35]
  PIN SET_ICASN[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6210.675 1046.435 6210.955 1047.435 ;
    END
  END SET_ICASN[36]
  PIN SET_ICASN[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6350.675 1046.435 6350.955 1047.435 ;
    END
  END SET_ICASN[37]
  PIN SET_ICASN[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6490.675 1046.435 6490.955 1047.435 ;
    END
  END SET_ICASN[38]
  PIN SET_ICASN[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6630.675 1046.435 6630.955 1047.435 ;
    END
  END SET_ICASN[39]
  PIN SET_ICASN[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6770.675 1046.435 6770.955 1047.435 ;
    END
  END SET_ICASN[40]
  PIN SET_ICASN[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6910.675 1046.435 6910.955 1047.435 ;
    END
  END SET_ICASN[41]
  PIN SET_ICASN[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7050.675 1046.435 7050.955 1047.435 ;
    END
  END SET_ICASN[42]
  PIN SET_ICASN[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7190.675 1046.435 7190.955 1047.435 ;
    END
  END SET_ICASN[43]
  PIN SET_ICASN[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7330.675 1046.435 7330.955 1047.435 ;
    END
  END SET_ICASN[44]
  PIN SET_ICASN[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7470.675 1046.435 7470.955 1047.435 ;
    END
  END SET_ICASN[45]
  PIN SET_ICASN[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7610.675 1046.435 7610.955 1047.435 ;
    END
  END SET_ICASN[46]
  PIN SET_ICASN[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7750.675 1046.435 7750.955 1047.435 ;
    END
  END SET_ICASN[47]
  PIN SET_ICASN[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7890.675 1046.435 7890.955 1047.435 ;
    END
  END SET_ICASN[48]
  PIN SET_ICASN[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8030.675 1046.435 8030.955 1047.435 ;
    END
  END SET_ICASN[49]
  PIN SET_ICASN[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8170.675 1046.435 8170.955 1047.435 ;
    END
  END SET_ICASN[50]
  PIN SET_ICASN[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8310.675 1046.435 8310.955 1047.435 ;
    END
  END SET_ICASN[51]
  PIN SET_ICASN[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8450.675 1046.435 8450.955 1047.435 ;
    END
  END SET_ICASN[52]
  PIN SET_ICASN[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8590.675 1046.435 8590.955 1047.435 ;
    END
  END SET_ICASN[53]
  PIN SET_ICASN[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8730.675 1046.435 8730.955 1047.435 ;
    END
  END SET_ICASN[54]
  PIN SET_ICASN[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8870.675 1046.435 8870.955 1047.435 ;
    END
  END SET_ICASN[55]
  PIN SET_ICASN[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9010.675 1046.435 9010.955 1047.435 ;
    END
  END SET_ICASN[56]
  PIN SET_ICASN[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9150.675 1046.435 9150.955 1047.435 ;
    END
  END SET_ICASN[57]
  PIN SET_ICASN[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9290.675 1046.435 9290.955 1047.435 ;
    END
  END SET_ICASN[58]
  PIN SET_ICASN[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9430.675 1046.435 9430.955 1047.435 ;
    END
  END SET_ICASN[59]
  PIN SET_ICASN[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9570.675 1046.435 9570.955 1047.435 ;
    END
  END SET_ICASN[60]
  PIN SET_ICASN[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9710.675 1046.435 9710.955 1047.435 ;
    END
  END SET_ICASN[61]
  PIN SET_ICASN[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9850.675 1046.435 9850.955 1047.435 ;
    END
  END SET_ICASN[62]
  PIN SET_ICASN[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9990.675 1046.435 9990.955 1047.435 ;
    END
  END SET_ICASN[63]
  PIN SET_ICASN[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10130.675 1046.435 10130.955 1047.435 ;
    END
  END SET_ICASN[64]
  PIN SET_ICASN[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10270.675 1046.435 10270.955 1047.435 ;
    END
  END SET_ICASN[65]
  PIN SET_ICASN[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10410.675 1046.435 10410.955 1047.435 ;
    END
  END SET_ICASN[66]
  PIN SET_ICASN[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10550.675 1046.435 10550.955 1047.435 ;
    END
  END SET_ICASN[67]
  PIN SET_ICASN[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10690.675 1046.435 10690.955 1047.435 ;
    END
  END SET_ICASN[68]
  PIN SET_ICASN[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10830.675 1046.435 10830.955 1047.435 ;
    END
  END SET_ICASN[69]
  PIN SET_ICASN[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10970.675 1046.435 10970.955 1047.435 ;
    END
  END SET_ICASN[70]
  PIN SET_ICASN[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11110.675 1046.435 11110.955 1047.435 ;
    END
  END SET_ICASN[71]
  PIN SET_ICASN[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11250.675 1046.435 11250.955 1047.435 ;
    END
  END SET_ICASN[72]
  PIN SET_ICASN[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11390.675 1046.435 11390.955 1047.435 ;
    END
  END SET_ICASN[73]
  PIN SET_ICASN[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11530.675 1046.435 11530.955 1047.435 ;
    END
  END SET_ICASN[74]
  PIN SET_ICASN[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11670.675 1046.435 11670.955 1047.435 ;
    END
  END SET_ICASN[75]
  PIN SET_ICASN[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11810.675 1046.435 11810.955 1047.435 ;
    END
  END SET_ICASN[76]
  PIN SET_ICASN[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11950.675 1046.435 11950.955 1047.435 ;
    END
  END SET_ICASN[77]
  PIN SET_ICASN[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12090.675 1046.435 12090.955 1047.435 ;
    END
  END SET_ICASN[78]
  PIN SET_ICASN[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12230.675 1046.435 12230.955 1047.435 ;
    END
  END SET_ICASN[79]
  PIN SET_ICASN[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12370.675 1046.435 12370.955 1047.435 ;
    END
  END SET_ICASN[80]
  PIN SET_ICASN[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12510.675 1046.435 12510.955 1047.435 ;
    END
  END SET_ICASN[81]
  PIN SET_ICASN[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12650.675 1046.435 12650.955 1047.435 ;
    END
  END SET_ICASN[82]
  PIN SET_ICASN[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12790.675 1046.435 12790.955 1047.435 ;
    END
  END SET_ICASN[83]
  PIN SET_ICASN[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12930.675 1046.435 12930.955 1047.435 ;
    END
  END SET_ICASN[84]
  PIN SET_ICASN[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13070.675 1046.435 13070.955 1047.435 ;
    END
  END SET_ICASN[85]
  PIN SET_ICASN[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13210.675 1046.435 13210.955 1047.435 ;
    END
  END SET_ICASN[86]
  PIN SET_ICASN[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13350.675 1046.435 13350.955 1047.435 ;
    END
  END SET_ICASN[87]
  PIN SET_ICASN[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13490.675 1046.435 13490.955 1047.435 ;
    END
  END SET_ICASN[88]
  PIN SET_ICASN[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13630.675 1046.435 13630.955 1047.435 ;
    END
  END SET_ICASN[89]
  PIN SET_ICASN[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13770.675 1046.435 13770.955 1047.435 ;
    END
  END SET_ICASN[90]
  PIN SET_ICASN[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13910.675 1046.435 13910.955 1047.435 ;
    END
  END SET_ICASN[91]
  PIN SET_ICASN[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14050.675 1046.435 14050.955 1047.435 ;
    END
  END SET_ICASN[92]
  PIN SET_ICASN[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14190.675 1046.435 14190.955 1047.435 ;
    END
  END SET_ICASN[93]
  PIN SET_ICASN[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14330.675 1046.435 14330.955 1047.435 ;
    END
  END SET_ICASN[94]
  PIN SET_ICASN[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14470.675 1046.435 14470.955 1047.435 ;
    END
  END SET_ICASN[95]
  PIN SET_ICASN[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14610.675 1046.435 14610.955 1047.435 ;
    END
  END SET_ICASN[96]
  PIN SET_ICASN[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14750.675 1046.435 14750.955 1047.435 ;
    END
  END SET_ICASN[97]
  PIN SET_ICASN[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14890.675 1046.435 14890.955 1047.435 ;
    END
  END SET_ICASN[98]
  PIN SET_ICASN[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15030.675 1046.435 15030.955 1047.435 ;
    END
  END SET_ICASN[99]
  PIN SET_ICASN[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15170.675 1046.435 15170.955 1047.435 ;
    END
  END SET_ICASN[100]
  PIN SET_ICASN[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15310.675 1046.435 15310.955 1047.435 ;
    END
  END SET_ICASN[101]
  PIN SET_ICASN[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15450.675 1046.435 15450.955 1047.435 ;
    END
  END SET_ICASN[102]
  PIN SET_ICASN[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15590.675 1046.435 15590.955 1047.435 ;
    END
  END SET_ICASN[103]
  PIN SET_ICASN[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15730.675 1046.435 15730.955 1047.435 ;
    END
  END SET_ICASN[104]
  PIN SET_ICASN[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15870.675 1046.435 15870.955 1047.435 ;
    END
  END SET_ICASN[105]
  PIN SET_ICASN[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16010.675 1046.435 16010.955 1047.435 ;
    END
  END SET_ICASN[106]
  PIN SET_ICASN[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16150.675 1046.435 16150.955 1047.435 ;
    END
  END SET_ICASN[107]
  PIN SET_ICASN[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16290.675 1046.435 16290.955 1047.435 ;
    END
  END SET_ICASN[108]
  PIN SET_ICASN[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16430.675 1046.435 16430.955 1047.435 ;
    END
  END SET_ICASN[109]
  PIN SET_ICASN[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16570.675 1046.435 16570.955 1047.435 ;
    END
  END SET_ICASN[110]
  PIN SET_ICASN[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16710.675 1046.435 16710.955 1047.435 ;
    END
  END SET_ICASN[111]
  PIN SET_ICASN[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16850.675 1046.435 16850.955 1047.435 ;
    END
  END SET_ICASN[112]
  PIN SET_ICASN[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16990.675 1046.435 16990.955 1047.435 ;
    END
  END SET_ICASN[113]
  PIN SET_ICASN[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17130.675 1046.435 17130.955 1047.435 ;
    END
  END SET_ICASN[114]
  PIN SET_ICASN[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17270.675 1046.435 17270.955 1047.435 ;
    END
  END SET_ICASN[115]
  PIN SET_ICASN[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17410.675 1046.435 17410.955 1047.435 ;
    END
  END SET_ICASN[116]
  PIN SET_ICASN[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17550.675 1046.435 17550.955 1047.435 ;
    END
  END SET_ICASN[117]
  PIN SET_ICASN[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17690.675 1046.435 17690.955 1047.435 ;
    END
  END SET_ICASN[118]
  PIN SET_ICASN[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17830.675 1046.435 17830.955 1047.435 ;
    END
  END SET_ICASN[119]
  PIN SET_ICASN[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17970.675 1046.435 17970.955 1047.435 ;
    END
  END SET_ICASN[120]
  PIN SET_ICASN[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18110.675 1046.435 18110.955 1047.435 ;
    END
  END SET_ICASN[121]
  PIN SET_ICASN[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18250.675 1046.435 18250.955 1047.435 ;
    END
  END SET_ICASN[122]
  PIN SET_ICASN[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18390.675 1046.435 18390.955 1047.435 ;
    END
  END SET_ICASN[123]
  PIN SET_ICASN[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18530.675 1046.435 18530.955 1047.435 ;
    END
  END SET_ICASN[124]
  PIN SET_ICASN[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18670.675 1046.435 18670.955 1047.435 ;
    END
  END SET_ICASN[125]
  PIN SET_ICASN[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18810.675 1046.435 18810.955 1047.435 ;
    END
  END SET_ICASN[126]
  PIN SET_VRESET_P[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15100.675 1046.435 15100.955 1047.435 ;
    END
  END SET_VRESET_P[99]
  PIN SET_VRESET_P[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15240.675 1046.435 15240.955 1047.435 ;
    END
  END SET_VRESET_P[100]
  PIN SET_VRESET_P[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15380.675 1046.435 15380.955 1047.435 ;
    END
  END SET_VRESET_P[101]
  PIN SET_VRESET_P[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15520.675 1046.435 15520.955 1047.435 ;
    END
  END SET_VRESET_P[102]
  PIN SET_VRESET_P[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15660.675 1046.435 15660.955 1047.435 ;
    END
  END SET_VRESET_P[103]
  PIN SET_VRESET_P[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15800.675 1046.435 15800.955 1047.435 ;
    END
  END SET_VRESET_P[104]
  PIN SET_VRESET_P[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15940.675 1046.435 15940.955 1047.435 ;
    END
  END SET_VRESET_P[105]
  PIN SET_VRESET_P[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16080.675 1046.435 16080.955 1047.435 ;
    END
  END SET_VRESET_P[106]
  PIN SET_VRESET_P[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16220.675 1046.435 16220.955 1047.435 ;
    END
  END SET_VRESET_P[107]
  PIN SET_VRESET_P[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16360.675 1046.435 16360.955 1047.435 ;
    END
  END SET_VRESET_P[108]
  PIN SET_VRESET_P[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16500.675 1046.435 16500.955 1047.435 ;
    END
  END SET_VRESET_P[109]
  PIN SET_VRESET_P[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16640.675 1046.435 16640.955 1047.435 ;
    END
  END SET_VRESET_P[110]
  PIN SET_VRESET_P[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16780.675 1046.435 16780.955 1047.435 ;
    END
  END SET_VRESET_P[111]
  PIN SET_VRESET_P[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16920.675 1046.435 16920.955 1047.435 ;
    END
  END SET_VRESET_P[112]
  PIN SET_VRESET_P[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17060.675 1046.435 17060.955 1047.435 ;
    END
  END SET_VRESET_P[113]
  PIN SET_VRESET_P[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17200.675 1046.435 17200.955 1047.435 ;
    END
  END SET_VRESET_P[114]
  PIN SET_VRESET_P[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17340.675 1046.435 17340.955 1047.435 ;
    END
  END SET_VRESET_P[115]
  PIN SET_VRESET_P[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17480.675 1046.435 17480.955 1047.435 ;
    END
  END SET_VRESET_P[116]
  PIN SET_VRESET_P[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17620.675 1046.435 17620.955 1047.435 ;
    END
  END SET_VRESET_P[117]
  PIN SET_VRESET_P[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17760.675 1046.435 17760.955 1047.435 ;
    END
  END SET_VRESET_P[118]
  PIN SET_VRESET_P[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17900.675 1046.435 17900.955 1047.435 ;
    END
  END SET_VRESET_P[119]
  PIN SET_VRESET_P[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18040.675 1046.435 18040.955 1047.435 ;
    END
  END SET_VRESET_P[120]
  PIN SET_VRESET_P[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18180.675 1046.435 18180.955 1047.435 ;
    END
  END SET_VRESET_P[121]
  PIN SET_VRESET_P[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18320.675 1046.435 18320.955 1047.435 ;
    END
  END SET_VRESET_P[122]
  PIN SET_VRESET_P[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18460.675 1046.435 18460.955 1047.435 ;
    END
  END SET_VRESET_P[123]
  PIN SET_VRESET_P[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18600.675 1046.435 18600.955 1047.435 ;
    END
  END SET_VRESET_P[124]
  PIN SET_VRESET_P[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18740.675 1046.435 18740.955 1047.435 ;
    END
  END SET_VRESET_P[125]
  PIN SET_VRESET_P[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18880.675 1046.435 18880.955 1047.435 ;
    END
  END SET_VRESET_P[126]
  PIN SET_VRESET_P[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19020.675 1046.435 19020.955 1047.435 ;
    END
  END SET_VRESET_P[127]
  PIN SET_VCLIP[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1244.315 1046.435 1244.595 1047.435 ;
    END
  END SET_VCLIP[0]
  PIN SET_VCLIP[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1384.315 1046.435 1384.595 1047.435 ;
    END
  END SET_VCLIP[1]
  PIN SET_VCLIP[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1524.315 1046.435 1524.595 1047.435 ;
    END
  END SET_VCLIP[2]
  PIN SET_VCLIP[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1664.315 1046.435 1664.595 1047.435 ;
    END
  END SET_VCLIP[3]
  PIN SET_VCLIP[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1804.315 1046.435 1804.595 1047.435 ;
    END
  END SET_VCLIP[4]
  PIN SET_VCLIP[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1944.315 1046.435 1944.595 1047.435 ;
    END
  END SET_VCLIP[5]
  PIN SET_VCLIP[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2084.315 1046.435 2084.595 1047.435 ;
    END
  END SET_VCLIP[6]
  PIN SET_VCLIP[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2224.315 1046.435 2224.595 1047.435 ;
    END
  END SET_VCLIP[7]
  PIN SET_VCLIP[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2364.315 1046.435 2364.595 1047.435 ;
    END
  END SET_VCLIP[8]
  PIN SET_VCLIP[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2504.315 1046.435 2504.595 1047.435 ;
    END
  END SET_VCLIP[9]
  PIN SET_VCLIP[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2644.315 1046.435 2644.595 1047.435 ;
    END
  END SET_VCLIP[10]
  PIN SET_VCLIP[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2784.315 1046.435 2784.595 1047.435 ;
    END
  END SET_VCLIP[11]
  PIN SET_VCLIP[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2924.315 1046.435 2924.595 1047.435 ;
    END
  END SET_VCLIP[12]
  PIN SET_VCLIP[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3064.315 1046.435 3064.595 1047.435 ;
    END
  END SET_VCLIP[13]
  PIN SET_VCLIP[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3204.315 1046.435 3204.595 1047.435 ;
    END
  END SET_VCLIP[14]
  PIN SET_VCLIP[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3344.315 1046.435 3344.595 1047.435 ;
    END
  END SET_VCLIP[15]
  PIN SET_VCLIP[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3484.315 1046.435 3484.595 1047.435 ;
    END
  END SET_VCLIP[16]
  PIN SET_VCLIP[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3624.315 1046.435 3624.595 1047.435 ;
    END
  END SET_VCLIP[17]
  PIN SET_VCLIP[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3764.315 1046.435 3764.595 1047.435 ;
    END
  END SET_VCLIP[18]
  PIN SET_VCLIP[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3904.315 1046.435 3904.595 1047.435 ;
    END
  END SET_VCLIP[19]
  PIN SET_VCLIP[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4044.315 1046.435 4044.595 1047.435 ;
    END
  END SET_VCLIP[20]
  PIN SET_VCLIP[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4184.315 1046.435 4184.595 1047.435 ;
    END
  END SET_VCLIP[21]
  PIN SET_VCLIP[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4324.315 1046.435 4324.595 1047.435 ;
    END
  END SET_VCLIP[22]
  PIN SET_VCLIP[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4464.315 1046.435 4464.595 1047.435 ;
    END
  END SET_VCLIP[23]
  PIN SET_VCLIP[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4604.315 1046.435 4604.595 1047.435 ;
    END
  END SET_VCLIP[24]
  PIN SET_VCLIP[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4744.315 1046.435 4744.595 1047.435 ;
    END
  END SET_VCLIP[25]
  PIN SET_VCLIP[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4884.315 1046.435 4884.595 1047.435 ;
    END
  END SET_VCLIP[26]
  PIN SET_VCLIP[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5024.315 1046.435 5024.595 1047.435 ;
    END
  END SET_VCLIP[27]
  PIN SET_VCLIP[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5164.315 1046.435 5164.595 1047.435 ;
    END
  END SET_VCLIP[28]
  PIN SET_VCLIP[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5304.315 1046.435 5304.595 1047.435 ;
    END
  END SET_VCLIP[29]
  PIN SET_VCLIP[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5444.315 1046.435 5444.595 1047.435 ;
    END
  END SET_VCLIP[30]
  PIN SET_VCLIP[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5584.315 1046.435 5584.595 1047.435 ;
    END
  END SET_VCLIP[31]
  PIN SET_VCLIP[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5724.315 1046.435 5724.595 1047.435 ;
    END
  END SET_VCLIP[32]
  PIN SET_VCLIP[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5864.315 1046.435 5864.595 1047.435 ;
    END
  END SET_VCLIP[33]
  PIN SET_VCLIP[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6004.315 1046.435 6004.595 1047.435 ;
    END
  END SET_VCLIP[34]
  PIN SET_VCLIP[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6144.315 1046.435 6144.595 1047.435 ;
    END
  END SET_VCLIP[35]
  PIN SET_VCLIP[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6284.315 1046.435 6284.595 1047.435 ;
    END
  END SET_VCLIP[36]
  PIN SET_VCLIP[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6424.315 1046.435 6424.595 1047.435 ;
    END
  END SET_VCLIP[37]
  PIN SET_VCLIP[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6564.315 1046.435 6564.595 1047.435 ;
    END
  END SET_VCLIP[38]
  PIN SET_VCLIP[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6704.315 1046.435 6704.595 1047.435 ;
    END
  END SET_VCLIP[39]
  PIN SET_VCLIP[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6844.315 1046.435 6844.595 1047.435 ;
    END
  END SET_VCLIP[40]
  PIN SET_VCLIP[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6984.315 1046.435 6984.595 1047.435 ;
    END
  END SET_VCLIP[41]
  PIN SET_VCLIP[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7124.315 1046.435 7124.595 1047.435 ;
    END
  END SET_VCLIP[42]
  PIN SET_VCLIP[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7264.315 1046.435 7264.595 1047.435 ;
    END
  END SET_VCLIP[43]
  PIN SET_VCLIP[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7404.315 1046.435 7404.595 1047.435 ;
    END
  END SET_VCLIP[44]
  PIN SET_VCLIP[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7544.315 1046.435 7544.595 1047.435 ;
    END
  END SET_VCLIP[45]
  PIN SET_VCLIP[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7684.315 1046.435 7684.595 1047.435 ;
    END
  END SET_VCLIP[46]
  PIN SET_VCLIP[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7824.315 1046.435 7824.595 1047.435 ;
    END
  END SET_VCLIP[47]
  PIN SET_VCLIP[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7964.315 1046.435 7964.595 1047.435 ;
    END
  END SET_VCLIP[48]
  PIN SET_VCLIP[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8104.315 1046.435 8104.595 1047.435 ;
    END
  END SET_VCLIP[49]
  PIN SET_VCLIP[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8244.315 1046.435 8244.595 1047.435 ;
    END
  END SET_VCLIP[50]
  PIN SET_VCLIP[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8384.315 1046.435 8384.595 1047.435 ;
    END
  END SET_VCLIP[51]
  PIN SET_VCLIP[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8524.315 1046.435 8524.595 1047.435 ;
    END
  END SET_VCLIP[52]
  PIN SET_VCLIP[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8664.315 1046.435 8664.595 1047.435 ;
    END
  END SET_VCLIP[53]
  PIN SET_VCLIP[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8804.315 1046.435 8804.595 1047.435 ;
    END
  END SET_VCLIP[54]
  PIN SET_VCLIP[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8944.315 1046.435 8944.595 1047.435 ;
    END
  END SET_VCLIP[55]
  PIN SET_VCLIP[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9084.315 1046.435 9084.595 1047.435 ;
    END
  END SET_VCLIP[56]
  PIN SET_VCLIP[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9224.315 1046.435 9224.595 1047.435 ;
    END
  END SET_VCLIP[57]
  PIN SET_VCLIP[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9364.315 1046.435 9364.595 1047.435 ;
    END
  END SET_VCLIP[58]
  PIN SET_VCLIP[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9504.315 1046.435 9504.595 1047.435 ;
    END
  END SET_VCLIP[59]
  PIN SET_VCLIP[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9644.315 1046.435 9644.595 1047.435 ;
    END
  END SET_VCLIP[60]
  PIN SET_VCLIP[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9784.315 1046.435 9784.595 1047.435 ;
    END
  END SET_VCLIP[61]
  PIN SET_VCLIP[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9924.315 1046.435 9924.595 1047.435 ;
    END
  END SET_VCLIP[62]
  PIN SET_VCLIP[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10064.315 1046.435 10064.595 1047.435 ;
    END
  END SET_VCLIP[63]
  PIN SET_VCLIP[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10204.315 1046.435 10204.595 1047.435 ;
    END
  END SET_VCLIP[64]
  PIN SET_VCLIP[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10344.315 1046.435 10344.595 1047.435 ;
    END
  END SET_VCLIP[65]
  PIN SET_VCLIP[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10484.315 1046.435 10484.595 1047.435 ;
    END
  END SET_VCLIP[66]
  PIN SET_VCLIP[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10624.315 1046.435 10624.595 1047.435 ;
    END
  END SET_VCLIP[67]
  PIN SET_VCLIP[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10764.315 1046.435 10764.595 1047.435 ;
    END
  END SET_VCLIP[68]
  PIN SET_VCLIP[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10904.315 1046.435 10904.595 1047.435 ;
    END
  END SET_VCLIP[69]
  PIN SET_VCLIP[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11044.315 1046.435 11044.595 1047.435 ;
    END
  END SET_VCLIP[70]
  PIN SET_VCLIP[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11184.315 1046.435 11184.595 1047.435 ;
    END
  END SET_VCLIP[71]
  PIN SET_VCLIP[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11324.315 1046.435 11324.595 1047.435 ;
    END
  END SET_VCLIP[72]
  PIN nRST[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10808.905 1046.435 10809.185 1047.435 ;
    END
  END nRST[121]
  PIN nRST[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10248.905 1046.435 10249.185 1047.435 ;
    END
  END nRST[114]
  PIN nRST[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5208.905 1046.435 5209.185 1047.435 ;
    END
  END nRST[51]
  PIN nRST[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4648.905 1046.435 4649.185 1047.435 ;
    END
  END nRST[44]
  PIN nRST[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10738.905 1046.435 10739.185 1047.435 ;
    END
  END nRST[120]
  PIN nRST[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10178.905 1046.435 10179.185 1047.435 ;
    END
  END nRST[113]
  PIN nRST[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9618.905 1046.435 9619.185 1047.435 ;
    END
  END nRST[106]
  PIN nRST[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1288.905 1046.435 1289.185 1047.435 ;
    END
  END nRST[2]
  PIN nRST[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4088.905 1046.435 4089.185 1047.435 ;
    END
  END nRST[37]
  PIN nRST[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3528.905 1046.435 3529.185 1047.435 ;
    END
  END nRST[30]
  PIN Data_COMP[341]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11438.345 1046.435 11438.625 1047.435 ;
    END
  END Data_COMP[341]
  PIN Data_COMP[342]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11435.545 1046.435 11435.825 1047.435 ;
    END
  END Data_COMP[342]
  PIN INJ_IN[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11434.425 1046.435 11434.705 1047.435 ;
    END
  END INJ_IN[257]
  PIN BcidMtx[772]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11392.425 1046.435 11392.705 1047.435 ;
    END
  END BcidMtx[772]
  PIN Read_COMP[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11390.745 1046.435 11391.025 1047.435 ;
    END
  END Read_COMP[16]
  PIN BcidMtx[769]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11389.625 1046.435 11389.905 1047.435 ;
    END
  END BcidMtx[769]
  PIN INJ_IN[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11387.945 1046.435 11388.225 1047.435 ;
    END
  END INJ_IN[256]
  PIN Data_COMP[346]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11384.585 1046.435 11384.865 1047.435 ;
    END
  END Data_COMP[346]
  PIN Data_COMP[340]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11384.025 1046.435 11384.305 1047.435 ;
    END
  END Data_COMP[340]
  PIN Data_COMP[337]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11382.345 1046.435 11382.625 1047.435 ;
    END
  END Data_COMP[337]
  PIN MASKD[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11371.145 1046.435 11371.425 1047.435 ;
    END
  END MASKD[256]
  PIN DIG_MON_COMP[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11370.025 1046.435 11370.305 1047.435 ;
    END
  END DIG_MON_COMP[32]
  PIN DIG_MON_SEL[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11367.785 1046.435 11368.065 1047.435 ;
    END
  END DIG_MON_SEL[255]
  PIN Data_COMP[333]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11361.345 1046.435 11361.625 1047.435 ;
    END
  END Data_COMP[333]
  PIN Data_COMP[323]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11360.785 1046.435 11361.065 1047.435 ;
    END
  END Data_COMP[323]
  PIN Data_COMP[320]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11359.105 1046.435 11359.385 1047.435 ;
    END
  END Data_COMP[320]
  PIN Data_COMP[321]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11330.825 1046.435 11331.105 1047.435 ;
    END
  END Data_COMP[321]
  PIN INJ_IN[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11329.705 1046.435 11329.985 1047.435 ;
    END
  END INJ_IN[255]
  PIN BcidMtx[766]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11326.905 1046.435 11327.185 1047.435 ;
    END
  END BcidMtx[766]
  PIN BcidMtx[763]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11324.105 1046.435 11324.385 1047.435 ;
    END
  END BcidMtx[763]
  PIN BcidMtx[762]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11323.545 1046.435 11323.825 1047.435 ;
    END
  END BcidMtx[762]
  PIN Data_COMP[318]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11321.305 1046.435 11321.585 1047.435 ;
    END
  END Data_COMP[318]
  PIN Data_COMP[319]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11305.625 1046.435 11305.905 1047.435 ;
    END
  END Data_COMP[319]
  PIN Data_COMP[331]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11305.065 1046.435 11305.345 1047.435 ;
    END
  END Data_COMP[331]
  PIN Data_COMP[315]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11303.385 1046.435 11303.665 1047.435 ;
    END
  END Data_COMP[315]
  PIN MASKH[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11301.705 1046.435 11301.985 1047.435 ;
    END
  END MASKH[127]
  PIN MASKD[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11296.665 1046.435 11296.945 1047.435 ;
    END
  END MASKD[253]
  PIN MASKV[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11293.865 1046.435 11294.145 1047.435 ;
    END
  END MASKV[253]
  PIN Data_COMP[306]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11252.425 1046.435 11252.705 1047.435 ;
    END
  END Data_COMP[306]
  PIN Data_COMP[307]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11250.745 1046.435 11251.025 1047.435 ;
    END
  END Data_COMP[307]
  PIN Data_COMP[301]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11249.065 1046.435 11249.345 1047.435 ;
    END
  END Data_COMP[301]
  PIN nTOK_COMP[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11246.265 1046.435 11246.545 1047.435 ;
    END
  END nTOK_COMP[14]
  PIN BcidMtx[759]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11244.025 1046.435 11244.305 1047.435 ;
    END
  END BcidMtx[759]
  PIN BcidMtx[758]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11242.345 1046.435 11242.625 1047.435 ;
    END
  END BcidMtx[758]
  PIN BcidMtx[756]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11241.225 1046.435 11241.505 1047.435 ;
    END
  END BcidMtx[756]
  PIN Data_COMP[296]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11230.025 1046.435 11230.305 1047.435 ;
    END
  END Data_COMP[296]
  PIN Data_COMP[304]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11228.345 1046.435 11228.625 1047.435 ;
    END
  END Data_COMP[304]
  PIN Data_COMP[305]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11226.665 1046.435 11226.945 1047.435 ;
    END
  END Data_COMP[305]
  PIN Data_COMP[311]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11224.985 1046.435 11225.265 1047.435 ;
    END
  END Data_COMP[311]
  PIN MASKD[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11221.345 1046.435 11221.625 1047.435 ;
    END
  END MASKD[252]
  PIN DIG_MON_SEL[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11218.545 1046.435 11218.825 1047.435 ;
    END
  END DIG_MON_SEL[252]
  PIN MASKD[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12310.825 1046.435 12311.105 1047.435 ;
    END
  END MASKD[279]
  PIN MASKV[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12308.025 1046.435 12308.305 1047.435 ;
    END
  END MASKV[279]
  PIN Data_COMP[579]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12306.345 1046.435 12306.625 1047.435 ;
    END
  END Data_COMP[579]
  PIN Data_COMP[580]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12304.665 1046.435 12304.945 1047.435 ;
    END
  END Data_COMP[580]
  PIN Data_COMP[574]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12302.985 1046.435 12303.265 1047.435 ;
    END
  END Data_COMP[574]
  PIN nTOK_COMP[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12300.185 1046.435 12300.465 1047.435 ;
    END
  END nTOK_COMP[27]
  PIN BcidMtx[837]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12284.505 1046.435 12284.785 1047.435 ;
    END
  END BcidMtx[837]
  PIN BcidMtx[836]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12282.825 1046.435 12283.105 1047.435 ;
    END
  END BcidMtx[836]
  PIN Read_HV[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18752.505 1046.435 18752.785 1047.435 ;
    END
  END Read_HV[52]
  PIN Data_COMP[570]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12279.465 1046.435 12279.745 1047.435 ;
    END
  END Data_COMP[570]
  PIN Data_COMP[582]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12277.785 1046.435 12278.065 1047.435 ;
    END
  END Data_COMP[582]
  PIN Data_COMP[578]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12275.545 1046.435 12275.825 1047.435 ;
    END
  END Data_COMP[578]
  PIN Data_COMP[567]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12274.425 1046.435 12274.705 1047.435 ;
    END
  END Data_COMP[567]
  PIN MASKH[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12234.105 1046.435 12234.385 1047.435 ;
    END
  END MASKH[139]
  PIN DIG_MON_SEL[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12230.745 1046.435 12231.025 1047.435 ;
    END
  END DIG_MON_SEL[278]
  PIN DIG_MON_COMP[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12227.945 1046.435 12228.225 1047.435 ;
    END
  END DIG_MON_COMP[53]
  PIN Data_COMP[564]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12225.705 1046.435 12225.985 1047.435 ;
    END
  END Data_COMP[564]
  PIN Data_COMP[558]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12224.585 1046.435 12224.865 1047.435 ;
    END
  END Data_COMP[558]
  PIN Data_COMP[566]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12222.345 1046.435 12222.625 1047.435 ;
    END
  END Data_COMP[566]
  PIN Data_COMP[552]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12212.265 1046.435 12212.545 1047.435 ;
    END
  END Data_COMP[552]
  PIN nTOK_COMP[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12210.025 1046.435 12210.305 1047.435 ;
    END
  END nTOK_COMP[26]
  PIN FREEZE_COMP[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12207.225 1046.435 12207.505 1047.435 ;
    END
  END FREEZE_COMP[26]
  PIN BcidMtx[829]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12205.545 1046.435 12205.825 1047.435 ;
    END
  END BcidMtx[829]
  PIN INJ_IN[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12201.905 1046.435 12202.185 1047.435 ;
    END
  END INJ_IN[276]
  PIN Data_COMP[561]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12199.105 1046.435 12199.385 1047.435 ;
    END
  END Data_COMP[561]
  PIN Data_COMP[562]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12171.945 1046.435 12172.225 1047.435 ;
    END
  END Data_COMP[562]
  PIN Data_COMP[547]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12170.825 1046.435 12171.105 1047.435 ;
    END
  END Data_COMP[547]
  PIN MASKH[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12168.585 1046.435 12168.865 1047.435 ;
    END
  END MASKH[138]
  PIN DIG_MON_SEL[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12164.665 1046.435 12164.945 1047.435 ;
    END
  END DIG_MON_SEL[275]
  PIN MASKV[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12160.745 1046.435 12161.025 1047.435 ;
    END
  END MASKV[275]
  PIN Data_COMP[537]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12146.185 1046.435 12146.465 1047.435 ;
    END
  END Data_COMP[537]
  PIN Data_COMP[530]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12145.065 1046.435 12145.345 1047.435 ;
    END
  END Data_COMP[530]
  PIN Data_COMP[545]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12143.945 1046.435 12144.225 1047.435 ;
    END
  END Data_COMP[545]
  PIN nTOK_COMP[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12140.025 1046.435 12140.305 1047.435 ;
    END
  END nTOK_COMP[25]
  PIN BcidMtx[825]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12137.785 1046.435 12138.065 1047.435 ;
    END
  END BcidMtx[825]
  PIN BcidMtx[824]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12136.105 1046.435 12136.385 1047.435 ;
    END
  END BcidMtx[824]
  PIN Data_COMP[528]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12094.105 1046.435 12094.385 1047.435 ;
    END
  END Data_COMP[528]
  PIN Data_COMP[534]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12092.985 1046.435 12093.265 1047.435 ;
    END
  END Data_COMP[534]
  PIN Data_COMP[529]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12091.305 1046.435 12091.585 1047.435 ;
    END
  END Data_COMP[529]
  PIN Data_COMP[525]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12089.065 1046.435 12089.345 1047.435 ;
    END
  END Data_COMP[525]
  PIN MASKV[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12087.945 1046.435 12088.225 1047.435 ;
    END
  END MASKV[274]
  PIN DIG_MON_COMP[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12085.705 1046.435 12085.985 1047.435 ;
    END
  END DIG_MON_COMP[50]
  PIN MASKD[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12082.345 1046.435 12082.625 1047.435 ;
    END
  END MASKD[273]
  PIN INJ_ROW[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12071.705 1046.435 12071.985 1047.435 ;
    END
  END INJ_ROW[136]
  PIN Data_COMP[512]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12070.025 1046.435 12070.305 1047.435 ;
    END
  END Data_COMP[512]
  PIN Data_COMP[517]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12067.785 1046.435 12068.065 1047.435 ;
    END
  END Data_COMP[517]
  PIN Data_COMP[518]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12066.665 1046.435 12066.945 1047.435 ;
    END
  END Data_COMP[518]
  PIN Data_COMP[510]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12065.545 1046.435 12065.825 1047.435 ;
    END
  END Data_COMP[510]
  PIN BcidMtx[820]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12059.665 1046.435 12059.945 1047.435 ;
    END
  END BcidMtx[820]
  PIN Read_COMP[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12032.505 1046.435 12032.785 1047.435 ;
    END
  END Read_COMP[24]
  PIN BcidMtx[816]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12030.825 1046.435 12031.105 1047.435 ;
    END
  END BcidMtx[816]
  PIN Data_COMP[506]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12028.025 1046.435 12028.305 1047.435 ;
    END
  END Data_COMP[506]
  PIN Data_COMP[514]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12026.345 1046.435 12026.625 1047.435 ;
    END
  END Data_COMP[514]
  PIN Data_COMP[515]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12024.665 1046.435 12024.945 1047.435 ;
    END
  END Data_COMP[515]
  PIN Data_COMP[521]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12022.985 1046.435 12023.265 1047.435 ;
    END
  END Data_COMP[521]
  PIN MASKH[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12021.865 1046.435 12022.145 1047.435 ;
    END
  END MASKH[136]
  PIN DIG_MON_COMP[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12020.185 1046.435 12020.465 1047.435 ;
    END
  END DIG_MON_COMP[48]
  PIN DIG_MON_SEL[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12005.065 1046.435 12005.345 1047.435 ;
    END
  END DIG_MON_SEL[271]
  PIN MASKV[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12001.145 1046.435 12001.425 1047.435 ;
    END
  END MASKV[271]
  PIN Data_COMP[491]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12000.025 1046.435 12000.305 1047.435 ;
    END
  END Data_COMP[491]
  PIN Data_COMP[488]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11998.345 1046.435 11998.625 1047.435 ;
    END
  END Data_COMP[488]
  PIN Data_COMP[490]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11996.105 1046.435 11996.385 1047.435 ;
    END
  END Data_COMP[490]
  PIN INJ_IN[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11994.425 1046.435 11994.705 1047.435 ;
    END
  END INJ_IN[271]
  PIN BcidMtx[815]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11952.985 1046.435 11953.265 1047.435 ;
    END
  END BcidMtx[815]
  PIN Read_COMP[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11950.745 1046.435 11951.025 1047.435 ;
    END
  END Read_COMP[23]
  PIN BcidMtx[811]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11949.625 1046.435 11949.905 1047.435 ;
    END
  END BcidMtx[811]
  PIN Data_COMP[486]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11946.825 1046.435 11947.105 1047.435 ;
    END
  END Data_COMP[486]
  PIN Data_COMP[493]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11944.585 1046.435 11944.865 1047.435 ;
    END
  END Data_COMP[493]
  PIN Data_COMP[499]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11943.465 1046.435 11943.745 1047.435 ;
    END
  END Data_COMP[499]
  PIN Data_COMP[483]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11941.785 1046.435 11942.065 1047.435 ;
    END
  END Data_COMP[483]
  PIN MASKD[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11931.145 1046.435 11931.425 1047.435 ;
    END
  END MASKD[270]
  PIN MASKD[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11926.665 1046.435 11926.945 1047.435 ;
    END
  END MASKD[269]
  PIN Data_COMP[480]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11921.345 1046.435 11921.625 1047.435 ;
    END
  END Data_COMP[480]
  PIN Data_COMP[481]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11919.665 1046.435 11919.945 1047.435 ;
    END
  END Data_COMP[481]
  PIN Data_COMP[475]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11893.065 1046.435 11893.345 1047.435 ;
    END
  END Data_COMP[475]
  PIN Data_COMP[469]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11891.385 1046.435 11891.665 1047.435 ;
    END
  END Data_COMP[469]
  PIN INJ_IN[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11889.705 1046.435 11889.985 1047.435 ;
    END
  END INJ_IN[269]
  PIN FREEZE_COMP[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11885.785 1046.435 11886.065 1047.435 ;
    END
  END FREEZE_COMP[22]
  PIN Read_COMP[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11885.225 1046.435 11885.505 1047.435 ;
    END
  END Read_COMP[22]
  PIN INJ_IN[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11882.425 1046.435 11882.705 1047.435 ;
    END
  END INJ_IN[268]
  PIN Data_COMP[471]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11880.185 1046.435 11880.465 1047.435 ;
    END
  END Data_COMP[471]
  PIN Data_COMP[472]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11866.185 1046.435 11866.465 1047.435 ;
    END
  END Data_COMP[472]
  PIN Data_COMP[463]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11863.945 1046.435 11864.225 1047.435 ;
    END
  END Data_COMP[463]
  PIN MASKV[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11862.265 1046.435 11862.545 1047.435 ;
    END
  END MASKV[268]
  PIN MASKD[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11861.145 1046.435 11861.425 1047.435 ;
    END
  END MASKD[268]
  PIN DIG_MON_SEL[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11857.785 1046.435 11858.065 1047.435 ;
    END
  END DIG_MON_SEL[267]
  PIN INJ_ROW[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11854.425 1046.435 11854.705 1047.435 ;
    END
  END INJ_ROW[133]
  PIN Data_COMP[459]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11813.545 1046.435 11813.825 1047.435 ;
    END
  END Data_COMP[459]
  PIN Data_COMP[454]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11810.745 1046.435 11811.025 1047.435 ;
    END
  END Data_COMP[454]
  PIN Data_COMP[448]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11809.065 1046.435 11809.345 1047.435 ;
    END
  END Data_COMP[448]
  PIN Data_COMP[447]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11808.505 1046.435 11808.785 1047.435 ;
    END
  END Data_COMP[447]
  PIN BcidMtx[801]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11804.025 1046.435 11804.305 1047.435 ;
    END
  END BcidMtx[801]
  PIN Read_COMP[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11802.905 1046.435 11803.185 1047.435 ;
    END
  END Read_COMP[21]
  PIN BcidMtx[798]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11801.225 1046.435 11801.505 1047.435 ;
    END
  END BcidMtx[798]
  PIN Data_COMP[450]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11789.465 1046.435 11789.745 1047.435 ;
    END
  END Data_COMP[450]
  PIN Data_COMP[445]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11787.785 1046.435 11788.065 1047.435 ;
    END
  END Data_COMP[445]
  PIN Data_COMP[452]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11786.665 1046.435 11786.945 1047.435 ;
    END
  END Data_COMP[452]
  PIN MASKV[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11782.465 1046.435 11782.745 1047.435 ;
    END
  END MASKV[266]
  PIN MASKD[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11781.345 1046.435 11781.625 1047.435 ;
    END
  END MASKD[266]
  PIN DIG_MON_SEL[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11778.545 1046.435 11778.825 1047.435 ;
    END
  END DIG_MON_SEL[266]
  PIN INJ_ROW[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12868.585 1046.435 12868.865 1047.435 ;
    END
  END INJ_ROW[146]
  PIN MASKV[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12868.025 1046.435 12868.305 1047.435 ;
    END
  END MASKV[293]
  PIN Data_COMP[726]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12866.345 1046.435 12866.625 1047.435 ;
    END
  END Data_COMP[726]
  PIN Data_COMP[728]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12863.545 1046.435 12863.825 1047.435 ;
    END
  END Data_COMP[728]
  PIN Data_COMP[720]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12862.425 1046.435 12862.705 1047.435 ;
    END
  END Data_COMP[720]
  PIN nTOK_COMP[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12860.185 1046.435 12860.465 1047.435 ;
    END
  END nTOK_COMP[34]
  PIN FREEZE_COMP[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12843.945 1046.435 12844.225 1047.435 ;
    END
  END FREEZE_COMP[34]
  PIN BcidMtx[877]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12842.265 1046.435 12842.545 1047.435 ;
    END
  END BcidMtx[877]
  PIN BcidMtx[876]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12841.705 1046.435 12841.985 1047.435 ;
    END
  END BcidMtx[876]
  PIN Data_COMP[729]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12837.785 1046.435 12838.065 1047.435 ;
    END
  END Data_COMP[729]
  PIN Data_COMP[730]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12836.105 1046.435 12836.385 1047.435 ;
    END
  END Data_COMP[730]
  PIN Data_COMP[715]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12834.985 1046.435 12835.265 1047.435 ;
    END
  END Data_COMP[715]
  PIN MASKH[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12794.105 1046.435 12794.385 1047.435 ;
    END
  END MASKH[146]
  PIN DIG_MON_SEL[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12790.185 1046.435 12790.465 1047.435 ;
    END
  END DIG_MON_SEL[291]
  PIN Data_COMP[711]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12785.705 1046.435 12785.985 1047.435 ;
    END
  END Data_COMP[711]
  PIN Data_COMP[705]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12784.585 1046.435 12784.865 1047.435 ;
    END
  END Data_COMP[705]
  PIN Data_COMP[698]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12783.465 1046.435 12783.745 1047.435 ;
    END
  END Data_COMP[698]
  PIN Data_COMP[700]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12781.225 1046.435 12781.505 1047.435 ;
    END
  END Data_COMP[700]
  PIN nTOK_COMP[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12770.025 1046.435 12770.305 1047.435 ;
    END
  END nTOK_COMP[33]
  PIN BcidMtx[874]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12768.345 1046.435 12768.625 1047.435 ;
    END
  END BcidMtx[874]
  PIN BcidMtx[871]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12765.545 1046.435 12765.825 1047.435 ;
    END
  END BcidMtx[871]
  PIN INJ_IN[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12761.905 1046.435 12762.185 1047.435 ;
    END
  END INJ_IN[290]
  PIN Data_COMP[702]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12759.665 1046.435 12759.945 1047.435 ;
    END
  END Data_COMP[702]
  PIN Data_COMP[709]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12731.945 1046.435 12732.225 1047.435 ;
    END
  END Data_COMP[709]
  PIN Data_COMP[704]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12731.385 1046.435 12731.665 1047.435 ;
    END
  END Data_COMP[704]
  PIN Data_COMP[710]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12729.705 1046.435 12729.985 1047.435 ;
    END
  END Data_COMP[710]
  PIN MASKD[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12728.025 1046.435 12728.305 1047.435 ;
    END
  END MASKD[290]
  PIN DIG_MON_SEL[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12725.225 1046.435 12725.505 1047.435 ;
    END
  END DIG_MON_SEL[290]
  PIN DIG_MON_COMP[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12722.425 1046.435 12722.705 1047.435 ;
    END
  END DIG_MON_COMP[65]
  PIN Data_COMP[690]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12720.185 1046.435 12720.465 1047.435 ;
    END
  END Data_COMP[690]
  PIN Data_COMP[691]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12705.625 1046.435 12705.905 1047.435 ;
    END
  END Data_COMP[691]
  PIN Data_COMP[692]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12703.945 1046.435 12704.225 1047.435 ;
    END
  END Data_COMP[692]
  PIN INJ_IN[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12701.145 1046.435 12701.425 1047.435 ;
    END
  END INJ_IN[289]
  PIN BcidMtx[869]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12698.905 1046.435 12699.185 1047.435 ;
    END
  END BcidMtx[869]
  PIN FREEZE_COMP[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12697.225 1046.435 12697.505 1047.435 ;
    END
  END FREEZE_COMP[32]
  PIN BcidMtx[864]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12694.985 1046.435 12695.265 1047.435 ;
    END
  END BcidMtx[864]
  PIN Data_COMP[675]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12654.105 1046.435 12654.385 1047.435 ;
    END
  END Data_COMP[675]
  PIN Data_COMP[687]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12652.425 1046.435 12652.705 1047.435 ;
    END
  END Data_COMP[687]
  PIN Data_COMP[688]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12650.745 1046.435 12651.025 1047.435 ;
    END
  END Data_COMP[688]
  PIN Data_COMP[672]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12649.065 1046.435 12649.345 1047.435 ;
    END
  END Data_COMP[672]
  PIN MASKH[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12647.385 1046.435 12647.665 1047.435 ;
    END
  END MASKH[144]
  PIN MASKD[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12642.345 1046.435 12642.625 1047.435 ;
    END
  END MASKD[287]
  PIN MASKV[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12631.145 1046.435 12631.425 1047.435 ;
    END
  END MASKV[287]
  PIN Data_COMP[663]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12629.465 1046.435 12629.745 1047.435 ;
    END
  END Data_COMP[663]
  PIN Data_COMP[656]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12628.345 1046.435 12628.625 1047.435 ;
    END
  END Data_COMP[656]
  PIN Data_COMP[665]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12626.665 1046.435 12626.945 1047.435 ;
    END
  END Data_COMP[665]
  PIN nTOK_COMP[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12621.345 1046.435 12621.625 1047.435 ;
    END
  END nTOK_COMP[31]
  PIN BcidMtx[862]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12619.665 1046.435 12619.945 1047.435 ;
    END
  END BcidMtx[862]
  PIN BcidMtx[860]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12591.945 1046.435 12592.225 1047.435 ;
    END
  END BcidMtx[860]
  PIN INJ_IN[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12589.705 1046.435 12589.985 1047.435 ;
    END
  END INJ_IN[286]
  PIN Data_COMP[660]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12587.465 1046.435 12587.745 1047.435 ;
    END
  END Data_COMP[660]
  PIN Data_COMP[655]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12585.785 1046.435 12586.065 1047.435 ;
    END
  END Data_COMP[655]
  PIN Data_COMP[652]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12584.105 1046.435 12584.385 1047.435 ;
    END
  END Data_COMP[652]
  PIN MASKV[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12582.425 1046.435 12582.705 1047.435 ;
    END
  END MASKV[286]
  PIN DIG_MON_COMP[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12580.185 1046.435 12580.465 1047.435 ;
    END
  END DIG_MON_COMP[62]
  PIN DIG_MON_SEL[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12565.065 1046.435 12565.345 1047.435 ;
    END
  END DIG_MON_SEL[285]
  PIN INJ_ROW[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12561.705 1046.435 12561.985 1047.435 ;
    END
  END INJ_ROW[142]
  PIN Data_COMP[638]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12560.025 1046.435 12560.305 1047.435 ;
    END
  END Data_COMP[638]
  PIN nRST[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2968.905 1046.435 2969.185 1047.435 ;
    END
  END nRST[23]
  PIN nRST[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 2408.905 1046.435 2409.185 1047.435 ;
    END
  END nRST[16]
  PIN nRST[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1848.905 1046.435 1849.185 1047.435 ;
    END
  END nRST[9]
  PIN Data_PMOS_NOSF[1020]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5026.345 1046.435 5026.625 1047.435 ;
    END
  END Data_PMOS_NOSF[1020]
  PIN Data_HV[1125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18866.185 1046.435 18866.465 1047.435 ;
    END
  END Data_HV[1125]
  PIN Data_PMOS_NOSF[1022]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5023.545 1046.435 5023.825 1047.435 ;
    END
  END Data_PMOS_NOSF[1022]
  PIN INJ_IN[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5021.305 1046.435 5021.585 1047.435 ;
    END
  END INJ_IN[97]
  PIN nTOK_PMOS_NOSF[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5020.185 1046.435 5020.465 1047.435 ;
    END
  END nTOK_PMOS_NOSF[48]
  PIN BcidMtx[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5004.505 1046.435 5004.785 1047.435 ;
    END
  END BcidMtx[291]
  PIN BcidMtx[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5002.825 1046.435 5003.105 1047.435 ;
    END
  END BcidMtx[290]
  PIN INJ_IN[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5000.585 1046.435 5000.865 1047.435 ;
    END
  END INJ_IN[96]
  PIN Data_PMOS_NOSF[1017]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4998.345 1046.435 4998.625 1047.435 ;
    END
  END Data_PMOS_NOSF[1017]
  PIN Data_PMOS_NOSF[1012]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4996.665 1046.435 4996.945 1047.435 ;
    END
  END Data_PMOS_NOSF[1012]
  PIN Data_PMOS_NOSF[1009]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4994.985 1046.435 4995.265 1047.435 ;
    END
  END Data_PMOS_NOSF[1009]
  PIN MASKV[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4954.665 1046.435 4954.945 1047.435 ;
    END
  END MASKV[96]
  PIN DIG_MON_PMOS_NOSF[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4952.425 1046.435 4952.705 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[96]
  PIN DIG_MON_SEL[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4950.745 1046.435 4951.025 1047.435 ;
    END
  END DIG_MON_SEL[96]
  PIN Data_PMOS_NOSF[1005]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4945.705 1046.435 4945.985 1047.435 ;
    END
  END Data_PMOS_NOSF[1005]
  PIN Data_PMOS_NOSF[1006]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4944.025 1046.435 4944.305 1047.435 ;
    END
  END Data_PMOS_NOSF[1006]
  PIN Data_PMOS_NOSF[1007]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4942.345 1046.435 4942.625 1047.435 ;
    END
  END Data_PMOS_NOSF[1007]
  PIN Data_PMOS_NOSF[994]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4941.225 1046.435 4941.505 1047.435 ;
    END
  END Data_PMOS_NOSF[994]
  PIN INJ_IN[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4931.145 1046.435 4931.425 1047.435 ;
    END
  END INJ_IN[95]
  PIN BcidMtx[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4927.785 1046.435 4928.065 1047.435 ;
    END
  END BcidMtx[285]
  PIN BcidMtx[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4926.105 1046.435 4926.385 1047.435 ;
    END
  END BcidMtx[284]
  PIN BcidMtx[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4924.985 1046.435 4925.265 1047.435 ;
    END
  END BcidMtx[282]
  PIN Data_PMOS_NOSF[996]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4919.665 1046.435 4919.945 1047.435 ;
    END
  END Data_PMOS_NOSF[996]
  PIN Data_PMOS_NOSF[991]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4892.505 1046.435 4892.785 1047.435 ;
    END
  END Data_PMOS_NOSF[991]
  PIN Data_PMOS_NOSF[998]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4891.385 1046.435 4891.665 1047.435 ;
    END
  END Data_PMOS_NOSF[998]
  PIN MASKV[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4889.145 1046.435 4889.425 1047.435 ;
    END
  END MASKV[94]
  PIN DIG_MON_PMOS_NOSF[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4886.905 1046.435 4887.185 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[94]
  PIN DIG_MON_SEL[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4885.225 1046.435 4885.505 1047.435 ;
    END
  END DIG_MON_SEL[94]
  PIN INJ_ROW[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4881.305 1046.435 4881.585 1047.435 ;
    END
  END INJ_ROW[46]
  PIN Data_PMOS_NOSF[974]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4879.625 1046.435 4879.905 1047.435 ;
    END
  END Data_PMOS_NOSF[974]
  PIN Data_PMOS_NOSF[985]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4865.625 1046.435 4865.905 1047.435 ;
    END
  END Data_PMOS_NOSF[985]
  PIN Data_PMOS_NOSF[980]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4863.385 1046.435 4863.665 1047.435 ;
    END
  END Data_PMOS_NOSF[980]
  PIN INJ_IN[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4861.145 1046.435 4861.425 1047.435 ;
    END
  END INJ_IN[93]
  PIN BcidMtx[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4858.905 1046.435 4859.185 1047.435 ;
    END
  END BcidMtx[281]
  PIN Read_PMOS_NOSF[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4856.665 1046.435 4856.945 1047.435 ;
    END
  END Read_PMOS_NOSF[46]
  PIN BcidMtx[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4854.985 1046.435 4855.265 1047.435 ;
    END
  END BcidMtx[276]
  PIN Data_PMOS_NOSF[969]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4814.105 1046.435 4814.385 1047.435 ;
    END
  END Data_PMOS_NOSF[969]
  PIN Data_PMOS_NOSF[976]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4811.865 1046.435 4812.145 1047.435 ;
    END
  END Data_PMOS_NOSF[976]
  PIN Data_PMOS_NOSF[977]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4810.185 1046.435 4810.465 1047.435 ;
    END
  END Data_PMOS_NOSF[977]
  PIN Data_PMOS_NOSF[966]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4809.065 1046.435 4809.345 1047.435 ;
    END
  END Data_PMOS_NOSF[966]
  PIN MASKD[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4806.825 1046.435 4807.105 1047.435 ;
    END
  END MASKD[92]
  PIN DIG_MON_SEL[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4804.025 1046.435 4804.305 1047.435 ;
    END
  END DIG_MON_SEL[92]
  PIN DIG_MON_SEL[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4803.465 1046.435 4803.745 1047.435 ;
    END
  END DIG_MON_SEL[91]
  PIN MASKV[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4791.145 1046.435 4791.425 1047.435 ;
    END
  END MASKV[91]
  PIN Data_PMOS_NOSF[957]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4789.465 1046.435 4789.745 1047.435 ;
    END
  END Data_PMOS_NOSF[957]
  PIN Data_PMOS_NOSF[950]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4788.345 1046.435 4788.625 1047.435 ;
    END
  END Data_PMOS_NOSF[950]
  PIN Data_PMOS_NOSF[952]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4786.105 1046.435 4786.385 1047.435 ;
    END
  END Data_PMOS_NOSF[952]
  PIN nTOK_PMOS_NOSF[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4781.345 1046.435 4781.625 1047.435 ;
    END
  END nTOK_PMOS_NOSF[45]
  PIN BcidMtx[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4779.665 1046.435 4779.945 1047.435 ;
    END
  END BcidMtx[274]
  PIN BcidMtx[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4751.385 1046.435 4751.665 1047.435 ;
    END
  END BcidMtx[271]
  PIN Data_PMOS_NOSF[948]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4748.585 1046.435 4748.865 1047.435 ;
    END
  END Data_PMOS_NOSF[948]
  PIN Data_PMOS_NOSF[954]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4747.465 1046.435 4747.745 1047.435 ;
    END
  END Data_PMOS_NOSF[954]
  PIN Data_PMOS_NOSF[961]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4745.225 1046.435 4745.505 1047.435 ;
    END
  END Data_PMOS_NOSF[961]
  PIN Data_PMOS_NOSF[945]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4743.545 1046.435 4743.825 1047.435 ;
    END
  END Data_PMOS_NOSF[945]
  PIN MASKV[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4742.425 1046.435 4742.705 1047.435 ;
    END
  END MASKV[90]
  PIN MASKD[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4723.945 1046.435 4724.225 1047.435 ;
    END
  END MASKD[89]
  PIN INJ_ROW[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4721.705 1046.435 4721.985 1047.435 ;
    END
  END INJ_ROW[44]
  PIN Data_PMOS_NOSF[936]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4719.465 1046.435 4719.745 1047.435 ;
    END
  END Data_PMOS_NOSF[936]
  PIN Data_PMOS_NOSF[937]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4717.785 1046.435 4718.065 1047.435 ;
    END
  END Data_PMOS_NOSF[937]
  PIN Data_PMOS_NOSF[938]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4716.665 1046.435 4716.945 1047.435 ;
    END
  END Data_PMOS_NOSF[938]
  PIN nTOK_PMOS_NOSF[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4674.105 1046.435 4674.385 1047.435 ;
    END
  END nTOK_PMOS_NOSF[44]
  PIN BcidMtx[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4671.865 1046.435 4672.145 1047.435 ;
    END
  END BcidMtx[267]
  PIN Read_PMOS_NOSF[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4670.745 1046.435 4671.025 1047.435 ;
    END
  END Read_PMOS_NOSF[44]
  PIN INJ_IN[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4667.945 1046.435 4668.225 1047.435 ;
    END
  END INJ_IN[88]
  PIN Data_PMOS_NOSF[933]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4665.705 1046.435 4665.985 1047.435 ;
    END
  END Data_PMOS_NOSF[933]
  PIN Data_PMOS_NOSF[934]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4664.585 1046.435 4664.865 1047.435 ;
    END
  END Data_PMOS_NOSF[934]
  PIN Data_PMOS_NOSF[925]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4662.345 1046.435 4662.625 1047.435 ;
    END
  END Data_PMOS_NOSF[925]
  PIN MASKV[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4652.265 1046.435 4652.545 1047.435 ;
    END
  END MASKV[88]
  PIN MASKD[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4651.145 1046.435 4651.425 1047.435 ;
    END
  END MASKD[88]
  PIN DIG_MON_SEL[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4647.785 1046.435 4648.065 1047.435 ;
    END
  END DIG_MON_SEL[87]
  PIN INJ_ROW[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4642.465 1046.435 4642.745 1047.435 ;
    END
  END INJ_ROW[43]
  PIN Data_PMOS_NOSF[921]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4641.345 1046.435 4641.625 1047.435 ;
    END
  END Data_PMOS_NOSF[921]
  PIN Data_PMOS_NOSF[908]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4639.105 1046.435 4639.385 1047.435 ;
    END
  END Data_PMOS_NOSF[908]
  PIN Data_PMOS_NOSF[917]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4611.945 1046.435 4612.225 1047.435 ;
    END
  END Data_PMOS_NOSF[917]
  PIN Data_PMOS_NOSF[909]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4610.825 1046.435 4611.105 1047.435 ;
    END
  END Data_PMOS_NOSF[909]
  PIN BcidMtx[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4606.905 1046.435 4607.185 1047.435 ;
    END
  END BcidMtx[262]
  PIN Read_PMOS_NOSF[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4605.225 1046.435 4605.505 1047.435 ;
    END
  END Read_PMOS_NOSF[43]
  PIN BcidMtx[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4604.105 1046.435 4604.385 1047.435 ;
    END
  END BcidMtx[259]
  PIN Data_PMOS_NOSF[905]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4600.745 1046.435 4601.025 1047.435 ;
    END
  END Data_PMOS_NOSF[905]
  PIN Data_PMOS_NOSF[913]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4586.185 1046.435 4586.465 1047.435 ;
    END
  END Data_PMOS_NOSF[913]
  PIN Data_PMOS_NOSF[919]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4585.065 1046.435 4585.345 1047.435 ;
    END
  END Data_PMOS_NOSF[919]
  PIN Data_PMOS_NOSF[920]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4582.825 1046.435 4583.105 1047.435 ;
    END
  END Data_PMOS_NOSF[920]
  PIN MASKD[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4581.145 1046.435 4581.425 1047.435 ;
    END
  END MASKD[86]
  PIN DIG_MON_PMOS_NOSF[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4575.545 1046.435 4575.825 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[85]
  PIN Data_HV[1133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18863.945 1046.435 18864.225 1047.435 ;
    END
  END Data_HV[1133]
  PIN Data_PMOS_NOSF[890]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4532.985 1046.435 4533.265 1047.435 ;
    END
  END Data_PMOS_NOSF[890]
  PIN Data_PMOS_NOSF[887]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4531.305 1046.435 4531.585 1047.435 ;
    END
  END Data_PMOS_NOSF[887]
  PIN Data_PMOS_NOSF[896]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4529.625 1046.435 4529.905 1047.435 ;
    END
  END Data_PMOS_NOSF[896]
  PIN Data_PMOS_NOSF[888]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4528.505 1046.435 4528.785 1047.435 ;
    END
  END Data_PMOS_NOSF[888]
  PIN BcidMtx[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4524.585 1046.435 4524.865 1047.435 ;
    END
  END BcidMtx[256]
  PIN FREEZE_PMOS_NOSF[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4523.465 1046.435 4523.745 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[42]
  PIN BcidMtx[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4522.345 1046.435 4522.625 1047.435 ;
    END
  END BcidMtx[254]
  PIN Data_PMOS_NOSF[885]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4510.585 1046.435 4510.865 1047.435 ;
    END
  END Data_PMOS_NOSF[885]
  PIN Data_PMOS_NOSF[897]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4508.905 1046.435 4509.185 1047.435 ;
    END
  END Data_PMOS_NOSF[897]
  PIN Data_PMOS_NOSF[886]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4507.785 1046.435 4508.065 1047.435 ;
    END
  END Data_PMOS_NOSF[886]
  PIN Data_PMOS_NOSF[882]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4505.545 1046.435 4505.825 1047.435 ;
    END
  END Data_PMOS_NOSF[882]
  PIN MASKH[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4501.905 1046.435 4502.185 1047.435 ;
    END
  END MASKH[42]
  PIN DIG_MON_PMOS_NOSF[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4500.225 1046.435 4500.505 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[84]
  PIN DIG_MON_SEL[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5591.945 1046.435 5592.225 1047.435 ;
    END
  END DIG_MON_SEL[111]
  PIN INJ_ROW[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5588.585 1046.435 5588.865 1047.435 ;
    END
  END INJ_ROW[55]
  PIN Data_PMOS_NOSF[869]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4466.905 1046.435 4467.185 1047.435 ;
    END
  END Data_PMOS_NOSF[869]
  PIN Data_PMOS_NOSF[880]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4465.785 1046.435 4466.065 1047.435 ;
    END
  END Data_PMOS_NOSF[880]
  PIN Data_PMOS_NOSF[874]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4464.665 1046.435 4464.945 1047.435 ;
    END
  END Data_PMOS_NOSF[874]
  PIN INJ_IN[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4461.305 1046.435 4461.585 1047.435 ;
    END
  END INJ_IN[83]
  PIN BcidMtx[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4445.625 1046.435 4445.905 1047.435 ;
    END
  END BcidMtx[251]
  PIN BcidMtx[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4444.505 1046.435 4444.785 1047.435 ;
    END
  END BcidMtx[249]
  PIN BcidMtx[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4442.265 1046.435 4442.545 1047.435 ;
    END
  END BcidMtx[247]
  PIN INJ_IN[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4440.585 1046.435 4440.865 1047.435 ;
    END
  END INJ_IN[82]
  PIN Data_PMOS_NOSF[863]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4438.905 1046.435 4439.185 1047.435 ;
    END
  END Data_PMOS_NOSF[863]
  PIN Data_PMOS_NOSF[877]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4436.105 1046.435 4436.385 1047.435 ;
    END
  END Data_PMOS_NOSF[877]
  PIN Data_PMOS_NOSF[862]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4434.985 1046.435 4435.265 1047.435 ;
    END
  END Data_PMOS_NOSF[862]
  PIN Data_PMOS_NOSF[878]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4433.865 1046.435 4434.145 1047.435 ;
    END
  END Data_PMOS_NOSF[878]
  PIN DIG_MON_SEL[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4390.185 1046.435 4390.465 1047.435 ;
    END
  END DIG_MON_SEL[81]
  PIN DIG_MON_PMOS_NOSF[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4387.945 1046.435 4388.225 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[81]
  PIN Data_PMOS_NOSF[852]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4384.585 1046.435 4384.865 1047.435 ;
    END
  END Data_PMOS_NOSF[852]
  PIN Data_PMOS_NOSF[845]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4383.465 1046.435 4383.745 1047.435 ;
    END
  END Data_PMOS_NOSF[845]
  PIN Data_PMOS_NOSF[860]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4382.345 1046.435 4382.625 1047.435 ;
    END
  END Data_PMOS_NOSF[860]
  PIN nTOK_PMOS_NOSF[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4370.025 1046.435 4370.305 1047.435 ;
    END
  END nTOK_PMOS_NOSF[40]
  PIN BcidMtx[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4368.345 1046.435 4368.625 1047.435 ;
    END
  END BcidMtx[244]
  PIN FREEZE_PMOS_NOSF[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4367.225 1046.435 4367.505 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[40]
  PIN INJ_IN[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4361.905 1046.435 4362.185 1047.435 ;
    END
  END INJ_IN[80]
  PIN Data_PMOS_NOSF[842]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4360.225 1046.435 4360.505 1047.435 ;
    END
  END Data_PMOS_NOSF[842]
  PIN Data_PMOS_NOSF[855]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4359.105 1046.435 4359.385 1047.435 ;
    END
  END Data_PMOS_NOSF[855]
  PIN Data_PMOS_NOSF[841]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4330.825 1046.435 4331.105 1047.435 ;
    END
  END Data_PMOS_NOSF[841]
  PIN Data_PMOS_NOSF[857]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4329.705 1046.435 4329.985 1047.435 ;
    END
  END Data_PMOS_NOSF[857]
  PIN MASKH[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4328.585 1046.435 4328.865 1047.435 ;
    END
  END MASKH[40]
  PIN DIG_MON_SEL[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4324.665 1046.435 4324.945 1047.435 ;
    END
  END DIG_MON_SEL[79]
  PIN INJ_ROW[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4321.305 1046.435 4321.585 1047.435 ;
    END
  END INJ_ROW[39]
  PIN Data_PMOS_NOSF[837]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4320.185 1046.435 4320.465 1047.435 ;
    END
  END Data_PMOS_NOSF[837]
  PIN Data_PMOS_NOSF[824]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4305.065 1046.435 4305.345 1047.435 ;
    END
  END Data_PMOS_NOSF[824]
  PIN Data_PMOS_NOSF[833]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4303.385 1046.435 4303.665 1047.435 ;
    END
  END Data_PMOS_NOSF[833]
  PIN Data_PMOS_NOSF[825]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4302.265 1046.435 4302.545 1047.435 ;
    END
  END Data_PMOS_NOSF[825]
  PIN BcidMtx[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4297.785 1046.435 4298.065 1047.435 ;
    END
  END BcidMtx[237]
  PIN Read_PMOS_NOSF[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4296.665 1046.435 4296.945 1047.435 ;
    END
  END Read_PMOS_NOSF[39]
  PIN BcidMtx[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4296.105 1046.435 4296.385 1047.435 ;
    END
  END BcidMtx[236]
  PIN Data_PMOS_NOSF[821]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4253.545 1046.435 4253.825 1047.435 ;
    END
  END Data_PMOS_NOSF[821]
  PIN Data_PMOS_NOSF[834]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4252.425 1046.435 4252.705 1047.435 ;
    END
  END Data_PMOS_NOSF[834]
  PIN Data_PMOS_NOSF[823]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4251.305 1046.435 4251.585 1047.435 ;
    END
  END Data_PMOS_NOSF[823]
  PIN Data_PMOS_NOSF[836]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4248.505 1046.435 4248.785 1047.435 ;
    END
  END Data_PMOS_NOSF[836]
  PIN MASKH[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4247.385 1046.435 4247.665 1047.435 ;
    END
  END MASKH[39]
  PIN DIG_MON_PMOS_NOSF[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4245.705 1046.435 4245.985 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[78]
  PIN DIG_MON_PMOS_NOSF[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4241.225 1046.435 4241.505 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[77]
  PIN Data_PMOS_NOSF[816]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4230.585 1046.435 4230.865 1047.435 ;
    END
  END Data_PMOS_NOSF[816]
  PIN Data_PMOS_NOSF[817]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4228.905 1046.435 4229.185 1047.435 ;
    END
  END Data_PMOS_NOSF[817]
  PIN Data_PMOS_NOSF[818]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4227.225 1046.435 4227.505 1047.435 ;
    END
  END Data_PMOS_NOSF[818]
  PIN Data_PMOS_NOSF[804]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4225.545 1046.435 4225.825 1047.435 ;
    END
  END Data_PMOS_NOSF[804]
  PIN BcidMtx[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4220.225 1046.435 4220.505 1047.435 ;
    END
  END BcidMtx[233]
  PIN Read_PMOS_NOSF[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4192.505 1046.435 4192.785 1047.435 ;
    END
  END Read_PMOS_NOSF[38]
  PIN BcidMtx[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4190.825 1046.435 4191.105 1047.435 ;
    END
  END BcidMtx[228]
  PIN Data_PMOS_NOSF[800]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4188.025 1046.435 4188.305 1047.435 ;
    END
  END Data_PMOS_NOSF[800]
  PIN Data_PMOS_NOSF[808]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4186.345 1046.435 4186.625 1047.435 ;
    END
  END Data_PMOS_NOSF[808]
  PIN Data_PMOS_NOSF[809]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4184.665 1046.435 4184.945 1047.435 ;
    END
  END Data_PMOS_NOSF[809]
  PIN Data_PMOS_NOSF[815]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4182.985 1046.435 4183.265 1047.435 ;
    END
  END Data_PMOS_NOSF[815]
  PIN MASKD[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4181.305 1046.435 4181.585 1047.435 ;
    END
  END MASKD[76]
  PIN MASKD[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4163.945 1046.435 4164.225 1047.435 ;
    END
  END MASKD[75]
  PIN MASKV[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4161.145 1046.435 4161.425 1047.435 ;
    END
  END MASKV[75]
  PIN Data_PMOS_NOSF[785]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4160.025 1046.435 4160.305 1047.435 ;
    END
  END Data_PMOS_NOSF[785]
  PIN Data_PMOS_NOSF[790]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4157.785 1046.435 4158.065 1047.435 ;
    END
  END Data_PMOS_NOSF[790]
  PIN Data_PMOS_NOSF[784]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4156.105 1046.435 4156.385 1047.435 ;
    END
  END Data_PMOS_NOSF[784]
  PIN INJ_IN[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4154.425 1046.435 4154.705 1047.435 ;
    END
  END INJ_IN[75]
  PIN BcidMtx[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4111.865 1046.435 4112.145 1047.435 ;
    END
  END BcidMtx[225]
  PIN BcidMtx[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4110.185 1046.435 4110.465 1047.435 ;
    END
  END BcidMtx[224]
  PIN BcidMtx[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4109.065 1046.435 4109.345 1047.435 ;
    END
  END BcidMtx[222]
  PIN Data_PMOS_NOSF[786]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4105.705 1046.435 4105.985 1047.435 ;
    END
  END Data_PMOS_NOSF[786]
  PIN Data_PMOS_NOSF[781]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4104.025 1046.435 4104.305 1047.435 ;
    END
  END Data_PMOS_NOSF[781]
  PIN Data_PMOS_NOSF[788]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4102.905 1046.435 4103.185 1047.435 ;
    END
  END Data_PMOS_NOSF[788]
  PIN MASKV[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4092.265 1046.435 4092.545 1047.435 ;
    END
  END MASKV[74]
  PIN DIG_MON_PMOS_NOSF[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4090.025 1046.435 4090.305 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[74]
  PIN DIG_MON_SEL[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4088.345 1046.435 4088.625 1047.435 ;
    END
  END DIG_MON_SEL[74]
  PIN MASKD[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4086.665 1046.435 4086.945 1047.435 ;
    END
  END MASKD[73]
  PIN MASKV[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4081.905 1046.435 4082.185 1047.435 ;
    END
  END MASKV[73]
  PIN Data_PMOS_NOSF[768]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4080.225 1046.435 4080.505 1047.435 ;
    END
  END Data_PMOS_NOSF[768]
  PIN Data_PMOS_NOSF[769]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4053.065 1046.435 4053.345 1047.435 ;
    END
  END Data_PMOS_NOSF[769]
  PIN Data_PMOS_NOSF[763]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4051.385 1046.435 4051.665 1047.435 ;
    END
  END Data_PMOS_NOSF[763]
  PIN nTOK_PMOS_NOSF[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4048.585 1046.435 4048.865 1047.435 ;
    END
  END nTOK_PMOS_NOSF[36]
  PIN BcidMtx[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4046.345 1046.435 4046.625 1047.435 ;
    END
  END BcidMtx[219]
  PIN BcidMtx[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4044.665 1046.435 4044.945 1047.435 ;
    END
  END BcidMtx[218]
  PIN INJ_IN[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4042.425 1046.435 4042.705 1047.435 ;
    END
  END INJ_IN[72]
  PIN Data_PMOS_NOSF[765]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4040.185 1046.435 4040.465 1047.435 ;
    END
  END Data_PMOS_NOSF[765]
  PIN Data_PMOS_NOSF[760]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4025.625 1046.435 4025.905 1047.435 ;
    END
  END Data_PMOS_NOSF[760]
  PIN Data_PMOS_NOSF[757]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4023.945 1046.435 4024.225 1047.435 ;
    END
  END Data_PMOS_NOSF[757]
  PIN MASKV[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4022.265 1046.435 4022.545 1047.435 ;
    END
  END MASKV[72]
  PIN DIG_MON_PMOS_NOSF[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4020.025 1046.435 4020.305 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[72]
  PIN DIG_MON_SEL[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4017.785 1046.435 4018.065 1047.435 ;
    END
  END DIG_MON_SEL[71]
  PIN INJ_ROW[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 4014.425 1046.435 4014.705 1047.435 ;
    END
  END INJ_ROW[35]
  PIN Data_PMOS_NOSF[743]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3972.985 1046.435 3973.265 1047.435 ;
    END
  END Data_PMOS_NOSF[743]
  PIN Data_PMOS_NOSF[740]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3971.305 1046.435 3971.585 1047.435 ;
    END
  END Data_PMOS_NOSF[740]
  PIN DIG_MON_HV[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18650.025 1046.435 18650.305 1047.435 ;
    END
  END DIG_MON_HV[102]
  PIN Data_PMOS_NOSF[742]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3969.065 1046.435 3969.345 1047.435 ;
    END
  END Data_PMOS_NOSF[742]
  PIN INJ_IN[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3967.385 1046.435 3967.665 1047.435 ;
    END
  END INJ_IN[71]
  PIN BcidMtx[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3964.585 1046.435 3964.865 1047.435 ;
    END
  END BcidMtx[214]
  PIN Read_PMOS_NOSF[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3962.905 1046.435 3963.185 1047.435 ;
    END
  END Read_PMOS_NOSF[35]
  PIN INJ_IN[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3951.705 1046.435 3951.985 1047.435 ;
    END
  END INJ_IN[70]
  PIN Data_PMOS_NOSF[737]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3950.025 1046.435 3950.305 1047.435 ;
    END
  END Data_PMOS_NOSF[737]
  PIN Data_PMOS_NOSF[745]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3948.345 1046.435 3948.625 1047.435 ;
    END
  END Data_PMOS_NOSF[745]
  PIN Data_PMOS_NOSF[746]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3946.665 1046.435 3946.945 1047.435 ;
    END
  END Data_PMOS_NOSF[746]
  PIN Data_PMOS_NOSF[752]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3944.985 1046.435 3945.265 1047.435 ;
    END
  END Data_PMOS_NOSF[752]
  PIN MASKD[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3941.345 1046.435 3941.625 1047.435 ;
    END
  END MASKD[70]
  PIN DIG_MON_SEL[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3938.545 1046.435 3938.825 1047.435 ;
    END
  END DIG_MON_SEL[70]
  PIN MASKD[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5030.825 1046.435 5031.105 1047.435 ;
    END
  END MASKD[97]
  PIN MASKV[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5028.025 1046.435 5028.305 1047.435 ;
    END
  END MASKV[97]
  PIN DIG_MON_PMOS[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6149.705 1046.435 6149.985 1047.435 ;
    END
  END DIG_MON_PMOS[13]
  PIN MASKV[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6148.025 1046.435 6148.305 1047.435 ;
    END
  END MASKV[125]
  PIN Data_PMOS[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6145.785 1046.435 6146.065 1047.435 ;
    END
  END Data_PMOS[145]
  PIN Data_PMOS[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6144.105 1046.435 6144.385 1047.435 ;
    END
  END Data_PMOS[146]
  PIN Data_PMOS[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6142.985 1046.435 6143.265 1047.435 ;
    END
  END Data_PMOS[133]
  PIN BcidMtx[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6125.625 1046.435 6125.905 1047.435 ;
    END
  END BcidMtx[377]
  PIN FREEZE_PMOS[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6123.945 1046.435 6124.225 1047.435 ;
    END
  END FREEZE_PMOS[6]
  PIN BcidMtx[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6122.825 1046.435 6123.105 1047.435 ;
    END
  END BcidMtx[374]
  PIN Data_PMOS[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6119.465 1046.435 6119.745 1047.435 ;
    END
  END Data_PMOS[129]
  PIN Data_PMOS[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6117.785 1046.435 6118.065 1047.435 ;
    END
  END Data_PMOS[141]
  PIN Data_PMOS[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6116.665 1046.435 6116.945 1047.435 ;
    END
  END Data_PMOS[130]
  PIN Data_PMOS[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6113.865 1046.435 6114.145 1047.435 ;
    END
  END Data_PMOS[143]
  PIN MASKH[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6074.105 1046.435 6074.385 1047.435 ;
    END
  END MASKH[62]
  PIN DIG_MON_PMOS[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6072.425 1046.435 6072.705 1047.435 ;
    END
  END DIG_MON_PMOS[12]
  PIN MASKD[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6069.065 1046.435 6069.345 1047.435 ;
    END
  END MASKD[123]
  PIN MASKV[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6066.265 1046.435 6066.545 1047.435 ;
    END
  END MASKV[123]
  PIN Data_PMOS[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6065.705 1046.435 6065.985 1047.435 ;
    END
  END Data_PMOS[123]
  PIN Data_PMOS[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6062.905 1046.435 6063.185 1047.435 ;
    END
  END Data_PMOS[118]
  PIN Data_PMOS[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6061.225 1046.435 6061.505 1047.435 ;
    END
  END Data_PMOS[112]
  PIN Data_PMOS[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6052.265 1046.435 6052.545 1047.435 ;
    END
  END Data_PMOS[111]
  PIN BcidMtx[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6047.785 1046.435 6048.065 1047.435 ;
    END
  END BcidMtx[369]
  PIN BcidMtx[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6046.105 1046.435 6046.385 1047.435 ;
    END
  END BcidMtx[368]
  PIN BcidMtx[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6045.545 1046.435 6045.825 1047.435 ;
    END
  END BcidMtx[367]
  PIN Data_PMOS[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6039.665 1046.435 6039.945 1047.435 ;
    END
  END Data_PMOS[114]
  PIN Data_PMOS[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6012.505 1046.435 6012.785 1047.435 ;
    END
  END Data_PMOS[109]
  PIN Data_PMOS[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6011.945 1046.435 6012.225 1047.435 ;
    END
  END Data_PMOS[121]
  PIN MASKV[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6009.145 1046.435 6009.425 1047.435 ;
    END
  END MASKV[122]
  PIN DIG_MON_PMOS[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6006.905 1046.435 6007.185 1047.435 ;
    END
  END DIG_MON_PMOS[10]
  PIN INJ_ROW[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6001.305 1046.435 6001.585 1047.435 ;
    END
  END INJ_ROW[60]
  PIN Data_PMOS[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6000.185 1046.435 6000.465 1047.435 ;
    END
  END Data_PMOS[102]
  PIN Data_PMOS[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5999.625 1046.435 5999.905 1047.435 ;
    END
  END Data_PMOS[92]
  PIN Data_PMOS[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5983.945 1046.435 5984.225 1047.435 ;
    END
  END Data_PMOS[104]
  PIN Data_PMOS[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5982.265 1046.435 5982.545 1047.435 ;
    END
  END Data_PMOS[90]
  PIN INJ_IN[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5981.145 1046.435 5981.425 1047.435 ;
    END
  END INJ_IN[121]
  PIN FREEZE_PMOS[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5977.225 1046.435 5977.505 1047.435 ;
    END
  END FREEZE_PMOS[4]
  PIN BcidMtx[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5975.545 1046.435 5975.825 1047.435 ;
    END
  END BcidMtx[361]
  PIN BcidMtx[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5974.985 1046.435 5975.265 1047.435 ;
    END
  END BcidMtx[360]
  PIN Data_PMOS[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5932.425 1046.435 5932.705 1047.435 ;
    END
  END Data_PMOS[99]
  PIN Data_PMOS[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5930.745 1046.435 5931.025 1047.435 ;
    END
  END Data_PMOS[100]
  PIN Data_PMOS[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5930.185 1046.435 5930.465 1047.435 ;
    END
  END Data_PMOS[95]
  PIN MASKH[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5927.385 1046.435 5927.665 1047.435 ;
    END
  END MASKH[60]
  PIN DIG_MON_SEL[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5924.025 1046.435 5924.305 1047.435 ;
    END
  END DIG_MON_SEL[120]
  PIN MASKV[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5911.145 1046.435 5911.425 1047.435 ;
    END
  END MASKV[119]
  PIN Data_PMOS[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5909.465 1046.435 5909.745 1047.435 ;
    END
  END Data_PMOS[75]
  PIN Data_PMOS[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5908.905 1046.435 5909.185 1047.435 ;
    END
  END Data_PMOS[82]
  PIN Data_PMOS[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5906.105 1046.435 5906.385 1047.435 ;
    END
  END Data_PMOS[70]
  PIN nTOK_PMOS[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5901.345 1046.435 5901.625 1047.435 ;
    END
  END nTOK_PMOS[3]
  PIN BcidMtx[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5900.225 1046.435 5900.505 1047.435 ;
    END
  END BcidMtx[359]
  PIN BcidMtx[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5871.385 1046.435 5871.665 1047.435 ;
    END
  END BcidMtx[355]
  PIN Data_PMOS[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5868.585 1046.435 5868.865 1047.435 ;
    END
  END Data_PMOS[66]
  PIN Data_PMOS[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5868.025 1046.435 5868.305 1047.435 ;
    END
  END Data_PMOS[65]
  PIN Data_PMOS[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5866.345 1046.435 5866.625 1047.435 ;
    END
  END Data_PMOS[73]
  PIN Data_PMOS[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5863.545 1046.435 5863.825 1047.435 ;
    END
  END Data_PMOS[63]
  PIN MASKV[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5862.425 1046.435 5862.705 1047.435 ;
    END
  END MASKV[118]
  PIN MASKD[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5861.305 1046.435 5861.585 1047.435 ;
    END
  END MASKD[118]
  PIN DIG_MON_SEL[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5845.625 1046.435 5845.905 1047.435 ;
    END
  END DIG_MON_SEL[118]
  PIN DIG_MON_PMOS[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5842.825 1046.435 5843.105 1047.435 ;
    END
  END DIG_MON_PMOS[5]
  PIN Data_PMOS[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5840.585 1046.435 5840.865 1047.435 ;
    END
  END Data_PMOS[60]
  PIN Data_PMOS[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5838.905 1046.435 5839.185 1047.435 ;
    END
  END Data_PMOS[61]
  PIN Data_PMOS[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5837.225 1046.435 5837.505 1047.435 ;
    END
  END Data_PMOS[62]
  PIN Data_PMOS[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5835.545 1046.435 5835.825 1047.435 ;
    END
  END Data_PMOS[48]
  PIN BcidMtx[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5792.985 1046.435 5793.265 1047.435 ;
    END
  END BcidMtx[353]
  PIN FREEZE_PMOS[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5791.305 1046.435 5791.585 1047.435 ;
    END
  END FREEZE_PMOS[2]
  PIN BcidMtx[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5789.625 1046.435 5789.905 1047.435 ;
    END
  END BcidMtx[349]
  PIN Data_PMOS[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5786.825 1046.435 5787.105 1047.435 ;
    END
  END Data_PMOS[45]
  PIN Data_PMOS[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5784.585 1046.435 5784.865 1047.435 ;
    END
  END Data_PMOS[52]
  PIN Data_PMOS[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5782.905 1046.435 5783.185 1047.435 ;
    END
  END Data_PMOS[53]
  PIN Data_PMOS[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5781.225 1046.435 5781.505 1047.435 ;
    END
  END Data_PMOS[59]
  PIN MASKD[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5771.145 1046.435 5771.425 1047.435 ;
    END
  END MASKD[116]
  PIN DIG_MON_SEL[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5768.345 1046.435 5768.625 1047.435 ;
    END
  END DIG_MON_SEL[116]
  PIN MASKV[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5761.905 1046.435 5762.185 1047.435 ;
    END
  END MASKV[115]
  PIN Data_PMOS[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5761.345 1046.435 5761.625 1047.435 ;
    END
  END Data_PMOS[39]
  PIN Data_PMOS[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5759.665 1046.435 5759.945 1047.435 ;
    END
  END Data_PMOS[40]
  PIN Data_PMOS[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5732.505 1046.435 5732.785 1047.435 ;
    END
  END Data_PMOS[41]
  PIN nTOK_PMOS[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5728.585 1046.435 5728.865 1047.435 ;
    END
  END nTOK_PMOS[1]
  PIN BcidMtx[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5727.465 1046.435 5727.745 1047.435 ;
    END
  END BcidMtx[347]
  PIN Read_PMOS[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5725.225 1046.435 5725.505 1047.435 ;
    END
  END Read_PMOS[1]
  PIN BcidMtx[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5724.105 1046.435 5724.385 1047.435 ;
    END
  END BcidMtx[343]
  PIN Data_PMOS[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5721.305 1046.435 5721.585 1047.435 ;
    END
  END Data_PMOS[24]
  PIN Data_PMOS[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5706.185 1046.435 5706.465 1047.435 ;
    END
  END Data_PMOS[31]
  PIN Data_PMOS[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5704.505 1046.435 5704.785 1047.435 ;
    END
  END Data_PMOS[32]
  PIN Data_PMOS[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5703.385 1046.435 5703.665 1047.435 ;
    END
  END Data_PMOS[21]
  PIN MASKH[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5701.705 1046.435 5701.985 1047.435 ;
    END
  END MASKH[57]
  PIN FREEZE_HV[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18857.225 1046.435 18857.505 1047.435 ;
    END
  END FREEZE_HV[53]
  PIN DIG_MON_SEL[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5698.345 1046.435 5698.625 1047.435 ;
    END
  END DIG_MON_SEL[114]
  PIN DIG_MON_PMOS[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5695.545 1046.435 5695.825 1047.435 ;
    END
  END DIG_MON_PMOS[1]
  PIN Data_PMOS[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5652.985 1046.435 5653.265 1047.435 ;
    END
  END Data_PMOS[8]
  PIN Data_PMOS[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5651.865 1046.435 5652.145 1047.435 ;
    END
  END Data_PMOS[19]
  PIN Data_PMOS[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5650.185 1046.435 5650.465 1047.435 ;
    END
  END Data_PMOS[20]
  PIN INJ_IN[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5647.385 1046.435 5647.665 1047.435 ;
    END
  END INJ_IN[113]
  PIN BcidMtx[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5645.145 1046.435 5645.425 1047.435 ;
    END
  END BcidMtx[341]
  PIN FREEZE_PMOS[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5643.465 1046.435 5643.745 1047.435 ;
    END
  END FREEZE_PMOS[0]
  PIN INJ_IN[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5631.705 1046.435 5631.985 1047.435 ;
    END
  END INJ_IN[112]
  PIN Data_PMOS[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5630.025 1046.435 5630.305 1047.435 ;
    END
  END Data_PMOS[2]
  PIN Data_PMOS[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5628.905 1046.435 5629.185 1047.435 ;
    END
  END Data_PMOS[15]
  PIN Data_PMOS[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5626.105 1046.435 5626.385 1047.435 ;
    END
  END Data_PMOS[1]
  PIN Data_PMOS[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5625.545 1046.435 5625.825 1047.435 ;
    END
  END Data_PMOS[0]
  PIN BcidMtx[1329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18857.785 1046.435 18858.065 1047.435 ;
    END
  END BcidMtx[1329]
  PIN Read_HV[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18856.665 1046.435 18856.945 1047.435 ;
    END
  END Read_HV[53]
  PIN FREEZE_PMOS[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5873.065 1046.435 5873.345 1047.435 ;
    END
  END FREEZE_PMOS[3]
  PIN Data_PMOS_NOSF[1173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5587.465 1046.435 5587.745 1047.435 ;
    END
  END Data_PMOS_NOSF[1173]
  PIN Data_PMOS_NOSF[1160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5585.225 1046.435 5585.505 1047.435 ;
    END
  END Data_PMOS_NOSF[1160]
  PIN Data_PMOS_NOSF[1175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5584.105 1046.435 5584.385 1047.435 ;
    END
  END Data_PMOS_NOSF[1175]
  PIN Data_PMOS_NOSF[1162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5582.985 1046.435 5583.265 1047.435 ;
    END
  END Data_PMOS_NOSF[1162]
  PIN BcidMtx[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5565.625 1046.435 5565.905 1047.435 ;
    END
  END BcidMtx[335]
  PIN FREEZE_PMOS_NOSF[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5563.945 1046.435 5564.225 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[55]
  PIN BcidMtx[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5562.825 1046.435 5563.105 1047.435 ;
    END
  END BcidMtx[332]
  PIN Data_PMOS_NOSF[1158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5559.465 1046.435 5559.745 1047.435 ;
    END
  END Data_PMOS_NOSF[1158]
  PIN Data_PMOS_NOSF[1170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5557.785 1046.435 5558.065 1047.435 ;
    END
  END Data_PMOS_NOSF[1170]
  PIN Data_PMOS_NOSF[1159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5556.665 1046.435 5556.945 1047.435 ;
    END
  END Data_PMOS_NOSF[1159]
  PIN Data_PMOS_NOSF[1155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5554.425 1046.435 5554.705 1047.435 ;
    END
  END Data_PMOS_NOSF[1155]
  PIN MASKH[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5514.105 1046.435 5514.385 1047.435 ;
    END
  END MASKH[55]
  PIN DIG_MON_PMOS_NOSF[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5512.425 1046.435 5512.705 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[110]
  PIN MASKD[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5509.065 1046.435 5509.345 1047.435 ;
    END
  END MASKD[109]
  PIN MASKV[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5506.265 1046.435 5506.545 1047.435 ;
    END
  END MASKV[109]
  PIN Data_PMOS_NOSF[1142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5505.145 1046.435 5505.425 1047.435 ;
    END
  END Data_PMOS_NOSF[1142]
  PIN Data_PMOS_NOSF[1147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5502.905 1046.435 5503.185 1047.435 ;
    END
  END Data_PMOS_NOSF[1147]
  PIN Data_PMOS_NOSF[1141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5501.225 1046.435 5501.505 1047.435 ;
    END
  END Data_PMOS_NOSF[1141]
  PIN INJ_IN[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5491.145 1046.435 5491.425 1047.435 ;
    END
  END INJ_IN[109]
  PIN BcidMtx[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5487.785 1046.435 5488.065 1047.435 ;
    END
  END BcidMtx[327]
  PIN BcidMtx[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5486.105 1046.435 5486.385 1047.435 ;
    END
  END BcidMtx[326]
  PIN BcidMtx[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5484.985 1046.435 5485.265 1047.435 ;
    END
  END BcidMtx[324]
  PIN Data_PMOS_NOSF[1143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5479.665 1046.435 5479.945 1047.435 ;
    END
  END Data_PMOS_NOSF[1143]
  PIN Data_PMOS_NOSF[1138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5452.505 1046.435 5452.785 1047.435 ;
    END
  END Data_PMOS_NOSF[1138]
  PIN Data_PMOS_NOSF[1145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5451.385 1046.435 5451.665 1047.435 ;
    END
  END Data_PMOS_NOSF[1145]
  PIN MASKV[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5449.145 1046.435 5449.425 1047.435 ;
    END
  END MASKV[108]
  PIN DIG_MON_PMOS_NOSF[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5446.905 1046.435 5447.185 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[108]
  PIN DIG_MON_SEL[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5445.225 1046.435 5445.505 1047.435 ;
    END
  END DIG_MON_SEL[108]
  PIN INJ_ROW[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5441.305 1046.435 5441.585 1047.435 ;
    END
  END INJ_ROW[53]
  PIN Data_PMOS_NOSF[1121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5439.625 1046.435 5439.905 1047.435 ;
    END
  END Data_PMOS_NOSF[1121]
  PIN Data_PMOS_NOSF[1132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5425.625 1046.435 5425.905 1047.435 ;
    END
  END Data_PMOS_NOSF[1132]
  PIN DIG_MON_SEL[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18648.345 1046.435 18648.625 1047.435 ;
    END
  END DIG_MON_SEL[438]
  PIN Data_PMOS_NOSF[1120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5422.825 1046.435 5423.105 1047.435 ;
    END
  END Data_PMOS_NOSF[1120]
  PIN INJ_IN[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5421.145 1046.435 5421.425 1047.435 ;
    END
  END INJ_IN[107]
  PIN BcidMtx[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5417.785 1046.435 5418.065 1047.435 ;
    END
  END BcidMtx[321]
  PIN BcidMtx[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5416.105 1046.435 5416.385 1047.435 ;
    END
  END BcidMtx[320]
  PIN BcidMtx[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5414.985 1046.435 5415.265 1047.435 ;
    END
  END BcidMtx[318]
  PIN Data_PMOS_NOSF[1122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5372.985 1046.435 5373.265 1047.435 ;
    END
  END Data_PMOS_NOSF[1122]
  PIN Data_PMOS_NOSF[1117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5371.305 1046.435 5371.585 1047.435 ;
    END
  END Data_PMOS_NOSF[1117]
  PIN Data_PMOS_NOSF[1124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5370.185 1046.435 5370.465 1047.435 ;
    END
  END Data_PMOS_NOSF[1124]
  PIN MASKV[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5367.945 1046.435 5368.225 1047.435 ;
    END
  END MASKV[106]
  PIN DIG_MON_PMOS_NOSF[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5365.705 1046.435 5365.985 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[106]
  PIN DIG_MON_SEL[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5364.025 1046.435 5364.305 1047.435 ;
    END
  END DIG_MON_SEL[106]
  PIN INJ_ROW[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5351.705 1046.435 5351.985 1047.435 ;
    END
  END INJ_ROW[52]
  PIN Data_PMOS_NOSF[1100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5350.025 1046.435 5350.305 1047.435 ;
    END
  END Data_PMOS_NOSF[1100]
  PIN Data_PMOS_NOSF[1111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5348.905 1046.435 5349.185 1047.435 ;
    END
  END Data_PMOS_NOSF[1111]
  PIN Data_PMOS_NOSF[1106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5346.665 1046.435 5346.945 1047.435 ;
    END
  END Data_PMOS_NOSF[1106]
  PIN INJ_IN[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5342.465 1046.435 5342.745 1047.435 ;
    END
  END INJ_IN[105]
  PIN BcidMtx[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5340.225 1046.435 5340.505 1047.435 ;
    END
  END BcidMtx[317]
  PIN BcidMtx[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5311.945 1046.435 5312.225 1047.435 ;
    END
  END BcidMtx[314]
  PIN INJ_IN[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5309.705 1046.435 5309.985 1047.435 ;
    END
  END INJ_IN[104]
  PIN Data_PMOS_NOSF[1094]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5308.025 1046.435 5308.305 1047.435 ;
    END
  END Data_PMOS_NOSF[1094]
  PIN Data_PMOS_NOSF[1096]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5305.785 1046.435 5306.065 1047.435 ;
    END
  END Data_PMOS_NOSF[1096]
  PIN Data_PMOS_NOSF[1093]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5304.105 1046.435 5304.385 1047.435 ;
    END
  END Data_PMOS_NOSF[1093]
  PIN Data_PMOS_NOSF[1109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5302.985 1046.435 5303.265 1047.435 ;
    END
  END Data_PMOS_NOSF[1109]
  PIN DIG_MON_PMOS_NOSF[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5300.185 1046.435 5300.465 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[104]
  PIN DIG_MON_SEL[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5285.065 1046.435 5285.345 1047.435 ;
    END
  END DIG_MON_SEL[103]
  PIN DIG_MON_PMOS_NOSF[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5282.825 1046.435 5283.105 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[103]
  PIN Data_PMOS_NOSF[1079]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5280.025 1046.435 5280.305 1047.435 ;
    END
  END Data_PMOS_NOSF[1079]
  PIN Data_PMOS_NOSF[1076]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5278.345 1046.435 5278.625 1047.435 ;
    END
  END Data_PMOS_NOSF[1076]
  PIN Data_PMOS_NOSF[1091]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5277.225 1046.435 5277.505 1047.435 ;
    END
  END Data_PMOS_NOSF[1091]
  PIN INJ_IN[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5274.425 1046.435 5274.705 1047.435 ;
    END
  END INJ_IN[103]
  PIN BcidMtx[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5232.425 1046.435 5232.705 1047.435 ;
    END
  END BcidMtx[310]
  PIN Read_PMOS_NOSF[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5230.745 1046.435 5231.025 1047.435 ;
    END
  END Read_PMOS_NOSF[51]
  PIN BcidMtx[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5230.185 1046.435 5230.465 1047.435 ;
    END
  END BcidMtx[308]
  PIN INJ_IN[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5227.945 1046.435 5228.225 1047.435 ;
    END
  END INJ_IN[102]
  PIN Data_PMOS_NOSF[1080]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5225.705 1046.435 5225.985 1047.435 ;
    END
  END Data_PMOS_NOSF[1080]
  PIN Data_PMOS_NOSF[1075]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5224.025 1046.435 5224.305 1047.435 ;
    END
  END Data_PMOS_NOSF[1075]
  PIN Data_PMOS_NOSF[1072]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5222.345 1046.435 5222.625 1047.435 ;
    END
  END Data_PMOS_NOSF[1072]
  PIN MASKV[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5212.265 1046.435 5212.545 1047.435 ;
    END
  END MASKV[102]
  PIN DIG_MON_PMOS_NOSF[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5210.025 1046.435 5210.305 1047.435 ;
    END
  END DIG_MON_PMOS_NOSF[102]
  PIN Data_HV[1081]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18664.585 1046.435 18664.865 1047.435 ;
    END
  END Data_HV[1081]
  PIN DIG_MON_SEL[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5207.785 1046.435 5208.065 1047.435 ;
    END
  END DIG_MON_SEL[101]
  PIN INJ_ROW[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5202.465 1046.435 5202.745 1047.435 ;
    END
  END INJ_ROW[50]
  PIN Data_PMOS_NOSF[1058]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5200.785 1046.435 5201.065 1047.435 ;
    END
  END Data_PMOS_NOSF[1058]
  PIN Data_PMOS_NOSF[1055]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5199.105 1046.435 5199.385 1047.435 ;
    END
  END Data_PMOS_NOSF[1055]
  PIN Data_PMOS_NOSF[1064]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5171.945 1046.435 5172.225 1047.435 ;
    END
  END Data_PMOS_NOSF[1064]
  PIN INJ_IN[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5169.705 1046.435 5169.985 1047.435 ;
    END
  END INJ_IN[101]
  PIN BcidMtx[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5166.905 1046.435 5167.185 1047.435 ;
    END
  END BcidMtx[304]
  PIN Read_PMOS_NOSF[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5165.225 1046.435 5165.505 1047.435 ;
    END
  END Read_PMOS_NOSF[50]
  PIN BcidMtx[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5163.545 1046.435 5163.825 1047.435 ;
    END
  END BcidMtx[300]
  PIN Data_PMOS_NOSF[1052]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5160.745 1046.435 5161.025 1047.435 ;
    END
  END Data_PMOS_NOSF[1052]
  PIN Data_PMOS_NOSF[1060]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5146.185 1046.435 5146.465 1047.435 ;
    END
  END Data_PMOS_NOSF[1060]
  PIN Data_PMOS_NOSF[1061]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5144.505 1046.435 5144.785 1047.435 ;
    END
  END Data_PMOS_NOSF[1061]
  PIN Data_PMOS_NOSF[1067]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5142.825 1046.435 5143.105 1047.435 ;
    END
  END Data_PMOS_NOSF[1067]
  PIN MASKD[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5141.145 1046.435 5141.425 1047.435 ;
    END
  END MASKD[100]
  PIN DIG_MON_SEL[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5138.345 1046.435 5138.625 1047.435 ;
    END
  END DIG_MON_SEL[100]
  PIN nTOK_HV[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18860.025 1046.435 18860.305 1047.435 ;
    END
  END nTOK_HV[53]
  PIN INJ_ROW[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5134.425 1046.435 5134.705 1047.435 ;
    END
  END INJ_ROW[49]
  PIN Data_PMOS_NOSF[1037]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5092.985 1046.435 5093.265 1047.435 ;
    END
  END Data_PMOS_NOSF[1037]
  PIN Data_PMOS_NOSF[1034]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5091.305 1046.435 5091.585 1047.435 ;
    END
  END Data_PMOS_NOSF[1034]
  PIN Data_PMOS_NOSF[1043]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5089.625 1046.435 5089.905 1047.435 ;
    END
  END Data_PMOS_NOSF[1043]
  PIN INJ_IN[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5087.385 1046.435 5087.665 1047.435 ;
    END
  END INJ_IN[99]
  PIN BcidMtx[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5084.585 1046.435 5084.865 1047.435 ;
    END
  END BcidMtx[298]
  PIN Read_PMOS_NOSF[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5082.905 1046.435 5083.185 1047.435 ;
    END
  END Read_PMOS_NOSF[49]
  PIN INJ_IN[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5071.705 1046.435 5071.985 1047.435 ;
    END
  END INJ_IN[98]
  PIN Data_PMOS_NOSF[1038]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5069.465 1046.435 5069.745 1047.435 ;
    END
  END Data_PMOS_NOSF[1038]
  PIN Data_PMOS_NOSF[1039]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5068.345 1046.435 5068.625 1047.435 ;
    END
  END Data_PMOS_NOSF[1039]
  PIN Data_PMOS_NOSF[1030]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5066.105 1046.435 5066.385 1047.435 ;
    END
  END Data_PMOS_NOSF[1030]
  PIN MASKV[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5062.465 1046.435 5062.745 1047.435 ;
    END
  END MASKV[98]
  PIN MASKD[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5061.345 1046.435 5061.625 1047.435 ;
    END
  END MASKD[98]
  PIN FREEZE_PMOS_NOSF[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5313.065 1046.435 5313.345 1047.435 ;
    END
  END FREEZE_PMOS_NOSF[52]
  PIN INJ_ROW[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7268.585 1046.435 7268.865 1047.435 ;
    END
  END INJ_ROW[76]
  PIN Data_PMOS[428]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7266.905 1046.435 7267.185 1047.435 ;
    END
  END Data_PMOS[428]
  PIN Data_PMOS[425]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7265.225 1046.435 7265.505 1047.435 ;
    END
  END Data_PMOS[425]
  PIN Data_PMOS[434]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7263.545 1046.435 7263.825 1047.435 ;
    END
  END Data_PMOS[434]
  PIN INJ_IN[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7261.305 1046.435 7261.585 1047.435 ;
    END
  END INJ_IN[153]
  PIN BcidMtx[460]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7245.065 1046.435 7245.345 1047.435 ;
    END
  END BcidMtx[460]
  PIN Read_PMOS[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7243.385 1046.435 7243.665 1047.435 ;
    END
  END Read_PMOS[20]
  PIN BcidMtx[456]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7241.705 1046.435 7241.985 1047.435 ;
    END
  END BcidMtx[456]
  PIN Data_PMOS[422]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7238.905 1046.435 7239.185 1047.435 ;
    END
  END Data_PMOS[422]
  PIN Data_PMOS[430]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7237.225 1046.435 7237.505 1047.435 ;
    END
  END Data_PMOS[430]
  PIN Data_PMOS[431]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7235.545 1046.435 7235.825 1047.435 ;
    END
  END Data_PMOS[431]
  PIN Data_PMOS[437]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7233.865 1046.435 7234.145 1047.435 ;
    END
  END Data_PMOS[437]
  PIN MASKD[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7193.545 1046.435 7193.825 1047.435 ;
    END
  END MASKD[152]
  PIN DIG_MON_SEL[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7190.745 1046.435 7191.025 1047.435 ;
    END
  END DIG_MON_SEL[152]
  PIN DIG_MON_PMOS[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7187.945 1046.435 7188.225 1047.435 ;
    END
  END DIG_MON_PMOS[39]
  PIN Data_PMOS[417]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7185.705 1046.435 7185.985 1047.435 ;
    END
  END Data_PMOS[417]
  PIN Data_PMOS[418]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7184.025 1046.435 7184.305 1047.435 ;
    END
  END Data_PMOS[418]
  PIN Data_PMOS[419]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7182.345 1046.435 7182.625 1047.435 ;
    END
  END Data_PMOS[419]
  PIN Data_PMOS[405]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7172.265 1046.435 7172.545 1047.435 ;
    END
  END Data_PMOS[405]
  PIN BcidMtx[455]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7168.905 1046.435 7169.185 1047.435 ;
    END
  END BcidMtx[455]
  PIN FREEZE_PMOS[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7167.225 1046.435 7167.505 1047.435 ;
    END
  END FREEZE_PMOS[19]
  PIN BcidMtx[451]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7165.545 1046.435 7165.825 1047.435 ;
    END
  END BcidMtx[451]
  PIN Data_PMOS[402]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7160.785 1046.435 7161.065 1047.435 ;
    END
  END Data_PMOS[402]
  PIN Data_PMOS[414]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7159.105 1046.435 7159.385 1047.435 ;
    END
  END Data_PMOS[414]
  PIN Data_PMOS[415]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7131.945 1046.435 7132.225 1047.435 ;
    END
  END Data_PMOS[415]
  PIN Data_PMOS[400]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7130.825 1046.435 7131.105 1047.435 ;
    END
  END Data_PMOS[400]
  PIN MASKV[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7129.145 1046.435 7129.425 1047.435 ;
    END
  END MASKV[150]
  PIN DIG_MON_PMOS[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7126.905 1046.435 7127.185 1047.435 ;
    END
  END DIG_MON_PMOS[38]
  PIN DIG_MON_SEL[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7124.665 1046.435 7124.945 1047.435 ;
    END
  END DIG_MON_SEL[149]
  PIN INJ_ROW[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7121.305 1046.435 7121.585 1047.435 ;
    END
  END INJ_ROW[74]
  PIN Data_PMOS[386]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7119.625 1046.435 7119.905 1047.435 ;
    END
  END Data_PMOS[386]
  PIN Data_PMOS[383]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7105.065 1046.435 7105.345 1047.435 ;
    END
  END Data_PMOS[383]
  PIN Data_PMOS[392]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7103.385 1046.435 7103.665 1047.435 ;
    END
  END Data_PMOS[392]
  PIN INJ_IN[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7101.145 1046.435 7101.425 1047.435 ;
    END
  END INJ_IN[149]
  PIN BcidMtx[448]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7098.345 1046.435 7098.625 1047.435 ;
    END
  END BcidMtx[448]
  PIN Read_PMOS[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7096.665 1046.435 7096.945 1047.435 ;
    END
  END Read_PMOS[18]
  PIN BcidMtx[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7094.985 1046.435 7095.265 1047.435 ;
    END
  END BcidMtx[444]
  PIN Data_PMOS[380]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7053.545 1046.435 7053.825 1047.435 ;
    END
  END Data_PMOS[380]
  PIN Data_PMOS[388]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7051.865 1046.435 7052.145 1047.435 ;
    END
  END Data_PMOS[388]
  PIN Data_PMOS[389]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7050.185 1046.435 7050.465 1047.435 ;
    END
  END Data_PMOS[389]
  PIN Data_PMOS[395]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7048.505 1046.435 7048.785 1047.435 ;
    END
  END Data_PMOS[395]
  PIN MASKD[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7046.825 1046.435 7047.105 1047.435 ;
    END
  END MASKD[148]
  PIN DIG_MON_SEL[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7044.025 1046.435 7044.305 1047.435 ;
    END
  END DIG_MON_SEL[148]
  PIN DIG_MON_PMOS[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7041.225 1046.435 7041.505 1047.435 ;
    END
  END DIG_MON_PMOS[35]
  PIN Data_PMOS[375]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7030.585 1046.435 7030.865 1047.435 ;
    END
  END Data_PMOS[375]
  PIN Data_PMOS[376]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7028.905 1046.435 7029.185 1047.435 ;
    END
  END Data_PMOS[376]
  PIN Data_PMOS[377]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7027.225 1046.435 7027.505 1047.435 ;
    END
  END Data_PMOS[377]
  PIN Data_PMOS[363]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7025.545 1046.435 7025.825 1047.435 ;
    END
  END Data_PMOS[363]
  PIN BcidMtx[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7020.225 1046.435 7020.505 1047.435 ;
    END
  END BcidMtx[443]
  PIN Read_PMOS[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6992.505 1046.435 6992.785 1047.435 ;
    END
  END Read_PMOS[17]
  PIN BcidMtx[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6990.825 1046.435 6991.105 1047.435 ;
    END
  END BcidMtx[438]
  PIN Data_PMOS[359]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6988.025 1046.435 6988.305 1047.435 ;
    END
  END Data_PMOS[359]
  PIN Data_PMOS[367]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6986.345 1046.435 6986.625 1047.435 ;
    END
  END Data_PMOS[367]
  PIN Data_PMOS[368]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6984.665 1046.435 6984.945 1047.435 ;
    END
  END Data_PMOS[368]
  PIN Data_PMOS[374]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6982.985 1046.435 6983.265 1047.435 ;
    END
  END Data_PMOS[374]
  PIN MASKD[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6981.305 1046.435 6981.585 1047.435 ;
    END
  END MASKD[146]
  PIN DIG_MON_SEL[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6965.625 1046.435 6965.905 1047.435 ;
    END
  END DIG_MON_SEL[146]
  PIN DIG_MON_PMOS[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6962.825 1046.435 6963.105 1047.435 ;
    END
  END DIG_MON_PMOS[33]
  PIN Data_PMOS[354]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6960.585 1046.435 6960.865 1047.435 ;
    END
  END Data_PMOS[354]
  PIN Data_PMOS[355]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6958.905 1046.435 6959.185 1047.435 ;
    END
  END Data_PMOS[355]
  PIN Data_PMOS[356]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6957.225 1046.435 6957.505 1047.435 ;
    END
  END Data_PMOS[356]
  PIN Data_PMOS[342]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6955.545 1046.435 6955.825 1047.435 ;
    END
  END Data_PMOS[342]
  PIN BcidMtx[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6912.985 1046.435 6913.265 1047.435 ;
    END
  END BcidMtx[437]
  PIN FREEZE_PMOS[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6911.305 1046.435 6911.585 1047.435 ;
    END
  END FREEZE_PMOS[16]
  PIN BcidMtx[1326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18854.985 1046.435 18855.265 1047.435 ;
    END
  END BcidMtx[1326]
  PIN INJ_IN[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6907.945 1046.435 6908.225 1047.435 ;
    END
  END INJ_IN[144]
  PIN Data_PMOS[345]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6905.705 1046.435 6905.985 1047.435 ;
    END
  END Data_PMOS[345]
  PIN Data_PMOS[340]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6904.025 1046.435 6904.305 1047.435 ;
    END
  END Data_PMOS[340]
  PIN Data_PMOS[337]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6902.345 1046.435 6902.625 1047.435 ;
    END
  END Data_PMOS[337]
  PIN MASKV[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6892.265 1046.435 6892.545 1047.435 ;
    END
  END MASKV[144]
  PIN DIG_MON_PMOS[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6890.025 1046.435 6890.305 1047.435 ;
    END
  END DIG_MON_PMOS[32]
  PIN DIG_MON_SEL[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6887.785 1046.435 6888.065 1047.435 ;
    END
  END DIG_MON_SEL[143]
  PIN DIG_MON_PMOS[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6885.545 1046.435 6885.825 1047.435 ;
    END
  END DIG_MON_PMOS[31]
  PIN Data_PMOS[333]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6881.345 1046.435 6881.625 1047.435 ;
    END
  END Data_PMOS[333]
  PIN Data_PMOS[320]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6879.105 1046.435 6879.385 1047.435 ;
    END
  END Data_PMOS[320]
  PIN Data_PMOS[329]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6851.945 1046.435 6852.225 1047.435 ;
    END
  END Data_PMOS[329]
  PIN INJ_IN[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6849.705 1046.435 6849.985 1047.435 ;
    END
  END INJ_IN[143]
  PIN BcidMtx[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6847.465 1046.435 6847.745 1047.435 ;
    END
  END BcidMtx[431]
  PIN FREEZE_PMOS[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6845.785 1046.435 6846.065 1047.435 ;
    END
  END FREEZE_PMOS[15]
  PIN BcidMtx[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6844.105 1046.435 6844.385 1047.435 ;
    END
  END BcidMtx[427]
  PIN Data_PMOS[318]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6841.305 1046.435 6841.585 1047.435 ;
    END
  END Data_PMOS[318]
  PIN Data_PMOS[330]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6826.745 1046.435 6827.025 1047.435 ;
    END
  END Data_PMOS[330]
  PIN Data_PMOS[331]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6825.065 1046.435 6825.345 1047.435 ;
    END
  END Data_PMOS[331]
  PIN Data_PMOS[315]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6823.385 1046.435 6823.665 1047.435 ;
    END
  END Data_PMOS[315]
  PIN MASKH[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6821.705 1046.435 6821.985 1047.435 ;
    END
  END MASKH[71]
  PIN MASKD[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6816.665 1046.435 6816.945 1047.435 ;
    END
  END MASKD[141]
  PIN MASKV[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6813.865 1046.435 6814.145 1047.435 ;
    END
  END MASKV[141]
  PIN Data_PMOS[306]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6772.425 1046.435 6772.705 1047.435 ;
    END
  END Data_PMOS[306]
  PIN Data_PMOS[307]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6770.745 1046.435 6771.025 1047.435 ;
    END
  END Data_PMOS[307]
  PIN Data_PMOS[301]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6769.065 1046.435 6769.345 1047.435 ;
    END
  END Data_PMOS[301]
  PIN nTOK_PMOS[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6766.265 1046.435 6766.545 1047.435 ;
    END
  END nTOK_PMOS[14]
  PIN BcidMtx[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6764.025 1046.435 6764.305 1047.435 ;
    END
  END BcidMtx[423]
  PIN BcidMtx[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6762.345 1046.435 6762.625 1047.435 ;
    END
  END BcidMtx[422]
  PIN Data_HV[1122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18812.985 1046.435 18813.265 1047.435 ;
    END
  END Data_HV[1122]
  PIN Data_PMOS[296]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6750.025 1046.435 6750.305 1047.435 ;
    END
  END Data_PMOS[296]
  PIN Data_PMOS[304]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6748.345 1046.435 6748.625 1047.435 ;
    END
  END Data_PMOS[304]
  PIN Data_PMOS[310]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6747.225 1046.435 6747.505 1047.435 ;
    END
  END Data_PMOS[310]
  PIN Data_PMOS[294]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6745.545 1046.435 6745.825 1047.435 ;
    END
  END Data_PMOS[294]
  PIN MASKH[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6741.905 1046.435 6742.185 1047.435 ;
    END
  END MASKH[70]
  PIN DIG_MON_SEL[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7831.945 1046.435 7832.225 1047.435 ;
    END
  END DIG_MON_SEL[167]
  PIN Data_COMP[194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10878.345 1046.435 10878.625 1047.435 ;
    END
  END Data_COMP[194]
  PIN Data_COMP[195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10875.545 1046.435 10875.825 1047.435 ;
    END
  END Data_COMP[195]
  PIN INJ_IN[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10874.425 1046.435 10874.705 1047.435 ;
    END
  END INJ_IN[243]
  PIN BcidMtx[730]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10832.425 1046.435 10832.705 1047.435 ;
    END
  END BcidMtx[730]
  PIN BcidMtx[727]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10829.625 1046.435 10829.905 1047.435 ;
    END
  END BcidMtx[727]
  PIN BcidMtx[726]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10829.065 1046.435 10829.345 1047.435 ;
    END
  END BcidMtx[726]
  PIN Data_COMP[192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10826.825 1046.435 10827.105 1047.435 ;
    END
  END Data_COMP[192]
  PIN Data_COMP[199]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10824.585 1046.435 10824.865 1047.435 ;
    END
  END Data_COMP[199]
  PIN Data_COMP[193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10824.025 1046.435 10824.305 1047.435 ;
    END
  END Data_COMP[193]
  PIN Data_COMP[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10822.345 1046.435 10822.625 1047.435 ;
    END
  END Data_COMP[190]
  PIN MASKD[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10811.145 1046.435 10811.425 1047.435 ;
    END
  END MASKD[242]
  PIN DIG_MON_COMP[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10810.025 1046.435 10810.305 1047.435 ;
    END
  END DIG_MON_COMP[18]
  PIN DIG_MON_SEL[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10807.785 1046.435 10808.065 1047.435 ;
    END
  END DIG_MON_SEL[241]
  PIN Data_COMP[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10801.345 1046.435 10801.625 1047.435 ;
    END
  END Data_COMP[186]
  PIN Data_COMP[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10800.785 1046.435 10801.065 1047.435 ;
    END
  END Data_COMP[176]
  PIN Data_COMP[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10799.105 1046.435 10799.385 1047.435 ;
    END
  END Data_COMP[173]
  PIN Data_COMP[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10770.825 1046.435 10771.105 1047.435 ;
    END
  END Data_COMP[174]
  PIN INJ_IN[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10769.705 1046.435 10769.985 1047.435 ;
    END
  END INJ_IN[241]
  PIN BcidMtx[724]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10766.905 1046.435 10767.185 1047.435 ;
    END
  END BcidMtx[724]
  PIN BcidMtx[721]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10764.105 1046.435 10764.385 1047.435 ;
    END
  END BcidMtx[721]
  PIN BcidMtx[720]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10763.545 1046.435 10763.825 1047.435 ;
    END
  END BcidMtx[720]
  PIN Data_COMP[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10761.305 1046.435 10761.585 1047.435 ;
    END
  END Data_COMP[171]
  PIN Data_COMP[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10745.625 1046.435 10745.905 1047.435 ;
    END
  END Data_COMP[172]
  PIN Data_COMP[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10745.065 1046.435 10745.345 1047.435 ;
    END
  END Data_COMP[184]
  PIN Data_COMP[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10744.505 1046.435 10744.785 1047.435 ;
    END
  END Data_COMP[179]
  PIN MASKH[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10741.705 1046.435 10741.985 1047.435 ;
    END
  END MASKH[120]
  PIN MASKD[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10741.145 1046.435 10741.425 1047.435 ;
    END
  END MASKD[240]
  PIN DIG_MON_SEL[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10738.345 1046.435 10738.625 1047.435 ;
    END
  END DIG_MON_SEL[240]
  PIN MASKV[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10733.865 1046.435 10734.145 1047.435 ;
    END
  END MASKV[239]
  PIN Data_COMP[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10693.545 1046.435 10693.825 1047.435 ;
    END
  END Data_COMP[165]
  PIN Data_COMP[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10691.865 1046.435 10692.145 1047.435 ;
    END
  END Data_COMP[166]
  PIN Data_COMP[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10689.065 1046.435 10689.345 1047.435 ;
    END
  END Data_COMP[154]
  PIN Data_COMP[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10688.505 1046.435 10688.785 1047.435 ;
    END
  END Data_COMP[153]
  PIN BcidMtx[719]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10685.145 1046.435 10685.425 1047.435 ;
    END
  END BcidMtx[719]
  PIN BcidMtx[716]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10682.345 1046.435 10682.625 1047.435 ;
    END
  END BcidMtx[716]
  PIN BcidMtx[715]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10681.785 1046.435 10682.065 1047.435 ;
    END
  END BcidMtx[715]
  PIN Data_COMP[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10670.585 1046.435 10670.865 1047.435 ;
    END
  END Data_COMP[150]
  PIN Data_COMP[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10667.785 1046.435 10668.065 1047.435 ;
    END
  END Data_COMP[151]
  PIN Data_COMP[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10667.225 1046.435 10667.505 1047.435 ;
    END
  END Data_COMP[163]
  PIN Data_COMP[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10665.545 1046.435 10665.825 1047.435 ;
    END
  END Data_COMP[147]
  PIN DIG_MON_COMP[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10660.225 1046.435 10660.505 1047.435 ;
    END
  END DIG_MON_COMP[14]
  PIN DIG_MON_SEL[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11751.945 1046.435 11752.225 1047.435 ;
    END
  END DIG_MON_SEL[265]
  PIN Data_COMP[438]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11747.465 1046.435 11747.745 1047.435 ;
    END
  END Data_COMP[438]
  PIN Data_COMP[428]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11746.905 1046.435 11747.185 1047.435 ;
    END
  END Data_COMP[428]
  PIN Data_COMP[425]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11745.225 1046.435 11745.505 1047.435 ;
    END
  END Data_COMP[425]
  PIN Data_COMP[426]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11742.425 1046.435 11742.705 1047.435 ;
    END
  END Data_COMP[426]
  PIN INJ_IN[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11741.305 1046.435 11741.585 1047.435 ;
    END
  END INJ_IN[265]
  PIN BcidMtx[796]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11725.065 1046.435 11725.345 1047.435 ;
    END
  END BcidMtx[796]
  PIN BcidMtx[793]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11722.265 1046.435 11722.545 1047.435 ;
    END
  END BcidMtx[793]
  PIN BcidMtx[792]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11721.705 1046.435 11721.985 1047.435 ;
    END
  END BcidMtx[792]
  PIN Data_COMP[422]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11718.905 1046.435 11719.185 1047.435 ;
    END
  END Data_COMP[422]
  PIN Data_COMP[436]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11716.105 1046.435 11716.385 1047.435 ;
    END
  END Data_COMP[436]
  PIN Data_COMP[431]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11715.545 1046.435 11715.825 1047.435 ;
    END
  END Data_COMP[431]
  PIN Data_COMP[437]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11713.865 1046.435 11714.145 1047.435 ;
    END
  END Data_COMP[437]
  PIN DIG_MON_SEL[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11670.745 1046.435 11671.025 1047.435 ;
    END
  END DIG_MON_SEL[264]
  PIN DIG_MON_COMP[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11667.945 1046.435 11668.225 1047.435 ;
    END
  END DIG_MON_COMP[39]
  PIN Data_COMP[411]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11664.585 1046.435 11664.865 1047.435 ;
    END
  END Data_COMP[411]
  PIN Data_COMP[418]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11664.025 1046.435 11664.305 1047.435 ;
    END
  END Data_COMP[418]
  PIN Data_COMP[419]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11662.345 1046.435 11662.625 1047.435 ;
    END
  END Data_COMP[419]
  PIN nTOK_COMP[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11650.025 1046.435 11650.305 1047.435 ;
    END
  END nTOK_COMP[19]
  PIN BcidMtx[791]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11648.905 1046.435 11649.185 1047.435 ;
    END
  END BcidMtx[791]
  PIN FREEZE_COMP[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11647.225 1046.435 11647.505 1047.435 ;
    END
  END FREEZE_COMP[19]
  PIN INJ_IN[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11641.905 1046.435 11642.185 1047.435 ;
    END
  END INJ_IN[262]
  PIN Data_COMP[402]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11640.785 1046.435 11641.065 1047.435 ;
    END
  END Data_COMP[402]
  PIN Data_COMP[414]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11639.105 1046.435 11639.385 1047.435 ;
    END
  END Data_COMP[414]
  PIN Data_COMP[400]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11610.825 1046.435 11611.105 1047.435 ;
    END
  END Data_COMP[400]
  PIN Data_COMP[399]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11610.265 1046.435 11610.545 1047.435 ;
    END
  END Data_COMP[399]
  PIN MASKH[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11608.585 1046.435 11608.865 1047.435 ;
    END
  END MASKH[131]
  PIN DIG_MON_SEL[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11604.665 1046.435 11604.945 1047.435 ;
    END
  END DIG_MON_SEL[261]
  PIN MASKD[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11603.545 1046.435 11603.825 1047.435 ;
    END
  END MASKD[261]
  PIN MASKV[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11600.745 1046.435 11601.025 1047.435 ;
    END
  END MASKV[261]
  PIN Data_COMP[383]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11585.065 1046.435 11585.345 1047.435 ;
    END
  END Data_COMP[383]
  PIN Data_COMP[391]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11584.505 1046.435 11584.785 1047.435 ;
    END
  END Data_COMP[391]
  PIN Data_COMP[385]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11582.825 1046.435 11583.105 1047.435 ;
    END
  END Data_COMP[385]
  PIN BcidMtx[784]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11578.345 1046.435 11578.625 1047.435 ;
    END
  END BcidMtx[784]
  PIN BcidMtx[783]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11577.785 1046.435 11578.065 1047.435 ;
    END
  END BcidMtx[783]
  PIN BcidMtx[782]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11576.105 1046.435 11576.385 1047.435 ;
    END
  END BcidMtx[782]
  PIN Data_COMP[380]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11533.545 1046.435 11533.825 1047.435 ;
    END
  END Data_COMP[380]
  PIN Data_COMP[387]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11532.985 1046.435 11533.265 1047.435 ;
    END
  END Data_COMP[387]
  PIN Data_COMP[382]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11531.305 1046.435 11531.585 1047.435 ;
    END
  END Data_COMP[382]
  PIN Data_COMP[395]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11528.505 1046.435 11528.785 1047.435 ;
    END
  END Data_COMP[395]
  PIN MASKV[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11527.945 1046.435 11528.225 1047.435 ;
    END
  END MASKV[260]
  PIN DIG_MON_COMP[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11525.705 1046.435 11525.985 1047.435 ;
    END
  END DIG_MON_COMP[36]
  PIN DIG_MON_COMP[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11521.225 1046.435 11521.505 1047.435 ;
    END
  END DIG_MON_COMP[35]
  PIN INJ_ROW[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11511.705 1046.435 11511.985 1047.435 ;
    END
  END INJ_ROW[129]
  PIN Data_COMP[365]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11510.025 1046.435 11510.305 1047.435 ;
    END
  END Data_COMP[365]
  PIN Data_COMP[377]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11507.225 1046.435 11507.505 1047.435 ;
    END
  END Data_COMP[377]
  PIN Data_COMP[371]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11506.665 1046.435 11506.945 1047.435 ;
    END
  END Data_COMP[371]
  PIN INJ_IN[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11502.465 1046.435 11502.745 1047.435 ;
    END
  END INJ_IN[259]
  PIN Read_COMP[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11472.505 1046.435 11472.785 1047.435 ;
    END
  END Read_COMP[17]
  PIN BcidMtx[776]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11471.945 1046.435 11472.225 1047.435 ;
    END
  END BcidMtx[776]
  PIN INJ_IN[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11469.705 1046.435 11469.985 1047.435 ;
    END
  END INJ_IN[258]
  PIN Data_COMP[367]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11466.345 1046.435 11466.625 1047.435 ;
    END
  END Data_COMP[367]
  PIN Data_COMP[361]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11465.785 1046.435 11466.065 1047.435 ;
    END
  END Data_COMP[361]
  PIN Data_COMP[358]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11464.105 1046.435 11464.385 1047.435 ;
    END
  END Data_COMP[358]
  PIN MASKD[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11461.305 1046.435 11461.585 1047.435 ;
    END
  END MASKD[258]
  PIN DIG_MON_COMP[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11460.185 1046.435 11460.465 1047.435 ;
    END
  END DIG_MON_COMP[34]
  PIN DIG_MON_SEL[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11445.065 1046.435 11445.345 1047.435 ;
    END
  END DIG_MON_SEL[257]
  PIN Data_COMP[354]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11440.585 1046.435 11440.865 1047.435 ;
    END
  END Data_COMP[354]
  PIN Data_COMP[344]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11440.025 1046.435 11440.305 1047.435 ;
    END
  END Data_COMP[344]
  PIN nRST[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 12418.905 1046.435 12419.185 1047.435 ;
    END
  END nRST[141]
  PIN nRST[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11858.905 1046.435 11859.185 1047.435 ;
    END
  END nRST[134]
  PIN nRST[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17458.905 1046.435 17459.185 1047.435 ;
    END
  END nRST[204]
  PIN nRST[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16898.905 1046.435 16899.185 1047.435 ;
    END
  END nRST[197]
  PIN nRST[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 9058.905 1046.435 9059.185 1047.435 ;
    END
  END nRST[99]
  PIN nRST[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 8498.905 1046.435 8499.185 1047.435 ;
    END
  END nRST[92]
  PIN nRST[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 11298.905 1046.435 11299.185 1047.435 ;
    END
  END nRST[127]
  PIN MASKD[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6710.825 1046.435 6711.105 1047.435 ;
    END
  END MASKD[139]
  PIN MASKV[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6708.025 1046.435 6708.305 1047.435 ;
    END
  END MASKV[139]
  PIN Data_PMOS[292]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6705.785 1046.435 6706.065 1047.435 ;
    END
  END Data_PMOS[292]
  PIN Data_PMOS[287]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6703.545 1046.435 6703.825 1047.435 ;
    END
  END Data_PMOS[287]
  PIN INJ_IN[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6701.305 1046.435 6701.585 1047.435 ;
    END
  END INJ_IN[139]
  PIN BcidMtx[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6685.065 1046.435 6685.345 1047.435 ;
    END
  END BcidMtx[418]
  PIN Read_PMOS[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6683.385 1046.435 6683.665 1047.435 ;
    END
  END Read_PMOS[13]
  PIN BcidMtx[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6681.705 1046.435 6681.985 1047.435 ;
    END
  END BcidMtx[414]
  PIN Data_PMOS[275]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6678.905 1046.435 6679.185 1047.435 ;
    END
  END Data_PMOS[275]
  PIN Data_PMOS[283]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6677.225 1046.435 6677.505 1047.435 ;
    END
  END Data_PMOS[283]
  PIN Data_PMOS[284]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6675.545 1046.435 6675.825 1047.435 ;
    END
  END Data_PMOS[284]
  PIN Data_PMOS[290]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6673.865 1046.435 6674.145 1047.435 ;
    END
  END Data_PMOS[290]
  PIN BcidMtx[1328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18856.105 1046.435 18856.385 1047.435 ;
    END
  END BcidMtx[1328]
  PIN MASKD[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6629.065 1046.435 6629.345 1047.435 ;
    END
  END MASKD[137]
  PIN MASKV[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6626.265 1046.435 6626.545 1047.435 ;
    END
  END MASKV[137]
  PIN Data_PMOS[264]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6624.585 1046.435 6624.865 1047.435 ;
    END
  END Data_PMOS[264]
  PIN Data_PMOS[265]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6622.905 1046.435 6623.185 1047.435 ;
    END
  END Data_PMOS[265]
  PIN Data_PMOS[259]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6621.225 1046.435 6621.505 1047.435 ;
    END
  END Data_PMOS[259]
  PIN nTOK_PMOS[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6610.025 1046.435 6610.305 1047.435 ;
    END
  END nTOK_PMOS[12]
  PIN BcidMtx[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6607.785 1046.435 6608.065 1047.435 ;
    END
  END BcidMtx[411]
  PIN BcidMtx[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6606.105 1046.435 6606.385 1047.435 ;
    END
  END BcidMtx[410]
  PIN INJ_IN[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6601.905 1046.435 6602.185 1047.435 ;
    END
  END INJ_IN[136]
  PIN Data_PMOS[261]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6599.665 1046.435 6599.945 1047.435 ;
    END
  END Data_PMOS[261]
  PIN Data_PMOS[256]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6572.505 1046.435 6572.785 1047.435 ;
    END
  END Data_PMOS[256]
  PIN Data_PMOS[253]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6570.825 1046.435 6571.105 1047.435 ;
    END
  END Data_PMOS[253]
  PIN MASKV[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6569.145 1046.435 6569.425 1047.435 ;
    END
  END MASKV[136]
  PIN DIG_MON_PMOS[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6566.905 1046.435 6567.185 1047.435 ;
    END
  END DIG_MON_PMOS[24]
  PIN DIG_MON_SEL[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6565.225 1046.435 6565.505 1047.435 ;
    END
  END DIG_MON_SEL[136]
  PIN DIG_MON_PMOS[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6562.425 1046.435 6562.705 1047.435 ;
    END
  END DIG_MON_PMOS[23]
  PIN Data_PMOS[249]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6560.185 1046.435 6560.465 1047.435 ;
    END
  END Data_PMOS[249]
  PIN Data_PMOS[250]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6545.625 1046.435 6545.905 1047.435 ;
    END
  END Data_PMOS[250]
  PIN Data_PMOS[251]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6543.945 1046.435 6544.225 1047.435 ;
    END
  END Data_PMOS[251]
  PIN Data_PMOS[237]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6542.265 1046.435 6542.545 1047.435 ;
    END
  END Data_PMOS[237]
  PIN BcidMtx[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6538.905 1046.435 6539.185 1047.435 ;
    END
  END BcidMtx[407]
  PIN BcidMtx[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6538.345 1046.435 6538.625 1047.435 ;
    END
  END BcidMtx[406]
  PIN BcidMtx[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6535.545 1046.435 6535.825 1047.435 ;
    END
  END BcidMtx[403]
  PIN Data_PMOS[234]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6494.105 1046.435 6494.385 1047.435 ;
    END
  END Data_PMOS[234]
  PIN Data_PMOS[246]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6492.425 1046.435 6492.705 1047.435 ;
    END
  END Data_PMOS[246]
  PIN Data_PMOS[247]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6490.745 1046.435 6491.025 1047.435 ;
    END
  END Data_PMOS[247]
  PIN Data_PMOS[231]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6489.065 1046.435 6489.345 1047.435 ;
    END
  END Data_PMOS[231]
  PIN MASKH[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6487.385 1046.435 6487.665 1047.435 ;
    END
  END MASKH[67]
  PIN MASKD[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6482.345 1046.435 6482.625 1047.435 ;
    END
  END MASKD[133]
  PIN MASKV[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6471.145 1046.435 6471.425 1047.435 ;
    END
  END MASKV[133]
  PIN Data_PMOS[222]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6469.465 1046.435 6469.745 1047.435 ;
    END
  END Data_PMOS[222]
  PIN Data_PMOS[223]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6467.785 1046.435 6468.065 1047.435 ;
    END
  END Data_PMOS[223]
  PIN Data_PMOS[217]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6466.105 1046.435 6466.385 1047.435 ;
    END
  END Data_PMOS[217]
  PIN nTOK_PMOS[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6461.345 1046.435 6461.625 1047.435 ;
    END
  END nTOK_PMOS[10]
  PIN BcidMtx[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6459.105 1046.435 6459.385 1047.435 ;
    END
  END BcidMtx[399]
  PIN BcidMtx[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6431.385 1046.435 6431.665 1047.435 ;
    END
  END BcidMtx[397]
  PIN Data_PMOS[213]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6428.585 1046.435 6428.865 1047.435 ;
    END
  END Data_PMOS[213]
  PIN Data_PMOS[225]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6426.905 1046.435 6427.185 1047.435 ;
    END
  END Data_PMOS[225]
  PIN Data_PMOS[226]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6425.225 1046.435 6425.505 1047.435 ;
    END
  END Data_PMOS[226]
  PIN Data_PMOS[210]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6423.545 1046.435 6423.825 1047.435 ;
    END
  END Data_PMOS[210]
  PIN MASKH[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6421.865 1046.435 6422.145 1047.435 ;
    END
  END MASKH[66]
  PIN MASKD[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6403.945 1046.435 6404.225 1047.435 ;
    END
  END MASKD[131]
  PIN MASKV[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6401.145 1046.435 6401.425 1047.435 ;
    END
  END MASKV[131]
  PIN Data_PMOS[201]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6399.465 1046.435 6399.745 1047.435 ;
    END
  END Data_PMOS[201]
  PIN Data_PMOS[202]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6397.785 1046.435 6398.065 1047.435 ;
    END
  END Data_PMOS[202]
  PIN Data_PMOS[196]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6396.105 1046.435 6396.385 1047.435 ;
    END
  END Data_PMOS[196]
  PIN nTOK_PMOS[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6354.105 1046.435 6354.385 1047.435 ;
    END
  END nTOK_PMOS[9]
  PIN BcidMtx[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6351.865 1046.435 6352.145 1047.435 ;
    END
  END BcidMtx[393]
  PIN BcidMtx[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6350.185 1046.435 6350.465 1047.435 ;
    END
  END BcidMtx[392]
  PIN INJ_IN[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6347.945 1046.435 6348.225 1047.435 ;
    END
  END INJ_IN[130]
  PIN Data_PMOS[198]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6345.705 1046.435 6345.985 1047.435 ;
    END
  END Data_PMOS[198]
  PIN Data_PMOS[193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6344.025 1046.435 6344.305 1047.435 ;
    END
  END Data_PMOS[193]
  PIN Data_PMOS[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6342.345 1046.435 6342.625 1047.435 ;
    END
  END Data_PMOS[190]
  PIN MASKV[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6332.265 1046.435 6332.545 1047.435 ;
    END
  END MASKV[130]
  PIN DIG_MON_PMOS[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6330.025 1046.435 6330.305 1047.435 ;
    END
  END DIG_MON_PMOS[18]
  PIN DIG_MON_SEL[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6327.785 1046.435 6328.065 1047.435 ;
    END
  END DIG_MON_SEL[129]
  PIN INJ_ROW[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6322.465 1046.435 6322.745 1047.435 ;
    END
  END INJ_ROW[64]
  PIN Data_PMOS[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6320.785 1046.435 6321.065 1047.435 ;
    END
  END Data_PMOS[176]
  PIN Data_PMOS[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6319.105 1046.435 6319.385 1047.435 ;
    END
  END Data_PMOS[173]
  PIN Data_PMOS[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6291.945 1046.435 6292.225 1047.435 ;
    END
  END Data_PMOS[182]
  PIN INJ_IN[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6289.705 1046.435 6289.985 1047.435 ;
    END
  END INJ_IN[129]
  PIN BcidMtx[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6286.905 1046.435 6287.185 1047.435 ;
    END
  END BcidMtx[388]
  PIN Read_PMOS[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6285.225 1046.435 6285.505 1047.435 ;
    END
  END Read_PMOS[8]
  PIN BcidMtx[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6283.545 1046.435 6283.825 1047.435 ;
    END
  END BcidMtx[384]
  PIN Data_PMOS[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6280.745 1046.435 6281.025 1047.435 ;
    END
  END Data_PMOS[170]
  PIN Data_PMOS[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6266.185 1046.435 6266.465 1047.435 ;
    END
  END Data_PMOS[178]
  PIN Data_PMOS[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6265.065 1046.435 6265.345 1047.435 ;
    END
  END Data_PMOS[184]
  PIN Data_PMOS[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6263.385 1046.435 6263.665 1047.435 ;
    END
  END Data_PMOS[168]
  PIN MASKH[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6261.705 1046.435 6261.985 1047.435 ;
    END
  END MASKH[64]
  PIN MASKD[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6256.665 1046.435 6256.945 1047.435 ;
    END
  END MASKD[127]
  PIN MASKV[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6253.865 1046.435 6254.145 1047.435 ;
    END
  END MASKV[127]
  PIN Data_PMOS[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6212.425 1046.435 6212.705 1047.435 ;
    END
  END Data_PMOS[159]
  PIN Data_PMOS[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6210.745 1046.435 6211.025 1047.435 ;
    END
  END Data_PMOS[160]
  PIN Data_PMOS[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6209.065 1046.435 6209.345 1047.435 ;
    END
  END Data_PMOS[154]
  PIN nTOK_PMOS[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6206.265 1046.435 6206.545 1047.435 ;
    END
  END nTOK_PMOS[7]
  PIN BcidMtx[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6204.025 1046.435 6204.305 1047.435 ;
    END
  END BcidMtx[381]
  PIN BcidMtx[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6202.345 1046.435 6202.625 1047.435 ;
    END
  END BcidMtx[380]
  PIN INJ_IN[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6191.705 1046.435 6191.985 1047.435 ;
    END
  END INJ_IN[126]
  PIN Data_PMOS[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6189.465 1046.435 6189.745 1047.435 ;
    END
  END Data_PMOS[156]
  PIN Data_PMOS[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6187.785 1046.435 6188.065 1047.435 ;
    END
  END Data_PMOS[151]
  PIN Data_PMOS[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6186.105 1046.435 6186.385 1047.435 ;
    END
  END Data_PMOS[148]
  PIN MASKV[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6182.465 1046.435 6182.745 1047.435 ;
    END
  END MASKV[126]
  PIN MASKH[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6181.905 1046.435 6182.185 1047.435 ;
    END
  END MASKH[63]
  PIN DIG_MON_SEL[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7271.945 1046.435 7272.225 1047.435 ;
    END
  END DIG_MON_SEL[153]
  PIN INJ_ROW[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7828.585 1046.435 7828.865 1047.435 ;
    END
  END INJ_ROW[83]
  PIN Data_PMOS[575]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7826.905 1046.435 7827.185 1047.435 ;
    END
  END Data_PMOS[575]
  PIN Data_PMOS[572]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7825.225 1046.435 7825.505 1047.435 ;
    END
  END Data_PMOS[572]
  PIN Data_PMOS[581]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7823.545 1046.435 7823.825 1047.435 ;
    END
  END Data_PMOS[581]
  PIN INJ_IN[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7821.305 1046.435 7821.585 1047.435 ;
    END
  END INJ_IN[167]
  PIN BcidMtx[502]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7805.065 1046.435 7805.345 1047.435 ;
    END
  END BcidMtx[502]
  PIN Read_PMOS[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7803.385 1046.435 7803.665 1047.435 ;
    END
  END Read_PMOS[27]
  PIN BcidMtx[498]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7801.705 1046.435 7801.985 1047.435 ;
    END
  END BcidMtx[498]
  PIN Data_PMOS[570]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7799.465 1046.435 7799.745 1047.435 ;
    END
  END Data_PMOS[570]
  PIN Data_PMOS[582]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7797.785 1046.435 7798.065 1047.435 ;
    END
  END Data_PMOS[582]
  PIN Data_PMOS[583]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7796.105 1046.435 7796.385 1047.435 ;
    END
  END Data_PMOS[583]
  PIN Data_PMOS[567]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7794.425 1046.435 7794.705 1047.435 ;
    END
  END Data_PMOS[567]
  PIN MASKH[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7754.105 1046.435 7754.385 1047.435 ;
    END
  END MASKH[83]
  PIN MASKD[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7749.065 1046.435 7749.345 1047.435 ;
    END
  END MASKD[165]
  PIN MASKV[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7746.265 1046.435 7746.545 1047.435 ;
    END
  END MASKV[165]
  PIN Data_PMOS[558]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7744.585 1046.435 7744.865 1047.435 ;
    END
  END Data_PMOS[558]
  PIN Data_PMOS[559]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7742.905 1046.435 7743.185 1047.435 ;
    END
  END Data_PMOS[559]
  PIN Data_PMOS[553]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7741.225 1046.435 7741.505 1047.435 ;
    END
  END Data_PMOS[553]
  PIN nTOK_PMOS[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7730.025 1046.435 7730.305 1047.435 ;
    END
  END nTOK_PMOS[26]
  PIN BcidMtx[495]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7727.785 1046.435 7728.065 1047.435 ;
    END
  END BcidMtx[495]
  PIN BcidMtx[494]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7726.105 1046.435 7726.385 1047.435 ;
    END
  END BcidMtx[494]
  PIN INJ_IN[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7721.905 1046.435 7722.185 1047.435 ;
    END
  END INJ_IN[164]
  PIN Data_PMOS[555]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7719.665 1046.435 7719.945 1047.435 ;
    END
  END Data_PMOS[555]
  PIN Data_PMOS[556]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7718.545 1046.435 7718.825 1047.435 ;
    END
  END Data_PMOS[556]
  PIN Data_PMOS[557]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7691.385 1046.435 7691.665 1047.435 ;
    END
  END Data_PMOS[557]
  PIN Data_PMOS[563]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7689.705 1046.435 7689.985 1047.435 ;
    END
  END Data_PMOS[563]
  PIN MASKD[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7688.025 1046.435 7688.305 1047.435 ;
    END
  END MASKD[164]
  PIN DIG_MON_SEL[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7685.225 1046.435 7685.505 1047.435 ;
    END
  END DIG_MON_SEL[164]
  PIN DIG_MON_PMOS[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7682.425 1046.435 7682.705 1047.435 ;
    END
  END DIG_MON_PMOS[51]
  PIN Data_PMOS[543]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7680.185 1046.435 7680.465 1047.435 ;
    END
  END Data_PMOS[543]
  PIN Data_PMOS[544]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7665.625 1046.435 7665.905 1047.435 ;
    END
  END Data_PMOS[544]
  PIN Data_PMOS[545]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7663.945 1046.435 7664.225 1047.435 ;
    END
  END Data_PMOS[545]
  PIN Data_PMOS[531]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7662.265 1046.435 7662.545 1047.435 ;
    END
  END Data_PMOS[531]
  PIN BcidMtx[491]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7658.905 1046.435 7659.185 1047.435 ;
    END
  END BcidMtx[491]
  PIN FREEZE_PMOS[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7657.225 1046.435 7657.505 1047.435 ;
    END
  END FREEZE_PMOS[25]
  PIN BcidMtx[487]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7655.545 1046.435 7655.825 1047.435 ;
    END
  END BcidMtx[487]
  PIN Data_PMOS[528]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7614.105 1046.435 7614.385 1047.435 ;
    END
  END Data_PMOS[528]
  PIN Data_PMOS[540]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7612.425 1046.435 7612.705 1047.435 ;
    END
  END Data_PMOS[540]
  PIN Data_PMOS[541]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7610.745 1046.435 7611.025 1047.435 ;
    END
  END Data_PMOS[541]
  PIN Data_PMOS[525]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7609.065 1046.435 7609.345 1047.435 ;
    END
  END Data_PMOS[525]
  PIN MASKH[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7607.385 1046.435 7607.665 1047.435 ;
    END
  END MASKH[81]
  PIN MASKD[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7602.345 1046.435 7602.625 1047.435 ;
    END
  END MASKD[161]
  PIN MASKV[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7591.145 1046.435 7591.425 1047.435 ;
    END
  END MASKV[161]
  PIN Data_PMOS[516]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7589.465 1046.435 7589.745 1047.435 ;
    END
  END Data_PMOS[516]
  PIN Data_PMOS[517]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7587.785 1046.435 7588.065 1047.435 ;
    END
  END Data_PMOS[517]
  PIN Data_PMOS[511]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7586.105 1046.435 7586.385 1047.435 ;
    END
  END Data_PMOS[511]
  PIN nTOK_PMOS[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7581.345 1046.435 7581.625 1047.435 ;
    END
  END nTOK_PMOS[24]
  PIN BcidMtx[483]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7579.105 1046.435 7579.385 1047.435 ;
    END
  END BcidMtx[483]
  PIN BcidMtx[481]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7551.385 1046.435 7551.665 1047.435 ;
    END
  END BcidMtx[481]
  PIN Data_PMOS[507]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7548.585 1046.435 7548.865 1047.435 ;
    END
  END Data_PMOS[507]
  PIN Data_PMOS[519]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7546.905 1046.435 7547.185 1047.435 ;
    END
  END Data_PMOS[519]
  PIN Data_PMOS[520]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7545.225 1046.435 7545.505 1047.435 ;
    END
  END Data_PMOS[520]
  PIN Data_PMOS[504]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7543.545 1046.435 7543.825 1047.435 ;
    END
  END Data_PMOS[504]
  PIN MASKH[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7541.865 1046.435 7542.145 1047.435 ;
    END
  END MASKH[80]
  PIN MASKD[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7523.945 1046.435 7524.225 1047.435 ;
    END
  END MASKD[159]
  PIN MASKV[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7521.145 1046.435 7521.425 1047.435 ;
    END
  END MASKV[159]
  PIN Data_PMOS[495]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7519.465 1046.435 7519.745 1047.435 ;
    END
  END Data_PMOS[495]
  PIN Data_PMOS[496]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7517.785 1046.435 7518.065 1047.435 ;
    END
  END Data_PMOS[496]
  PIN Data_PMOS[490]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7516.105 1046.435 7516.385 1047.435 ;
    END
  END Data_PMOS[490]
  PIN nTOK_PMOS[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7474.105 1046.435 7474.385 1047.435 ;
    END
  END nTOK_PMOS[23]
  PIN DIG_MON_HV[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18645.545 1046.435 18645.825 1047.435 ;
    END
  END DIG_MON_HV[101]
  PIN BcidMtx[477]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7471.865 1046.435 7472.145 1047.435 ;
    END
  END BcidMtx[477]
  PIN BcidMtx[476]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7470.185 1046.435 7470.465 1047.435 ;
    END
  END BcidMtx[476]
  PIN INJ_IN[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7467.945 1046.435 7468.225 1047.435 ;
    END
  END INJ_IN[158]
  PIN Data_PMOS[492]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7465.705 1046.435 7465.985 1047.435 ;
    END
  END Data_PMOS[492]
  PIN Data_PMOS[487]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7464.025 1046.435 7464.305 1047.435 ;
    END
  END Data_PMOS[487]
  PIN Data_PMOS[484]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7462.345 1046.435 7462.625 1047.435 ;
    END
  END Data_PMOS[484]
  PIN MASKV[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7452.265 1046.435 7452.545 1047.435 ;
    END
  END MASKV[158]
  PIN DIG_MON_PMOS[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7450.025 1046.435 7450.305 1047.435 ;
    END
  END DIG_MON_PMOS[46]
  PIN DIG_MON_SEL[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7447.785 1046.435 7448.065 1047.435 ;
    END
  END DIG_MON_SEL[157]
  PIN DIG_MON_PMOS[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7445.545 1046.435 7445.825 1047.435 ;
    END
  END DIG_MON_PMOS[45]
  PIN Data_PMOS[470]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7440.785 1046.435 7441.065 1047.435 ;
    END
  END Data_PMOS[470]
  PIN Data_PMOS[467]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7439.105 1046.435 7439.385 1047.435 ;
    END
  END Data_PMOS[467]
  PIN Data_PMOS[482]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7412.505 1046.435 7412.785 1047.435 ;
    END
  END Data_PMOS[482]
  PIN INJ_IN[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7409.705 1046.435 7409.985 1047.435 ;
    END
  END INJ_IN[157]
  PIN Data_HV[1129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18810.745 1046.435 18811.025 1047.435 ;
    END
  END Data_HV[1129]
  PIN BcidMtx[471]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7406.345 1046.435 7406.625 1047.435 ;
    END
  END BcidMtx[471]
  PIN INJ_ROW[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18642.465 1046.435 18642.745 1047.435 ;
    END
  END INJ_ROW[218]
  PIN BcidMtx[468]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7403.545 1046.435 7403.825 1047.435 ;
    END
  END BcidMtx[468]
  PIN Data_PMOS[465]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7401.305 1046.435 7401.585 1047.435 ;
    END
  END Data_PMOS[465]
  PIN Data_PMOS[472]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7386.185 1046.435 7386.465 1047.435 ;
    END
  END Data_PMOS[472]
  PIN Data_PMOS[473]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7384.505 1046.435 7384.785 1047.435 ;
    END
  END Data_PMOS[473]
  PIN Data_PMOS[462]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7383.385 1046.435 7383.665 1047.435 ;
    END
  END Data_PMOS[462]
  PIN MASKH[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7381.705 1046.435 7381.985 1047.435 ;
    END
  END MASKH[78]
  PIN MASKD[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7376.665 1046.435 7376.945 1047.435 ;
    END
  END MASKD[155]
  PIN MASKV[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7373.865 1046.435 7374.145 1047.435 ;
    END
  END MASKV[155]
  PIN Data_PMOS[453]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7332.425 1046.435 7332.705 1047.435 ;
    END
  END Data_PMOS[453]
  PIN Data_PMOS[454]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7330.745 1046.435 7331.025 1047.435 ;
    END
  END Data_PMOS[454]
  PIN Data_PMOS[448]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7329.065 1046.435 7329.345 1047.435 ;
    END
  END Data_PMOS[448]
  PIN nTOK_PMOS[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7326.265 1046.435 7326.545 1047.435 ;
    END
  END nTOK_PMOS[21]
  PIN BcidMtx[466]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7324.585 1046.435 7324.865 1047.435 ;
    END
  END BcidMtx[466]
  PIN Read_PMOS[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7322.905 1046.435 7323.185 1047.435 ;
    END
  END Read_PMOS[21]
  PIN BcidMtx[462]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7321.225 1046.435 7321.505 1047.435 ;
    END
  END BcidMtx[462]
  PIN Data_PMOS[444]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7310.585 1046.435 7310.865 1047.435 ;
    END
  END Data_PMOS[444]
  PIN Data_PMOS[451]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7308.345 1046.435 7308.625 1047.435 ;
    END
  END Data_PMOS[451]
  PIN Data_PMOS[452]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7306.665 1046.435 7306.945 1047.435 ;
    END
  END Data_PMOS[452]
  PIN Data_PMOS[458]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 7304.985 1046.435 7305.265 1047.435 ;
    END
  END Data_PMOS[458]
  PIN Data_HV[841]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17770.825 1046.435 17771.105 1047.435 ;
    END
  END Data_HV[841]
  PIN MASKV[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17769.145 1046.435 17769.425 1047.435 ;
    END
  END MASKV[416]
  PIN MASKD[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17768.025 1046.435 17768.305 1047.435 ;
    END
  END MASKD[416]
  PIN Data_HV[1088]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18661.225 1046.435 18661.505 1047.435 ;
    END
  END Data_HV[1088]
  PIN DIG_MON_HV[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17762.425 1046.435 17762.705 1047.435 ;
    END
  END DIG_MON_HV[79]
  PIN MASKV[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17760.745 1046.435 17761.025 1047.435 ;
    END
  END MASKV[415]
  PIN Data_HV[838]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17745.625 1046.435 17745.905 1047.435 ;
    END
  END Data_HV[838]
  PIN Data_HV[839]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17743.945 1046.435 17744.225 1047.435 ;
    END
  END Data_HV[839]
  PIN Data_HV[826]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17742.825 1046.435 17743.105 1047.435 ;
    END
  END Data_HV[826]
  PIN BcidMtx[1247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17738.905 1046.435 17739.185 1047.435 ;
    END
  END BcidMtx[1247]
  PIN FREEZE_HV[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17737.225 1046.435 17737.505 1047.435 ;
    END
  END FREEZE_HV[39]
  PIN BcidMtx[1244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17736.105 1046.435 17736.385 1047.435 ;
    END
  END BcidMtx[1244]
  PIN Data_HV[822]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17694.105 1046.435 17694.385 1047.435 ;
    END
  END Data_HV[822]
  PIN Data_HV[834]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17692.425 1046.435 17692.705 1047.435 ;
    END
  END Data_HV[834]
  PIN Data_HV[823]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17691.305 1046.435 17691.585 1047.435 ;
    END
  END Data_HV[823]
  PIN Data_HV[819]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17689.065 1046.435 17689.345 1047.435 ;
    END
  END Data_HV[819]
  PIN MASKH[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17687.385 1046.435 17687.665 1047.435 ;
    END
  END MASKH[207]
  PIN DIG_MON_HV[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17685.705 1046.435 17685.985 1047.435 ;
    END
  END DIG_MON_HV[78]
  PIN DIG_MON_SEL[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17683.465 1046.435 17683.745 1047.435 ;
    END
  END DIG_MON_SEL[413]
  PIN DIG_MON_HV[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17681.225 1046.435 17681.505 1047.435 ;
    END
  END DIG_MON_HV[77]
  PIN MASKV[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17671.145 1046.435 17671.425 1047.435 ;
    END
  END MASKV[413]
  PIN Data_HV[817]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17668.905 1046.435 17669.185 1047.435 ;
    END
  END Data_HV[817]
  PIN Data_HV[818]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17667.225 1046.435 17667.505 1047.435 ;
    END
  END Data_HV[818]
  PIN Data_HV[805]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17666.105 1046.435 17666.385 1047.435 ;
    END
  END Data_HV[805]
  PIN BcidMtx[1241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17660.225 1046.435 17660.505 1047.435 ;
    END
  END BcidMtx[1241]
  PIN Read_HV[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17632.505 1046.435 17632.785 1047.435 ;
    END
  END Read_HV[38]
  PIN BcidMtx[1237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17631.385 1046.435 17631.665 1047.435 ;
    END
  END BcidMtx[1237]
  PIN Data_HV[800]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17628.025 1046.435 17628.305 1047.435 ;
    END
  END Data_HV[800]
  PIN Data_HV[808]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17626.345 1046.435 17626.625 1047.435 ;
    END
  END Data_HV[808]
  PIN Data_HV[814]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17625.225 1046.435 17625.505 1047.435 ;
    END
  END Data_HV[814]
  PIN Data_HV[815]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17622.985 1046.435 17623.265 1047.435 ;
    END
  END Data_HV[815]
  PIN MASKD[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17621.305 1046.435 17621.585 1047.435 ;
    END
  END MASKD[412]
  PIN MASKD[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17603.945 1046.435 17604.225 1047.435 ;
    END
  END MASKD[411]
  PIN Data_HV[1051]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18583.945 1046.435 18584.225 1047.435 ;
    END
  END Data_HV[1051]
  PIN MASKV[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17601.145 1046.435 17601.425 1047.435 ;
    END
  END MASKV[411]
  PIN Data_HV[796]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17598.905 1046.435 17599.185 1047.435 ;
    END
  END Data_HV[796]
  PIN Data_HV[797]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17597.225 1046.435 17597.505 1047.435 ;
    END
  END Data_HV[797]
  PIN Data_HV[784]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17596.105 1046.435 17596.385 1047.435 ;
    END
  END Data_HV[784]
  PIN BcidMtx[1235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17552.985 1046.435 17553.265 1047.435 ;
    END
  END BcidMtx[1235]
  PIN FREEZE_HV[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17551.305 1046.435 17551.585 1047.435 ;
    END
  END FREEZE_HV[37]
  PIN BcidMtx[1232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17550.185 1046.435 17550.465 1047.435 ;
    END
  END BcidMtx[1232]
  PIN Data_HV[780]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17546.825 1046.435 17547.105 1047.435 ;
    END
  END Data_HV[780]
  PIN Data_HV[792]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17545.145 1046.435 17545.425 1047.435 ;
    END
  END Data_HV[792]
  PIN Data_HV[781]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17544.025 1046.435 17544.305 1047.435 ;
    END
  END Data_HV[781]
  PIN Data_HV[777]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17541.785 1046.435 17542.065 1047.435 ;
    END
  END Data_HV[777]
  PIN MASKH[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17531.705 1046.435 17531.985 1047.435 ;
    END
  END MASKH[205]
  PIN DIG_MON_HV[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17530.025 1046.435 17530.305 1047.435 ;
    END
  END DIG_MON_HV[74]
  PIN MASKD[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17526.665 1046.435 17526.945 1047.435 ;
    END
  END MASKD[409]
  PIN MASKV[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17521.905 1046.435 17522.185 1047.435 ;
    END
  END MASKV[409]
  PIN Data_HV[764]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17520.785 1046.435 17521.065 1047.435 ;
    END
  END Data_HV[764]
  PIN Data_HV[769]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17493.065 1046.435 17493.345 1047.435 ;
    END
  END Data_HV[769]
  PIN Data_HV[763]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17491.385 1046.435 17491.665 1047.435 ;
    END
  END Data_HV[763]
  PIN INJ_IN[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17489.705 1046.435 17489.985 1047.435 ;
    END
  END INJ_IN[409]
  PIN BcidMtx[1227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17486.345 1046.435 17486.625 1047.435 ;
    END
  END BcidMtx[1227]
  PIN BcidMtx[1226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17484.665 1046.435 17484.945 1047.435 ;
    END
  END BcidMtx[1226]
  PIN BcidMtx[1224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17483.545 1046.435 17483.825 1047.435 ;
    END
  END BcidMtx[1224]
  PIN Data_HV[765]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17480.185 1046.435 17480.465 1047.435 ;
    END
  END Data_HV[765]
  PIN Data_HV[760]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17465.625 1046.435 17465.905 1047.435 ;
    END
  END Data_HV[760]
  PIN Data_HV[767]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17464.505 1046.435 17464.785 1047.435 ;
    END
  END Data_HV[767]
  PIN MASKV[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17462.265 1046.435 17462.545 1047.435 ;
    END
  END MASKV[408]
  PIN DIG_MON_HV[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17460.025 1046.435 17460.305 1047.435 ;
    END
  END DIG_MON_HV[72]
  PIN DIG_MON_SEL[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17458.345 1046.435 17458.625 1047.435 ;
    END
  END DIG_MON_SEL[408]
  PIN INJ_ROW[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17454.425 1046.435 17454.705 1047.435 ;
    END
  END INJ_ROW[203]
  PIN Data_HV[743]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17412.985 1046.435 17413.265 1047.435 ;
    END
  END Data_HV[743]
  PIN Data_HV[754]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17411.865 1046.435 17412.145 1047.435 ;
    END
  END Data_HV[754]
  PIN Data_HV[749]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17409.625 1046.435 17409.905 1047.435 ;
    END
  END Data_HV[749]
  PIN INJ_IN[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17407.385 1046.435 17407.665 1047.435 ;
    END
  END INJ_IN[407]
  PIN BcidMtx[1223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17405.145 1046.435 17405.425 1047.435 ;
    END
  END BcidMtx[1223]
  PIN Read_HV[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17402.905 1046.435 17403.185 1047.435 ;
    END
  END Read_HV[35]
  PIN BcidMtx[1218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17401.225 1046.435 17401.505 1047.435 ;
    END
  END BcidMtx[1218]
  PIN Data_HV[738]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17390.585 1046.435 17390.865 1047.435 ;
    END
  END Data_HV[738]
  PIN Data_HV[745]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17388.345 1046.435 17388.625 1047.435 ;
    END
  END Data_HV[745]
  PIN Data_HV[746]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17386.665 1046.435 17386.945 1047.435 ;
    END
  END Data_HV[746]
  PIN Data_HV[735]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17385.545 1046.435 17385.825 1047.435 ;
    END
  END Data_HV[735]
  PIN MASKD[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17381.345 1046.435 17381.625 1047.435 ;
    END
  END MASKD[406]
  PIN DIG_MON_SEL[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17378.545 1046.435 17378.825 1047.435 ;
    END
  END DIG_MON_SEL[406]
  PIN DIG_MON_SEL[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18471.945 1046.435 18472.225 1047.435 ;
    END
  END DIG_MON_SEL[433]
  PIN MASKV[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18468.025 1046.435 18468.305 1047.435 ;
    END
  END MASKV[433]
  PIN Data_HV[1020]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18466.345 1046.435 18466.625 1047.435 ;
    END
  END Data_HV[1020]
  PIN Data_HV[1021]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18464.665 1046.435 18464.945 1047.435 ;
    END
  END Data_HV[1021]
  PIN Data_HV[1015]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18462.985 1046.435 18463.265 1047.435 ;
    END
  END Data_HV[1015]
  PIN nTOK_HV[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18460.185 1046.435 18460.465 1047.435 ;
    END
  END nTOK_HV[48]
  PIN BcidMtx[1299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18444.505 1046.435 18444.785 1047.435 ;
    END
  END BcidMtx[1299]
  PIN BcidMtx[1298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18442.825 1046.435 18443.105 1047.435 ;
    END
  END BcidMtx[1298]
  PIN INJ_IN[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18440.585 1046.435 18440.865 1047.435 ;
    END
  END INJ_IN[432]
  PIN Data_HV[1017]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18438.345 1046.435 18438.625 1047.435 ;
    END
  END Data_HV[1017]
  PIN Data_HV[1012]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18436.665 1046.435 18436.945 1047.435 ;
    END
  END Data_HV[1012]
  PIN Data_HV[1009]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18434.985 1046.435 18435.265 1047.435 ;
    END
  END Data_HV[1009]
  PIN MASKV[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18394.665 1046.435 18394.945 1047.435 ;
    END
  END MASKV[432]
  PIN DIG_MON_HV[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18392.425 1046.435 18392.705 1047.435 ;
    END
  END DIG_MON_HV[96]
  PIN DIG_MON_SEL[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18390.185 1046.435 18390.465 1047.435 ;
    END
  END DIG_MON_SEL[431]
  PIN INJ_ROW[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18386.825 1046.435 18387.105 1047.435 ;
    END
  END INJ_ROW[215]
  PIN Data_HV[995]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18385.145 1046.435 18385.425 1047.435 ;
    END
  END Data_HV[995]
  PIN Data_HV[992]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18383.465 1046.435 18383.745 1047.435 ;
    END
  END Data_HV[992]
  PIN Data_HV[1001]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18381.785 1046.435 18382.065 1047.435 ;
    END
  END Data_HV[1001]
  PIN INJ_IN[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18371.145 1046.435 18371.425 1047.435 ;
    END
  END INJ_IN[431]
  PIN BcidMtx[1294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18368.345 1046.435 18368.625 1047.435 ;
    END
  END BcidMtx[1294]
  PIN Read_HV[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18366.665 1046.435 18366.945 1047.435 ;
    END
  END Read_HV[47]
  PIN BcidMtx[1290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18364.985 1046.435 18365.265 1047.435 ;
    END
  END BcidMtx[1290]
  PIN Data_HV[989]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18360.225 1046.435 18360.505 1047.435 ;
    END
  END Data_HV[989]
  PIN Data_HV[997]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 18358.545 1046.435 18358.825 1047.435 ;
    END
  END Data_HV[997]
  PIN OUTA_MON_L_PAD[0]
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 616.1 8960.155 618.1 8995.155 ;
    END
  END OUTA_MON_L_PAD[0]
  PIN VCASN_DAC_MON_L_PAD
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 616.1 8720.15 618.1 8755.15 ;
    END
  END VCASN_DAC_MON_L_PAD
  PIN VCASN_MON_L_PAD
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 616.1 8840.155 618.1 8875.155 ;
    END
  END VCASN_MON_L_PAD
  PIN DACMON_ICASN_PAD
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 616.1 680.155 618.1 715.155 ;
    END
  END DACMON_ICASN_PAD
  PIN DACMON_IRESET_PAD
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 616.1 800.155 618.1 835.155 ;
    END
  END DACMON_IRESET_PAD
  PIN DACMON_IDB_PAD
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 616.1 920.155 618.1 955.155 ;
    END
  END DACMON_IDB_PAD
  PIN DACMON_ITHR_PAD
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 616.1 1040.155 618.1 1075.155 ;
    END
  END DACMON_ITHR_PAD
  PIN DACMON_IBIAS_PAD
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 616.1 1160.155 618.1 1195.155 ;
    END
  END DACMON_IBIAS_PAD
  PIN PSUB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER TOP_M ;
        RECT 746.1 9398.18 748.1 9448.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 638.18 748.1 688.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 9398.18 19453.9 9448.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 638.18 19453.9 688.18 ;
    END
  END PSUB
  PIN PWELL
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 746.1 9278.18 748.1 9328.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 5438.18 748.1 5488.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 1478.18 748.1 1528.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 9278.18 19453.9 9328.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 5438.18 19453.9 5488.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 1478.18 19453.9 1528.18 ;
    END
  END PWELL
  PIN VDDA
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 746.1 9158.18 748.1 9208.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 8678.18 748.1 8728.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 8198.18 748.1 8248.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 7718.18 748.1 7768.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 7238.18 748.1 7288.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 6758.18 748.1 6808.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 6278.18 748.1 6328.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 5798.18 748.1 5848.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 5318.18 748.1 5368.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 4838.18 748.1 4888.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 4358.18 748.1 4408.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 3878.18 748.1 3928.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 3398.18 748.1 3448.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 2918.18 748.1 2968.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 2438.18 748.1 2488.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 1958.18 748.1 2008.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 9158.18 19453.9 9208.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 8678.18 19453.9 8728.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 8198.18 19453.9 8248.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 7718.18 19453.9 7768.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 7238.18 19453.9 7288.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 6758.18 19453.9 6808.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 6278.18 19453.9 6328.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 5798.18 19453.9 5848.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 5318.18 19453.9 5368.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 4838.18 19453.9 4888.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 4358.18 19453.9 4408.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 3878.18 19453.9 3928.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 3398.18 19453.9 3448.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 2918.18 19453.9 2968.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 2438.18 19453.9 2488.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 1958.18 19453.9 2008.18 ;
    END
  END VDDA
  PIN GNDA
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 746.1 9038.18 748.1 9088.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 8558.18 748.1 8608.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 8078.18 748.1 8128.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 7598.18 748.1 7648.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 7118.18 748.1 7168.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 6638.18 748.1 6688.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 6158.18 748.1 6208.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 5678.18 748.1 5728.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 5198.18 748.1 5248.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 4718.18 748.1 4768.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 4238.18 748.1 4288.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 3758.18 748.1 3808.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 3278.18 748.1 3328.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 2798.18 748.1 2848.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 2318.18 748.1 2368.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 1838.18 748.1 1888.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 9038.18 19453.9 9088.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 8558.18 19453.9 8608.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 8078.18 19453.9 8128.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 7598.18 19453.9 7648.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 7118.18 19453.9 7168.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 6638.18 19453.9 6688.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 6158.18 19453.9 6208.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 5678.18 19453.9 5728.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 5198.18 19453.9 5248.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 4718.18 19453.9 4768.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 4238.18 19453.9 4288.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 3758.18 19453.9 3808.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 3278.18 19453.9 3328.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 2798.18 19453.9 2848.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 2318.18 19453.9 2368.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 1838.18 19453.9 1888.18 ;
    END
  END GNDA
  PIN VDDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER TOP_M ;
        RECT 746.1 8918.18 748.1 8968.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 8438.18 748.1 8488.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 7958.18 748.1 8008.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 7478.18 748.1 7528.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 6998.18 748.1 7048.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 6518.18 748.1 6568.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 6038.18 748.1 6088.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 5558.18 748.1 5608.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 5078.18 748.1 5128.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 4598.18 748.1 4648.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 4118.18 748.1 4168.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 3638.18 748.1 3688.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 3158.18 748.1 3208.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 2678.18 748.1 2728.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 2198.18 748.1 2248.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 1718.18 748.1 1768.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 8918.18 19453.9 8968.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 8438.18 19453.9 8488.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 7958.18 19453.9 8008.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 7478.18 19453.9 7528.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 6998.18 19453.9 7048.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 6518.18 19453.9 6568.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 6038.18 19453.9 6088.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 5078.18 19453.9 5128.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 4598.18 19453.9 4648.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 4118.18 19453.9 4168.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 3638.18 19453.9 3688.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 3158.18 19453.9 3208.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 2678.18 19453.9 2728.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 2198.18 19453.9 2248.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 1718.18 19453.9 1768.18 ;
    END
  END VDDD
  PIN GNDD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER TOP_M ;
        RECT 746.1 8798.18 748.1 8848.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 8318.18 748.1 8368.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 7838.18 748.1 7888.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 7358.18 748.1 7408.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 6878.18 748.1 6928.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 6398.18 748.1 6448.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 5918.18 748.1 5968.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 4958.18 748.1 5008.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 4478.18 748.1 4528.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 3998.18 748.1 4048.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 3518.18 748.1 3568.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 3038.18 748.1 3088.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 2558.18 748.1 2608.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 2078.18 748.1 2128.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 1598.18 748.1 1648.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 8798.18 19453.9 8848.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 8318.18 19453.9 8368.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 7838.18 19453.9 7888.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 7358.18 19453.9 7408.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 6878.18 19453.9 6928.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 6398.18 19453.9 6448.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 5918.18 19453.9 5968.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 4958.18 19453.9 5008.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 4478.18 19453.9 4528.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 3998.18 19453.9 4048.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 3518.18 19453.9 3568.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 3038.18 19453.9 3088.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 2558.18 19453.9 2608.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 2078.18 19453.9 2128.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 1598.18 19453.9 1648.18 ;
    END
  END GNDD
  PIN GNDA_DAC
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 746.1 998.18 748.1 1048.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 758.18 748.1 808.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 998.18 19453.9 1048.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 758.18 19453.9 808.18 ;
    END
  END GNDA_DAC
  PIN VDDA_DAC
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 746.1 1118.18 748.1 1168.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 746.1 878.18 748.1 928.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 1118.18 19453.9 1168.18 ;
    END
    PORT
      LAYER TOP_M ;
        RECT 19451.9 878.18 19453.9 928.18 ;
    END
  END VDDA_DAC
  PIN VPCNOSF
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 616.1 1298.18 618.1 1348.18 ;
    END
  END VPCNOSF
  PIN OUTA_MON_L_PAD[1]
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 616.1 9080.155 618.1 9115.155 ;
    END
  END OUTA_MON_L_PAD[1]
  PIN OUTA_MON_L_PAD[2]
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 616.1 9200.155 618.1 9235.155 ;
    END
  END OUTA_MON_L_PAD[2]
  PIN OUTA_MON_L_PAD[3]
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 616.1 9320.155 618.1 9355.155 ;
    END
  END OUTA_MON_L_PAD[3]
  PIN OUTA_MON_R_PAD[3]
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 19581.9 9320.155 19583.9 9355.155 ;
    END
  END OUTA_MON_R_PAD[3]
  PIN OUTA_MON_R_PAD[2]
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 19581.9 9200.155 19583.9 9235.155 ;
    END
  END OUTA_MON_R_PAD[2]
  PIN OUTA_MON_R_PAD[1]
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 19581.9 9080.155 19583.9 9115.155 ;
    END
  END OUTA_MON_R_PAD[1]
  PIN OUTA_MON_R_PAD[0]
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 19581.9 8960.155 19583.9 8995.155 ;
    END
  END OUTA_MON_R_PAD[0]
  PIN VCASN_MON_R_PAD
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 19581.9 8840.155 19583.9 8875.155 ;
    END
  END VCASN_MON_R_PAD
  PIN VCASN_DAC_MON_R_PAD
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 19581.9 8720.15 19583.9 8755.15 ;
    END
  END VCASN_DAC_MON_R_PAD
  PIN HV_DIODE
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 19451.9 5558.18 19453.9 5608.18 ;
    END
  END HV_DIODE
  PIN DACMON_VL_PAD
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 19581.9 1040.155 19583.9 1075.155 ;
    END
  END DACMON_VL_PAD
  PIN DACMON_VH_PAD
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 19581.9 920.155 19583.9 955.155 ;
    END
  END DACMON_VH_PAD
  PIN DACMON_VRESET_P_PAD
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 19581.9 800.155 19583.9 835.155 ;
    END
  END DACMON_VRESET_P_PAD
  PIN VPC_PAD
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 19581.9 1280.155 19583.9 1315.155 ;
    END
  END VPC_PAD
  PIN BiasSF_PAD
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 19581.9 1400.155 19583.9 1435.155 ;
    END
  END BiasSF_PAD
  PIN DACMON_VCASN_DAC_PAD
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER TOP_M ;
        RECT 19581.9 680.155 19583.9 715.155 ;
    END
  END DACMON_VCASN_DAC_PAD
  OBS
    LAYER M1 ;
      RECT 4.1 9985 20195.9 9995.9 ;
      RECT 20190 4.1 20195.9 9995.9 ;
      RECT 19150 9953.14 19170 9995.9 ;
      RECT 990 9953.14 1010 9995.9 ;
      RECT 4.1 4.1 10 9995.9 ;
      RECT 4.1 9974.53 20195.9 9979.53 ;
      RECT 4.1 9964.31 20195.9 9969.31 ;
      RECT 4.1 9953.565 20195.9 9958.565 ;
      RECT 30 9953.56 20170 9958.565 ;
      RECT 19150.42 9952.8 19169.58 9995.9 ;
      RECT 19169.24 9472.58 19169.58 9995.9 ;
      RECT 990.42 9952.8 1009.58 9995.9 ;
      RECT 1009.24 9473.18 1009.58 9995.9 ;
      RECT 19150.42 9473.18 19150.76 9995.9 ;
      RECT 990.42 9472.58 990.76 9995.9 ;
      RECT 19150.42 9832.8 19169.58 9834.32 ;
      RECT 990.42 9832.8 1009.58 9834.32 ;
      RECT 19150 9833.14 19170 9833.98 ;
      RECT 990 9833.14 1010 9833.98 ;
      RECT 19150.42 9712.8 19169.58 9714.32 ;
      RECT 990.42 9712.8 1009.58 9714.32 ;
      RECT 19150 9713.14 19170 9713.98 ;
      RECT 990 9713.14 1010 9713.98 ;
      RECT 19150.42 9592.8 19169.58 9594.32 ;
      RECT 990.42 9592.8 1009.58 9594.32 ;
      RECT 19150 9593.14 19170 9593.98 ;
      RECT 990 9593.14 1010 9593.98 ;
      RECT 19150.42 9473.18 19169.58 9474.32 ;
      RECT 990.42 9473.18 1009.58 9474.32 ;
      RECT 19150 9473.18 19170 9473.98 ;
      RECT 990 9473.18 1010 9473.98 ;
      RECT 19432.99 1042.86 19433.99 9473.58 ;
      RECT 766.01 9472.58 1001.04 9473.58 ;
      RECT 4.1 9473.18 20195.9 9473.56 ;
      RECT 19158.96 9472.58 19433.99 9473.58 ;
      RECT 19158.96 1042.86 19159.96 9474.32 ;
      RECT 1000.04 1042.86 1001.04 9474.32 ;
      RECT 766.01 1042.86 767.01 9473.58 ;
      RECT 19158.96 9422.7 19433.99 9423.7 ;
      RECT 766.01 9422.7 1001.04 9423.7 ;
      RECT 19158.96 9372.82 19433.99 9373.82 ;
      RECT 766.01 9372.82 1001.04 9373.82 ;
      RECT 19158.96 9322.94 19433.99 9323.94 ;
      RECT 766.01 9322.94 1001.04 9323.94 ;
      RECT 19158.96 9273.06 19433.99 9274.06 ;
      RECT 766.01 9273.06 1001.04 9274.06 ;
      RECT 19158.96 9223.18 19433.99 9224.18 ;
      RECT 766.01 9223.18 1001.04 9224.18 ;
      RECT 19158.96 9173.3 19433.99 9174.3 ;
      RECT 766.01 9173.3 1001.04 9174.3 ;
      RECT 19158.96 9123.42 19433.99 9124.42 ;
      RECT 766.01 9123.42 1001.04 9124.42 ;
      RECT 19158.96 9073.54 19433.99 9074.54 ;
      RECT 766.01 9073.54 1001.04 9074.54 ;
      RECT 19158.96 9023.66 19433.99 9024.66 ;
      RECT 766.01 9023.66 1001.04 9024.66 ;
      RECT 19158.96 8973.78 19433.99 8974.78 ;
      RECT 766.01 8973.78 1001.04 8974.78 ;
      RECT 19158.96 8923.9 19433.99 8924.9 ;
      RECT 766.01 8923.9 1001.04 8924.9 ;
      RECT 19158.96 8874.02 19433.99 8875.02 ;
      RECT 766.01 8874.02 1001.04 8875.02 ;
      RECT 19158.96 8824.14 19433.99 8825.14 ;
      RECT 766.01 8824.14 1001.04 8825.14 ;
      RECT 19158.96 8774.26 19433.99 8775.26 ;
      RECT 766.01 8774.26 1001.04 8775.26 ;
      RECT 19158.96 8724.38 19433.99 8725.38 ;
      RECT 766.01 8724.38 1001.04 8725.38 ;
      RECT 19158.96 8674.5 19433.99 8675.5 ;
      RECT 766.01 8674.5 1001.04 8675.5 ;
      RECT 19158.96 8624.62 19433.99 8625.62 ;
      RECT 766.01 8624.62 1001.04 8625.62 ;
      RECT 19158.96 8574.74 19433.99 8575.74 ;
      RECT 766.01 8574.74 1001.04 8575.74 ;
      RECT 19158.96 8524.86 19433.99 8525.86 ;
      RECT 766.01 8524.86 1001.04 8525.86 ;
      RECT 19158.96 8474.98 19433.99 8475.98 ;
      RECT 766.01 8474.98 1001.04 8475.98 ;
      RECT 19158.96 8425.1 19433.99 8426.1 ;
      RECT 766.01 8425.1 1001.04 8426.1 ;
      RECT 19158.96 8375.22 19433.99 8376.22 ;
      RECT 766.01 8375.22 1001.04 8376.22 ;
      RECT 19158.96 8325.34 19433.99 8326.34 ;
      RECT 766.01 8325.34 1001.04 8326.34 ;
      RECT 19158.96 8275.46 19433.99 8276.46 ;
      RECT 766.01 8275.46 1001.04 8276.46 ;
      RECT 19158.96 8225.58 19433.99 8226.58 ;
      RECT 766.01 8225.58 1001.04 8226.58 ;
      RECT 19158.96 8175.7 19433.99 8176.7 ;
      RECT 766.01 8175.7 1001.04 8176.7 ;
      RECT 19158.96 8125.82 19433.99 8126.82 ;
      RECT 766.01 8125.82 1001.04 8126.82 ;
      RECT 19158.96 8075.94 19433.99 8076.94 ;
      RECT 766.01 8075.94 1001.04 8076.94 ;
      RECT 19158.96 8026.06 19433.99 8027.06 ;
      RECT 766.01 8026.06 1001.04 8027.06 ;
      RECT 19158.96 7976.18 19433.99 7977.18 ;
      RECT 766.01 7976.18 1001.04 7977.18 ;
      RECT 19158.96 7926.3 19433.99 7927.3 ;
      RECT 766.01 7926.3 1001.04 7927.3 ;
      RECT 19158.96 7876.42 19433.99 7877.42 ;
      RECT 766.01 7876.42 1001.04 7877.42 ;
      RECT 19158.96 7826.54 19433.99 7827.54 ;
      RECT 766.01 7826.54 1001.04 7827.54 ;
      RECT 19158.96 7776.66 19433.99 7777.66 ;
      RECT 766.01 7776.66 1001.04 7777.66 ;
      RECT 19158.96 7726.78 19433.99 7727.78 ;
      RECT 766.01 7726.78 1001.04 7727.78 ;
      RECT 19158.96 7676.9 19433.99 7677.9 ;
      RECT 766.01 7676.9 1001.04 7677.9 ;
      RECT 19158.96 7627.02 19433.99 7628.02 ;
      RECT 766.01 7627.02 1001.04 7628.02 ;
      RECT 19158.96 7577.14 19433.99 7578.14 ;
      RECT 766.01 7577.14 1001.04 7578.14 ;
      RECT 19158.96 7527.26 19433.99 7528.26 ;
      RECT 766.01 7527.26 1001.04 7528.26 ;
      RECT 19158.96 7477.38 19433.99 7478.38 ;
      RECT 766.01 7477.38 1001.04 7478.38 ;
      RECT 19158.96 7427.5 19433.99 7428.5 ;
      RECT 766.01 7427.5 1001.04 7428.5 ;
      RECT 19158.96 7377.62 19433.99 7378.62 ;
      RECT 766.01 7377.62 1001.04 7378.62 ;
      RECT 19158.96 7327.74 19433.99 7328.74 ;
      RECT 766.01 7327.74 1001.04 7328.74 ;
      RECT 19158.96 7277.86 19433.99 7278.86 ;
      RECT 766.01 7277.86 1001.04 7278.86 ;
      RECT 19158.96 7227.98 19433.99 7228.98 ;
      RECT 766.01 7227.98 1001.04 7228.98 ;
      RECT 19158.96 7178.1 19433.99 7179.1 ;
      RECT 766.01 7178.1 1001.04 7179.1 ;
      RECT 19158.96 7128.22 19433.99 7129.22 ;
      RECT 766.01 7128.22 1001.04 7129.22 ;
      RECT 19158.96 7078.34 19433.99 7079.34 ;
      RECT 766.01 7078.34 1001.04 7079.34 ;
      RECT 19158.96 7028.46 19433.99 7029.46 ;
      RECT 766.01 7028.46 1001.04 7029.46 ;
      RECT 19158.96 6978.58 19433.99 6979.58 ;
      RECT 766.01 6978.58 1001.04 6979.58 ;
      RECT 19158.96 6928.7 19433.99 6929.7 ;
      RECT 766.01 6928.7 1001.04 6929.7 ;
      RECT 19158.96 6878.82 19433.99 6879.82 ;
      RECT 766.01 6878.82 1001.04 6879.82 ;
      RECT 19158.96 6828.94 19433.99 6829.94 ;
      RECT 766.01 6828.94 1001.04 6829.94 ;
      RECT 19158.96 6779.06 19433.99 6780.06 ;
      RECT 766.01 6779.06 1001.04 6780.06 ;
      RECT 19158.96 6729.18 19433.99 6730.18 ;
      RECT 766.01 6729.18 1001.04 6730.18 ;
      RECT 19158.96 6679.3 19433.99 6680.3 ;
      RECT 766.01 6679.3 1001.04 6680.3 ;
      RECT 19158.96 6629.42 19433.99 6630.42 ;
      RECT 766.01 6629.42 1001.04 6630.42 ;
      RECT 19158.96 6579.54 19433.99 6580.54 ;
      RECT 766.01 6579.54 1001.04 6580.54 ;
      RECT 19158.96 6529.66 19433.99 6530.66 ;
      RECT 766.01 6529.66 1001.04 6530.66 ;
      RECT 19158.96 6479.78 19433.99 6480.78 ;
      RECT 766.01 6479.78 1001.04 6480.78 ;
      RECT 19158.96 6429.9 19433.99 6430.9 ;
      RECT 766.01 6429.9 1001.04 6430.9 ;
      RECT 19158.96 6380.02 19433.99 6381.02 ;
      RECT 766.01 6380.02 1001.04 6381.02 ;
      RECT 19158.96 6330.14 19433.99 6331.14 ;
      RECT 766.01 6330.14 1001.04 6331.14 ;
      RECT 19158.96 6280.26 19433.99 6281.26 ;
      RECT 766.01 6280.26 1001.04 6281.26 ;
      RECT 19158.96 6230.38 19433.99 6231.38 ;
      RECT 766.01 6230.38 1001.04 6231.38 ;
      RECT 19158.96 6180.5 19433.99 6181.5 ;
      RECT 766.01 6180.5 1001.04 6181.5 ;
      RECT 19158.96 6130.62 19433.99 6131.62 ;
      RECT 766.01 6130.62 1001.04 6131.62 ;
      RECT 19158.96 6080.74 19433.99 6081.74 ;
      RECT 766.01 6080.74 1001.04 6081.74 ;
      RECT 19158.96 6030.86 19433.99 6031.86 ;
      RECT 766.01 6030.86 1001.04 6031.86 ;
      RECT 19158.96 5980.98 19433.99 5981.98 ;
      RECT 766.01 5980.98 1001.04 5981.98 ;
      RECT 19158.96 5931.1 19433.99 5932.1 ;
      RECT 766.01 5931.1 1001.04 5932.1 ;
      RECT 19158.96 5881.22 19433.99 5882.22 ;
      RECT 766.01 5881.22 1001.04 5882.22 ;
      RECT 19158.96 5831.34 19433.99 5832.34 ;
      RECT 766.01 5831.34 1001.04 5832.34 ;
      RECT 19158.96 5781.46 19433.99 5782.46 ;
      RECT 766.01 5781.46 1001.04 5782.46 ;
      RECT 19158.96 5731.58 19433.99 5732.58 ;
      RECT 766.01 5731.58 1001.04 5732.58 ;
      RECT 19158.96 5681.7 19433.99 5682.7 ;
      RECT 766.01 5681.7 1001.04 5682.7 ;
      RECT 19158.96 5631.82 19433.99 5632.82 ;
      RECT 766.01 5631.82 1001.04 5632.82 ;
      RECT 19158.96 5581.94 19433.99 5582.94 ;
      RECT 766.01 5581.94 1001.04 5582.94 ;
      RECT 19158.96 5532.06 19433.99 5533.06 ;
      RECT 766.01 5532.06 1001.04 5533.06 ;
      RECT 19158.96 5482.18 19433.99 5483.18 ;
      RECT 766.01 5482.18 1001.04 5483.18 ;
      RECT 19158.96 5432.3 19433.99 5433.3 ;
      RECT 766.01 5432.3 1001.04 5433.3 ;
      RECT 19158.96 5382.42 19433.99 5383.42 ;
      RECT 766.01 5382.42 1001.04 5383.42 ;
      RECT 19158.96 5332.54 19433.99 5333.54 ;
      RECT 766.01 5332.54 1001.04 5333.54 ;
      RECT 19158.96 5282.66 19433.99 5283.66 ;
      RECT 766.01 5282.66 1001.04 5283.66 ;
      RECT 19158.96 5232.78 19433.99 5233.78 ;
      RECT 766.01 5232.78 1001.04 5233.78 ;
      RECT 19158.96 5182.9 19433.99 5183.9 ;
      RECT 766.01 5182.9 1001.04 5183.9 ;
      RECT 19158.96 5133.02 19433.99 5134.02 ;
      RECT 766.01 5133.02 1001.04 5134.02 ;
      RECT 19158.96 5083.14 19433.99 5084.14 ;
      RECT 766.01 5083.14 1001.04 5084.14 ;
      RECT 19158.96 5033.26 19433.99 5034.26 ;
      RECT 766.01 5033.26 1001.04 5034.26 ;
      RECT 19158.96 4983.38 19433.99 4984.38 ;
      RECT 766.01 4983.38 1001.04 4984.38 ;
      RECT 19158.96 4933.5 19433.99 4934.5 ;
      RECT 766.01 4933.5 1001.04 4934.5 ;
      RECT 19158.96 4883.62 19433.99 4884.62 ;
      RECT 766.01 4883.62 1001.04 4884.62 ;
      RECT 19158.96 4833.74 19433.99 4834.74 ;
      RECT 766.01 4833.74 1001.04 4834.74 ;
      RECT 19158.96 4783.86 19433.99 4784.86 ;
      RECT 766.01 4783.86 1001.04 4784.86 ;
      RECT 19158.96 4733.98 19433.99 4734.98 ;
      RECT 766.01 4733.98 1001.04 4734.98 ;
      RECT 19158.96 4684.1 19433.99 4685.1 ;
      RECT 766.01 4684.1 1001.04 4685.1 ;
      RECT 19158.96 4634.22 19433.99 4635.22 ;
      RECT 766.01 4634.22 1001.04 4635.22 ;
      RECT 19158.96 4584.34 19433.99 4585.34 ;
      RECT 766.01 4584.34 1001.04 4585.34 ;
      RECT 19158.96 4534.46 19433.99 4535.46 ;
      RECT 766.01 4534.46 1001.04 4535.46 ;
      RECT 19158.96 4484.58 19433.99 4485.58 ;
      RECT 766.01 4484.58 1001.04 4485.58 ;
      RECT 19158.96 4434.7 19433.99 4435.7 ;
      RECT 766.01 4434.7 1001.04 4435.7 ;
      RECT 19158.96 4384.82 19433.99 4385.82 ;
      RECT 766.01 4384.82 1001.04 4385.82 ;
      RECT 19158.96 4334.94 19433.99 4335.94 ;
      RECT 766.01 4334.94 1001.04 4335.94 ;
      RECT 19158.96 4285.06 19433.99 4286.06 ;
      RECT 766.01 4285.06 1001.04 4286.06 ;
      RECT 19158.96 4235.18 19433.99 4236.18 ;
      RECT 766.01 4235.18 1001.04 4236.18 ;
      RECT 19158.96 4185.3 19433.99 4186.3 ;
      RECT 766.01 4185.3 1001.04 4186.3 ;
      RECT 19158.96 4135.42 19433.99 4136.42 ;
      RECT 766.01 4135.42 1001.04 4136.42 ;
      RECT 19158.96 4085.54 19433.99 4086.54 ;
      RECT 766.01 4085.54 1001.04 4086.54 ;
      RECT 19158.96 4035.66 19433.99 4036.66 ;
      RECT 766.01 4035.66 1001.04 4036.66 ;
      RECT 19158.96 3985.78 19433.99 3986.78 ;
      RECT 766.01 3985.78 1001.04 3986.78 ;
      RECT 19158.96 3935.9 19433.99 3936.9 ;
      RECT 766.01 3935.9 1001.04 3936.9 ;
      RECT 19158.96 3886.02 19433.99 3887.02 ;
      RECT 766.01 3886.02 1001.04 3887.02 ;
      RECT 19158.96 3836.14 19433.99 3837.14 ;
      RECT 766.01 3836.14 1001.04 3837.14 ;
      RECT 19158.96 3786.26 19433.99 3787.26 ;
      RECT 766.01 3786.26 1001.04 3787.26 ;
      RECT 19158.96 3736.38 19433.99 3737.38 ;
      RECT 766.01 3736.38 1001.04 3737.38 ;
      RECT 19158.96 3686.5 19433.99 3687.5 ;
      RECT 766.01 3686.5 1001.04 3687.5 ;
      RECT 19158.96 3636.62 19433.99 3637.62 ;
      RECT 766.01 3636.62 1001.04 3637.62 ;
      RECT 19158.96 3586.74 19433.99 3587.74 ;
      RECT 766.01 3586.74 1001.04 3587.74 ;
      RECT 19158.96 3536.86 19433.99 3537.86 ;
      RECT 766.01 3536.86 1001.04 3537.86 ;
      RECT 19158.96 3486.98 19433.99 3487.98 ;
      RECT 766.01 3486.98 1001.04 3487.98 ;
      RECT 19158.96 3437.1 19433.99 3438.1 ;
      RECT 766.01 3437.1 1001.04 3438.1 ;
      RECT 19158.96 3387.22 19433.99 3388.22 ;
      RECT 766.01 3387.22 1001.04 3388.22 ;
      RECT 19158.96 3337.34 19433.99 3338.34 ;
      RECT 766.01 3337.34 1001.04 3338.34 ;
      RECT 19158.96 3287.46 19433.99 3288.46 ;
      RECT 766.01 3287.46 1001.04 3288.46 ;
      RECT 19158.96 3237.58 19433.99 3238.58 ;
      RECT 766.01 3237.58 1001.04 3238.58 ;
      RECT 19158.96 3187.7 19433.99 3188.7 ;
      RECT 766.01 3187.7 1001.04 3188.7 ;
      RECT 19158.96 3137.82 19433.99 3138.82 ;
      RECT 766.01 3137.82 1001.04 3138.82 ;
      RECT 19158.96 3087.94 19433.99 3088.94 ;
      RECT 766.01 3087.94 1001.04 3088.94 ;
      RECT 19158.96 3038.06 19433.99 3039.06 ;
      RECT 766.01 3038.06 1001.04 3039.06 ;
      RECT 19158.96 2988.18 19433.99 2989.18 ;
      RECT 766.01 2988.18 1001.04 2989.18 ;
      RECT 19158.96 2938.3 19433.99 2939.3 ;
      RECT 766.01 2938.3 1001.04 2939.3 ;
      RECT 19158.96 2888.42 19433.99 2889.42 ;
      RECT 766.01 2888.42 1001.04 2889.42 ;
      RECT 19158.96 2838.54 19433.99 2839.54 ;
      RECT 766.01 2838.54 1001.04 2839.54 ;
      RECT 19158.96 2788.66 19433.99 2789.66 ;
      RECT 766.01 2788.66 1001.04 2789.66 ;
      RECT 19158.96 2738.78 19433.99 2739.78 ;
      RECT 766.01 2738.78 1001.04 2739.78 ;
      RECT 19158.96 2688.9 19433.99 2689.9 ;
      RECT 766.01 2688.9 1001.04 2689.9 ;
      RECT 19158.96 2639.02 19433.99 2640.02 ;
      RECT 766.01 2639.02 1001.04 2640.02 ;
      RECT 19158.96 2589.14 19433.99 2590.14 ;
      RECT 766.01 2589.14 1001.04 2590.14 ;
      RECT 19158.96 2539.26 19433.99 2540.26 ;
      RECT 766.01 2539.26 1001.04 2540.26 ;
      RECT 19158.96 2489.38 19433.99 2490.38 ;
      RECT 766.01 2489.38 1001.04 2490.38 ;
      RECT 19158.96 2439.5 19433.99 2440.5 ;
      RECT 766.01 2439.5 1001.04 2440.5 ;
      RECT 19158.96 2389.62 19433.99 2390.62 ;
      RECT 766.01 2389.62 1001.04 2390.62 ;
      RECT 19158.96 2339.74 19433.99 2340.74 ;
      RECT 766.01 2339.74 1001.04 2340.74 ;
      RECT 19158.96 2289.86 19433.99 2290.86 ;
      RECT 766.01 2289.86 1001.04 2290.86 ;
      RECT 19158.96 2239.98 19433.99 2240.98 ;
      RECT 766.01 2239.98 1001.04 2240.98 ;
      RECT 19158.96 2190.1 19433.99 2191.1 ;
      RECT 766.01 2190.1 1001.04 2191.1 ;
      RECT 19158.96 2140.22 19433.99 2141.22 ;
      RECT 766.01 2140.22 1001.04 2141.22 ;
      RECT 19158.96 2090.34 19433.99 2091.34 ;
      RECT 766.01 2090.34 1001.04 2091.34 ;
      RECT 19158.96 2040.46 19433.99 2041.46 ;
      RECT 766.01 2040.46 1001.04 2041.46 ;
      RECT 19158.96 1990.58 19433.99 1991.58 ;
      RECT 766.01 1990.58 1001.04 1991.58 ;
      RECT 19158.96 1940.7 19433.99 1941.7 ;
      RECT 766.01 1940.7 1001.04 1941.7 ;
      RECT 19158.96 1890.82 19433.99 1891.82 ;
      RECT 766.01 1890.82 1001.04 1891.82 ;
      RECT 19158.96 1840.94 19433.99 1841.94 ;
      RECT 766.01 1840.94 1001.04 1841.94 ;
      RECT 19158.96 1791.06 19433.99 1792.06 ;
      RECT 766.01 1791.06 1001.04 1792.06 ;
      RECT 19158.96 1741.18 19433.99 1742.18 ;
      RECT 766.01 1741.18 1001.04 1742.18 ;
      RECT 19158.96 1691.3 19433.99 1692.3 ;
      RECT 766.01 1691.3 1001.04 1692.3 ;
      RECT 19158.96 1641.42 19433.99 1642.42 ;
      RECT 766.01 1641.42 1001.04 1642.42 ;
      RECT 19158.96 1591.54 19433.99 1592.54 ;
      RECT 766.01 1591.54 1001.04 1592.54 ;
      RECT 19158.96 1541.66 19433.99 1542.66 ;
      RECT 766.01 1541.66 1001.04 1542.66 ;
      RECT 19158.96 1491.78 19433.99 1492.78 ;
      RECT 766.01 1491.78 1001.04 1492.78 ;
      RECT 19158.96 1441.9 19433.99 1442.9 ;
      RECT 766.01 1441.9 1001.04 1442.9 ;
      RECT 19158.96 1392.02 19433.99 1393.02 ;
      RECT 766.01 1392.02 1001.04 1393.02 ;
      RECT 19158.96 1342.14 19433.99 1343.14 ;
      RECT 766.01 1342.14 1001.04 1343.14 ;
      RECT 19158.96 1292.26 19433.99 1293.26 ;
      RECT 766.01 1292.26 1001.04 1293.26 ;
      RECT 19158.96 1242.38 19433.99 1243.38 ;
      RECT 766.01 1242.38 1001.04 1243.38 ;
      RECT 19158.96 1192.5 19433.99 1193.5 ;
      RECT 766.01 1192.5 1001.04 1193.5 ;
      RECT 19158.96 1142.62 19433.99 1143.62 ;
      RECT 766.01 1142.62 1001.04 1143.62 ;
      RECT 19158.96 1092.74 19433.99 1093.74 ;
      RECT 766.01 1092.74 1001.04 1093.74 ;
      RECT 19157.4 646.015 19158.96 1049.355 ;
      RECT 1001.04 650.935 1003.6 1049.355 ;
      RECT 19156.4 1042.86 19433.99 1043.86 ;
      RECT 766.01 1042.86 1003.6 1043.86 ;
      RECT 19156.4 650.935 19158.96 1049.355 ;
      RECT 1001.04 650.935 19158.96 651.935 ;
      RECT 1001.04 646.015 1002.6 1049.355 ;
      RECT 4.1 4.1 20195.9 10 ;
      RECT 19163.33 9478.7 19163.63 9479.91 ;
      RECT 19163.33 9478.7 19164.09 9479 ;
      RECT 19163.79 9476.66 19164.09 9479 ;
      RECT 19161.16 9476.66 19161.46 9479 ;
      RECT 19155.9 9476.66 19168 9477.66 ;
      RECT 19163.33 9490.08 19163.63 9491.29 ;
      RECT 19163.33 9490.08 19164.09 9490.38 ;
      RECT 19163.79 9485.79 19164.09 9490.38 ;
      RECT 19161.16 9485.79 19161.46 9490.38 ;
      RECT 19155.035 9487.585 19168 9488.585 ;
      RECT 19163.33 9485.79 19164.09 9486.09 ;
      RECT 19163.33 9484.88 19163.63 9486.09 ;
      RECT 19163.33 9501.46 19163.63 9502.67 ;
      RECT 19163.33 9501.46 19164.09 9501.76 ;
      RECT 19163.79 9497.17 19164.09 9501.76 ;
      RECT 19161.16 9497.17 19161.46 9501.76 ;
      RECT 19155.035 9498.965 19168 9499.965 ;
      RECT 19163.33 9497.17 19164.09 9497.47 ;
      RECT 19163.33 9496.26 19163.63 9497.47 ;
      RECT 19163.33 9512.84 19163.63 9514.05 ;
      RECT 19163.33 9512.84 19164.09 9513.14 ;
      RECT 19163.79 9508.55 19164.09 9513.14 ;
      RECT 19161.16 9508.55 19161.46 9513.14 ;
      RECT 19155.035 9510.345 19168 9511.345 ;
      RECT 19163.33 9508.55 19164.09 9508.85 ;
      RECT 19163.33 9507.64 19163.63 9508.85 ;
      RECT 19163.33 9524.22 19163.63 9525.43 ;
      RECT 19163.33 9524.22 19164.09 9524.52 ;
      RECT 19163.79 9519.93 19164.09 9524.52 ;
      RECT 19161.16 9519.93 19161.46 9524.52 ;
      RECT 19155.035 9521.725 19168 9522.725 ;
      RECT 19163.33 9519.93 19164.09 9520.23 ;
      RECT 19163.33 9519.02 19163.63 9520.23 ;
      RECT 19163.33 9535.6 19163.63 9536.81 ;
      RECT 19163.33 9535.6 19164.09 9535.9 ;
      RECT 19163.79 9531.31 19164.09 9535.9 ;
      RECT 19161.16 9531.31 19161.46 9535.9 ;
      RECT 19155.035 9533.105 19168 9534.105 ;
      RECT 19163.33 9531.31 19164.09 9531.61 ;
      RECT 19163.33 9530.4 19163.63 9531.61 ;
      RECT 19163.33 9546.98 19163.63 9548.19 ;
      RECT 19163.33 9546.98 19164.09 9547.28 ;
      RECT 19163.79 9542.69 19164.09 9547.28 ;
      RECT 19161.16 9542.69 19161.46 9547.28 ;
      RECT 19155.035 9544.485 19168 9545.485 ;
      RECT 19163.33 9542.69 19164.09 9542.99 ;
      RECT 19163.33 9541.78 19163.63 9542.99 ;
      RECT 19163.33 9558.36 19163.63 9559.57 ;
      RECT 19163.33 9558.36 19164.09 9558.66 ;
      RECT 19163.79 9554.07 19164.09 9558.66 ;
      RECT 19161.16 9554.07 19161.46 9558.66 ;
      RECT 19155.035 9555.865 19168 9556.865 ;
      RECT 19163.33 9554.07 19164.09 9554.37 ;
      RECT 19163.33 9553.16 19163.63 9554.37 ;
      RECT 19163.33 9569.74 19163.63 9570.95 ;
      RECT 19163.33 9569.74 19164.09 9570.04 ;
      RECT 19163.79 9565.45 19164.09 9570.04 ;
      RECT 19161.16 9565.45 19161.46 9570.04 ;
      RECT 19155.035 9567.245 19168 9568.245 ;
      RECT 19163.33 9565.45 19164.09 9565.75 ;
      RECT 19163.33 9564.54 19163.63 9565.75 ;
      RECT 19163.33 9581.12 19163.63 9582.33 ;
      RECT 19163.33 9581.12 19164.09 9581.42 ;
      RECT 19163.79 9576.83 19164.09 9581.42 ;
      RECT 19161.16 9576.83 19161.46 9581.42 ;
      RECT 19155.035 9578.625 19168 9579.625 ;
      RECT 19163.33 9576.83 19164.09 9577.13 ;
      RECT 19163.33 9575.92 19163.63 9577.13 ;
      RECT 19155.035 9590.005 19168 9591.005 ;
      RECT 19163.79 9588.21 19164.09 9591.005 ;
      RECT 19161.16 9588.21 19161.46 9591.005 ;
      RECT 19163.33 9588.21 19164.09 9588.51 ;
      RECT 19163.33 9587.3 19163.63 9588.51 ;
      RECT 19163.33 9598.7 19163.63 9599.91 ;
      RECT 19163.33 9598.7 19164.09 9599 ;
      RECT 19163.79 9596.66 19164.09 9599 ;
      RECT 19161.16 9596.66 19161.46 9599 ;
      RECT 19155.9 9596.66 19168 9597.66 ;
      RECT 19163.33 9610.08 19163.63 9611.29 ;
      RECT 19163.33 9610.08 19164.09 9610.38 ;
      RECT 19163.79 9605.79 19164.09 9610.38 ;
      RECT 19161.16 9605.79 19161.46 9610.38 ;
      RECT 19155.035 9607.585 19168 9608.585 ;
      RECT 19163.33 9605.79 19164.09 9606.09 ;
      RECT 19163.33 9604.88 19163.63 9606.09 ;
      RECT 19163.33 9621.46 19163.63 9622.67 ;
      RECT 19163.33 9621.46 19164.09 9621.76 ;
      RECT 19163.79 9617.17 19164.09 9621.76 ;
      RECT 19161.16 9617.17 19161.46 9621.76 ;
      RECT 19155.035 9618.965 19168 9619.965 ;
      RECT 19163.33 9617.17 19164.09 9617.47 ;
      RECT 19163.33 9616.26 19163.63 9617.47 ;
      RECT 19163.33 9632.84 19163.63 9634.05 ;
      RECT 19163.33 9632.84 19164.09 9633.14 ;
      RECT 19163.79 9628.55 19164.09 9633.14 ;
      RECT 19161.16 9628.55 19161.46 9633.14 ;
      RECT 19155.035 9630.345 19168 9631.345 ;
      RECT 19163.33 9628.55 19164.09 9628.85 ;
      RECT 19163.33 9627.64 19163.63 9628.85 ;
      RECT 19163.33 9644.22 19163.63 9645.43 ;
      RECT 19163.33 9644.22 19164.09 9644.52 ;
      RECT 19163.79 9639.93 19164.09 9644.52 ;
      RECT 19161.16 9639.93 19161.46 9644.52 ;
      RECT 19155.035 9641.725 19168 9642.725 ;
      RECT 19163.33 9639.93 19164.09 9640.23 ;
      RECT 19163.33 9639.02 19163.63 9640.23 ;
      RECT 19163.33 9655.6 19163.63 9656.81 ;
      RECT 19163.33 9655.6 19164.09 9655.9 ;
      RECT 19163.79 9651.31 19164.09 9655.9 ;
      RECT 19161.16 9651.31 19161.46 9655.9 ;
      RECT 19155.035 9653.105 19168 9654.105 ;
      RECT 19163.33 9651.31 19164.09 9651.61 ;
      RECT 19163.33 9650.4 19163.63 9651.61 ;
      RECT 19163.33 9666.98 19163.63 9668.19 ;
      RECT 19163.33 9666.98 19164.09 9667.28 ;
      RECT 19163.79 9662.69 19164.09 9667.28 ;
      RECT 19161.16 9662.69 19161.46 9667.28 ;
      RECT 19155.035 9664.485 19168 9665.485 ;
      RECT 19163.33 9662.69 19164.09 9662.99 ;
      RECT 19163.33 9661.78 19163.63 9662.99 ;
      RECT 19163.33 9678.36 19163.63 9679.57 ;
      RECT 19163.33 9678.36 19164.09 9678.66 ;
      RECT 19163.79 9674.07 19164.09 9678.66 ;
      RECT 19161.16 9674.07 19161.46 9678.66 ;
      RECT 19155.035 9675.865 19168 9676.865 ;
      RECT 19163.33 9674.07 19164.09 9674.37 ;
      RECT 19163.33 9673.16 19163.63 9674.37 ;
      RECT 19163.33 9689.74 19163.63 9690.95 ;
      RECT 19163.33 9689.74 19164.09 9690.04 ;
      RECT 19163.79 9685.45 19164.09 9690.04 ;
      RECT 19161.16 9685.45 19161.46 9690.04 ;
      RECT 19155.035 9687.245 19168 9688.245 ;
      RECT 19163.33 9685.45 19164.09 9685.75 ;
      RECT 19163.33 9684.54 19163.63 9685.75 ;
      RECT 19163.33 9701.12 19163.63 9702.33 ;
      RECT 19163.33 9701.12 19164.09 9701.42 ;
      RECT 19163.79 9696.83 19164.09 9701.42 ;
      RECT 19161.16 9696.83 19161.46 9701.42 ;
      RECT 19155.035 9698.625 19168 9699.625 ;
      RECT 19163.33 9696.83 19164.09 9697.13 ;
      RECT 19163.33 9695.92 19163.63 9697.13 ;
      RECT 19155.035 9710.005 19168 9711.005 ;
      RECT 19163.79 9708.21 19164.09 9711.005 ;
      RECT 19161.16 9708.21 19161.46 9711.005 ;
      RECT 19163.33 9708.21 19164.09 9708.51 ;
      RECT 19163.33 9707.3 19163.63 9708.51 ;
      RECT 19163.33 9718.7 19163.63 9719.91 ;
      RECT 19163.33 9718.7 19164.09 9719 ;
      RECT 19163.79 9716.66 19164.09 9719 ;
      RECT 19161.16 9716.66 19161.46 9719 ;
      RECT 19155.9 9716.66 19168 9717.66 ;
      RECT 19163.33 9730.08 19163.63 9731.29 ;
      RECT 19163.33 9730.08 19164.09 9730.38 ;
      RECT 19163.79 9725.79 19164.09 9730.38 ;
      RECT 19161.16 9725.79 19161.46 9730.38 ;
      RECT 19155.035 9727.585 19168 9728.585 ;
      RECT 19163.33 9725.79 19164.09 9726.09 ;
      RECT 19163.33 9724.88 19163.63 9726.09 ;
      RECT 19163.33 9741.46 19163.63 9742.67 ;
      RECT 19163.33 9741.46 19164.09 9741.76 ;
      RECT 19163.79 9737.17 19164.09 9741.76 ;
      RECT 19161.16 9737.17 19161.46 9741.76 ;
      RECT 19155.035 9738.965 19168 9739.965 ;
      RECT 19163.33 9737.17 19164.09 9737.47 ;
      RECT 19163.33 9736.26 19163.63 9737.47 ;
      RECT 19163.33 9752.84 19163.63 9754.05 ;
      RECT 19163.33 9752.84 19164.09 9753.14 ;
      RECT 19163.79 9748.55 19164.09 9753.14 ;
      RECT 19161.16 9748.55 19161.46 9753.14 ;
      RECT 19155.035 9750.345 19168 9751.345 ;
      RECT 19163.33 9748.55 19164.09 9748.85 ;
      RECT 19163.33 9747.64 19163.63 9748.85 ;
      RECT 19163.33 9764.22 19163.63 9765.43 ;
      RECT 19163.33 9764.22 19164.09 9764.52 ;
      RECT 19163.79 9759.93 19164.09 9764.52 ;
      RECT 19161.16 9759.93 19161.46 9764.52 ;
      RECT 19155.035 9761.725 19168 9762.725 ;
      RECT 19163.33 9759.93 19164.09 9760.23 ;
      RECT 19163.33 9759.02 19163.63 9760.23 ;
      RECT 19163.33 9775.6 19163.63 9776.81 ;
      RECT 19163.33 9775.6 19164.09 9775.9 ;
      RECT 19163.79 9771.31 19164.09 9775.9 ;
      RECT 19161.16 9771.31 19161.46 9775.9 ;
      RECT 19155.035 9773.105 19168 9774.105 ;
      RECT 19163.33 9771.31 19164.09 9771.61 ;
      RECT 19163.33 9770.4 19163.63 9771.61 ;
      RECT 19163.33 9786.98 19163.63 9788.19 ;
      RECT 19163.33 9786.98 19164.09 9787.28 ;
      RECT 19163.79 9782.69 19164.09 9787.28 ;
      RECT 19161.16 9782.69 19161.46 9787.28 ;
      RECT 19155.035 9784.485 19168 9785.485 ;
      RECT 19163.33 9782.69 19164.09 9782.99 ;
      RECT 19163.33 9781.78 19163.63 9782.99 ;
      RECT 19163.33 9798.36 19163.63 9799.57 ;
      RECT 19163.33 9798.36 19164.09 9798.66 ;
      RECT 19163.79 9794.07 19164.09 9798.66 ;
      RECT 19161.16 9794.07 19161.46 9798.66 ;
      RECT 19155.035 9795.865 19168 9796.865 ;
      RECT 19163.33 9794.07 19164.09 9794.37 ;
      RECT 19163.33 9793.16 19163.63 9794.37 ;
      RECT 19163.33 9809.74 19163.63 9810.95 ;
      RECT 19163.33 9809.74 19164.09 9810.04 ;
      RECT 19163.79 9805.45 19164.09 9810.04 ;
      RECT 19161.16 9805.45 19161.46 9810.04 ;
      RECT 19155.035 9807.245 19168 9808.245 ;
      RECT 19163.33 9805.45 19164.09 9805.75 ;
      RECT 19163.33 9804.54 19163.63 9805.75 ;
      RECT 19163.33 9821.12 19163.63 9822.33 ;
      RECT 19163.33 9821.12 19164.09 9821.42 ;
      RECT 19163.79 9816.83 19164.09 9821.42 ;
      RECT 19161.16 9816.83 19161.46 9821.42 ;
      RECT 19155.035 9818.625 19168 9819.625 ;
      RECT 19163.33 9816.83 19164.09 9817.13 ;
      RECT 19163.33 9815.92 19163.63 9817.13 ;
      RECT 19155.035 9830.005 19168 9831.005 ;
      RECT 19163.79 9828.21 19164.09 9831.005 ;
      RECT 19161.16 9828.21 19161.46 9831.005 ;
      RECT 19163.33 9828.21 19164.09 9828.51 ;
      RECT 19163.33 9827.3 19163.63 9828.51 ;
      RECT 19163.33 9838.7 19163.63 9839.91 ;
      RECT 19163.33 9838.7 19164.09 9839 ;
      RECT 19163.79 9836.66 19164.09 9839 ;
      RECT 19161.16 9836.66 19161.46 9839 ;
      RECT 19155.9 9836.66 19168 9837.66 ;
      RECT 19163.33 9850.08 19163.63 9851.29 ;
      RECT 19163.33 9850.08 19164.09 9850.38 ;
      RECT 19163.79 9845.79 19164.09 9850.38 ;
      RECT 19161.16 9845.79 19161.46 9850.38 ;
      RECT 19155.035 9847.585 19168 9848.585 ;
      RECT 19163.33 9845.79 19164.09 9846.09 ;
      RECT 19163.33 9844.88 19163.63 9846.09 ;
      RECT 19163.33 9861.46 19163.63 9862.67 ;
      RECT 19163.33 9861.46 19164.09 9861.76 ;
      RECT 19163.79 9857.17 19164.09 9861.76 ;
      RECT 19161.16 9857.17 19161.46 9861.76 ;
      RECT 19155.035 9858.965 19168 9859.965 ;
      RECT 19163.33 9857.17 19164.09 9857.47 ;
      RECT 19163.33 9856.26 19163.63 9857.47 ;
      RECT 19163.33 9872.84 19163.63 9874.05 ;
      RECT 19163.33 9872.84 19164.09 9873.14 ;
      RECT 19163.79 9868.55 19164.09 9873.14 ;
      RECT 19161.16 9868.55 19161.46 9873.14 ;
      RECT 19155.035 9870.345 19168 9871.345 ;
      RECT 19163.33 9868.55 19164.09 9868.85 ;
      RECT 19163.33 9867.64 19163.63 9868.85 ;
      RECT 19163.33 9884.22 19163.63 9885.43 ;
      RECT 19163.33 9884.22 19164.09 9884.52 ;
      RECT 19163.79 9879.93 19164.09 9884.52 ;
      RECT 19161.16 9879.93 19161.46 9884.52 ;
      RECT 19155.035 9881.725 19168 9882.725 ;
      RECT 19163.33 9879.93 19164.09 9880.23 ;
      RECT 19163.33 9879.02 19163.63 9880.23 ;
      RECT 19163.33 9895.6 19163.63 9896.81 ;
      RECT 19163.33 9895.6 19164.09 9895.9 ;
      RECT 19163.79 9891.31 19164.09 9895.9 ;
      RECT 19161.16 9891.31 19161.46 9895.9 ;
      RECT 19155.035 9893.105 19168 9894.105 ;
      RECT 19163.33 9891.31 19164.09 9891.61 ;
      RECT 19163.33 9890.4 19163.63 9891.61 ;
      RECT 19163.33 9906.98 19163.63 9908.19 ;
      RECT 19163.33 9906.98 19164.09 9907.28 ;
      RECT 19163.79 9902.69 19164.09 9907.28 ;
      RECT 19161.16 9902.69 19161.46 9907.28 ;
      RECT 19155.035 9904.485 19168 9905.485 ;
      RECT 19163.33 9902.69 19164.09 9902.99 ;
      RECT 19163.33 9901.78 19163.63 9902.99 ;
      RECT 19163.33 9918.36 19163.63 9919.57 ;
      RECT 19163.33 9918.36 19164.09 9918.66 ;
      RECT 19163.79 9914.07 19164.09 9918.66 ;
      RECT 19161.16 9914.07 19161.46 9918.66 ;
      RECT 19155.035 9915.865 19168 9916.865 ;
      RECT 19163.33 9914.07 19164.09 9914.37 ;
      RECT 19163.33 9913.16 19163.63 9914.37 ;
      RECT 19163.33 9929.74 19163.63 9930.95 ;
      RECT 19163.33 9929.74 19164.09 9930.04 ;
      RECT 19163.79 9925.45 19164.09 9930.04 ;
      RECT 19161.16 9925.45 19161.46 9930.04 ;
      RECT 19155.035 9927.245 19168 9928.245 ;
      RECT 19163.33 9925.45 19164.09 9925.75 ;
      RECT 19163.33 9924.54 19163.63 9925.75 ;
      RECT 19163.33 9941.12 19163.63 9942.33 ;
      RECT 19163.33 9941.12 19164.09 9941.42 ;
      RECT 19163.79 9936.83 19164.09 9941.42 ;
      RECT 19161.16 9936.83 19161.46 9941.42 ;
      RECT 19155.035 9938.625 19168 9939.625 ;
      RECT 19163.33 9936.83 19164.09 9937.13 ;
      RECT 19163.33 9935.92 19163.63 9937.13 ;
      RECT 19155.035 9950.005 19168 9951.005 ;
      RECT 19163.79 9948.21 19164.09 9951.005 ;
      RECT 19161.16 9948.21 19161.46 9951.005 ;
      RECT 19163.33 9948.21 19164.09 9948.51 ;
      RECT 19163.33 9947.3 19163.63 9948.51 ;
      RECT 19161.62 9485.15 19162.43 9485.49 ;
      RECT 19158.99 9484.23 19159.29 9485.44 ;
      RECT 19161.62 9484.23 19161.92 9485.49 ;
      RECT 19163.87 9480.26 19164.17 9484.53 ;
      RECT 19161.16 9484.23 19161.92 9484.53 ;
      RECT 19158.53 9484.23 19159.29 9484.53 ;
      RECT 19161.16 9480.26 19161.54 9484.53 ;
      RECT 19158.53 9480.26 19158.83 9484.53 ;
      RECT 19152 9481.895 19164.965 9482.895 ;
      RECT 19161.16 9480.26 19161.92 9480.56 ;
      RECT 19161.62 9479.3 19161.92 9480.56 ;
      RECT 19158.53 9480.26 19159.29 9480.56 ;
      RECT 19158.99 9479.35 19159.29 9480.56 ;
      RECT 19161.62 9479.3 19162.43 9479.64 ;
      RECT 19161.62 9496.53 19162.43 9496.87 ;
      RECT 19158.99 9495.61 19159.29 9496.82 ;
      RECT 19161.62 9495.61 19161.92 9496.87 ;
      RECT 19163.87 9491.64 19164.17 9495.91 ;
      RECT 19161.16 9495.61 19161.92 9495.91 ;
      RECT 19158.53 9495.61 19159.29 9495.91 ;
      RECT 19161.16 9491.64 19161.54 9495.91 ;
      RECT 19158.53 9491.64 19158.83 9495.91 ;
      RECT 19152 9493.275 19164.965 9494.275 ;
      RECT 19161.16 9491.64 19161.92 9491.94 ;
      RECT 19161.62 9490.68 19161.92 9491.94 ;
      RECT 19158.53 9491.64 19159.29 9491.94 ;
      RECT 19158.99 9490.73 19159.29 9491.94 ;
      RECT 19161.62 9490.68 19162.43 9491.02 ;
      RECT 19161.62 9507.91 19162.43 9508.25 ;
      RECT 19158.99 9506.99 19159.29 9508.2 ;
      RECT 19161.62 9506.99 19161.92 9508.25 ;
      RECT 19163.87 9503.02 19164.17 9507.29 ;
      RECT 19161.16 9506.99 19161.92 9507.29 ;
      RECT 19158.53 9506.99 19159.29 9507.29 ;
      RECT 19161.16 9503.02 19161.54 9507.29 ;
      RECT 19158.53 9503.02 19158.83 9507.29 ;
      RECT 19152 9504.655 19164.965 9505.655 ;
      RECT 19161.16 9503.02 19161.92 9503.32 ;
      RECT 19161.62 9502.06 19161.92 9503.32 ;
      RECT 19158.53 9503.02 19159.29 9503.32 ;
      RECT 19158.99 9502.11 19159.29 9503.32 ;
      RECT 19161.62 9502.06 19162.43 9502.4 ;
      RECT 19161.62 9519.29 19162.43 9519.63 ;
      RECT 19158.99 9518.37 19159.29 9519.58 ;
      RECT 19161.62 9518.37 19161.92 9519.63 ;
      RECT 19163.87 9514.4 19164.17 9518.67 ;
      RECT 19161.16 9518.37 19161.92 9518.67 ;
      RECT 19158.53 9518.37 19159.29 9518.67 ;
      RECT 19161.16 9514.4 19161.54 9518.67 ;
      RECT 19158.53 9514.4 19158.83 9518.67 ;
      RECT 19152 9516.035 19164.965 9517.035 ;
      RECT 19161.16 9514.4 19161.92 9514.7 ;
      RECT 19161.62 9513.44 19161.92 9514.7 ;
      RECT 19158.53 9514.4 19159.29 9514.7 ;
      RECT 19158.99 9513.49 19159.29 9514.7 ;
      RECT 19161.62 9513.44 19162.43 9513.78 ;
      RECT 19161.62 9530.67 19162.43 9531.01 ;
      RECT 19158.99 9529.75 19159.29 9530.96 ;
      RECT 19161.62 9529.75 19161.92 9531.01 ;
      RECT 19163.87 9525.78 19164.17 9530.05 ;
      RECT 19161.16 9529.75 19161.92 9530.05 ;
      RECT 19158.53 9529.75 19159.29 9530.05 ;
      RECT 19161.16 9525.78 19161.54 9530.05 ;
      RECT 19158.53 9525.78 19158.83 9530.05 ;
      RECT 19152 9527.415 19164.965 9528.415 ;
      RECT 19161.16 9525.78 19161.92 9526.08 ;
      RECT 19161.62 9524.82 19161.92 9526.08 ;
      RECT 19158.53 9525.78 19159.29 9526.08 ;
      RECT 19158.99 9524.87 19159.29 9526.08 ;
      RECT 19161.62 9524.82 19162.43 9525.16 ;
      RECT 19161.62 9542.05 19162.43 9542.39 ;
      RECT 19158.99 9541.13 19159.29 9542.34 ;
      RECT 19161.62 9541.13 19161.92 9542.39 ;
      RECT 19163.87 9537.16 19164.17 9541.43 ;
      RECT 19161.16 9541.13 19161.92 9541.43 ;
      RECT 19158.53 9541.13 19159.29 9541.43 ;
      RECT 19161.16 9537.16 19161.54 9541.43 ;
      RECT 19158.53 9537.16 19158.83 9541.43 ;
      RECT 19152 9538.795 19164.965 9539.795 ;
      RECT 19161.16 9537.16 19161.92 9537.46 ;
      RECT 19161.62 9536.2 19161.92 9537.46 ;
      RECT 19158.53 9537.16 19159.29 9537.46 ;
      RECT 19158.99 9536.25 19159.29 9537.46 ;
      RECT 19161.62 9536.2 19162.43 9536.54 ;
      RECT 19161.62 9553.43 19162.43 9553.77 ;
      RECT 19158.99 9552.51 19159.29 9553.72 ;
      RECT 19161.62 9552.51 19161.92 9553.77 ;
      RECT 19163.87 9548.54 19164.17 9552.81 ;
      RECT 19161.16 9552.51 19161.92 9552.81 ;
      RECT 19158.53 9552.51 19159.29 9552.81 ;
      RECT 19161.16 9548.54 19161.54 9552.81 ;
      RECT 19158.53 9548.54 19158.83 9552.81 ;
      RECT 19152 9550.175 19164.965 9551.175 ;
      RECT 19161.16 9548.54 19161.92 9548.84 ;
      RECT 19161.62 9547.58 19161.92 9548.84 ;
      RECT 19158.53 9548.54 19159.29 9548.84 ;
      RECT 19158.99 9547.63 19159.29 9548.84 ;
      RECT 19161.62 9547.58 19162.43 9547.92 ;
      RECT 19161.62 9564.81 19162.43 9565.15 ;
      RECT 19158.99 9563.89 19159.29 9565.1 ;
      RECT 19161.62 9563.89 19161.92 9565.15 ;
      RECT 19163.87 9559.92 19164.17 9564.19 ;
      RECT 19161.16 9563.89 19161.92 9564.19 ;
      RECT 19158.53 9563.89 19159.29 9564.19 ;
      RECT 19161.16 9559.92 19161.54 9564.19 ;
      RECT 19158.53 9559.92 19158.83 9564.19 ;
      RECT 19152 9561.555 19164.965 9562.555 ;
      RECT 19161.16 9559.92 19161.92 9560.22 ;
      RECT 19161.62 9558.96 19161.92 9560.22 ;
      RECT 19158.53 9559.92 19159.29 9560.22 ;
      RECT 19158.99 9559.01 19159.29 9560.22 ;
      RECT 19161.62 9558.96 19162.43 9559.3 ;
      RECT 19161.62 9576.19 19162.43 9576.53 ;
      RECT 19158.99 9575.27 19159.29 9576.48 ;
      RECT 19161.62 9575.27 19161.92 9576.53 ;
      RECT 19163.87 9571.3 19164.17 9575.57 ;
      RECT 19161.16 9575.27 19161.92 9575.57 ;
      RECT 19158.53 9575.27 19159.29 9575.57 ;
      RECT 19161.16 9571.3 19161.54 9575.57 ;
      RECT 19158.53 9571.3 19158.83 9575.57 ;
      RECT 19152 9572.935 19164.965 9573.935 ;
      RECT 19161.16 9571.3 19161.92 9571.6 ;
      RECT 19161.62 9570.34 19161.92 9571.6 ;
      RECT 19158.53 9571.3 19159.29 9571.6 ;
      RECT 19158.99 9570.39 19159.29 9571.6 ;
      RECT 19161.62 9570.34 19162.43 9570.68 ;
      RECT 19161.62 9587.57 19162.43 9587.91 ;
      RECT 19158.99 9586.65 19159.29 9587.86 ;
      RECT 19161.62 9586.65 19161.92 9587.91 ;
      RECT 19163.87 9582.68 19164.17 9586.95 ;
      RECT 19161.16 9586.65 19161.92 9586.95 ;
      RECT 19158.53 9586.65 19159.29 9586.95 ;
      RECT 19161.16 9582.68 19161.54 9586.95 ;
      RECT 19158.53 9582.68 19158.83 9586.95 ;
      RECT 19152 9584.315 19164.965 9585.315 ;
      RECT 19161.16 9582.68 19161.92 9582.98 ;
      RECT 19161.62 9581.72 19161.92 9582.98 ;
      RECT 19158.53 9582.68 19159.29 9582.98 ;
      RECT 19158.99 9581.77 19159.29 9582.98 ;
      RECT 19161.62 9581.72 19162.43 9582.06 ;
      RECT 19161.62 9605.15 19162.43 9605.49 ;
      RECT 19158.99 9604.23 19159.29 9605.44 ;
      RECT 19161.62 9604.23 19161.92 9605.49 ;
      RECT 19163.87 9600.26 19164.17 9604.53 ;
      RECT 19161.16 9604.23 19161.92 9604.53 ;
      RECT 19158.53 9604.23 19159.29 9604.53 ;
      RECT 19161.16 9600.26 19161.54 9604.53 ;
      RECT 19158.53 9600.26 19158.83 9604.53 ;
      RECT 19152 9601.895 19164.965 9602.895 ;
      RECT 19161.16 9600.26 19161.92 9600.56 ;
      RECT 19161.62 9599.3 19161.92 9600.56 ;
      RECT 19158.53 9600.26 19159.29 9600.56 ;
      RECT 19158.99 9599.35 19159.29 9600.56 ;
      RECT 19161.62 9599.3 19162.43 9599.64 ;
      RECT 19161.62 9616.53 19162.43 9616.87 ;
      RECT 19158.99 9615.61 19159.29 9616.82 ;
      RECT 19161.62 9615.61 19161.92 9616.87 ;
      RECT 19163.87 9611.64 19164.17 9615.91 ;
      RECT 19161.16 9615.61 19161.92 9615.91 ;
      RECT 19158.53 9615.61 19159.29 9615.91 ;
      RECT 19161.16 9611.64 19161.54 9615.91 ;
      RECT 19158.53 9611.64 19158.83 9615.91 ;
      RECT 19152 9613.275 19164.965 9614.275 ;
      RECT 19161.16 9611.64 19161.92 9611.94 ;
      RECT 19161.62 9610.68 19161.92 9611.94 ;
      RECT 19158.53 9611.64 19159.29 9611.94 ;
      RECT 19158.99 9610.73 19159.29 9611.94 ;
      RECT 19161.62 9610.68 19162.43 9611.02 ;
      RECT 19161.62 9627.91 19162.43 9628.25 ;
      RECT 19158.99 9626.99 19159.29 9628.2 ;
      RECT 19161.62 9626.99 19161.92 9628.25 ;
      RECT 19163.87 9623.02 19164.17 9627.29 ;
      RECT 19161.16 9626.99 19161.92 9627.29 ;
      RECT 19158.53 9626.99 19159.29 9627.29 ;
      RECT 19161.16 9623.02 19161.54 9627.29 ;
      RECT 19158.53 9623.02 19158.83 9627.29 ;
      RECT 19152 9624.655 19164.965 9625.655 ;
      RECT 19161.16 9623.02 19161.92 9623.32 ;
      RECT 19161.62 9622.06 19161.92 9623.32 ;
      RECT 19158.53 9623.02 19159.29 9623.32 ;
      RECT 19158.99 9622.11 19159.29 9623.32 ;
      RECT 19161.62 9622.06 19162.43 9622.4 ;
      RECT 19161.62 9639.29 19162.43 9639.63 ;
      RECT 19158.99 9638.37 19159.29 9639.58 ;
      RECT 19161.62 9638.37 19161.92 9639.63 ;
      RECT 19163.87 9634.4 19164.17 9638.67 ;
      RECT 19161.16 9638.37 19161.92 9638.67 ;
      RECT 19158.53 9638.37 19159.29 9638.67 ;
      RECT 19161.16 9634.4 19161.54 9638.67 ;
      RECT 19158.53 9634.4 19158.83 9638.67 ;
      RECT 19152 9636.035 19164.965 9637.035 ;
      RECT 19161.16 9634.4 19161.92 9634.7 ;
      RECT 19161.62 9633.44 19161.92 9634.7 ;
      RECT 19158.53 9634.4 19159.29 9634.7 ;
      RECT 19158.99 9633.49 19159.29 9634.7 ;
      RECT 19161.62 9633.44 19162.43 9633.78 ;
      RECT 19161.62 9650.67 19162.43 9651.01 ;
      RECT 19158.99 9649.75 19159.29 9650.96 ;
      RECT 19161.62 9649.75 19161.92 9651.01 ;
      RECT 19163.87 9645.78 19164.17 9650.05 ;
      RECT 19161.16 9649.75 19161.92 9650.05 ;
      RECT 19158.53 9649.75 19159.29 9650.05 ;
      RECT 19161.16 9645.78 19161.54 9650.05 ;
      RECT 19158.53 9645.78 19158.83 9650.05 ;
      RECT 19152 9647.415 19164.965 9648.415 ;
      RECT 19161.16 9645.78 19161.92 9646.08 ;
      RECT 19161.62 9644.82 19161.92 9646.08 ;
      RECT 19158.53 9645.78 19159.29 9646.08 ;
      RECT 19158.99 9644.87 19159.29 9646.08 ;
      RECT 19161.62 9644.82 19162.43 9645.16 ;
      RECT 19161.62 9662.05 19162.43 9662.39 ;
      RECT 19158.99 9661.13 19159.29 9662.34 ;
      RECT 19161.62 9661.13 19161.92 9662.39 ;
      RECT 19163.87 9657.16 19164.17 9661.43 ;
      RECT 19161.16 9661.13 19161.92 9661.43 ;
      RECT 19158.53 9661.13 19159.29 9661.43 ;
      RECT 19161.16 9657.16 19161.54 9661.43 ;
      RECT 19158.53 9657.16 19158.83 9661.43 ;
      RECT 19152 9658.795 19164.965 9659.795 ;
      RECT 19161.16 9657.16 19161.92 9657.46 ;
      RECT 19161.62 9656.2 19161.92 9657.46 ;
      RECT 19158.53 9657.16 19159.29 9657.46 ;
      RECT 19158.99 9656.25 19159.29 9657.46 ;
      RECT 19161.62 9656.2 19162.43 9656.54 ;
      RECT 19161.62 9673.43 19162.43 9673.77 ;
      RECT 19158.99 9672.51 19159.29 9673.72 ;
      RECT 19161.62 9672.51 19161.92 9673.77 ;
      RECT 19163.87 9668.54 19164.17 9672.81 ;
      RECT 19161.16 9672.51 19161.92 9672.81 ;
      RECT 19158.53 9672.51 19159.29 9672.81 ;
      RECT 19161.16 9668.54 19161.54 9672.81 ;
      RECT 19158.53 9668.54 19158.83 9672.81 ;
      RECT 19152 9670.175 19164.965 9671.175 ;
      RECT 19161.16 9668.54 19161.92 9668.84 ;
      RECT 19161.62 9667.58 19161.92 9668.84 ;
      RECT 19158.53 9668.54 19159.29 9668.84 ;
      RECT 19158.99 9667.63 19159.29 9668.84 ;
      RECT 19161.62 9667.58 19162.43 9667.92 ;
      RECT 19161.62 9684.81 19162.43 9685.15 ;
      RECT 19158.99 9683.89 19159.29 9685.1 ;
      RECT 19161.62 9683.89 19161.92 9685.15 ;
      RECT 19163.87 9679.92 19164.17 9684.19 ;
      RECT 19161.16 9683.89 19161.92 9684.19 ;
      RECT 19158.53 9683.89 19159.29 9684.19 ;
      RECT 19161.16 9679.92 19161.54 9684.19 ;
      RECT 19158.53 9679.92 19158.83 9684.19 ;
      RECT 19152 9681.555 19164.965 9682.555 ;
      RECT 19161.16 9679.92 19161.92 9680.22 ;
      RECT 19161.62 9678.96 19161.92 9680.22 ;
      RECT 19158.53 9679.92 19159.29 9680.22 ;
      RECT 19158.99 9679.01 19159.29 9680.22 ;
      RECT 19161.62 9678.96 19162.43 9679.3 ;
      RECT 19161.62 9696.19 19162.43 9696.53 ;
      RECT 19158.99 9695.27 19159.29 9696.48 ;
      RECT 19161.62 9695.27 19161.92 9696.53 ;
      RECT 19163.87 9691.3 19164.17 9695.57 ;
      RECT 19161.16 9695.27 19161.92 9695.57 ;
      RECT 19158.53 9695.27 19159.29 9695.57 ;
      RECT 19161.16 9691.3 19161.54 9695.57 ;
      RECT 19158.53 9691.3 19158.83 9695.57 ;
      RECT 19152 9692.935 19164.965 9693.935 ;
      RECT 19161.16 9691.3 19161.92 9691.6 ;
      RECT 19161.62 9690.34 19161.92 9691.6 ;
      RECT 19158.53 9691.3 19159.29 9691.6 ;
      RECT 19158.99 9690.39 19159.29 9691.6 ;
      RECT 19161.62 9690.34 19162.43 9690.68 ;
      RECT 19161.62 9707.57 19162.43 9707.91 ;
      RECT 19158.99 9706.65 19159.29 9707.86 ;
      RECT 19161.62 9706.65 19161.92 9707.91 ;
      RECT 19163.87 9702.68 19164.17 9706.95 ;
      RECT 19161.16 9706.65 19161.92 9706.95 ;
      RECT 19158.53 9706.65 19159.29 9706.95 ;
      RECT 19161.16 9702.68 19161.54 9706.95 ;
      RECT 19158.53 9702.68 19158.83 9706.95 ;
      RECT 19152 9704.315 19164.965 9705.315 ;
      RECT 19161.16 9702.68 19161.92 9702.98 ;
      RECT 19161.62 9701.72 19161.92 9702.98 ;
      RECT 19158.53 9702.68 19159.29 9702.98 ;
      RECT 19158.99 9701.77 19159.29 9702.98 ;
      RECT 19161.62 9701.72 19162.43 9702.06 ;
      RECT 19161.62 9725.15 19162.43 9725.49 ;
      RECT 19158.99 9724.23 19159.29 9725.44 ;
      RECT 19161.62 9724.23 19161.92 9725.49 ;
      RECT 19163.87 9720.26 19164.17 9724.53 ;
      RECT 19161.16 9724.23 19161.92 9724.53 ;
      RECT 19158.53 9724.23 19159.29 9724.53 ;
      RECT 19161.16 9720.26 19161.54 9724.53 ;
      RECT 19158.53 9720.26 19158.83 9724.53 ;
      RECT 19152 9721.895 19164.965 9722.895 ;
      RECT 19161.16 9720.26 19161.92 9720.56 ;
      RECT 19161.62 9719.3 19161.92 9720.56 ;
      RECT 19158.53 9720.26 19159.29 9720.56 ;
      RECT 19158.99 9719.35 19159.29 9720.56 ;
      RECT 19161.62 9719.3 19162.43 9719.64 ;
      RECT 19161.62 9736.53 19162.43 9736.87 ;
      RECT 19158.99 9735.61 19159.29 9736.82 ;
      RECT 19161.62 9735.61 19161.92 9736.87 ;
      RECT 19163.87 9731.64 19164.17 9735.91 ;
      RECT 19161.16 9735.61 19161.92 9735.91 ;
      RECT 19158.53 9735.61 19159.29 9735.91 ;
      RECT 19161.16 9731.64 19161.54 9735.91 ;
      RECT 19158.53 9731.64 19158.83 9735.91 ;
      RECT 19152 9733.275 19164.965 9734.275 ;
      RECT 19161.16 9731.64 19161.92 9731.94 ;
      RECT 19161.62 9730.68 19161.92 9731.94 ;
      RECT 19158.53 9731.64 19159.29 9731.94 ;
      RECT 19158.99 9730.73 19159.29 9731.94 ;
      RECT 19161.62 9730.68 19162.43 9731.02 ;
      RECT 19161.62 9747.91 19162.43 9748.25 ;
      RECT 19158.99 9746.99 19159.29 9748.2 ;
      RECT 19161.62 9746.99 19161.92 9748.25 ;
      RECT 19163.87 9743.02 19164.17 9747.29 ;
      RECT 19161.16 9746.99 19161.92 9747.29 ;
      RECT 19158.53 9746.99 19159.29 9747.29 ;
      RECT 19161.16 9743.02 19161.54 9747.29 ;
      RECT 19158.53 9743.02 19158.83 9747.29 ;
      RECT 19152 9744.655 19164.965 9745.655 ;
      RECT 19161.16 9743.02 19161.92 9743.32 ;
      RECT 19161.62 9742.06 19161.92 9743.32 ;
      RECT 19158.53 9743.02 19159.29 9743.32 ;
      RECT 19158.99 9742.11 19159.29 9743.32 ;
      RECT 19161.62 9742.06 19162.43 9742.4 ;
      RECT 19161.62 9759.29 19162.43 9759.63 ;
      RECT 19158.99 9758.37 19159.29 9759.58 ;
      RECT 19161.62 9758.37 19161.92 9759.63 ;
      RECT 19163.87 9754.4 19164.17 9758.67 ;
      RECT 19161.16 9758.37 19161.92 9758.67 ;
      RECT 19158.53 9758.37 19159.29 9758.67 ;
      RECT 19161.16 9754.4 19161.54 9758.67 ;
      RECT 19158.53 9754.4 19158.83 9758.67 ;
      RECT 19152 9756.035 19164.965 9757.035 ;
      RECT 19161.16 9754.4 19161.92 9754.7 ;
      RECT 19161.62 9753.44 19161.92 9754.7 ;
      RECT 19158.53 9754.4 19159.29 9754.7 ;
      RECT 19158.99 9753.49 19159.29 9754.7 ;
      RECT 19161.62 9753.44 19162.43 9753.78 ;
      RECT 19161.62 9770.67 19162.43 9771.01 ;
      RECT 19158.99 9769.75 19159.29 9770.96 ;
      RECT 19161.62 9769.75 19161.92 9771.01 ;
      RECT 19163.87 9765.78 19164.17 9770.05 ;
      RECT 19161.16 9769.75 19161.92 9770.05 ;
      RECT 19158.53 9769.75 19159.29 9770.05 ;
      RECT 19161.16 9765.78 19161.54 9770.05 ;
      RECT 19158.53 9765.78 19158.83 9770.05 ;
      RECT 19152 9767.415 19164.965 9768.415 ;
      RECT 19161.16 9765.78 19161.92 9766.08 ;
      RECT 19161.62 9764.82 19161.92 9766.08 ;
      RECT 19158.53 9765.78 19159.29 9766.08 ;
      RECT 19158.99 9764.87 19159.29 9766.08 ;
      RECT 19161.62 9764.82 19162.43 9765.16 ;
      RECT 19161.62 9782.05 19162.43 9782.39 ;
      RECT 19158.99 9781.13 19159.29 9782.34 ;
      RECT 19161.62 9781.13 19161.92 9782.39 ;
      RECT 19163.87 9777.16 19164.17 9781.43 ;
      RECT 19161.16 9781.13 19161.92 9781.43 ;
      RECT 19158.53 9781.13 19159.29 9781.43 ;
      RECT 19161.16 9777.16 19161.54 9781.43 ;
      RECT 19158.53 9777.16 19158.83 9781.43 ;
      RECT 19152 9778.795 19164.965 9779.795 ;
      RECT 19161.16 9777.16 19161.92 9777.46 ;
      RECT 19161.62 9776.2 19161.92 9777.46 ;
      RECT 19158.53 9777.16 19159.29 9777.46 ;
      RECT 19158.99 9776.25 19159.29 9777.46 ;
      RECT 19161.62 9776.2 19162.43 9776.54 ;
      RECT 19161.62 9793.43 19162.43 9793.77 ;
      RECT 19158.99 9792.51 19159.29 9793.72 ;
      RECT 19161.62 9792.51 19161.92 9793.77 ;
      RECT 19163.87 9788.54 19164.17 9792.81 ;
      RECT 19161.16 9792.51 19161.92 9792.81 ;
      RECT 19158.53 9792.51 19159.29 9792.81 ;
      RECT 19161.16 9788.54 19161.54 9792.81 ;
      RECT 19158.53 9788.54 19158.83 9792.81 ;
      RECT 19152 9790.175 19164.965 9791.175 ;
      RECT 19161.16 9788.54 19161.92 9788.84 ;
      RECT 19161.62 9787.58 19161.92 9788.84 ;
      RECT 19158.53 9788.54 19159.29 9788.84 ;
      RECT 19158.99 9787.63 19159.29 9788.84 ;
      RECT 19161.62 9787.58 19162.43 9787.92 ;
      RECT 19161.62 9804.81 19162.43 9805.15 ;
      RECT 19158.99 9803.89 19159.29 9805.1 ;
      RECT 19161.62 9803.89 19161.92 9805.15 ;
      RECT 19163.87 9799.92 19164.17 9804.19 ;
      RECT 19161.16 9803.89 19161.92 9804.19 ;
      RECT 19158.53 9803.89 19159.29 9804.19 ;
      RECT 19161.16 9799.92 19161.54 9804.19 ;
      RECT 19158.53 9799.92 19158.83 9804.19 ;
      RECT 19152 9801.555 19164.965 9802.555 ;
      RECT 19161.16 9799.92 19161.92 9800.22 ;
      RECT 19161.62 9798.96 19161.92 9800.22 ;
      RECT 19158.53 9799.92 19159.29 9800.22 ;
      RECT 19158.99 9799.01 19159.29 9800.22 ;
      RECT 19161.62 9798.96 19162.43 9799.3 ;
      RECT 19161.62 9816.19 19162.43 9816.53 ;
      RECT 19158.99 9815.27 19159.29 9816.48 ;
      RECT 19161.62 9815.27 19161.92 9816.53 ;
      RECT 19163.87 9811.3 19164.17 9815.57 ;
      RECT 19161.16 9815.27 19161.92 9815.57 ;
      RECT 19158.53 9815.27 19159.29 9815.57 ;
      RECT 19161.16 9811.3 19161.54 9815.57 ;
      RECT 19158.53 9811.3 19158.83 9815.57 ;
      RECT 19152 9812.935 19164.965 9813.935 ;
      RECT 19161.16 9811.3 19161.92 9811.6 ;
      RECT 19161.62 9810.34 19161.92 9811.6 ;
      RECT 19158.53 9811.3 19159.29 9811.6 ;
      RECT 19158.99 9810.39 19159.29 9811.6 ;
      RECT 19161.62 9810.34 19162.43 9810.68 ;
      RECT 19161.62 9827.57 19162.43 9827.91 ;
      RECT 19158.99 9826.65 19159.29 9827.86 ;
      RECT 19161.62 9826.65 19161.92 9827.91 ;
      RECT 19163.87 9822.68 19164.17 9826.95 ;
      RECT 19161.16 9826.65 19161.92 9826.95 ;
      RECT 19158.53 9826.65 19159.29 9826.95 ;
      RECT 19161.16 9822.68 19161.54 9826.95 ;
      RECT 19158.53 9822.68 19158.83 9826.95 ;
      RECT 19152 9824.315 19164.965 9825.315 ;
      RECT 19161.16 9822.68 19161.92 9822.98 ;
      RECT 19161.62 9821.72 19161.92 9822.98 ;
      RECT 19158.53 9822.68 19159.29 9822.98 ;
      RECT 19158.99 9821.77 19159.29 9822.98 ;
      RECT 19161.62 9821.72 19162.43 9822.06 ;
      RECT 19161.62 9845.15 19162.43 9845.49 ;
      RECT 19158.99 9844.23 19159.29 9845.44 ;
      RECT 19161.62 9844.23 19161.92 9845.49 ;
      RECT 19163.87 9840.26 19164.17 9844.53 ;
      RECT 19161.16 9844.23 19161.92 9844.53 ;
      RECT 19158.53 9844.23 19159.29 9844.53 ;
      RECT 19161.16 9840.26 19161.54 9844.53 ;
      RECT 19158.53 9840.26 19158.83 9844.53 ;
      RECT 19152 9841.895 19164.965 9842.895 ;
      RECT 19161.16 9840.26 19161.92 9840.56 ;
      RECT 19161.62 9839.3 19161.92 9840.56 ;
      RECT 19158.53 9840.26 19159.29 9840.56 ;
      RECT 19158.99 9839.35 19159.29 9840.56 ;
      RECT 19161.62 9839.3 19162.43 9839.64 ;
      RECT 19161.62 9856.53 19162.43 9856.87 ;
      RECT 19158.99 9855.61 19159.29 9856.82 ;
      RECT 19161.62 9855.61 19161.92 9856.87 ;
      RECT 19163.87 9851.64 19164.17 9855.91 ;
      RECT 19161.16 9855.61 19161.92 9855.91 ;
      RECT 19158.53 9855.61 19159.29 9855.91 ;
      RECT 19161.16 9851.64 19161.54 9855.91 ;
      RECT 19158.53 9851.64 19158.83 9855.91 ;
      RECT 19152 9853.275 19164.965 9854.275 ;
      RECT 19161.16 9851.64 19161.92 9851.94 ;
      RECT 19161.62 9850.68 19161.92 9851.94 ;
      RECT 19158.53 9851.64 19159.29 9851.94 ;
      RECT 19158.99 9850.73 19159.29 9851.94 ;
      RECT 19161.62 9850.68 19162.43 9851.02 ;
      RECT 19161.62 9867.91 19162.43 9868.25 ;
      RECT 19158.99 9866.99 19159.29 9868.2 ;
      RECT 19161.62 9866.99 19161.92 9868.25 ;
      RECT 19163.87 9863.02 19164.17 9867.29 ;
      RECT 19161.16 9866.99 19161.92 9867.29 ;
      RECT 19158.53 9866.99 19159.29 9867.29 ;
      RECT 19161.16 9863.02 19161.54 9867.29 ;
      RECT 19158.53 9863.02 19158.83 9867.29 ;
      RECT 19152 9864.655 19164.965 9865.655 ;
      RECT 19161.16 9863.02 19161.92 9863.32 ;
      RECT 19161.62 9862.06 19161.92 9863.32 ;
      RECT 19158.53 9863.02 19159.29 9863.32 ;
      RECT 19158.99 9862.11 19159.29 9863.32 ;
      RECT 19161.62 9862.06 19162.43 9862.4 ;
      RECT 19161.62 9879.29 19162.43 9879.63 ;
      RECT 19158.99 9878.37 19159.29 9879.58 ;
      RECT 19161.62 9878.37 19161.92 9879.63 ;
      RECT 19163.87 9874.4 19164.17 9878.67 ;
      RECT 19161.16 9878.37 19161.92 9878.67 ;
      RECT 19158.53 9878.37 19159.29 9878.67 ;
      RECT 19161.16 9874.4 19161.54 9878.67 ;
      RECT 19158.53 9874.4 19158.83 9878.67 ;
      RECT 19152 9876.035 19164.965 9877.035 ;
      RECT 19161.16 9874.4 19161.92 9874.7 ;
      RECT 19161.62 9873.44 19161.92 9874.7 ;
      RECT 19158.53 9874.4 19159.29 9874.7 ;
      RECT 19158.99 9873.49 19159.29 9874.7 ;
      RECT 19161.62 9873.44 19162.43 9873.78 ;
      RECT 19161.62 9890.67 19162.43 9891.01 ;
      RECT 19158.99 9889.75 19159.29 9890.96 ;
      RECT 19161.62 9889.75 19161.92 9891.01 ;
      RECT 19163.87 9885.78 19164.17 9890.05 ;
      RECT 19161.16 9889.75 19161.92 9890.05 ;
      RECT 19158.53 9889.75 19159.29 9890.05 ;
      RECT 19161.16 9885.78 19161.54 9890.05 ;
      RECT 19158.53 9885.78 19158.83 9890.05 ;
      RECT 19152 9887.415 19164.965 9888.415 ;
      RECT 19161.16 9885.78 19161.92 9886.08 ;
      RECT 19161.62 9884.82 19161.92 9886.08 ;
      RECT 19158.53 9885.78 19159.29 9886.08 ;
      RECT 19158.99 9884.87 19159.29 9886.08 ;
      RECT 19161.62 9884.82 19162.43 9885.16 ;
      RECT 19161.62 9902.05 19162.43 9902.39 ;
      RECT 19158.99 9901.13 19159.29 9902.34 ;
      RECT 19161.62 9901.13 19161.92 9902.39 ;
      RECT 19163.87 9897.16 19164.17 9901.43 ;
      RECT 19161.16 9901.13 19161.92 9901.43 ;
      RECT 19158.53 9901.13 19159.29 9901.43 ;
      RECT 19161.16 9897.16 19161.54 9901.43 ;
      RECT 19158.53 9897.16 19158.83 9901.43 ;
      RECT 19152 9898.795 19164.965 9899.795 ;
      RECT 19161.16 9897.16 19161.92 9897.46 ;
      RECT 19161.62 9896.2 19161.92 9897.46 ;
      RECT 19158.53 9897.16 19159.29 9897.46 ;
      RECT 19158.99 9896.25 19159.29 9897.46 ;
      RECT 19161.62 9896.2 19162.43 9896.54 ;
      RECT 19161.62 9913.43 19162.43 9913.77 ;
      RECT 19158.99 9912.51 19159.29 9913.72 ;
      RECT 19161.62 9912.51 19161.92 9913.77 ;
      RECT 19163.87 9908.54 19164.17 9912.81 ;
      RECT 19161.16 9912.51 19161.92 9912.81 ;
      RECT 19158.53 9912.51 19159.29 9912.81 ;
      RECT 19161.16 9908.54 19161.54 9912.81 ;
      RECT 19158.53 9908.54 19158.83 9912.81 ;
      RECT 19152 9910.175 19164.965 9911.175 ;
      RECT 19161.16 9908.54 19161.92 9908.84 ;
      RECT 19161.62 9907.58 19161.92 9908.84 ;
      RECT 19158.53 9908.54 19159.29 9908.84 ;
      RECT 19158.99 9907.63 19159.29 9908.84 ;
      RECT 19161.62 9907.58 19162.43 9907.92 ;
      RECT 19161.62 9924.81 19162.43 9925.15 ;
      RECT 19158.99 9923.89 19159.29 9925.1 ;
      RECT 19161.62 9923.89 19161.92 9925.15 ;
      RECT 19163.87 9919.92 19164.17 9924.19 ;
      RECT 19161.16 9923.89 19161.92 9924.19 ;
      RECT 19158.53 9923.89 19159.29 9924.19 ;
      RECT 19161.16 9919.92 19161.54 9924.19 ;
      RECT 19158.53 9919.92 19158.83 9924.19 ;
      RECT 19152 9921.555 19164.965 9922.555 ;
      RECT 19161.16 9919.92 19161.92 9920.22 ;
      RECT 19161.62 9918.96 19161.92 9920.22 ;
      RECT 19158.53 9919.92 19159.29 9920.22 ;
      RECT 19158.99 9919.01 19159.29 9920.22 ;
      RECT 19161.62 9918.96 19162.43 9919.3 ;
      RECT 19161.62 9936.19 19162.43 9936.53 ;
      RECT 19158.99 9935.27 19159.29 9936.48 ;
      RECT 19161.62 9935.27 19161.92 9936.53 ;
      RECT 19163.87 9931.3 19164.17 9935.57 ;
      RECT 19161.16 9935.27 19161.92 9935.57 ;
      RECT 19158.53 9935.27 19159.29 9935.57 ;
      RECT 19161.16 9931.3 19161.54 9935.57 ;
      RECT 19158.53 9931.3 19158.83 9935.57 ;
      RECT 19152 9932.935 19164.965 9933.935 ;
      RECT 19161.16 9931.3 19161.92 9931.6 ;
      RECT 19161.62 9930.34 19161.92 9931.6 ;
      RECT 19158.53 9931.3 19159.29 9931.6 ;
      RECT 19158.99 9930.39 19159.29 9931.6 ;
      RECT 19161.62 9930.34 19162.43 9930.68 ;
      RECT 19161.62 9947.57 19162.43 9947.91 ;
      RECT 19158.99 9946.65 19159.29 9947.86 ;
      RECT 19161.62 9946.65 19161.92 9947.91 ;
      RECT 19163.87 9942.68 19164.17 9946.95 ;
      RECT 19161.16 9946.65 19161.92 9946.95 ;
      RECT 19158.53 9946.65 19159.29 9946.95 ;
      RECT 19161.16 9942.68 19161.54 9946.95 ;
      RECT 19158.53 9942.68 19158.83 9946.95 ;
      RECT 19152 9944.315 19164.965 9945.315 ;
      RECT 19161.16 9942.68 19161.92 9942.98 ;
      RECT 19161.62 9941.72 19161.92 9942.98 ;
      RECT 19158.53 9942.68 19159.29 9942.98 ;
      RECT 19158.99 9941.77 19159.29 9942.98 ;
      RECT 19161.62 9941.72 19162.43 9942.06 ;
      RECT 997.56 9479.62 998.37 9479.96 ;
      RECT 998.07 9478.7 998.37 9479.96 ;
      RECT 998.07 9478.7 998.83 9479 ;
      RECT 998.53 9476.66 998.83 9479 ;
      RECT 995.9 9476.66 996.2 9479 ;
      RECT 995.9 9476.66 1008 9477.66 ;
      RECT 997.56 9491 998.37 9491.34 ;
      RECT 998.07 9490.08 998.37 9491.34 ;
      RECT 998.07 9490.08 998.83 9490.38 ;
      RECT 998.53 9485.79 998.83 9490.38 ;
      RECT 995.9 9485.79 996.2 9490.38 ;
      RECT 995.035 9487.585 1008 9488.585 ;
      RECT 998.07 9485.79 998.83 9486.09 ;
      RECT 998.07 9484.83 998.37 9486.09 ;
      RECT 997.56 9484.83 998.37 9485.17 ;
      RECT 997.56 9502.38 998.37 9502.72 ;
      RECT 998.07 9501.46 998.37 9502.72 ;
      RECT 998.07 9501.46 998.83 9501.76 ;
      RECT 998.53 9497.17 998.83 9501.76 ;
      RECT 995.9 9497.17 996.2 9501.76 ;
      RECT 995.035 9498.965 1008 9499.965 ;
      RECT 998.07 9497.17 998.83 9497.47 ;
      RECT 998.07 9496.21 998.37 9497.47 ;
      RECT 997.56 9496.21 998.37 9496.55 ;
      RECT 997.56 9513.76 998.37 9514.1 ;
      RECT 998.07 9512.84 998.37 9514.1 ;
      RECT 998.07 9512.84 998.83 9513.14 ;
      RECT 998.53 9508.55 998.83 9513.14 ;
      RECT 995.9 9508.55 996.2 9513.14 ;
      RECT 995.035 9510.345 1008 9511.345 ;
      RECT 998.07 9508.55 998.83 9508.85 ;
      RECT 998.07 9507.59 998.37 9508.85 ;
      RECT 997.56 9507.59 998.37 9507.93 ;
      RECT 997.56 9525.14 998.37 9525.48 ;
      RECT 998.07 9524.22 998.37 9525.48 ;
      RECT 998.07 9524.22 998.83 9524.52 ;
      RECT 998.53 9519.93 998.83 9524.52 ;
      RECT 995.9 9519.93 996.2 9524.52 ;
      RECT 995.035 9521.725 1008 9522.725 ;
      RECT 998.07 9519.93 998.83 9520.23 ;
      RECT 998.07 9518.97 998.37 9520.23 ;
      RECT 997.56 9518.97 998.37 9519.31 ;
      RECT 997.56 9536.52 998.37 9536.86 ;
      RECT 998.07 9535.6 998.37 9536.86 ;
      RECT 998.07 9535.6 998.83 9535.9 ;
      RECT 998.53 9531.31 998.83 9535.9 ;
      RECT 995.9 9531.31 996.2 9535.9 ;
      RECT 995.035 9533.105 1008 9534.105 ;
      RECT 998.07 9531.31 998.83 9531.61 ;
      RECT 998.07 9530.35 998.37 9531.61 ;
      RECT 997.56 9530.35 998.37 9530.69 ;
      RECT 997.56 9547.9 998.37 9548.24 ;
      RECT 998.07 9546.98 998.37 9548.24 ;
      RECT 998.07 9546.98 998.83 9547.28 ;
      RECT 998.53 9542.69 998.83 9547.28 ;
      RECT 995.9 9542.69 996.2 9547.28 ;
      RECT 995.035 9544.485 1008 9545.485 ;
      RECT 998.07 9542.69 998.83 9542.99 ;
      RECT 998.07 9541.73 998.37 9542.99 ;
      RECT 997.56 9541.73 998.37 9542.07 ;
      RECT 997.56 9559.28 998.37 9559.62 ;
      RECT 998.07 9558.36 998.37 9559.62 ;
      RECT 998.07 9558.36 998.83 9558.66 ;
      RECT 998.53 9554.07 998.83 9558.66 ;
      RECT 995.9 9554.07 996.2 9558.66 ;
      RECT 995.035 9555.865 1008 9556.865 ;
      RECT 998.07 9554.07 998.83 9554.37 ;
      RECT 998.07 9553.11 998.37 9554.37 ;
      RECT 997.56 9553.11 998.37 9553.45 ;
      RECT 997.56 9570.66 998.37 9571 ;
      RECT 998.07 9569.74 998.37 9571 ;
      RECT 998.07 9569.74 998.83 9570.04 ;
      RECT 998.53 9565.45 998.83 9570.04 ;
      RECT 995.9 9565.45 996.2 9570.04 ;
      RECT 995.035 9567.245 1008 9568.245 ;
      RECT 998.07 9565.45 998.83 9565.75 ;
      RECT 998.07 9564.49 998.37 9565.75 ;
      RECT 997.56 9564.49 998.37 9564.83 ;
      RECT 997.56 9582.04 998.37 9582.38 ;
      RECT 998.07 9581.12 998.37 9582.38 ;
      RECT 998.07 9581.12 998.83 9581.42 ;
      RECT 998.53 9576.83 998.83 9581.42 ;
      RECT 995.9 9576.83 996.2 9581.42 ;
      RECT 995.035 9578.625 1008 9579.625 ;
      RECT 998.07 9576.83 998.83 9577.13 ;
      RECT 998.07 9575.87 998.37 9577.13 ;
      RECT 997.56 9575.87 998.37 9576.21 ;
      RECT 995.035 9590.005 1008 9591.005 ;
      RECT 998.53 9588.21 998.83 9591.005 ;
      RECT 995.9 9588.21 996.2 9591.005 ;
      RECT 998.07 9588.21 998.83 9588.51 ;
      RECT 998.07 9587.25 998.37 9588.51 ;
      RECT 997.56 9587.25 998.37 9587.59 ;
      RECT 997.56 9599.62 998.37 9599.96 ;
      RECT 998.07 9598.7 998.37 9599.96 ;
      RECT 998.07 9598.7 998.83 9599 ;
      RECT 998.53 9596.66 998.83 9599 ;
      RECT 995.9 9596.66 996.2 9599 ;
      RECT 995.9 9596.66 1008 9597.66 ;
      RECT 997.56 9611 998.37 9611.34 ;
      RECT 998.07 9610.08 998.37 9611.34 ;
      RECT 998.07 9610.08 998.83 9610.38 ;
      RECT 998.53 9605.79 998.83 9610.38 ;
      RECT 995.9 9605.79 996.2 9610.38 ;
      RECT 995.035 9607.585 1008 9608.585 ;
      RECT 998.07 9605.79 998.83 9606.09 ;
      RECT 998.07 9604.83 998.37 9606.09 ;
      RECT 997.56 9604.83 998.37 9605.17 ;
      RECT 997.56 9622.38 998.37 9622.72 ;
      RECT 998.07 9621.46 998.37 9622.72 ;
      RECT 998.07 9621.46 998.83 9621.76 ;
      RECT 998.53 9617.17 998.83 9621.76 ;
      RECT 995.9 9617.17 996.2 9621.76 ;
      RECT 995.035 9618.965 1008 9619.965 ;
      RECT 998.07 9617.17 998.83 9617.47 ;
      RECT 998.07 9616.21 998.37 9617.47 ;
      RECT 997.56 9616.21 998.37 9616.55 ;
      RECT 997.56 9633.76 998.37 9634.1 ;
      RECT 998.07 9632.84 998.37 9634.1 ;
      RECT 998.07 9632.84 998.83 9633.14 ;
      RECT 998.53 9628.55 998.83 9633.14 ;
      RECT 995.9 9628.55 996.2 9633.14 ;
      RECT 995.035 9630.345 1008 9631.345 ;
      RECT 998.07 9628.55 998.83 9628.85 ;
      RECT 998.07 9627.59 998.37 9628.85 ;
      RECT 997.56 9627.59 998.37 9627.93 ;
      RECT 997.56 9645.14 998.37 9645.48 ;
      RECT 998.07 9644.22 998.37 9645.48 ;
      RECT 998.07 9644.22 998.83 9644.52 ;
      RECT 998.53 9639.93 998.83 9644.52 ;
      RECT 995.9 9639.93 996.2 9644.52 ;
      RECT 995.035 9641.725 1008 9642.725 ;
      RECT 998.07 9639.93 998.83 9640.23 ;
      RECT 998.07 9638.97 998.37 9640.23 ;
      RECT 997.56 9638.97 998.37 9639.31 ;
      RECT 997.56 9656.52 998.37 9656.86 ;
      RECT 998.07 9655.6 998.37 9656.86 ;
      RECT 998.07 9655.6 998.83 9655.9 ;
      RECT 998.53 9651.31 998.83 9655.9 ;
      RECT 995.9 9651.31 996.2 9655.9 ;
      RECT 995.035 9653.105 1008 9654.105 ;
      RECT 998.07 9651.31 998.83 9651.61 ;
      RECT 998.07 9650.35 998.37 9651.61 ;
      RECT 997.56 9650.35 998.37 9650.69 ;
      RECT 997.56 9667.9 998.37 9668.24 ;
      RECT 998.07 9666.98 998.37 9668.24 ;
      RECT 998.07 9666.98 998.83 9667.28 ;
      RECT 998.53 9662.69 998.83 9667.28 ;
      RECT 995.9 9662.69 996.2 9667.28 ;
      RECT 995.035 9664.485 1008 9665.485 ;
      RECT 998.07 9662.69 998.83 9662.99 ;
      RECT 998.07 9661.73 998.37 9662.99 ;
      RECT 997.56 9661.73 998.37 9662.07 ;
      RECT 997.56 9679.28 998.37 9679.62 ;
      RECT 998.07 9678.36 998.37 9679.62 ;
      RECT 998.07 9678.36 998.83 9678.66 ;
      RECT 998.53 9674.07 998.83 9678.66 ;
      RECT 995.9 9674.07 996.2 9678.66 ;
      RECT 995.035 9675.865 1008 9676.865 ;
      RECT 998.07 9674.07 998.83 9674.37 ;
      RECT 998.07 9673.11 998.37 9674.37 ;
      RECT 997.56 9673.11 998.37 9673.45 ;
      RECT 997.56 9690.66 998.37 9691 ;
      RECT 998.07 9689.74 998.37 9691 ;
      RECT 998.07 9689.74 998.83 9690.04 ;
      RECT 998.53 9685.45 998.83 9690.04 ;
      RECT 995.9 9685.45 996.2 9690.04 ;
      RECT 995.035 9687.245 1008 9688.245 ;
      RECT 998.07 9685.45 998.83 9685.75 ;
      RECT 998.07 9684.49 998.37 9685.75 ;
      RECT 997.56 9684.49 998.37 9684.83 ;
      RECT 997.56 9702.04 998.37 9702.38 ;
      RECT 998.07 9701.12 998.37 9702.38 ;
      RECT 998.07 9701.12 998.83 9701.42 ;
      RECT 998.53 9696.83 998.83 9701.42 ;
      RECT 995.9 9696.83 996.2 9701.42 ;
      RECT 995.035 9698.625 1008 9699.625 ;
      RECT 998.07 9696.83 998.83 9697.13 ;
      RECT 998.07 9695.87 998.37 9697.13 ;
      RECT 997.56 9695.87 998.37 9696.21 ;
      RECT 995.035 9710.005 1008 9711.005 ;
      RECT 998.53 9708.21 998.83 9711.005 ;
      RECT 995.9 9708.21 996.2 9711.005 ;
      RECT 998.07 9708.21 998.83 9708.51 ;
      RECT 998.07 9707.25 998.37 9708.51 ;
      RECT 997.56 9707.25 998.37 9707.59 ;
      RECT 997.56 9719.62 998.37 9719.96 ;
      RECT 998.07 9718.7 998.37 9719.96 ;
      RECT 998.07 9718.7 998.83 9719 ;
      RECT 998.53 9716.66 998.83 9719 ;
      RECT 995.9 9716.66 996.2 9719 ;
      RECT 995.9 9716.66 1008 9717.66 ;
      RECT 997.56 9731 998.37 9731.34 ;
      RECT 998.07 9730.08 998.37 9731.34 ;
      RECT 998.07 9730.08 998.83 9730.38 ;
      RECT 998.53 9725.79 998.83 9730.38 ;
      RECT 995.9 9725.79 996.2 9730.38 ;
      RECT 995.035 9727.585 1008 9728.585 ;
      RECT 998.07 9725.79 998.83 9726.09 ;
      RECT 998.07 9724.83 998.37 9726.09 ;
      RECT 997.56 9724.83 998.37 9725.17 ;
      RECT 997.56 9742.38 998.37 9742.72 ;
      RECT 998.07 9741.46 998.37 9742.72 ;
      RECT 998.07 9741.46 998.83 9741.76 ;
      RECT 998.53 9737.17 998.83 9741.76 ;
      RECT 995.9 9737.17 996.2 9741.76 ;
      RECT 995.035 9738.965 1008 9739.965 ;
      RECT 998.07 9737.17 998.83 9737.47 ;
      RECT 998.07 9736.21 998.37 9737.47 ;
      RECT 997.56 9736.21 998.37 9736.55 ;
      RECT 997.56 9753.76 998.37 9754.1 ;
      RECT 998.07 9752.84 998.37 9754.1 ;
      RECT 998.07 9752.84 998.83 9753.14 ;
      RECT 998.53 9748.55 998.83 9753.14 ;
      RECT 995.9 9748.55 996.2 9753.14 ;
      RECT 995.035 9750.345 1008 9751.345 ;
      RECT 998.07 9748.55 998.83 9748.85 ;
      RECT 998.07 9747.59 998.37 9748.85 ;
      RECT 997.56 9747.59 998.37 9747.93 ;
      RECT 997.56 9765.14 998.37 9765.48 ;
      RECT 998.07 9764.22 998.37 9765.48 ;
      RECT 998.07 9764.22 998.83 9764.52 ;
      RECT 998.53 9759.93 998.83 9764.52 ;
      RECT 995.9 9759.93 996.2 9764.52 ;
      RECT 995.035 9761.725 1008 9762.725 ;
      RECT 998.07 9759.93 998.83 9760.23 ;
      RECT 998.07 9758.97 998.37 9760.23 ;
      RECT 997.56 9758.97 998.37 9759.31 ;
      RECT 997.56 9776.52 998.37 9776.86 ;
      RECT 998.07 9775.6 998.37 9776.86 ;
      RECT 998.07 9775.6 998.83 9775.9 ;
      RECT 998.53 9771.31 998.83 9775.9 ;
      RECT 995.9 9771.31 996.2 9775.9 ;
      RECT 995.035 9773.105 1008 9774.105 ;
      RECT 998.07 9771.31 998.83 9771.61 ;
      RECT 998.07 9770.35 998.37 9771.61 ;
      RECT 997.56 9770.35 998.37 9770.69 ;
      RECT 997.56 9787.9 998.37 9788.24 ;
      RECT 998.07 9786.98 998.37 9788.24 ;
      RECT 998.07 9786.98 998.83 9787.28 ;
      RECT 998.53 9782.69 998.83 9787.28 ;
      RECT 995.9 9782.69 996.2 9787.28 ;
      RECT 995.035 9784.485 1008 9785.485 ;
      RECT 998.07 9782.69 998.83 9782.99 ;
      RECT 998.07 9781.73 998.37 9782.99 ;
      RECT 997.56 9781.73 998.37 9782.07 ;
      RECT 997.56 9799.28 998.37 9799.62 ;
      RECT 998.07 9798.36 998.37 9799.62 ;
      RECT 998.07 9798.36 998.83 9798.66 ;
      RECT 998.53 9794.07 998.83 9798.66 ;
      RECT 995.9 9794.07 996.2 9798.66 ;
      RECT 995.035 9795.865 1008 9796.865 ;
      RECT 998.07 9794.07 998.83 9794.37 ;
      RECT 998.07 9793.11 998.37 9794.37 ;
      RECT 997.56 9793.11 998.37 9793.45 ;
      RECT 997.56 9810.66 998.37 9811 ;
      RECT 998.07 9809.74 998.37 9811 ;
      RECT 998.07 9809.74 998.83 9810.04 ;
      RECT 998.53 9805.45 998.83 9810.04 ;
      RECT 995.9 9805.45 996.2 9810.04 ;
      RECT 995.035 9807.245 1008 9808.245 ;
      RECT 998.07 9805.45 998.83 9805.75 ;
      RECT 998.07 9804.49 998.37 9805.75 ;
      RECT 997.56 9804.49 998.37 9804.83 ;
      RECT 997.56 9822.04 998.37 9822.38 ;
      RECT 998.07 9821.12 998.37 9822.38 ;
      RECT 998.07 9821.12 998.83 9821.42 ;
      RECT 998.53 9816.83 998.83 9821.42 ;
      RECT 995.9 9816.83 996.2 9821.42 ;
      RECT 995.035 9818.625 1008 9819.625 ;
      RECT 998.07 9816.83 998.83 9817.13 ;
      RECT 998.07 9815.87 998.37 9817.13 ;
      RECT 997.56 9815.87 998.37 9816.21 ;
      RECT 995.035 9830.005 1008 9831.005 ;
      RECT 998.53 9828.21 998.83 9831.005 ;
      RECT 995.9 9828.21 996.2 9831.005 ;
      RECT 998.07 9828.21 998.83 9828.51 ;
      RECT 998.07 9827.25 998.37 9828.51 ;
      RECT 997.56 9827.25 998.37 9827.59 ;
      RECT 997.56 9839.62 998.37 9839.96 ;
      RECT 998.07 9838.7 998.37 9839.96 ;
      RECT 998.07 9838.7 998.83 9839 ;
      RECT 998.53 9836.66 998.83 9839 ;
      RECT 995.9 9836.66 996.2 9839 ;
      RECT 995.9 9836.66 1008 9837.66 ;
      RECT 997.56 9851 998.37 9851.34 ;
      RECT 998.07 9850.08 998.37 9851.34 ;
      RECT 998.07 9850.08 998.83 9850.38 ;
      RECT 998.53 9845.79 998.83 9850.38 ;
      RECT 995.9 9845.79 996.2 9850.38 ;
      RECT 995.035 9847.585 1008 9848.585 ;
      RECT 998.07 9845.79 998.83 9846.09 ;
      RECT 998.07 9844.83 998.37 9846.09 ;
      RECT 997.56 9844.83 998.37 9845.17 ;
      RECT 997.56 9862.38 998.37 9862.72 ;
      RECT 998.07 9861.46 998.37 9862.72 ;
      RECT 998.07 9861.46 998.83 9861.76 ;
      RECT 998.53 9857.17 998.83 9861.76 ;
      RECT 995.9 9857.17 996.2 9861.76 ;
      RECT 995.035 9858.965 1008 9859.965 ;
      RECT 998.07 9857.17 998.83 9857.47 ;
      RECT 998.07 9856.21 998.37 9857.47 ;
      RECT 997.56 9856.21 998.37 9856.55 ;
      RECT 997.56 9873.76 998.37 9874.1 ;
      RECT 998.07 9872.84 998.37 9874.1 ;
      RECT 998.07 9872.84 998.83 9873.14 ;
      RECT 998.53 9868.55 998.83 9873.14 ;
      RECT 995.9 9868.55 996.2 9873.14 ;
      RECT 995.035 9870.345 1008 9871.345 ;
      RECT 998.07 9868.55 998.83 9868.85 ;
      RECT 998.07 9867.59 998.37 9868.85 ;
      RECT 997.56 9867.59 998.37 9867.93 ;
      RECT 997.56 9885.14 998.37 9885.48 ;
      RECT 998.07 9884.22 998.37 9885.48 ;
      RECT 998.07 9884.22 998.83 9884.52 ;
      RECT 998.53 9879.93 998.83 9884.52 ;
      RECT 995.9 9879.93 996.2 9884.52 ;
      RECT 995.035 9881.725 1008 9882.725 ;
      RECT 998.07 9879.93 998.83 9880.23 ;
      RECT 998.07 9878.97 998.37 9880.23 ;
      RECT 997.56 9878.97 998.37 9879.31 ;
      RECT 997.56 9896.52 998.37 9896.86 ;
      RECT 998.07 9895.6 998.37 9896.86 ;
      RECT 998.07 9895.6 998.83 9895.9 ;
      RECT 998.53 9891.31 998.83 9895.9 ;
      RECT 995.9 9891.31 996.2 9895.9 ;
      RECT 995.035 9893.105 1008 9894.105 ;
      RECT 998.07 9891.31 998.83 9891.61 ;
      RECT 998.07 9890.35 998.37 9891.61 ;
      RECT 997.56 9890.35 998.37 9890.69 ;
      RECT 997.56 9907.9 998.37 9908.24 ;
      RECT 998.07 9906.98 998.37 9908.24 ;
      RECT 998.07 9906.98 998.83 9907.28 ;
      RECT 998.53 9902.69 998.83 9907.28 ;
      RECT 995.9 9902.69 996.2 9907.28 ;
      RECT 995.035 9904.485 1008 9905.485 ;
      RECT 998.07 9902.69 998.83 9902.99 ;
      RECT 998.07 9901.73 998.37 9902.99 ;
      RECT 997.56 9901.73 998.37 9902.07 ;
      RECT 997.56 9919.28 998.37 9919.62 ;
      RECT 998.07 9918.36 998.37 9919.62 ;
      RECT 998.07 9918.36 998.83 9918.66 ;
      RECT 998.53 9914.07 998.83 9918.66 ;
      RECT 995.9 9914.07 996.2 9918.66 ;
      RECT 995.035 9915.865 1008 9916.865 ;
      RECT 998.07 9914.07 998.83 9914.37 ;
      RECT 998.07 9913.11 998.37 9914.37 ;
      RECT 997.56 9913.11 998.37 9913.45 ;
      RECT 997.56 9930.66 998.37 9931 ;
      RECT 998.07 9929.74 998.37 9931 ;
      RECT 998.07 9929.74 998.83 9930.04 ;
      RECT 998.53 9925.45 998.83 9930.04 ;
      RECT 995.9 9925.45 996.2 9930.04 ;
      RECT 995.035 9927.245 1008 9928.245 ;
      RECT 998.07 9925.45 998.83 9925.75 ;
      RECT 998.07 9924.49 998.37 9925.75 ;
      RECT 997.56 9924.49 998.37 9924.83 ;
      RECT 997.56 9942.04 998.37 9942.38 ;
      RECT 998.07 9941.12 998.37 9942.38 ;
      RECT 998.07 9941.12 998.83 9941.42 ;
      RECT 998.53 9936.83 998.83 9941.42 ;
      RECT 995.9 9936.83 996.2 9941.42 ;
      RECT 995.035 9938.625 1008 9939.625 ;
      RECT 998.07 9936.83 998.83 9937.13 ;
      RECT 998.07 9935.87 998.37 9937.13 ;
      RECT 997.56 9935.87 998.37 9936.21 ;
      RECT 995.035 9950.005 1008 9951.005 ;
      RECT 998.53 9948.21 998.83 9951.005 ;
      RECT 995.9 9948.21 996.2 9951.005 ;
      RECT 998.07 9948.21 998.83 9948.51 ;
      RECT 998.07 9947.25 998.37 9948.51 ;
      RECT 997.56 9947.25 998.37 9947.59 ;
      RECT 996.36 9484.23 996.66 9485.44 ;
      RECT 998.61 9480.26 998.91 9484.53 ;
      RECT 995.9 9484.23 996.66 9484.53 ;
      RECT 995.9 9480.26 996.2 9484.53 ;
      RECT 992 9481.895 1004.965 9482.895 ;
      RECT 995.9 9480.26 996.66 9480.56 ;
      RECT 996.36 9479.35 996.66 9480.56 ;
      RECT 996.36 9495.61 996.66 9496.82 ;
      RECT 998.61 9491.64 998.91 9495.91 ;
      RECT 995.9 9495.61 996.66 9495.91 ;
      RECT 995.9 9491.64 996.2 9495.91 ;
      RECT 992 9493.275 1004.965 9494.275 ;
      RECT 995.9 9491.64 996.66 9491.94 ;
      RECT 996.36 9490.73 996.66 9491.94 ;
      RECT 996.36 9506.99 996.66 9508.2 ;
      RECT 998.61 9503.02 998.91 9507.29 ;
      RECT 995.9 9506.99 996.66 9507.29 ;
      RECT 995.9 9503.02 996.2 9507.29 ;
      RECT 992 9504.655 1004.965 9505.655 ;
      RECT 995.9 9503.02 996.66 9503.32 ;
      RECT 996.36 9502.11 996.66 9503.32 ;
      RECT 996.36 9518.37 996.66 9519.58 ;
      RECT 998.61 9514.4 998.91 9518.67 ;
      RECT 995.9 9518.37 996.66 9518.67 ;
      RECT 995.9 9514.4 996.2 9518.67 ;
      RECT 992 9516.035 1004.965 9517.035 ;
      RECT 995.9 9514.4 996.66 9514.7 ;
      RECT 996.36 9513.49 996.66 9514.7 ;
      RECT 996.36 9529.75 996.66 9530.96 ;
      RECT 998.61 9525.78 998.91 9530.05 ;
      RECT 995.9 9529.75 996.66 9530.05 ;
      RECT 995.9 9525.78 996.2 9530.05 ;
      RECT 992 9527.415 1004.965 9528.415 ;
      RECT 995.9 9525.78 996.66 9526.08 ;
      RECT 996.36 9524.87 996.66 9526.08 ;
      RECT 996.36 9541.13 996.66 9542.34 ;
      RECT 998.61 9537.16 998.91 9541.43 ;
      RECT 995.9 9541.13 996.66 9541.43 ;
      RECT 995.9 9537.16 996.2 9541.43 ;
      RECT 992 9538.795 1004.965 9539.795 ;
      RECT 995.9 9537.16 996.66 9537.46 ;
      RECT 996.36 9536.25 996.66 9537.46 ;
      RECT 996.36 9552.51 996.66 9553.72 ;
      RECT 998.61 9548.54 998.91 9552.81 ;
      RECT 995.9 9552.51 996.66 9552.81 ;
      RECT 995.9 9548.54 996.2 9552.81 ;
      RECT 992 9550.175 1004.965 9551.175 ;
      RECT 995.9 9548.54 996.66 9548.84 ;
      RECT 996.36 9547.63 996.66 9548.84 ;
      RECT 996.36 9563.89 996.66 9565.1 ;
      RECT 998.61 9559.92 998.91 9564.19 ;
      RECT 995.9 9563.89 996.66 9564.19 ;
      RECT 995.9 9559.92 996.2 9564.19 ;
      RECT 992 9561.555 1004.965 9562.555 ;
      RECT 995.9 9559.92 996.66 9560.22 ;
      RECT 996.36 9559.01 996.66 9560.22 ;
      RECT 996.36 9575.27 996.66 9576.48 ;
      RECT 998.61 9571.3 998.91 9575.57 ;
      RECT 995.9 9575.27 996.66 9575.57 ;
      RECT 995.9 9571.3 996.2 9575.57 ;
      RECT 992 9572.935 1004.965 9573.935 ;
      RECT 995.9 9571.3 996.66 9571.6 ;
      RECT 996.36 9570.39 996.66 9571.6 ;
      RECT 996.36 9586.65 996.66 9587.86 ;
      RECT 998.61 9582.68 998.91 9586.95 ;
      RECT 995.9 9586.65 996.66 9586.95 ;
      RECT 995.9 9582.68 996.2 9586.95 ;
      RECT 992 9584.315 1004.965 9585.315 ;
      RECT 995.9 9582.68 996.66 9582.98 ;
      RECT 996.36 9581.77 996.66 9582.98 ;
      RECT 996.36 9604.23 996.66 9605.44 ;
      RECT 998.61 9600.26 998.91 9604.53 ;
      RECT 995.9 9604.23 996.66 9604.53 ;
      RECT 995.9 9600.26 996.2 9604.53 ;
      RECT 992 9601.895 1004.965 9602.895 ;
      RECT 995.9 9600.26 996.66 9600.56 ;
      RECT 996.36 9599.35 996.66 9600.56 ;
      RECT 996.36 9615.61 996.66 9616.82 ;
      RECT 998.61 9611.64 998.91 9615.91 ;
      RECT 995.9 9615.61 996.66 9615.91 ;
      RECT 995.9 9611.64 996.2 9615.91 ;
      RECT 992 9613.275 1004.965 9614.275 ;
      RECT 995.9 9611.64 996.66 9611.94 ;
      RECT 996.36 9610.73 996.66 9611.94 ;
      RECT 996.36 9626.99 996.66 9628.2 ;
      RECT 998.61 9623.02 998.91 9627.29 ;
      RECT 995.9 9626.99 996.66 9627.29 ;
      RECT 995.9 9623.02 996.2 9627.29 ;
      RECT 992 9624.655 1004.965 9625.655 ;
      RECT 995.9 9623.02 996.66 9623.32 ;
      RECT 996.36 9622.11 996.66 9623.32 ;
      RECT 996.36 9638.37 996.66 9639.58 ;
      RECT 998.61 9634.4 998.91 9638.67 ;
      RECT 995.9 9638.37 996.66 9638.67 ;
      RECT 995.9 9634.4 996.2 9638.67 ;
      RECT 992 9636.035 1004.965 9637.035 ;
      RECT 995.9 9634.4 996.66 9634.7 ;
      RECT 996.36 9633.49 996.66 9634.7 ;
      RECT 996.36 9649.75 996.66 9650.96 ;
      RECT 998.61 9645.78 998.91 9650.05 ;
      RECT 995.9 9649.75 996.66 9650.05 ;
      RECT 995.9 9645.78 996.2 9650.05 ;
      RECT 992 9647.415 1004.965 9648.415 ;
      RECT 995.9 9645.78 996.66 9646.08 ;
      RECT 996.36 9644.87 996.66 9646.08 ;
      RECT 996.36 9661.13 996.66 9662.34 ;
      RECT 998.61 9657.16 998.91 9661.43 ;
      RECT 995.9 9661.13 996.66 9661.43 ;
      RECT 995.9 9657.16 996.2 9661.43 ;
      RECT 992 9658.795 1004.965 9659.795 ;
      RECT 995.9 9657.16 996.66 9657.46 ;
      RECT 996.36 9656.25 996.66 9657.46 ;
      RECT 996.36 9672.51 996.66 9673.72 ;
      RECT 998.61 9668.54 998.91 9672.81 ;
      RECT 995.9 9672.51 996.66 9672.81 ;
      RECT 995.9 9668.54 996.2 9672.81 ;
      RECT 992 9670.175 1004.965 9671.175 ;
      RECT 995.9 9668.54 996.66 9668.84 ;
      RECT 996.36 9667.63 996.66 9668.84 ;
      RECT 996.36 9683.89 996.66 9685.1 ;
      RECT 998.61 9679.92 998.91 9684.19 ;
      RECT 995.9 9683.89 996.66 9684.19 ;
      RECT 995.9 9679.92 996.2 9684.19 ;
      RECT 992 9681.555 1004.965 9682.555 ;
      RECT 995.9 9679.92 996.66 9680.22 ;
      RECT 996.36 9679.01 996.66 9680.22 ;
      RECT 996.36 9695.27 996.66 9696.48 ;
      RECT 998.61 9691.3 998.91 9695.57 ;
      RECT 995.9 9695.27 996.66 9695.57 ;
      RECT 995.9 9691.3 996.2 9695.57 ;
      RECT 992 9692.935 1004.965 9693.935 ;
      RECT 995.9 9691.3 996.66 9691.6 ;
      RECT 996.36 9690.39 996.66 9691.6 ;
      RECT 996.36 9706.65 996.66 9707.86 ;
      RECT 998.61 9702.68 998.91 9706.95 ;
      RECT 995.9 9706.65 996.66 9706.95 ;
      RECT 995.9 9702.68 996.2 9706.95 ;
      RECT 992 9704.315 1004.965 9705.315 ;
      RECT 995.9 9702.68 996.66 9702.98 ;
      RECT 996.36 9701.77 996.66 9702.98 ;
      RECT 996.36 9724.23 996.66 9725.44 ;
      RECT 998.61 9720.26 998.91 9724.53 ;
      RECT 995.9 9724.23 996.66 9724.53 ;
      RECT 995.9 9720.26 996.2 9724.53 ;
      RECT 992 9721.895 1004.965 9722.895 ;
      RECT 995.9 9720.26 996.66 9720.56 ;
      RECT 996.36 9719.35 996.66 9720.56 ;
      RECT 996.36 9735.61 996.66 9736.82 ;
      RECT 998.61 9731.64 998.91 9735.91 ;
      RECT 995.9 9735.61 996.66 9735.91 ;
      RECT 995.9 9731.64 996.2 9735.91 ;
      RECT 992 9733.275 1004.965 9734.275 ;
      RECT 995.9 9731.64 996.66 9731.94 ;
      RECT 996.36 9730.73 996.66 9731.94 ;
      RECT 996.36 9746.99 996.66 9748.2 ;
      RECT 998.61 9743.02 998.91 9747.29 ;
      RECT 995.9 9746.99 996.66 9747.29 ;
      RECT 995.9 9743.02 996.2 9747.29 ;
      RECT 992 9744.655 1004.965 9745.655 ;
      RECT 995.9 9743.02 996.66 9743.32 ;
      RECT 996.36 9742.11 996.66 9743.32 ;
      RECT 996.36 9758.37 996.66 9759.58 ;
      RECT 998.61 9754.4 998.91 9758.67 ;
      RECT 995.9 9758.37 996.66 9758.67 ;
      RECT 995.9 9754.4 996.2 9758.67 ;
      RECT 992 9756.035 1004.965 9757.035 ;
      RECT 995.9 9754.4 996.66 9754.7 ;
      RECT 996.36 9753.49 996.66 9754.7 ;
      RECT 996.36 9769.75 996.66 9770.96 ;
      RECT 998.61 9765.78 998.91 9770.05 ;
      RECT 995.9 9769.75 996.66 9770.05 ;
      RECT 995.9 9765.78 996.2 9770.05 ;
      RECT 992 9767.415 1004.965 9768.415 ;
      RECT 995.9 9765.78 996.66 9766.08 ;
      RECT 996.36 9764.87 996.66 9766.08 ;
      RECT 996.36 9781.13 996.66 9782.34 ;
      RECT 998.61 9777.16 998.91 9781.43 ;
      RECT 995.9 9781.13 996.66 9781.43 ;
      RECT 995.9 9777.16 996.2 9781.43 ;
      RECT 992 9778.795 1004.965 9779.795 ;
      RECT 995.9 9777.16 996.66 9777.46 ;
      RECT 996.36 9776.25 996.66 9777.46 ;
      RECT 996.36 9792.51 996.66 9793.72 ;
      RECT 998.61 9788.54 998.91 9792.81 ;
      RECT 995.9 9792.51 996.66 9792.81 ;
      RECT 995.9 9788.54 996.2 9792.81 ;
      RECT 992 9790.175 1004.965 9791.175 ;
      RECT 995.9 9788.54 996.66 9788.84 ;
      RECT 996.36 9787.63 996.66 9788.84 ;
      RECT 996.36 9803.89 996.66 9805.1 ;
      RECT 998.61 9799.92 998.91 9804.19 ;
      RECT 995.9 9803.89 996.66 9804.19 ;
      RECT 995.9 9799.92 996.2 9804.19 ;
      RECT 992 9801.555 1004.965 9802.555 ;
      RECT 995.9 9799.92 996.66 9800.22 ;
      RECT 996.36 9799.01 996.66 9800.22 ;
      RECT 996.36 9815.27 996.66 9816.48 ;
      RECT 998.61 9811.3 998.91 9815.57 ;
      RECT 995.9 9815.27 996.66 9815.57 ;
      RECT 995.9 9811.3 996.2 9815.57 ;
      RECT 992 9812.935 1004.965 9813.935 ;
      RECT 995.9 9811.3 996.66 9811.6 ;
      RECT 996.36 9810.39 996.66 9811.6 ;
      RECT 996.36 9826.65 996.66 9827.86 ;
      RECT 998.61 9822.68 998.91 9826.95 ;
      RECT 995.9 9826.65 996.66 9826.95 ;
      RECT 995.9 9822.68 996.2 9826.95 ;
      RECT 992 9824.315 1004.965 9825.315 ;
      RECT 995.9 9822.68 996.66 9822.98 ;
      RECT 996.36 9821.77 996.66 9822.98 ;
      RECT 996.36 9844.23 996.66 9845.44 ;
      RECT 998.61 9840.26 998.91 9844.53 ;
      RECT 995.9 9844.23 996.66 9844.53 ;
      RECT 995.9 9840.26 996.2 9844.53 ;
      RECT 992 9841.895 1004.965 9842.895 ;
      RECT 995.9 9840.26 996.66 9840.56 ;
      RECT 996.36 9839.35 996.66 9840.56 ;
      RECT 996.36 9855.61 996.66 9856.82 ;
      RECT 998.61 9851.64 998.91 9855.91 ;
      RECT 995.9 9855.61 996.66 9855.91 ;
      RECT 995.9 9851.64 996.2 9855.91 ;
      RECT 992 9853.275 1004.965 9854.275 ;
      RECT 995.9 9851.64 996.66 9851.94 ;
      RECT 996.36 9850.73 996.66 9851.94 ;
      RECT 996.36 9866.99 996.66 9868.2 ;
      RECT 998.61 9863.02 998.91 9867.29 ;
      RECT 995.9 9866.99 996.66 9867.29 ;
      RECT 995.9 9863.02 996.2 9867.29 ;
      RECT 992 9864.655 1004.965 9865.655 ;
      RECT 995.9 9863.02 996.66 9863.32 ;
      RECT 996.36 9862.11 996.66 9863.32 ;
      RECT 996.36 9878.37 996.66 9879.58 ;
      RECT 998.61 9874.4 998.91 9878.67 ;
      RECT 995.9 9878.37 996.66 9878.67 ;
      RECT 995.9 9874.4 996.2 9878.67 ;
      RECT 992 9876.035 1004.965 9877.035 ;
      RECT 995.9 9874.4 996.66 9874.7 ;
      RECT 996.36 9873.49 996.66 9874.7 ;
      RECT 996.36 9889.75 996.66 9890.96 ;
      RECT 998.61 9885.78 998.91 9890.05 ;
      RECT 995.9 9889.75 996.66 9890.05 ;
      RECT 995.9 9885.78 996.2 9890.05 ;
      RECT 992 9887.415 1004.965 9888.415 ;
      RECT 995.9 9885.78 996.66 9886.08 ;
      RECT 996.36 9884.87 996.66 9886.08 ;
      RECT 996.36 9901.13 996.66 9902.34 ;
      RECT 998.61 9897.16 998.91 9901.43 ;
      RECT 995.9 9901.13 996.66 9901.43 ;
      RECT 995.9 9897.16 996.2 9901.43 ;
      RECT 992 9898.795 1004.965 9899.795 ;
      RECT 995.9 9897.16 996.66 9897.46 ;
      RECT 996.36 9896.25 996.66 9897.46 ;
      RECT 996.36 9912.51 996.66 9913.72 ;
      RECT 998.61 9908.54 998.91 9912.81 ;
      RECT 995.9 9912.51 996.66 9912.81 ;
      RECT 995.9 9908.54 996.2 9912.81 ;
      RECT 992 9910.175 1004.965 9911.175 ;
      RECT 995.9 9908.54 996.66 9908.84 ;
      RECT 996.36 9907.63 996.66 9908.84 ;
      RECT 996.36 9923.89 996.66 9925.1 ;
      RECT 998.61 9919.92 998.91 9924.19 ;
      RECT 995.9 9923.89 996.66 9924.19 ;
      RECT 995.9 9919.92 996.2 9924.19 ;
      RECT 992 9921.555 1004.965 9922.555 ;
      RECT 995.9 9919.92 996.66 9920.22 ;
      RECT 996.36 9919.01 996.66 9920.22 ;
      RECT 996.36 9935.27 996.66 9936.48 ;
      RECT 998.61 9931.3 998.91 9935.57 ;
      RECT 995.9 9935.27 996.66 9935.57 ;
      RECT 995.9 9931.3 996.2 9935.57 ;
      RECT 992 9932.935 1004.965 9933.935 ;
      RECT 995.9 9931.3 996.66 9931.6 ;
      RECT 996.36 9930.39 996.66 9931.6 ;
      RECT 996.36 9946.65 996.66 9947.86 ;
      RECT 998.61 9942.68 998.91 9946.95 ;
      RECT 995.9 9946.65 996.66 9946.95 ;
      RECT 995.9 9942.68 996.2 9946.95 ;
      RECT 992 9944.315 1004.965 9945.315 ;
      RECT 995.9 9942.68 996.66 9942.98 ;
      RECT 996.36 9941.77 996.66 9942.98 ;
    LAYER M1 SPACING 0.23 ;
      RECT 998.1 1046.435 19161.9 10000 ;
    LAYER M2 ;
      RECT 0.5 9996.5 20199.5 9999.5 ;
      RECT 20196.5 0.5 20199.5 9999.5 ;
      RECT 0.5 0.5 3.5 9999.5 ;
      RECT 0.5 0.5 20199.5 3.5 ;
      RECT 4.1 9990 20195.9 9995.9 ;
      RECT 20190 4.1 20195.9 9995.9 ;
      RECT 19150 9953.565 19170 9995.9 ;
      RECT 990 9953.565 1010 9995.9 ;
      RECT 4.1 4.1 10 9995.9 ;
      RECT 4.1 4.1 20195.9 10 ;
      RECT 10100.705 1048.035 10102.645 1048.22 ;
      RECT 10102.555 1047.94 10102.645 1048.22 ;
      RECT 10100.705 1047.94 10100.795 1048.22 ;
      RECT 19157.85 1363.955 19429.88 1365.955 ;
      RECT 19157.85 1366.935 19429.88 1368.935 ;
      RECT 19146.565 9441.09 19352.21 9442.51 ;
      RECT 19146.565 9402.575 19335.79 9403.995 ;
      RECT 19146.565 9369.09 19319.37 9370.51 ;
      RECT 19146.565 9330.58 19302.95 9332 ;
      RECT 19146.565 9297.09 19286.53 9298.51 ;
      RECT 19158.16 1126.185 19277.57 1127.385 ;
      RECT 19146.565 9258.575 19270.11 9259.995 ;
      RECT 19158.16 1123.785 19261.37 1124.985 ;
      RECT 19158.16 1121.385 19245.17 1122.585 ;
      RECT 19158.16 1118.985 19228.97 1120.185 ;
      RECT 19150 9497.56 19170 9527.56 ;
      RECT 19150 9529.56 19170 9559.56 ;
      RECT 19150 9617.56 19170 9647.56 ;
      RECT 19150 9649.56 19170 9679.56 ;
      RECT 19150 9737.56 19170 9767.56 ;
      RECT 19150 9769.56 19170 9799.56 ;
      RECT 19150 9857.56 19170 9887.56 ;
      RECT 19150 9889.56 19170 9919.56 ;
      RECT 19155.875 1048.035 19156.155 1111.38 ;
      RECT 19155.315 1048.035 19155.595 1111.38 ;
      RECT 19154.755 1048.035 19155.035 1111.38 ;
      RECT 19154.195 1048.035 19154.475 1111.38 ;
      RECT 19153.635 1048.035 19153.915 1111.38 ;
      RECT 19153.075 1048.035 19153.355 1111.38 ;
      RECT 19152.515 1048.035 19152.795 1111.38 ;
      RECT 19151.955 1048.035 19152.235 1111.38 ;
      RECT 19027.955 1048.035 19028.235 1049.3 ;
      RECT 19024.315 1048.035 19024.595 1049.265 ;
      RECT 19020.675 1048.035 19020.955 1049.32 ;
      RECT 19017.035 1048.035 19017.315 1049.36 ;
      RECT 19013.395 1048.035 19013.675 1049.345 ;
      RECT 19009.755 1048.035 19010.035 1049.255 ;
      RECT 18950.675 1048.035 18950.955 1049.155 ;
      RECT 18946.755 1048.035 18947.035 1049.2 ;
      RECT 18942.835 1048.035 18943.115 1048.93 ;
      RECT 18938.915 1048.035 18939.195 1049.155 ;
      RECT 18934.995 1048.035 18935.275 1064.6 ;
      RECT 18887.955 1048.035 18888.235 1049.3 ;
      RECT 18884.315 1048.035 18884.595 1049.265 ;
      RECT 18880.675 1048.035 18880.955 1049.32 ;
      RECT 18877.035 1048.035 18877.315 1049.36 ;
      RECT 18873.395 1048.035 18873.675 1049.345 ;
      RECT 18869.755 1048.035 18870.035 1049.255 ;
      RECT 18810.675 1048.035 18810.955 1049.155 ;
      RECT 18806.755 1048.035 18807.035 1049.2 ;
      RECT 18802.835 1048.035 18803.115 1048.93 ;
      RECT 18798.915 1048.035 18799.195 1049.155 ;
      RECT 18794.995 1048.035 18795.275 1064.6 ;
      RECT 18747.955 1048.035 18748.235 1049.3 ;
      RECT 18744.315 1048.035 18744.595 1049.265 ;
      RECT 18740.675 1048.035 18740.955 1049.32 ;
      RECT 18737.035 1048.035 18737.315 1049.36 ;
      RECT 18733.395 1048.035 18733.675 1049.345 ;
      RECT 18729.755 1048.035 18730.035 1049.255 ;
      RECT 18670.675 1048.035 18670.955 1049.155 ;
      RECT 18666.755 1048.035 18667.035 1049.2 ;
      RECT 18662.835 1048.035 18663.115 1048.93 ;
      RECT 18658.915 1048.035 18659.195 1049.155 ;
      RECT 18654.995 1048.035 18655.275 1064.6 ;
      RECT 18607.955 1048.035 18608.235 1049.3 ;
      RECT 18604.315 1048.035 18604.595 1049.265 ;
      RECT 18600.675 1048.035 18600.955 1049.32 ;
      RECT 18597.035 1048.035 18597.315 1049.36 ;
      RECT 18593.395 1048.035 18593.675 1049.345 ;
      RECT 18589.755 1048.035 18590.035 1049.255 ;
      RECT 18530.675 1048.035 18530.955 1049.155 ;
      RECT 18526.755 1048.035 18527.035 1049.2 ;
      RECT 18522.835 1048.035 18523.115 1048.93 ;
      RECT 18518.915 1048.035 18519.195 1049.155 ;
      RECT 18514.995 1048.035 18515.275 1064.6 ;
      RECT 18467.955 1048.035 18468.235 1049.3 ;
      RECT 18464.315 1048.035 18464.595 1049.265 ;
      RECT 18460.675 1048.035 18460.955 1049.32 ;
      RECT 18457.035 1048.035 18457.315 1049.36 ;
      RECT 18453.395 1048.035 18453.675 1049.345 ;
      RECT 18449.755 1048.035 18450.035 1049.255 ;
      RECT 18390.675 1048.035 18390.955 1049.155 ;
      RECT 18386.755 1048.035 18387.035 1049.2 ;
      RECT 18382.835 1048.035 18383.115 1048.93 ;
      RECT 18378.915 1048.035 18379.195 1049.155 ;
      RECT 18374.995 1048.035 18375.275 1064.6 ;
      RECT 18327.955 1048.035 18328.235 1049.3 ;
      RECT 18324.315 1048.035 18324.595 1049.265 ;
      RECT 18320.675 1048.035 18320.955 1049.32 ;
      RECT 18317.035 1048.035 18317.315 1049.36 ;
      RECT 18313.395 1048.035 18313.675 1049.345 ;
      RECT 18309.755 1048.035 18310.035 1049.255 ;
      RECT 18250.675 1048.035 18250.955 1049.155 ;
      RECT 18246.755 1048.035 18247.035 1049.2 ;
      RECT 18242.835 1048.035 18243.115 1048.93 ;
      RECT 18238.915 1048.035 18239.195 1049.155 ;
      RECT 18234.995 1048.035 18235.275 1064.6 ;
      RECT 18187.955 1048.035 18188.235 1049.3 ;
      RECT 18184.315 1048.035 18184.595 1049.265 ;
      RECT 18180.675 1048.035 18180.955 1049.32 ;
      RECT 18177.035 1048.035 18177.315 1049.36 ;
      RECT 18173.395 1048.035 18173.675 1049.345 ;
      RECT 18169.755 1048.035 18170.035 1049.255 ;
      RECT 18110.675 1048.035 18110.955 1049.155 ;
      RECT 18106.755 1048.035 18107.035 1049.2 ;
      RECT 18102.835 1048.035 18103.115 1048.93 ;
      RECT 18098.915 1048.035 18099.195 1049.155 ;
      RECT 18094.995 1048.035 18095.275 1064.6 ;
      RECT 18047.955 1048.035 18048.235 1049.3 ;
      RECT 18044.315 1048.035 18044.595 1049.265 ;
      RECT 18040.675 1048.035 18040.955 1049.32 ;
      RECT 18037.035 1048.035 18037.315 1049.36 ;
      RECT 18033.395 1048.035 18033.675 1049.345 ;
      RECT 18029.755 1048.035 18030.035 1049.255 ;
      RECT 17970.675 1048.035 17970.955 1049.155 ;
      RECT 17966.755 1048.035 17967.035 1049.2 ;
      RECT 17962.835 1048.035 17963.115 1048.93 ;
      RECT 17958.915 1048.035 17959.195 1049.155 ;
      RECT 17954.995 1048.035 17955.275 1064.6 ;
      RECT 17907.955 1048.035 17908.235 1049.3 ;
      RECT 17904.315 1048.035 17904.595 1049.265 ;
      RECT 17900.675 1048.035 17900.955 1049.32 ;
      RECT 17897.035 1048.035 17897.315 1049.36 ;
      RECT 17893.395 1048.035 17893.675 1049.345 ;
      RECT 17889.755 1048.035 17890.035 1049.255 ;
      RECT 17830.675 1048.035 17830.955 1049.155 ;
      RECT 17826.755 1048.035 17827.035 1049.2 ;
      RECT 17822.835 1048.035 17823.115 1048.93 ;
      RECT 17818.915 1048.035 17819.195 1049.155 ;
      RECT 17814.995 1048.035 17815.275 1064.6 ;
      RECT 17767.955 1048.035 17768.235 1049.3 ;
      RECT 17764.315 1048.035 17764.595 1049.265 ;
      RECT 17760.675 1048.035 17760.955 1049.32 ;
      RECT 17757.035 1048.035 17757.315 1049.36 ;
      RECT 17753.395 1048.035 17753.675 1049.345 ;
      RECT 17749.755 1048.035 17750.035 1049.255 ;
      RECT 17690.675 1048.035 17690.955 1049.155 ;
      RECT 17686.755 1048.035 17687.035 1049.2 ;
      RECT 17682.835 1048.035 17683.115 1048.93 ;
      RECT 17678.915 1048.035 17679.195 1049.155 ;
      RECT 17674.995 1048.035 17675.275 1064.6 ;
      RECT 17627.955 1048.035 17628.235 1049.3 ;
      RECT 17624.315 1048.035 17624.595 1049.265 ;
      RECT 17620.675 1048.035 17620.955 1049.32 ;
      RECT 17617.035 1048.035 17617.315 1049.36 ;
      RECT 17613.395 1048.035 17613.675 1049.345 ;
      RECT 17609.755 1048.035 17610.035 1049.255 ;
      RECT 17550.675 1048.035 17550.955 1049.155 ;
      RECT 17546.755 1048.035 17547.035 1049.2 ;
      RECT 17542.835 1048.035 17543.115 1048.93 ;
      RECT 17538.915 1048.035 17539.195 1049.155 ;
      RECT 17534.995 1048.035 17535.275 1064.6 ;
      RECT 17487.955 1048.035 17488.235 1049.3 ;
      RECT 17484.315 1048.035 17484.595 1049.265 ;
      RECT 17480.675 1048.035 17480.955 1049.32 ;
      RECT 17477.035 1048.035 17477.315 1049.36 ;
      RECT 17473.395 1048.035 17473.675 1049.345 ;
      RECT 17469.755 1048.035 17470.035 1049.255 ;
      RECT 17410.675 1048.035 17410.955 1049.155 ;
      RECT 17406.755 1048.035 17407.035 1049.2 ;
      RECT 17402.835 1048.035 17403.115 1048.93 ;
      RECT 17398.915 1048.035 17399.195 1049.155 ;
      RECT 17394.995 1048.035 17395.275 1064.6 ;
      RECT 17347.955 1048.035 17348.235 1049.3 ;
      RECT 17344.315 1048.035 17344.595 1049.265 ;
      RECT 17340.675 1048.035 17340.955 1049.32 ;
      RECT 17337.035 1048.035 17337.315 1049.36 ;
      RECT 17333.395 1048.035 17333.675 1049.345 ;
      RECT 17329.755 1048.035 17330.035 1049.255 ;
      RECT 17270.675 1048.035 17270.955 1049.155 ;
      RECT 17266.755 1048.035 17267.035 1049.2 ;
      RECT 17262.835 1048.035 17263.115 1048.93 ;
      RECT 17258.915 1048.035 17259.195 1049.155 ;
      RECT 17254.995 1048.035 17255.275 1064.6 ;
      RECT 17207.955 1048.035 17208.235 1049.3 ;
      RECT 17204.315 1048.035 17204.595 1049.265 ;
      RECT 17200.675 1048.035 17200.955 1049.32 ;
      RECT 17197.035 1048.035 17197.315 1049.36 ;
      RECT 17193.395 1048.035 17193.675 1049.345 ;
      RECT 17189.755 1048.035 17190.035 1049.255 ;
      RECT 17130.675 1048.035 17130.955 1049.155 ;
      RECT 17126.755 1048.035 17127.035 1049.2 ;
      RECT 17122.835 1048.035 17123.115 1048.93 ;
      RECT 17118.915 1048.035 17119.195 1049.155 ;
      RECT 17114.995 1048.035 17115.275 1064.6 ;
      RECT 17067.955 1048.035 17068.235 1049.3 ;
      RECT 17064.315 1048.035 17064.595 1049.265 ;
      RECT 17060.675 1048.035 17060.955 1049.32 ;
      RECT 17057.035 1048.035 17057.315 1049.36 ;
      RECT 17053.395 1048.035 17053.675 1049.345 ;
      RECT 17049.755 1048.035 17050.035 1049.255 ;
      RECT 16990.675 1048.035 16990.955 1049.155 ;
      RECT 16986.755 1048.035 16987.035 1049.2 ;
      RECT 16982.835 1048.035 16983.115 1048.93 ;
      RECT 16978.915 1048.035 16979.195 1049.155 ;
      RECT 16974.995 1048.035 16975.275 1064.6 ;
      RECT 16927.955 1048.035 16928.235 1049.3 ;
      RECT 16924.315 1048.035 16924.595 1049.265 ;
      RECT 16920.675 1048.035 16920.955 1049.32 ;
      RECT 16917.035 1048.035 16917.315 1049.36 ;
      RECT 16913.395 1048.035 16913.675 1049.345 ;
      RECT 16909.755 1048.035 16910.035 1049.255 ;
      RECT 16850.675 1048.035 16850.955 1049.155 ;
      RECT 16846.755 1048.035 16847.035 1049.2 ;
      RECT 16842.835 1048.035 16843.115 1048.93 ;
      RECT 16838.915 1048.035 16839.195 1049.155 ;
      RECT 16834.995 1048.035 16835.275 1064.6 ;
      RECT 16787.955 1048.035 16788.235 1049.3 ;
      RECT 16784.315 1048.035 16784.595 1049.265 ;
      RECT 16780.675 1048.035 16780.955 1049.32 ;
      RECT 16777.035 1048.035 16777.315 1049.36 ;
      RECT 16773.395 1048.035 16773.675 1049.345 ;
      RECT 16769.755 1048.035 16770.035 1049.255 ;
      RECT 16710.675 1048.035 16710.955 1049.155 ;
      RECT 16706.755 1048.035 16707.035 1049.2 ;
      RECT 16702.835 1048.035 16703.115 1048.93 ;
      RECT 16698.915 1048.035 16699.195 1049.155 ;
      RECT 16694.995 1048.035 16695.275 1064.6 ;
      RECT 16647.955 1048.035 16648.235 1049.3 ;
      RECT 16644.315 1048.035 16644.595 1049.265 ;
      RECT 16640.675 1048.035 16640.955 1049.32 ;
      RECT 16637.035 1048.035 16637.315 1049.36 ;
      RECT 16633.395 1048.035 16633.675 1049.345 ;
      RECT 16629.755 1048.035 16630.035 1049.255 ;
      RECT 16570.675 1048.035 16570.955 1049.155 ;
      RECT 16566.755 1048.035 16567.035 1049.2 ;
      RECT 16562.835 1048.035 16563.115 1048.93 ;
      RECT 16558.915 1048.035 16559.195 1049.155 ;
      RECT 16554.995 1048.035 16555.275 1064.6 ;
      RECT 16507.955 1048.035 16508.235 1049.3 ;
      RECT 16504.315 1048.035 16504.595 1049.265 ;
      RECT 16500.675 1048.035 16500.955 1049.32 ;
      RECT 16497.035 1048.035 16497.315 1049.36 ;
      RECT 16493.395 1048.035 16493.675 1049.345 ;
      RECT 16489.755 1048.035 16490.035 1049.255 ;
      RECT 16430.675 1048.035 16430.955 1049.155 ;
      RECT 16426.755 1048.035 16427.035 1049.2 ;
      RECT 16422.835 1048.035 16423.115 1048.93 ;
      RECT 16418.915 1048.035 16419.195 1049.155 ;
      RECT 16414.995 1048.035 16415.275 1064.6 ;
      RECT 16367.955 1048.035 16368.235 1049.3 ;
      RECT 16364.315 1048.035 16364.595 1049.265 ;
      RECT 16360.675 1048.035 16360.955 1049.32 ;
      RECT 16357.035 1048.035 16357.315 1049.36 ;
      RECT 16353.395 1048.035 16353.675 1049.345 ;
      RECT 16349.755 1048.035 16350.035 1049.255 ;
      RECT 16290.675 1048.035 16290.955 1049.155 ;
      RECT 16286.755 1048.035 16287.035 1049.2 ;
      RECT 16282.835 1048.035 16283.115 1048.93 ;
      RECT 16278.915 1048.035 16279.195 1049.155 ;
      RECT 16274.995 1048.035 16275.275 1064.6 ;
      RECT 16227.955 1048.035 16228.235 1049.3 ;
      RECT 16224.315 1048.035 16224.595 1049.265 ;
      RECT 16220.675 1048.035 16220.955 1049.32 ;
      RECT 16217.035 1048.035 16217.315 1049.36 ;
      RECT 16213.395 1048.035 16213.675 1049.345 ;
      RECT 16209.755 1048.035 16210.035 1049.255 ;
      RECT 16150.675 1048.035 16150.955 1049.155 ;
      RECT 16146.755 1048.035 16147.035 1049.2 ;
      RECT 16142.835 1048.035 16143.115 1048.93 ;
      RECT 16138.915 1048.035 16139.195 1049.155 ;
      RECT 16134.995 1048.035 16135.275 1064.6 ;
      RECT 16087.955 1048.035 16088.235 1049.3 ;
      RECT 16084.315 1048.035 16084.595 1049.265 ;
      RECT 16080.675 1048.035 16080.955 1049.32 ;
      RECT 16077.035 1048.035 16077.315 1049.36 ;
      RECT 16073.395 1048.035 16073.675 1049.345 ;
      RECT 16069.755 1048.035 16070.035 1049.255 ;
      RECT 16010.675 1048.035 16010.955 1049.155 ;
      RECT 16006.755 1048.035 16007.035 1049.2 ;
      RECT 16002.835 1048.035 16003.115 1048.93 ;
      RECT 15998.915 1048.035 15999.195 1049.155 ;
      RECT 15994.995 1048.035 15995.275 1064.6 ;
      RECT 15947.955 1048.035 15948.235 1049.3 ;
      RECT 15944.315 1048.035 15944.595 1049.265 ;
      RECT 15940.675 1048.035 15940.955 1049.32 ;
      RECT 15937.035 1048.035 15937.315 1049.36 ;
      RECT 15933.395 1048.035 15933.675 1049.345 ;
      RECT 15929.755 1048.035 15930.035 1049.255 ;
      RECT 15870.675 1048.035 15870.955 1049.155 ;
      RECT 15866.755 1048.035 15867.035 1049.2 ;
      RECT 15862.835 1048.035 15863.115 1048.93 ;
      RECT 15858.915 1048.035 15859.195 1049.155 ;
      RECT 15854.995 1048.035 15855.275 1064.6 ;
      RECT 15807.955 1048.035 15808.235 1049.3 ;
      RECT 15804.315 1048.035 15804.595 1049.265 ;
      RECT 15800.675 1048.035 15800.955 1049.32 ;
      RECT 15797.035 1048.035 15797.315 1049.36 ;
      RECT 15793.395 1048.035 15793.675 1049.345 ;
      RECT 15789.755 1048.035 15790.035 1049.255 ;
      RECT 15730.675 1048.035 15730.955 1049.155 ;
      RECT 15726.755 1048.035 15727.035 1049.2 ;
      RECT 15722.835 1048.035 15723.115 1048.93 ;
      RECT 15718.915 1048.035 15719.195 1049.155 ;
      RECT 15714.995 1048.035 15715.275 1064.6 ;
      RECT 15667.955 1048.035 15668.235 1049.3 ;
      RECT 15664.315 1048.035 15664.595 1049.265 ;
      RECT 15660.675 1048.035 15660.955 1049.32 ;
      RECT 15657.035 1048.035 15657.315 1049.36 ;
      RECT 15653.395 1048.035 15653.675 1049.345 ;
      RECT 15649.755 1048.035 15650.035 1049.255 ;
      RECT 15590.675 1048.035 15590.955 1049.155 ;
      RECT 15586.755 1048.035 15587.035 1049.2 ;
      RECT 15582.835 1048.035 15583.115 1048.93 ;
      RECT 15578.915 1048.035 15579.195 1049.155 ;
      RECT 15574.995 1048.035 15575.275 1064.6 ;
      RECT 15527.955 1048.035 15528.235 1049.3 ;
      RECT 15524.315 1048.035 15524.595 1049.265 ;
      RECT 15520.675 1048.035 15520.955 1049.32 ;
      RECT 15517.035 1048.035 15517.315 1049.36 ;
      RECT 15513.395 1048.035 15513.675 1049.345 ;
      RECT 15509.755 1048.035 15510.035 1049.255 ;
      RECT 15450.675 1048.035 15450.955 1049.155 ;
      RECT 15446.755 1048.035 15447.035 1049.2 ;
      RECT 15442.835 1048.035 15443.115 1048.93 ;
      RECT 15438.915 1048.035 15439.195 1049.155 ;
      RECT 15434.995 1048.035 15435.275 1064.6 ;
      RECT 15387.955 1048.035 15388.235 1049.3 ;
      RECT 15384.315 1048.035 15384.595 1049.265 ;
      RECT 15380.675 1048.035 15380.955 1049.32 ;
      RECT 15377.035 1048.035 15377.315 1049.36 ;
      RECT 15373.395 1048.035 15373.675 1049.345 ;
      RECT 15369.755 1048.035 15370.035 1049.255 ;
      RECT 15310.675 1048.035 15310.955 1049.155 ;
      RECT 15306.755 1048.035 15307.035 1049.2 ;
      RECT 15302.835 1048.035 15303.115 1048.93 ;
      RECT 15298.915 1048.035 15299.195 1049.155 ;
      RECT 15294.995 1048.035 15295.275 1064.6 ;
      RECT 15247.955 1048.035 15248.235 1049.3 ;
      RECT 15244.315 1048.035 15244.595 1049.265 ;
      RECT 15240.675 1048.035 15240.955 1049.32 ;
      RECT 15237.035 1048.035 15237.315 1049.36 ;
      RECT 15233.395 1048.035 15233.675 1049.345 ;
      RECT 15229.755 1048.035 15230.035 1049.255 ;
      RECT 15170.675 1048.035 15170.955 1049.155 ;
      RECT 15166.755 1048.035 15167.035 1049.2 ;
      RECT 15162.835 1048.035 15163.115 1048.93 ;
      RECT 15158.915 1048.035 15159.195 1049.155 ;
      RECT 15154.995 1048.035 15155.275 1064.6 ;
      RECT 15107.955 1048.035 15108.235 1049.3 ;
      RECT 15104.315 1048.035 15104.595 1049.265 ;
      RECT 15100.675 1048.035 15100.955 1049.32 ;
      RECT 15097.035 1048.035 15097.315 1049.36 ;
      RECT 15093.395 1048.035 15093.675 1049.345 ;
      RECT 15089.755 1048.035 15090.035 1049.255 ;
      RECT 15030.675 1048.035 15030.955 1049.155 ;
      RECT 15026.755 1048.035 15027.035 1049.2 ;
      RECT 15022.835 1048.035 15023.115 1048.93 ;
      RECT 15018.915 1048.035 15019.195 1049.155 ;
      RECT 15014.995 1048.035 15015.275 1064.6 ;
      RECT 14967.955 1048.035 14968.235 1049.3 ;
      RECT 14964.315 1048.035 14964.595 1049.265 ;
      RECT 14960.675 1048.035 14960.955 1049.32 ;
      RECT 14957.035 1048.035 14957.315 1049.36 ;
      RECT 14953.395 1048.035 14953.675 1049.345 ;
      RECT 14949.755 1048.035 14950.035 1049.255 ;
      RECT 14890.675 1048.035 14890.955 1049.155 ;
      RECT 14886.755 1048.035 14887.035 1049.2 ;
      RECT 14882.835 1048.035 14883.115 1048.93 ;
      RECT 14878.915 1048.035 14879.195 1049.155 ;
      RECT 14874.995 1048.035 14875.275 1064.6 ;
      RECT 14827.955 1048.035 14828.235 1049.3 ;
      RECT 14824.315 1048.035 14824.595 1049.265 ;
      RECT 14820.675 1048.035 14820.955 1049.32 ;
      RECT 14817.035 1048.035 14817.315 1049.36 ;
      RECT 14813.395 1048.035 14813.675 1049.345 ;
      RECT 14809.755 1048.035 14810.035 1049.255 ;
      RECT 14750.675 1048.035 14750.955 1049.155 ;
      RECT 14746.755 1048.035 14747.035 1049.2 ;
      RECT 14742.835 1048.035 14743.115 1048.93 ;
      RECT 14738.915 1048.035 14739.195 1049.155 ;
      RECT 14734.995 1048.035 14735.275 1064.6 ;
      RECT 14687.955 1048.035 14688.235 1049.3 ;
      RECT 14684.315 1048.035 14684.595 1049.265 ;
      RECT 14680.675 1048.035 14680.955 1049.32 ;
      RECT 14677.035 1048.035 14677.315 1049.36 ;
      RECT 14673.395 1048.035 14673.675 1049.345 ;
      RECT 14669.755 1048.035 14670.035 1049.255 ;
      RECT 14610.675 1048.035 14610.955 1049.155 ;
      RECT 14606.755 1048.035 14607.035 1049.2 ;
      RECT 14602.835 1048.035 14603.115 1048.93 ;
      RECT 14598.915 1048.035 14599.195 1049.155 ;
      RECT 14594.995 1048.035 14595.275 1064.6 ;
      RECT 14547.955 1048.035 14548.235 1049.3 ;
      RECT 14544.315 1048.035 14544.595 1049.265 ;
      RECT 14540.675 1048.035 14540.955 1049.32 ;
      RECT 14537.035 1048.035 14537.315 1049.36 ;
      RECT 14533.395 1048.035 14533.675 1049.345 ;
      RECT 14529.755 1048.035 14530.035 1049.255 ;
      RECT 14470.675 1048.035 14470.955 1049.155 ;
      RECT 14466.755 1048.035 14467.035 1049.2 ;
      RECT 14462.835 1048.035 14463.115 1048.93 ;
      RECT 14458.915 1048.035 14459.195 1049.155 ;
      RECT 14454.995 1048.035 14455.275 1064.6 ;
      RECT 14407.955 1048.035 14408.235 1049.3 ;
      RECT 14404.315 1048.035 14404.595 1049.265 ;
      RECT 14400.675 1048.035 14400.955 1049.32 ;
      RECT 14397.035 1048.035 14397.315 1049.36 ;
      RECT 14393.395 1048.035 14393.675 1049.345 ;
      RECT 14389.755 1048.035 14390.035 1049.255 ;
      RECT 14330.675 1048.035 14330.955 1049.155 ;
      RECT 14326.755 1048.035 14327.035 1049.2 ;
      RECT 14322.835 1048.035 14323.115 1048.93 ;
      RECT 14318.915 1048.035 14319.195 1049.155 ;
      RECT 14314.995 1048.035 14315.275 1064.6 ;
      RECT 14267.955 1048.035 14268.235 1049.3 ;
      RECT 14264.315 1048.035 14264.595 1049.265 ;
      RECT 14260.675 1048.035 14260.955 1049.32 ;
      RECT 14257.035 1048.035 14257.315 1049.36 ;
      RECT 14253.395 1048.035 14253.675 1049.345 ;
      RECT 14249.755 1048.035 14250.035 1049.255 ;
      RECT 14190.675 1048.035 14190.955 1049.155 ;
      RECT 14186.755 1048.035 14187.035 1049.2 ;
      RECT 14182.835 1048.035 14183.115 1048.93 ;
      RECT 14178.915 1048.035 14179.195 1049.155 ;
      RECT 14174.995 1048.035 14175.275 1064.6 ;
      RECT 14127.955 1048.035 14128.235 1049.3 ;
      RECT 14124.315 1048.035 14124.595 1049.265 ;
      RECT 14120.675 1048.035 14120.955 1049.32 ;
      RECT 14117.035 1048.035 14117.315 1049.36 ;
      RECT 14113.395 1048.035 14113.675 1049.345 ;
      RECT 14109.755 1048.035 14110.035 1049.255 ;
      RECT 14050.675 1048.035 14050.955 1049.155 ;
      RECT 14046.755 1048.035 14047.035 1049.2 ;
      RECT 14042.835 1048.035 14043.115 1048.93 ;
      RECT 14038.915 1048.035 14039.195 1049.155 ;
      RECT 14034.995 1048.035 14035.275 1064.6 ;
      RECT 13987.955 1048.035 13988.235 1049.3 ;
      RECT 13984.315 1048.035 13984.595 1049.265 ;
      RECT 13980.675 1048.035 13980.955 1049.32 ;
      RECT 13977.035 1048.035 13977.315 1049.36 ;
      RECT 13973.395 1048.035 13973.675 1049.345 ;
      RECT 13969.755 1048.035 13970.035 1049.255 ;
      RECT 13910.675 1048.035 13910.955 1049.155 ;
      RECT 13906.755 1048.035 13907.035 1049.2 ;
      RECT 13902.835 1048.035 13903.115 1048.93 ;
      RECT 13898.915 1048.035 13899.195 1049.155 ;
      RECT 13894.995 1048.035 13895.275 1064.6 ;
      RECT 13847.955 1048.035 13848.235 1049.3 ;
      RECT 13844.315 1048.035 13844.595 1049.265 ;
      RECT 13840.675 1048.035 13840.955 1049.32 ;
      RECT 13837.035 1048.035 13837.315 1049.36 ;
      RECT 13833.395 1048.035 13833.675 1049.345 ;
      RECT 13829.755 1048.035 13830.035 1049.255 ;
      RECT 13770.675 1048.035 13770.955 1049.155 ;
      RECT 13766.755 1048.035 13767.035 1049.2 ;
      RECT 13762.835 1048.035 13763.115 1048.93 ;
      RECT 13758.915 1048.035 13759.195 1049.155 ;
      RECT 13754.995 1048.035 13755.275 1064.6 ;
      RECT 13707.955 1048.035 13708.235 1049.3 ;
      RECT 13704.315 1048.035 13704.595 1049.265 ;
      RECT 13700.675 1048.035 13700.955 1049.32 ;
      RECT 13697.035 1048.035 13697.315 1049.36 ;
      RECT 13693.395 1048.035 13693.675 1049.345 ;
      RECT 13689.755 1048.035 13690.035 1049.255 ;
      RECT 13630.675 1048.035 13630.955 1049.155 ;
      RECT 13626.755 1048.035 13627.035 1049.2 ;
      RECT 13622.835 1048.035 13623.115 1048.93 ;
      RECT 13618.915 1048.035 13619.195 1049.155 ;
      RECT 13614.995 1048.035 13615.275 1064.6 ;
      RECT 13567.955 1048.035 13568.235 1049.3 ;
      RECT 13564.315 1048.035 13564.595 1049.265 ;
      RECT 13560.675 1048.035 13560.955 1049.32 ;
      RECT 13557.035 1048.035 13557.315 1049.36 ;
      RECT 13553.395 1048.035 13553.675 1049.345 ;
      RECT 13549.755 1048.035 13550.035 1049.255 ;
      RECT 13490.675 1048.035 13490.955 1049.155 ;
      RECT 13486.755 1048.035 13487.035 1049.2 ;
      RECT 13482.835 1048.035 13483.115 1048.93 ;
      RECT 13478.915 1048.035 13479.195 1049.155 ;
      RECT 13474.995 1048.035 13475.275 1064.6 ;
      RECT 13427.955 1048.035 13428.235 1049.3 ;
      RECT 13424.315 1048.035 13424.595 1049.265 ;
      RECT 13420.675 1048.035 13420.955 1049.32 ;
      RECT 13417.035 1048.035 13417.315 1049.36 ;
      RECT 13413.395 1048.035 13413.675 1049.345 ;
      RECT 13409.755 1048.035 13410.035 1049.255 ;
      RECT 13350.675 1048.035 13350.955 1049.155 ;
      RECT 13346.755 1048.035 13347.035 1049.2 ;
      RECT 13342.835 1048.035 13343.115 1048.93 ;
      RECT 13338.915 1048.035 13339.195 1049.155 ;
      RECT 13334.995 1048.035 13335.275 1064.6 ;
      RECT 13287.955 1048.035 13288.235 1049.3 ;
      RECT 13284.315 1048.035 13284.595 1049.265 ;
      RECT 13280.675 1048.035 13280.955 1049.32 ;
      RECT 13277.035 1048.035 13277.315 1049.36 ;
      RECT 13273.395 1048.035 13273.675 1049.345 ;
      RECT 13269.755 1048.035 13270.035 1049.255 ;
      RECT 13210.675 1048.035 13210.955 1049.155 ;
      RECT 13206.755 1048.035 13207.035 1049.2 ;
      RECT 13202.835 1048.035 13203.115 1048.93 ;
      RECT 13198.915 1048.035 13199.195 1049.155 ;
      RECT 13194.995 1048.035 13195.275 1064.6 ;
      RECT 13147.955 1048.035 13148.235 1049.3 ;
      RECT 13144.315 1048.035 13144.595 1049.265 ;
      RECT 13140.675 1048.035 13140.955 1049.32 ;
      RECT 13137.035 1048.035 13137.315 1049.36 ;
      RECT 13133.395 1048.035 13133.675 1049.345 ;
      RECT 13129.755 1048.035 13130.035 1049.255 ;
      RECT 13070.675 1048.035 13070.955 1049.155 ;
      RECT 13066.755 1048.035 13067.035 1049.2 ;
      RECT 13062.835 1048.035 13063.115 1048.93 ;
      RECT 13058.915 1048.035 13059.195 1049.155 ;
      RECT 13054.995 1048.035 13055.275 1064.6 ;
      RECT 13007.955 1048.035 13008.235 1049.3 ;
      RECT 13004.315 1048.035 13004.595 1049.265 ;
      RECT 13000.675 1048.035 13000.955 1049.32 ;
      RECT 12997.035 1048.035 12997.315 1049.36 ;
      RECT 12993.395 1048.035 12993.675 1049.345 ;
      RECT 12989.755 1048.035 12990.035 1049.255 ;
      RECT 12930.675 1048.035 12930.955 1049.155 ;
      RECT 12926.755 1048.035 12927.035 1049.2 ;
      RECT 12922.835 1048.035 12923.115 1048.93 ;
      RECT 12918.915 1048.035 12919.195 1049.155 ;
      RECT 12914.995 1048.035 12915.275 1064.6 ;
      RECT 12867.955 1048.035 12868.235 1049.3 ;
      RECT 12864.315 1048.035 12864.595 1049.265 ;
      RECT 12860.675 1048.035 12860.955 1049.32 ;
      RECT 12857.035 1048.035 12857.315 1049.36 ;
      RECT 12853.395 1048.035 12853.675 1049.345 ;
      RECT 12849.755 1048.035 12850.035 1049.255 ;
      RECT 12790.675 1048.035 12790.955 1049.155 ;
      RECT 12786.755 1048.035 12787.035 1049.2 ;
      RECT 12782.835 1048.035 12783.115 1048.93 ;
      RECT 12778.915 1048.035 12779.195 1049.155 ;
      RECT 12774.995 1048.035 12775.275 1064.6 ;
      RECT 12727.955 1048.035 12728.235 1049.3 ;
      RECT 12724.315 1048.035 12724.595 1049.265 ;
      RECT 12720.675 1048.035 12720.955 1049.32 ;
      RECT 12717.035 1048.035 12717.315 1049.36 ;
      RECT 12713.395 1048.035 12713.675 1049.345 ;
      RECT 12709.755 1048.035 12710.035 1049.255 ;
      RECT 12650.675 1048.035 12650.955 1049.155 ;
      RECT 12646.755 1048.035 12647.035 1049.2 ;
      RECT 12642.835 1048.035 12643.115 1048.93 ;
      RECT 12638.915 1048.035 12639.195 1049.155 ;
      RECT 12634.995 1048.035 12635.275 1064.6 ;
      RECT 12587.955 1048.035 12588.235 1049.3 ;
      RECT 12584.315 1048.035 12584.595 1049.265 ;
      RECT 12580.675 1048.035 12580.955 1049.32 ;
      RECT 12577.035 1048.035 12577.315 1049.36 ;
      RECT 12573.395 1048.035 12573.675 1049.345 ;
      RECT 12569.755 1048.035 12570.035 1049.255 ;
      RECT 12510.675 1048.035 12510.955 1049.155 ;
      RECT 12506.755 1048.035 12507.035 1049.2 ;
      RECT 12502.835 1048.035 12503.115 1048.93 ;
      RECT 12498.915 1048.035 12499.195 1049.155 ;
      RECT 12494.995 1048.035 12495.275 1064.6 ;
      RECT 12447.955 1048.035 12448.235 1049.3 ;
      RECT 12444.315 1048.035 12444.595 1049.265 ;
      RECT 12440.675 1048.035 12440.955 1049.32 ;
      RECT 12437.035 1048.035 12437.315 1049.36 ;
      RECT 12433.395 1048.035 12433.675 1049.345 ;
      RECT 12429.755 1048.035 12430.035 1049.255 ;
      RECT 12370.675 1048.035 12370.955 1049.155 ;
      RECT 12366.755 1048.035 12367.035 1049.2 ;
      RECT 12362.835 1048.035 12363.115 1048.93 ;
      RECT 12358.915 1048.035 12359.195 1049.155 ;
      RECT 12354.995 1048.035 12355.275 1064.6 ;
      RECT 12307.955 1048.035 12308.235 1049.3 ;
      RECT 12304.315 1048.035 12304.595 1049.265 ;
      RECT 12300.675 1048.035 12300.955 1049.32 ;
      RECT 12297.035 1048.035 12297.315 1049.36 ;
      RECT 12293.395 1048.035 12293.675 1049.345 ;
      RECT 12289.755 1048.035 12290.035 1049.255 ;
      RECT 12230.675 1048.035 12230.955 1049.155 ;
      RECT 12226.755 1048.035 12227.035 1049.2 ;
      RECT 12222.835 1048.035 12223.115 1048.93 ;
      RECT 12218.915 1048.035 12219.195 1049.155 ;
      RECT 12214.995 1048.035 12215.275 1064.6 ;
      RECT 12167.955 1048.035 12168.235 1049.3 ;
      RECT 12164.315 1048.035 12164.595 1049.265 ;
      RECT 12160.675 1048.035 12160.955 1049.32 ;
      RECT 12157.035 1048.035 12157.315 1049.36 ;
      RECT 12153.395 1048.035 12153.675 1049.345 ;
      RECT 12149.755 1048.035 12150.035 1049.255 ;
      RECT 12090.675 1048.035 12090.955 1049.155 ;
      RECT 12086.755 1048.035 12087.035 1049.2 ;
      RECT 12082.835 1048.035 12083.115 1048.93 ;
      RECT 12078.915 1048.035 12079.195 1049.155 ;
      RECT 12074.995 1048.035 12075.275 1064.6 ;
      RECT 12027.955 1048.035 12028.235 1049.3 ;
      RECT 12024.315 1048.035 12024.595 1049.265 ;
      RECT 12020.675 1048.035 12020.955 1049.32 ;
      RECT 12017.035 1048.035 12017.315 1049.36 ;
      RECT 12013.395 1048.035 12013.675 1049.345 ;
      RECT 12009.755 1048.035 12010.035 1049.255 ;
      RECT 11950.675 1048.035 11950.955 1049.155 ;
      RECT 11946.755 1048.035 11947.035 1049.2 ;
      RECT 11942.835 1048.035 11943.115 1048.93 ;
      RECT 11938.915 1048.035 11939.195 1049.155 ;
      RECT 11934.995 1048.035 11935.275 1064.6 ;
      RECT 11887.955 1048.035 11888.235 1049.3 ;
      RECT 11884.315 1048.035 11884.595 1049.265 ;
      RECT 11880.675 1048.035 11880.955 1049.32 ;
      RECT 11877.035 1048.035 11877.315 1049.36 ;
      RECT 11873.395 1048.035 11873.675 1049.345 ;
      RECT 11869.755 1048.035 11870.035 1049.255 ;
      RECT 11810.675 1048.035 11810.955 1049.155 ;
      RECT 11806.755 1048.035 11807.035 1049.2 ;
      RECT 11802.835 1048.035 11803.115 1048.93 ;
      RECT 11798.915 1048.035 11799.195 1049.155 ;
      RECT 11794.995 1048.035 11795.275 1064.6 ;
      RECT 11747.955 1048.035 11748.235 1049.3 ;
      RECT 11744.315 1048.035 11744.595 1049.265 ;
      RECT 11740.675 1048.035 11740.955 1049.32 ;
      RECT 11737.035 1048.035 11737.315 1049.36 ;
      RECT 11733.395 1048.035 11733.675 1049.345 ;
      RECT 11729.755 1048.035 11730.035 1049.255 ;
      RECT 11670.675 1048.035 11670.955 1049.155 ;
      RECT 11666.755 1048.035 11667.035 1049.2 ;
      RECT 11662.835 1048.035 11663.115 1048.93 ;
      RECT 11658.915 1048.035 11659.195 1049.155 ;
      RECT 11654.995 1048.035 11655.275 1064.6 ;
      RECT 11607.955 1048.035 11608.235 1049.3 ;
      RECT 11604.315 1048.035 11604.595 1049.265 ;
      RECT 11600.675 1048.035 11600.955 1049.32 ;
      RECT 11597.035 1048.035 11597.315 1049.36 ;
      RECT 11593.395 1048.035 11593.675 1049.345 ;
      RECT 11589.755 1048.035 11590.035 1049.255 ;
      RECT 11530.675 1048.035 11530.955 1049.155 ;
      RECT 11526.755 1048.035 11527.035 1049.2 ;
      RECT 11522.835 1048.035 11523.115 1048.93 ;
      RECT 11518.915 1048.035 11519.195 1049.155 ;
      RECT 11514.995 1048.035 11515.275 1064.6 ;
      RECT 11467.955 1048.035 11468.235 1049.3 ;
      RECT 11464.315 1048.035 11464.595 1049.265 ;
      RECT 11460.675 1048.035 11460.955 1049.32 ;
      RECT 11457.035 1048.035 11457.315 1049.36 ;
      RECT 11453.395 1048.035 11453.675 1049.345 ;
      RECT 11449.755 1048.035 11450.035 1049.255 ;
      RECT 11390.675 1048.035 11390.955 1049.155 ;
      RECT 11386.755 1048.035 11387.035 1049.2 ;
      RECT 11382.835 1048.035 11383.115 1048.93 ;
      RECT 11378.915 1048.035 11379.195 1049.155 ;
      RECT 11374.995 1048.035 11375.275 1064.6 ;
      RECT 11327.955 1048.035 11328.235 1049.3 ;
      RECT 11324.315 1048.035 11324.595 1049.265 ;
      RECT 11320.675 1048.035 11320.955 1049.32 ;
      RECT 11317.035 1048.035 11317.315 1049.36 ;
      RECT 11313.395 1048.035 11313.675 1049.345 ;
      RECT 11309.755 1048.035 11310.035 1049.255 ;
      RECT 11250.675 1048.035 11250.955 1049.155 ;
      RECT 11246.755 1048.035 11247.035 1049.2 ;
      RECT 11242.835 1048.035 11243.115 1048.93 ;
      RECT 11238.915 1048.035 11239.195 1049.155 ;
      RECT 11234.995 1048.035 11235.275 1064.6 ;
      RECT 11187.955 1048.035 11188.235 1049.3 ;
      RECT 11184.315 1048.035 11184.595 1049.265 ;
      RECT 11180.675 1048.035 11180.955 1049.32 ;
      RECT 11177.035 1048.035 11177.315 1049.36 ;
      RECT 11173.395 1048.035 11173.675 1049.345 ;
      RECT 11169.755 1048.035 11170.035 1049.255 ;
      RECT 11110.675 1048.035 11110.955 1049.155 ;
      RECT 11106.755 1048.035 11107.035 1049.2 ;
      RECT 11102.835 1048.035 11103.115 1048.93 ;
      RECT 11098.915 1048.035 11099.195 1049.155 ;
      RECT 11094.995 1048.035 11095.275 1064.6 ;
      RECT 11047.955 1048.035 11048.235 1049.3 ;
      RECT 11044.315 1048.035 11044.595 1049.265 ;
      RECT 11040.675 1048.035 11040.955 1049.32 ;
      RECT 11037.035 1048.035 11037.315 1049.36 ;
      RECT 11033.395 1048.035 11033.675 1049.345 ;
      RECT 11029.755 1048.035 11030.035 1049.255 ;
      RECT 10970.675 1048.035 10970.955 1049.155 ;
      RECT 10966.755 1048.035 10967.035 1049.2 ;
      RECT 10962.835 1048.035 10963.115 1048.93 ;
      RECT 10958.915 1048.035 10959.195 1049.155 ;
      RECT 10954.995 1048.035 10955.275 1064.6 ;
      RECT 10907.955 1048.035 10908.235 1049.3 ;
      RECT 10904.315 1048.035 10904.595 1049.265 ;
      RECT 10900.675 1048.035 10900.955 1049.32 ;
      RECT 10897.035 1048.035 10897.315 1049.36 ;
      RECT 10893.395 1048.035 10893.675 1049.345 ;
      RECT 10889.755 1048.035 10890.035 1049.255 ;
      RECT 10830.675 1048.035 10830.955 1049.155 ;
      RECT 10826.755 1048.035 10827.035 1049.2 ;
      RECT 10822.835 1048.035 10823.115 1048.93 ;
      RECT 10818.915 1048.035 10819.195 1049.155 ;
      RECT 10814.995 1048.035 10815.275 1064.6 ;
      RECT 10767.955 1048.035 10768.235 1049.3 ;
      RECT 10764.315 1048.035 10764.595 1049.265 ;
      RECT 10760.675 1048.035 10760.955 1049.32 ;
      RECT 10757.035 1048.035 10757.315 1049.36 ;
      RECT 10753.395 1048.035 10753.675 1049.345 ;
      RECT 10749.755 1048.035 10750.035 1049.255 ;
      RECT 10690.675 1048.035 10690.955 1049.155 ;
      RECT 10686.755 1048.035 10687.035 1049.2 ;
      RECT 10682.835 1048.035 10683.115 1048.93 ;
      RECT 10678.915 1048.035 10679.195 1049.155 ;
      RECT 10674.995 1048.035 10675.275 1064.6 ;
      RECT 10627.955 1048.035 10628.235 1049.3 ;
      RECT 10624.315 1048.035 10624.595 1049.265 ;
      RECT 10620.675 1048.035 10620.955 1049.32 ;
      RECT 10617.035 1048.035 10617.315 1049.36 ;
      RECT 10613.395 1048.035 10613.675 1049.345 ;
      RECT 10609.755 1048.035 10610.035 1049.255 ;
      RECT 10550.675 1048.035 10550.955 1049.155 ;
      RECT 10546.755 1048.035 10547.035 1049.2 ;
      RECT 10542.835 1048.035 10543.115 1048.93 ;
      RECT 10538.915 1048.035 10539.195 1049.155 ;
      RECT 10534.995 1048.035 10535.275 1064.6 ;
      RECT 10487.955 1048.035 10488.235 1049.3 ;
      RECT 10484.315 1048.035 10484.595 1049.265 ;
      RECT 10480.675 1048.035 10480.955 1049.32 ;
      RECT 10477.035 1048.035 10477.315 1049.36 ;
      RECT 10473.395 1048.035 10473.675 1049.345 ;
      RECT 10469.755 1048.035 10470.035 1049.255 ;
      RECT 10410.675 1048.035 10410.955 1049.155 ;
      RECT 10406.755 1048.035 10407.035 1049.2 ;
      RECT 10402.835 1048.035 10403.115 1048.93 ;
      RECT 10398.915 1048.035 10399.195 1049.155 ;
      RECT 10394.995 1048.035 10395.275 1064.6 ;
      RECT 10347.955 1048.035 10348.235 1049.3 ;
      RECT 10344.315 1048.035 10344.595 1049.265 ;
      RECT 10340.675 1048.035 10340.955 1049.32 ;
      RECT 10337.035 1048.035 10337.315 1049.36 ;
      RECT 10333.395 1048.035 10333.675 1049.345 ;
      RECT 10329.755 1048.035 10330.035 1049.255 ;
      RECT 10270.675 1048.035 10270.955 1049.155 ;
      RECT 10266.755 1048.035 10267.035 1049.2 ;
      RECT 10262.835 1048.035 10263.115 1048.93 ;
      RECT 10258.915 1048.035 10259.195 1049.155 ;
      RECT 10254.995 1048.035 10255.275 1064.6 ;
      RECT 10207.955 1048.035 10208.235 1049.3 ;
      RECT 10204.315 1048.035 10204.595 1049.265 ;
      RECT 10200.675 1048.035 10200.955 1049.32 ;
      RECT 10197.035 1048.035 10197.315 1049.36 ;
      RECT 10193.395 1048.035 10193.675 1049.345 ;
      RECT 10189.755 1048.035 10190.035 1049.255 ;
      RECT 10130.675 1048.035 10130.955 1049.155 ;
      RECT 10126.755 1048.035 10127.035 1049.2 ;
      RECT 10122.835 1048.035 10123.115 1048.93 ;
      RECT 10118.915 1048.035 10119.195 1049.155 ;
      RECT 10114.995 1048.035 10115.275 1064.6 ;
      RECT 10104.235 1047.01 10104.325 1047.29 ;
      RECT 10102.385 1047.01 10102.475 1047.29 ;
      RECT 10099.715 1048.035 10100.275 1049.01 ;
      RECT 10098.035 1048.035 10098.595 1049.94 ;
      RECT 10096.355 1048.035 10096.915 1050.87 ;
      RECT 10094.675 1048.035 10095.235 1051.8 ;
      RECT 10092.995 1048.035 10093.555 1052.73 ;
      RECT 10091.315 1048.035 10091.875 1053.66 ;
      RECT 10089.635 1048.035 10090.195 1054.59 ;
      RECT 10087.955 1048.035 10088.515 1055.51 ;
      RECT 10086.275 1048.035 10086.835 1056.44 ;
      RECT 10084.595 1048.035 10085.155 1057.37 ;
      RECT 10082.915 1048.035 10083.475 1058.3 ;
      RECT 10081.235 1048.035 10081.795 1059.23 ;
      RECT 10079.555 1048.035 10080.115 1060.16 ;
      RECT 10067.955 1048.035 10068.235 1049.3 ;
      RECT 10064.315 1048.035 10064.595 1049.265 ;
      RECT 10060.675 1048.035 10060.955 1049.32 ;
      RECT 10057.035 1048.035 10057.315 1049.36 ;
      RECT 10053.395 1048.035 10053.675 1049.345 ;
      RECT 10049.755 1048.035 10050.035 1049.255 ;
      RECT 9990.675 1048.035 9990.955 1049.155 ;
      RECT 9986.755 1048.035 9987.035 1049.2 ;
      RECT 9982.835 1048.035 9983.115 1048.93 ;
      RECT 9978.915 1048.035 9979.195 1049.155 ;
      RECT 9974.995 1048.035 9975.275 1064.6 ;
      RECT 9927.955 1048.035 9928.235 1049.3 ;
      RECT 9924.315 1048.035 9924.595 1049.265 ;
      RECT 9920.675 1048.035 9920.955 1049.32 ;
      RECT 9917.035 1048.035 9917.315 1049.36 ;
      RECT 9913.395 1048.035 9913.675 1049.345 ;
      RECT 9909.755 1048.035 9910.035 1049.255 ;
      RECT 9850.675 1048.035 9850.955 1049.155 ;
      RECT 9846.755 1048.035 9847.035 1049.2 ;
      RECT 9842.835 1048.035 9843.115 1048.93 ;
      RECT 9838.915 1048.035 9839.195 1049.155 ;
      RECT 9834.995 1048.035 9835.275 1064.6 ;
      RECT 9787.955 1048.035 9788.235 1049.3 ;
      RECT 9784.315 1048.035 9784.595 1049.265 ;
      RECT 9780.675 1048.035 9780.955 1049.32 ;
      RECT 9777.035 1048.035 9777.315 1049.36 ;
      RECT 9773.395 1048.035 9773.675 1049.345 ;
      RECT 9769.755 1048.035 9770.035 1049.255 ;
      RECT 9710.675 1048.035 9710.955 1049.155 ;
      RECT 9706.755 1048.035 9707.035 1049.2 ;
      RECT 9702.835 1048.035 9703.115 1048.93 ;
      RECT 9698.915 1048.035 9699.195 1049.155 ;
      RECT 9694.995 1048.035 9695.275 1064.6 ;
      RECT 9647.955 1048.035 9648.235 1049.3 ;
      RECT 9644.315 1048.035 9644.595 1049.265 ;
      RECT 9640.675 1048.035 9640.955 1049.32 ;
      RECT 9637.035 1048.035 9637.315 1049.36 ;
      RECT 9633.395 1048.035 9633.675 1049.345 ;
      RECT 9629.755 1048.035 9630.035 1049.255 ;
      RECT 9570.675 1048.035 9570.955 1049.155 ;
      RECT 9566.755 1048.035 9567.035 1049.2 ;
      RECT 9562.835 1048.035 9563.115 1048.93 ;
      RECT 9558.915 1048.035 9559.195 1049.155 ;
      RECT 9554.995 1048.035 9555.275 1064.6 ;
      RECT 9507.955 1048.035 9508.235 1049.3 ;
      RECT 9504.315 1048.035 9504.595 1049.265 ;
      RECT 9500.675 1048.035 9500.955 1049.32 ;
      RECT 9497.035 1048.035 9497.315 1049.36 ;
      RECT 9493.395 1048.035 9493.675 1049.345 ;
      RECT 9489.755 1048.035 9490.035 1049.255 ;
      RECT 9430.675 1048.035 9430.955 1049.155 ;
      RECT 9426.755 1048.035 9427.035 1049.2 ;
      RECT 9422.835 1048.035 9423.115 1048.93 ;
      RECT 9418.915 1048.035 9419.195 1049.155 ;
      RECT 9414.995 1048.035 9415.275 1064.6 ;
      RECT 9367.955 1048.035 9368.235 1049.3 ;
      RECT 9364.315 1048.035 9364.595 1049.265 ;
      RECT 9360.675 1048.035 9360.955 1049.32 ;
      RECT 9357.035 1048.035 9357.315 1049.36 ;
      RECT 9353.395 1048.035 9353.675 1049.345 ;
      RECT 9349.755 1048.035 9350.035 1049.255 ;
      RECT 9290.675 1048.035 9290.955 1049.155 ;
      RECT 9286.755 1048.035 9287.035 1049.2 ;
      RECT 9282.835 1048.035 9283.115 1048.93 ;
      RECT 9278.915 1048.035 9279.195 1049.155 ;
      RECT 9274.995 1048.035 9275.275 1064.6 ;
      RECT 9227.955 1048.035 9228.235 1049.3 ;
      RECT 9224.315 1048.035 9224.595 1049.265 ;
      RECT 9220.675 1048.035 9220.955 1049.32 ;
      RECT 9217.035 1048.035 9217.315 1049.36 ;
      RECT 9213.395 1048.035 9213.675 1049.345 ;
      RECT 9209.755 1048.035 9210.035 1049.255 ;
      RECT 9150.675 1048.035 9150.955 1049.155 ;
      RECT 9146.755 1048.035 9147.035 1049.2 ;
      RECT 9142.835 1048.035 9143.115 1048.93 ;
      RECT 9138.915 1048.035 9139.195 1049.155 ;
      RECT 9134.995 1048.035 9135.275 1064.6 ;
      RECT 9087.955 1048.035 9088.235 1049.3 ;
      RECT 9084.315 1048.035 9084.595 1049.265 ;
      RECT 9080.675 1048.035 9080.955 1049.32 ;
      RECT 9077.035 1048.035 9077.315 1049.36 ;
      RECT 9073.395 1048.035 9073.675 1049.345 ;
      RECT 9069.755 1048.035 9070.035 1049.255 ;
      RECT 9010.675 1048.035 9010.955 1049.155 ;
      RECT 9006.755 1048.035 9007.035 1049.2 ;
      RECT 9002.835 1048.035 9003.115 1048.93 ;
      RECT 8998.915 1048.035 8999.195 1049.155 ;
      RECT 8994.995 1048.035 8995.275 1064.6 ;
      RECT 8947.955 1048.035 8948.235 1049.3 ;
      RECT 8944.315 1048.035 8944.595 1049.265 ;
      RECT 8940.675 1048.035 8940.955 1049.32 ;
      RECT 8937.035 1048.035 8937.315 1049.36 ;
      RECT 8933.395 1048.035 8933.675 1049.345 ;
      RECT 8929.755 1048.035 8930.035 1049.255 ;
      RECT 8870.675 1048.035 8870.955 1049.155 ;
      RECT 8866.755 1048.035 8867.035 1049.2 ;
      RECT 8862.835 1048.035 8863.115 1048.93 ;
      RECT 8858.915 1048.035 8859.195 1049.155 ;
      RECT 8854.995 1048.035 8855.275 1064.6 ;
      RECT 8807.955 1048.035 8808.235 1049.3 ;
      RECT 8804.315 1048.035 8804.595 1049.265 ;
      RECT 8800.675 1048.035 8800.955 1049.32 ;
      RECT 8797.035 1048.035 8797.315 1049.36 ;
      RECT 8793.395 1048.035 8793.675 1049.345 ;
      RECT 8789.755 1048.035 8790.035 1049.255 ;
      RECT 8730.675 1048.035 8730.955 1049.155 ;
      RECT 8726.755 1048.035 8727.035 1049.2 ;
      RECT 8722.835 1048.035 8723.115 1048.93 ;
      RECT 8718.915 1048.035 8719.195 1049.155 ;
      RECT 8714.995 1048.035 8715.275 1064.6 ;
      RECT 8667.955 1048.035 8668.235 1049.3 ;
      RECT 8664.315 1048.035 8664.595 1049.265 ;
      RECT 8660.675 1048.035 8660.955 1049.32 ;
      RECT 8657.035 1048.035 8657.315 1049.36 ;
      RECT 8653.395 1048.035 8653.675 1049.345 ;
      RECT 8649.755 1048.035 8650.035 1049.255 ;
      RECT 8590.675 1048.035 8590.955 1049.155 ;
      RECT 8586.755 1048.035 8587.035 1049.2 ;
      RECT 8582.835 1048.035 8583.115 1048.93 ;
      RECT 8578.915 1048.035 8579.195 1049.155 ;
      RECT 8574.995 1048.035 8575.275 1064.6 ;
      RECT 8527.955 1048.035 8528.235 1049.3 ;
      RECT 8524.315 1048.035 8524.595 1049.265 ;
      RECT 8520.675 1048.035 8520.955 1049.32 ;
      RECT 8517.035 1048.035 8517.315 1049.36 ;
      RECT 8513.395 1048.035 8513.675 1049.345 ;
      RECT 8509.755 1048.035 8510.035 1049.255 ;
      RECT 8450.675 1048.035 8450.955 1049.155 ;
      RECT 8446.755 1048.035 8447.035 1049.2 ;
      RECT 8442.835 1048.035 8443.115 1048.93 ;
      RECT 8438.915 1048.035 8439.195 1049.155 ;
      RECT 8434.995 1048.035 8435.275 1064.6 ;
      RECT 8387.955 1048.035 8388.235 1049.3 ;
      RECT 8384.315 1048.035 8384.595 1049.265 ;
      RECT 8380.675 1048.035 8380.955 1049.32 ;
      RECT 8377.035 1048.035 8377.315 1049.36 ;
      RECT 8373.395 1048.035 8373.675 1049.345 ;
      RECT 8369.755 1048.035 8370.035 1049.255 ;
      RECT 8310.675 1048.035 8310.955 1049.155 ;
      RECT 8306.755 1048.035 8307.035 1049.2 ;
      RECT 8302.835 1048.035 8303.115 1048.93 ;
      RECT 8298.915 1048.035 8299.195 1049.155 ;
      RECT 8294.995 1048.035 8295.275 1064.6 ;
      RECT 8247.955 1048.035 8248.235 1049.3 ;
      RECT 8244.315 1048.035 8244.595 1049.265 ;
      RECT 8240.675 1048.035 8240.955 1049.32 ;
      RECT 8237.035 1048.035 8237.315 1049.36 ;
      RECT 8233.395 1048.035 8233.675 1049.345 ;
      RECT 8229.755 1048.035 8230.035 1049.255 ;
      RECT 8170.675 1048.035 8170.955 1049.155 ;
      RECT 8166.755 1048.035 8167.035 1049.2 ;
      RECT 8162.835 1048.035 8163.115 1048.93 ;
      RECT 8158.915 1048.035 8159.195 1049.155 ;
      RECT 8154.995 1048.035 8155.275 1064.6 ;
      RECT 8107.955 1048.035 8108.235 1049.3 ;
      RECT 8104.315 1048.035 8104.595 1049.265 ;
      RECT 8100.675 1048.035 8100.955 1049.32 ;
      RECT 8097.035 1048.035 8097.315 1049.36 ;
      RECT 8093.395 1048.035 8093.675 1049.345 ;
      RECT 8089.755 1048.035 8090.035 1049.255 ;
      RECT 8030.675 1048.035 8030.955 1049.155 ;
      RECT 8026.755 1048.035 8027.035 1049.2 ;
      RECT 8022.835 1048.035 8023.115 1048.93 ;
      RECT 8018.915 1048.035 8019.195 1049.155 ;
      RECT 8014.995 1048.035 8015.275 1064.6 ;
      RECT 7967.955 1048.035 7968.235 1049.3 ;
      RECT 7964.315 1048.035 7964.595 1049.265 ;
      RECT 7960.675 1048.035 7960.955 1049.32 ;
      RECT 7957.035 1048.035 7957.315 1049.36 ;
      RECT 7953.395 1048.035 7953.675 1049.345 ;
      RECT 7949.755 1048.035 7950.035 1049.255 ;
      RECT 7890.675 1048.035 7890.955 1049.155 ;
      RECT 7886.755 1048.035 7887.035 1049.2 ;
      RECT 7882.835 1048.035 7883.115 1048.93 ;
      RECT 7878.915 1048.035 7879.195 1049.155 ;
      RECT 7874.995 1048.035 7875.275 1064.6 ;
      RECT 7827.955 1048.035 7828.235 1049.3 ;
      RECT 7824.315 1048.035 7824.595 1049.265 ;
      RECT 7820.675 1048.035 7820.955 1049.32 ;
      RECT 7817.035 1048.035 7817.315 1049.36 ;
      RECT 7813.395 1048.035 7813.675 1049.345 ;
      RECT 7809.755 1048.035 7810.035 1049.255 ;
      RECT 7750.675 1048.035 7750.955 1049.155 ;
      RECT 7746.755 1048.035 7747.035 1049.2 ;
      RECT 7742.835 1048.035 7743.115 1048.93 ;
      RECT 7738.915 1048.035 7739.195 1049.155 ;
      RECT 7734.995 1048.035 7735.275 1064.6 ;
      RECT 7687.955 1048.035 7688.235 1049.3 ;
      RECT 7684.315 1048.035 7684.595 1049.265 ;
      RECT 7680.675 1048.035 7680.955 1049.32 ;
      RECT 7677.035 1048.035 7677.315 1049.36 ;
      RECT 7673.395 1048.035 7673.675 1049.345 ;
      RECT 7669.755 1048.035 7670.035 1049.255 ;
      RECT 7610.675 1048.035 7610.955 1049.155 ;
      RECT 7606.755 1048.035 7607.035 1049.2 ;
      RECT 7602.835 1048.035 7603.115 1048.93 ;
      RECT 7598.915 1048.035 7599.195 1049.155 ;
      RECT 7594.995 1048.035 7595.275 1064.6 ;
      RECT 7547.955 1048.035 7548.235 1049.3 ;
      RECT 7544.315 1048.035 7544.595 1049.265 ;
      RECT 7540.675 1048.035 7540.955 1049.32 ;
      RECT 7537.035 1048.035 7537.315 1049.36 ;
      RECT 7533.395 1048.035 7533.675 1049.345 ;
      RECT 7529.755 1048.035 7530.035 1049.255 ;
      RECT 7470.675 1048.035 7470.955 1049.155 ;
      RECT 7466.755 1048.035 7467.035 1049.2 ;
      RECT 7462.835 1048.035 7463.115 1048.93 ;
      RECT 7458.915 1048.035 7459.195 1049.155 ;
      RECT 7454.995 1048.035 7455.275 1064.6 ;
      RECT 7407.955 1048.035 7408.235 1049.3 ;
      RECT 7404.315 1048.035 7404.595 1049.265 ;
      RECT 7400.675 1048.035 7400.955 1049.32 ;
      RECT 7397.035 1048.035 7397.315 1049.36 ;
      RECT 7393.395 1048.035 7393.675 1049.345 ;
      RECT 7389.755 1048.035 7390.035 1049.255 ;
      RECT 7330.675 1048.035 7330.955 1049.155 ;
      RECT 7326.755 1048.035 7327.035 1049.2 ;
      RECT 7322.835 1048.035 7323.115 1048.93 ;
      RECT 7318.915 1048.035 7319.195 1049.155 ;
      RECT 7314.995 1048.035 7315.275 1064.6 ;
      RECT 7267.955 1048.035 7268.235 1049.3 ;
      RECT 7264.315 1048.035 7264.595 1049.265 ;
      RECT 7260.675 1048.035 7260.955 1049.32 ;
      RECT 7257.035 1048.035 7257.315 1049.36 ;
      RECT 7253.395 1048.035 7253.675 1049.345 ;
      RECT 7249.755 1048.035 7250.035 1049.255 ;
      RECT 7190.675 1048.035 7190.955 1049.155 ;
      RECT 7186.755 1048.035 7187.035 1049.2 ;
      RECT 7182.835 1048.035 7183.115 1048.93 ;
      RECT 7178.915 1048.035 7179.195 1049.155 ;
      RECT 7174.995 1048.035 7175.275 1064.6 ;
      RECT 7127.955 1048.035 7128.235 1049.3 ;
      RECT 7124.315 1048.035 7124.595 1049.265 ;
      RECT 7120.675 1048.035 7120.955 1049.32 ;
      RECT 7117.035 1048.035 7117.315 1049.36 ;
      RECT 7113.395 1048.035 7113.675 1049.345 ;
      RECT 7109.755 1048.035 7110.035 1049.255 ;
      RECT 7050.675 1048.035 7050.955 1049.155 ;
      RECT 7046.755 1048.035 7047.035 1049.2 ;
      RECT 7042.835 1048.035 7043.115 1048.93 ;
      RECT 7038.915 1048.035 7039.195 1049.155 ;
      RECT 7034.995 1048.035 7035.275 1064.6 ;
      RECT 6987.955 1048.035 6988.235 1049.3 ;
      RECT 6984.315 1048.035 6984.595 1049.265 ;
      RECT 6980.675 1048.035 6980.955 1049.32 ;
      RECT 6977.035 1048.035 6977.315 1049.36 ;
      RECT 6973.395 1048.035 6973.675 1049.345 ;
      RECT 6969.755 1048.035 6970.035 1049.255 ;
      RECT 6910.675 1048.035 6910.955 1049.155 ;
      RECT 6906.755 1048.035 6907.035 1049.2 ;
      RECT 6902.835 1048.035 6903.115 1048.93 ;
      RECT 6898.915 1048.035 6899.195 1049.155 ;
      RECT 6894.995 1048.035 6895.275 1064.6 ;
      RECT 6847.955 1048.035 6848.235 1049.3 ;
      RECT 6844.315 1048.035 6844.595 1049.265 ;
      RECT 6840.675 1048.035 6840.955 1049.32 ;
      RECT 6837.035 1048.035 6837.315 1049.36 ;
      RECT 6833.395 1048.035 6833.675 1049.345 ;
      RECT 6829.755 1048.035 6830.035 1049.255 ;
      RECT 6770.675 1048.035 6770.955 1049.155 ;
      RECT 6766.755 1048.035 6767.035 1049.2 ;
      RECT 6762.835 1048.035 6763.115 1048.93 ;
      RECT 6758.915 1048.035 6759.195 1049.155 ;
      RECT 6754.995 1048.035 6755.275 1064.6 ;
      RECT 6707.955 1048.035 6708.235 1049.3 ;
      RECT 6704.315 1048.035 6704.595 1049.265 ;
      RECT 6700.675 1048.035 6700.955 1049.32 ;
      RECT 6697.035 1048.035 6697.315 1049.36 ;
      RECT 6693.395 1048.035 6693.675 1049.345 ;
      RECT 6689.755 1048.035 6690.035 1049.255 ;
      RECT 6630.675 1048.035 6630.955 1049.155 ;
      RECT 6626.755 1048.035 6627.035 1049.2 ;
      RECT 6622.835 1048.035 6623.115 1048.93 ;
      RECT 6618.915 1048.035 6619.195 1049.155 ;
      RECT 6614.995 1048.035 6615.275 1064.6 ;
      RECT 6567.955 1048.035 6568.235 1049.3 ;
      RECT 6564.315 1048.035 6564.595 1049.265 ;
      RECT 6560.675 1048.035 6560.955 1049.32 ;
      RECT 6557.035 1048.035 6557.315 1049.36 ;
      RECT 6553.395 1048.035 6553.675 1049.345 ;
      RECT 6549.755 1048.035 6550.035 1049.255 ;
      RECT 6490.675 1048.035 6490.955 1049.155 ;
      RECT 6486.755 1048.035 6487.035 1049.2 ;
      RECT 6482.835 1048.035 6483.115 1048.93 ;
      RECT 6478.915 1048.035 6479.195 1049.155 ;
      RECT 6474.995 1048.035 6475.275 1064.6 ;
      RECT 6427.955 1048.035 6428.235 1049.3 ;
      RECT 6424.315 1048.035 6424.595 1049.265 ;
      RECT 6420.675 1048.035 6420.955 1049.32 ;
      RECT 6417.035 1048.035 6417.315 1049.36 ;
      RECT 6413.395 1048.035 6413.675 1049.345 ;
      RECT 6409.755 1048.035 6410.035 1049.255 ;
      RECT 6350.675 1048.035 6350.955 1049.155 ;
      RECT 6346.755 1048.035 6347.035 1049.2 ;
      RECT 6342.835 1048.035 6343.115 1048.93 ;
      RECT 6338.915 1048.035 6339.195 1049.155 ;
      RECT 6334.995 1048.035 6335.275 1064.6 ;
      RECT 6287.955 1048.035 6288.235 1049.3 ;
      RECT 6284.315 1048.035 6284.595 1049.265 ;
      RECT 6280.675 1048.035 6280.955 1049.32 ;
      RECT 6277.035 1048.035 6277.315 1049.36 ;
      RECT 6273.395 1048.035 6273.675 1049.345 ;
      RECT 6269.755 1048.035 6270.035 1049.255 ;
      RECT 6210.675 1048.035 6210.955 1049.155 ;
      RECT 6206.755 1048.035 6207.035 1049.2 ;
      RECT 6202.835 1048.035 6203.115 1048.93 ;
      RECT 6198.915 1048.035 6199.195 1049.155 ;
      RECT 6194.995 1048.035 6195.275 1064.6 ;
      RECT 6147.955 1048.035 6148.235 1049.3 ;
      RECT 6144.315 1048.035 6144.595 1049.265 ;
      RECT 6140.675 1048.035 6140.955 1049.32 ;
      RECT 6137.035 1048.035 6137.315 1049.36 ;
      RECT 6133.395 1048.035 6133.675 1049.345 ;
      RECT 6129.755 1048.035 6130.035 1049.255 ;
      RECT 6070.675 1048.035 6070.955 1049.155 ;
      RECT 6066.755 1048.035 6067.035 1049.2 ;
      RECT 6062.835 1048.035 6063.115 1048.93 ;
      RECT 6058.915 1048.035 6059.195 1049.155 ;
      RECT 6054.995 1048.035 6055.275 1064.6 ;
      RECT 6007.955 1048.035 6008.235 1049.3 ;
      RECT 6004.315 1048.035 6004.595 1049.265 ;
      RECT 6000.675 1048.035 6000.955 1049.32 ;
      RECT 5997.035 1048.035 5997.315 1049.36 ;
      RECT 5993.395 1048.035 5993.675 1049.345 ;
      RECT 5989.755 1048.035 5990.035 1049.255 ;
      RECT 5930.675 1048.035 5930.955 1049.155 ;
      RECT 5926.755 1048.035 5927.035 1049.2 ;
      RECT 5922.835 1048.035 5923.115 1048.93 ;
      RECT 5918.915 1048.035 5919.195 1049.155 ;
      RECT 5914.995 1048.035 5915.275 1064.6 ;
      RECT 5867.955 1048.035 5868.235 1049.3 ;
      RECT 5864.315 1048.035 5864.595 1049.265 ;
      RECT 5860.675 1048.035 5860.955 1049.32 ;
      RECT 5857.035 1048.035 5857.315 1049.36 ;
      RECT 5853.395 1048.035 5853.675 1049.345 ;
      RECT 5849.755 1048.035 5850.035 1049.255 ;
      RECT 5790.675 1048.035 5790.955 1049.155 ;
      RECT 5786.755 1048.035 5787.035 1049.2 ;
      RECT 5782.835 1048.035 5783.115 1048.93 ;
      RECT 5778.915 1048.035 5779.195 1049.155 ;
      RECT 5774.995 1048.035 5775.275 1064.6 ;
      RECT 5727.955 1048.035 5728.235 1049.3 ;
      RECT 5724.315 1048.035 5724.595 1049.265 ;
      RECT 5720.675 1048.035 5720.955 1049.32 ;
      RECT 5717.035 1048.035 5717.315 1049.36 ;
      RECT 5713.395 1048.035 5713.675 1049.345 ;
      RECT 5709.755 1048.035 5710.035 1049.255 ;
      RECT 5650.675 1048.035 5650.955 1049.155 ;
      RECT 5646.755 1048.035 5647.035 1049.2 ;
      RECT 5642.835 1048.035 5643.115 1048.93 ;
      RECT 5638.915 1048.035 5639.195 1049.155 ;
      RECT 5634.995 1048.035 5635.275 1064.6 ;
      RECT 5587.955 1048.035 5588.235 1049.3 ;
      RECT 5584.315 1048.035 5584.595 1049.265 ;
      RECT 5580.675 1048.035 5580.955 1049.32 ;
      RECT 5577.035 1048.035 5577.315 1049.36 ;
      RECT 5573.395 1048.035 5573.675 1049.345 ;
      RECT 5569.755 1048.035 5570.035 1049.255 ;
      RECT 5510.675 1048.035 5510.955 1049.155 ;
      RECT 5506.755 1048.035 5507.035 1049.2 ;
      RECT 5502.835 1048.035 5503.115 1048.93 ;
      RECT 5498.915 1048.035 5499.195 1049.155 ;
      RECT 5494.995 1048.035 5495.275 1064.6 ;
      RECT 5447.955 1048.035 5448.235 1049.3 ;
      RECT 5444.315 1048.035 5444.595 1049.265 ;
      RECT 5440.675 1048.035 5440.955 1049.32 ;
      RECT 5437.035 1048.035 5437.315 1049.36 ;
      RECT 5433.395 1048.035 5433.675 1049.345 ;
      RECT 5429.755 1048.035 5430.035 1049.255 ;
      RECT 5370.675 1048.035 5370.955 1049.155 ;
      RECT 5366.755 1048.035 5367.035 1049.2 ;
      RECT 5362.835 1048.035 5363.115 1048.93 ;
      RECT 5358.915 1048.035 5359.195 1049.155 ;
      RECT 5354.995 1048.035 5355.275 1064.6 ;
      RECT 5307.955 1048.035 5308.235 1049.3 ;
      RECT 5304.315 1048.035 5304.595 1049.265 ;
      RECT 5300.675 1048.035 5300.955 1049.32 ;
      RECT 5297.035 1048.035 5297.315 1049.36 ;
      RECT 5293.395 1048.035 5293.675 1049.345 ;
      RECT 5289.755 1048.035 5290.035 1049.255 ;
      RECT 5230.675 1048.035 5230.955 1049.155 ;
      RECT 5226.755 1048.035 5227.035 1049.2 ;
      RECT 5222.835 1048.035 5223.115 1048.93 ;
      RECT 5218.915 1048.035 5219.195 1049.155 ;
      RECT 5214.995 1048.035 5215.275 1064.6 ;
      RECT 5167.955 1048.035 5168.235 1049.3 ;
      RECT 5164.315 1048.035 5164.595 1049.265 ;
      RECT 5160.675 1048.035 5160.955 1049.32 ;
      RECT 5157.035 1048.035 5157.315 1049.36 ;
      RECT 5153.395 1048.035 5153.675 1049.345 ;
      RECT 5149.755 1048.035 5150.035 1049.255 ;
      RECT 5090.675 1048.035 5090.955 1049.155 ;
      RECT 5086.755 1048.035 5087.035 1049.2 ;
      RECT 5082.835 1048.035 5083.115 1048.93 ;
      RECT 5078.915 1048.035 5079.195 1049.155 ;
      RECT 5074.995 1048.035 5075.275 1064.6 ;
      RECT 5027.955 1048.035 5028.235 1049.3 ;
      RECT 5024.315 1048.035 5024.595 1049.265 ;
      RECT 5020.675 1048.035 5020.955 1049.32 ;
      RECT 5017.035 1048.035 5017.315 1049.36 ;
      RECT 5013.395 1048.035 5013.675 1049.345 ;
      RECT 5009.755 1048.035 5010.035 1049.255 ;
      RECT 4950.675 1048.035 4950.955 1049.155 ;
      RECT 4946.755 1048.035 4947.035 1049.2 ;
      RECT 4942.835 1048.035 4943.115 1048.93 ;
      RECT 4938.915 1048.035 4939.195 1049.155 ;
      RECT 4934.995 1048.035 4935.275 1064.6 ;
      RECT 4887.955 1048.035 4888.235 1049.3 ;
      RECT 4884.315 1048.035 4884.595 1049.265 ;
      RECT 4880.675 1048.035 4880.955 1049.32 ;
      RECT 4877.035 1048.035 4877.315 1049.36 ;
      RECT 4873.395 1048.035 4873.675 1049.345 ;
      RECT 4869.755 1048.035 4870.035 1049.255 ;
      RECT 4810.675 1048.035 4810.955 1049.155 ;
      RECT 4806.755 1048.035 4807.035 1049.2 ;
      RECT 4802.835 1048.035 4803.115 1048.93 ;
      RECT 4798.915 1048.035 4799.195 1049.155 ;
      RECT 4794.995 1048.035 4795.275 1064.6 ;
      RECT 4747.955 1048.035 4748.235 1049.3 ;
      RECT 4744.315 1048.035 4744.595 1049.265 ;
      RECT 4740.675 1048.035 4740.955 1049.32 ;
      RECT 4737.035 1048.035 4737.315 1049.36 ;
      RECT 4733.395 1048.035 4733.675 1049.345 ;
      RECT 4729.755 1048.035 4730.035 1049.255 ;
      RECT 4670.675 1048.035 4670.955 1049.155 ;
      RECT 4666.755 1048.035 4667.035 1049.2 ;
      RECT 4662.835 1048.035 4663.115 1048.93 ;
      RECT 4658.915 1048.035 4659.195 1049.155 ;
      RECT 4654.995 1048.035 4655.275 1064.6 ;
      RECT 4607.955 1048.035 4608.235 1049.3 ;
      RECT 4604.315 1048.035 4604.595 1049.265 ;
      RECT 4600.675 1048.035 4600.955 1049.32 ;
      RECT 4597.035 1048.035 4597.315 1049.36 ;
      RECT 4593.395 1048.035 4593.675 1049.345 ;
      RECT 4589.755 1048.035 4590.035 1049.255 ;
      RECT 4530.675 1048.035 4530.955 1049.155 ;
      RECT 4526.755 1048.035 4527.035 1049.2 ;
      RECT 4522.835 1048.035 4523.115 1048.93 ;
      RECT 4518.915 1048.035 4519.195 1049.155 ;
      RECT 4514.995 1048.035 4515.275 1064.6 ;
      RECT 4467.955 1048.035 4468.235 1049.3 ;
      RECT 4464.315 1048.035 4464.595 1049.265 ;
      RECT 4460.675 1048.035 4460.955 1049.32 ;
      RECT 4457.035 1048.035 4457.315 1049.36 ;
      RECT 4453.395 1048.035 4453.675 1049.345 ;
      RECT 4449.755 1048.035 4450.035 1049.255 ;
      RECT 4390.675 1048.035 4390.955 1049.155 ;
      RECT 4386.755 1048.035 4387.035 1049.2 ;
      RECT 4382.835 1048.035 4383.115 1048.93 ;
      RECT 4378.915 1048.035 4379.195 1049.155 ;
      RECT 4374.995 1048.035 4375.275 1064.6 ;
      RECT 4327.955 1048.035 4328.235 1049.3 ;
      RECT 4324.315 1048.035 4324.595 1049.265 ;
      RECT 4320.675 1048.035 4320.955 1049.32 ;
      RECT 4317.035 1048.035 4317.315 1049.36 ;
      RECT 4313.395 1048.035 4313.675 1049.345 ;
      RECT 4309.755 1048.035 4310.035 1049.255 ;
      RECT 4250.675 1048.035 4250.955 1049.155 ;
      RECT 4246.755 1048.035 4247.035 1049.2 ;
      RECT 4242.835 1048.035 4243.115 1048.93 ;
      RECT 4238.915 1048.035 4239.195 1049.155 ;
      RECT 4234.995 1048.035 4235.275 1064.6 ;
      RECT 4187.955 1048.035 4188.235 1049.3 ;
      RECT 4184.315 1048.035 4184.595 1049.265 ;
      RECT 4180.675 1048.035 4180.955 1049.32 ;
      RECT 4177.035 1048.035 4177.315 1049.36 ;
      RECT 4173.395 1048.035 4173.675 1049.345 ;
      RECT 4169.755 1048.035 4170.035 1049.255 ;
      RECT 4110.675 1048.035 4110.955 1049.155 ;
      RECT 4106.755 1048.035 4107.035 1049.2 ;
      RECT 4102.835 1048.035 4103.115 1048.93 ;
      RECT 4098.915 1048.035 4099.195 1049.155 ;
      RECT 4094.995 1048.035 4095.275 1064.6 ;
      RECT 4047.955 1048.035 4048.235 1049.3 ;
      RECT 4044.315 1048.035 4044.595 1049.265 ;
      RECT 4040.675 1048.035 4040.955 1049.32 ;
      RECT 4037.035 1048.035 4037.315 1049.36 ;
      RECT 4033.395 1048.035 4033.675 1049.345 ;
      RECT 4029.755 1048.035 4030.035 1049.255 ;
      RECT 3970.675 1048.035 3970.955 1049.155 ;
      RECT 3966.755 1048.035 3967.035 1049.2 ;
      RECT 3962.835 1048.035 3963.115 1048.93 ;
      RECT 3958.915 1048.035 3959.195 1049.155 ;
      RECT 3954.995 1048.035 3955.275 1064.6 ;
      RECT 3907.955 1048.035 3908.235 1049.3 ;
      RECT 3904.315 1048.035 3904.595 1049.265 ;
      RECT 3900.675 1048.035 3900.955 1049.32 ;
      RECT 3897.035 1048.035 3897.315 1049.36 ;
      RECT 3893.395 1048.035 3893.675 1049.345 ;
      RECT 3889.755 1048.035 3890.035 1049.255 ;
      RECT 3830.675 1048.035 3830.955 1049.155 ;
      RECT 3826.755 1048.035 3827.035 1049.2 ;
      RECT 3822.835 1048.035 3823.115 1048.93 ;
      RECT 3818.915 1048.035 3819.195 1049.155 ;
      RECT 3814.995 1048.035 3815.275 1064.6 ;
      RECT 3767.955 1048.035 3768.235 1049.3 ;
      RECT 3764.315 1048.035 3764.595 1049.265 ;
      RECT 3760.675 1048.035 3760.955 1049.32 ;
      RECT 3757.035 1048.035 3757.315 1049.36 ;
      RECT 3753.395 1048.035 3753.675 1049.345 ;
      RECT 3749.755 1048.035 3750.035 1049.255 ;
      RECT 3690.675 1048.035 3690.955 1049.155 ;
      RECT 3686.755 1048.035 3687.035 1049.2 ;
      RECT 3682.835 1048.035 3683.115 1048.93 ;
      RECT 3678.915 1048.035 3679.195 1049.155 ;
      RECT 3674.995 1048.035 3675.275 1064.6 ;
      RECT 3627.955 1048.035 3628.235 1049.3 ;
      RECT 3624.315 1048.035 3624.595 1049.265 ;
      RECT 3620.675 1048.035 3620.955 1049.32 ;
      RECT 3617.035 1048.035 3617.315 1049.36 ;
      RECT 3613.395 1048.035 3613.675 1049.345 ;
      RECT 3609.755 1048.035 3610.035 1049.255 ;
      RECT 3550.675 1048.035 3550.955 1049.155 ;
      RECT 3546.755 1048.035 3547.035 1049.2 ;
      RECT 3542.835 1048.035 3543.115 1048.93 ;
      RECT 3538.915 1048.035 3539.195 1049.155 ;
      RECT 3534.995 1048.035 3535.275 1064.6 ;
      RECT 3487.955 1048.035 3488.235 1049.3 ;
      RECT 3484.315 1048.035 3484.595 1049.265 ;
      RECT 3480.675 1048.035 3480.955 1049.32 ;
      RECT 3477.035 1048.035 3477.315 1049.36 ;
      RECT 3473.395 1048.035 3473.675 1049.345 ;
      RECT 3469.755 1048.035 3470.035 1049.255 ;
      RECT 3410.675 1048.035 3410.955 1049.155 ;
      RECT 3406.755 1048.035 3407.035 1049.2 ;
      RECT 3402.835 1048.035 3403.115 1048.93 ;
      RECT 3398.915 1048.035 3399.195 1049.155 ;
      RECT 3394.995 1048.035 3395.275 1064.6 ;
      RECT 3347.955 1048.035 3348.235 1049.3 ;
      RECT 3344.315 1048.035 3344.595 1049.265 ;
      RECT 3340.675 1048.035 3340.955 1049.32 ;
      RECT 3337.035 1048.035 3337.315 1049.36 ;
      RECT 3333.395 1048.035 3333.675 1049.345 ;
      RECT 3329.755 1048.035 3330.035 1049.255 ;
      RECT 3270.675 1048.035 3270.955 1049.155 ;
      RECT 3266.755 1048.035 3267.035 1049.2 ;
      RECT 3262.835 1048.035 3263.115 1048.93 ;
      RECT 3258.915 1048.035 3259.195 1049.155 ;
      RECT 3254.995 1048.035 3255.275 1064.6 ;
      RECT 3207.955 1048.035 3208.235 1049.3 ;
      RECT 3204.315 1048.035 3204.595 1049.265 ;
      RECT 3200.675 1048.035 3200.955 1049.32 ;
      RECT 3197.035 1048.035 3197.315 1049.36 ;
      RECT 3193.395 1048.035 3193.675 1049.345 ;
      RECT 3189.755 1048.035 3190.035 1049.255 ;
      RECT 3130.675 1048.035 3130.955 1049.155 ;
      RECT 3126.755 1048.035 3127.035 1049.2 ;
      RECT 3122.835 1048.035 3123.115 1048.93 ;
      RECT 3118.915 1048.035 3119.195 1049.155 ;
      RECT 3114.995 1048.035 3115.275 1064.6 ;
      RECT 3067.955 1048.035 3068.235 1049.3 ;
      RECT 3064.315 1048.035 3064.595 1049.265 ;
      RECT 3060.675 1048.035 3060.955 1049.32 ;
      RECT 3057.035 1048.035 3057.315 1049.36 ;
      RECT 3053.395 1048.035 3053.675 1049.345 ;
      RECT 3049.755 1048.035 3050.035 1049.255 ;
      RECT 2990.675 1048.035 2990.955 1049.155 ;
      RECT 2986.755 1048.035 2987.035 1049.2 ;
      RECT 2982.835 1048.035 2983.115 1048.93 ;
      RECT 2978.915 1048.035 2979.195 1049.155 ;
      RECT 2974.995 1048.035 2975.275 1064.6 ;
      RECT 2927.955 1048.035 2928.235 1049.3 ;
      RECT 2924.315 1048.035 2924.595 1049.265 ;
      RECT 2920.675 1048.035 2920.955 1049.32 ;
      RECT 2917.035 1048.035 2917.315 1049.36 ;
      RECT 2913.395 1048.035 2913.675 1049.345 ;
      RECT 2909.755 1048.035 2910.035 1049.255 ;
      RECT 2850.675 1048.035 2850.955 1049.155 ;
      RECT 2846.755 1048.035 2847.035 1049.2 ;
      RECT 2842.835 1048.035 2843.115 1048.93 ;
      RECT 2838.915 1048.035 2839.195 1049.155 ;
      RECT 2834.995 1048.035 2835.275 1064.6 ;
      RECT 2787.955 1048.035 2788.235 1049.3 ;
      RECT 2784.315 1048.035 2784.595 1049.265 ;
      RECT 2780.675 1048.035 2780.955 1049.32 ;
      RECT 2777.035 1048.035 2777.315 1049.36 ;
      RECT 2773.395 1048.035 2773.675 1049.345 ;
      RECT 2769.755 1048.035 2770.035 1049.255 ;
      RECT 2710.675 1048.035 2710.955 1049.155 ;
      RECT 2706.755 1048.035 2707.035 1049.2 ;
      RECT 2702.835 1048.035 2703.115 1048.93 ;
      RECT 2698.915 1048.035 2699.195 1049.155 ;
      RECT 2694.995 1048.035 2695.275 1064.6 ;
      RECT 2647.955 1048.035 2648.235 1049.3 ;
      RECT 2644.315 1048.035 2644.595 1049.265 ;
      RECT 2640.675 1048.035 2640.955 1049.32 ;
      RECT 2637.035 1048.035 2637.315 1049.36 ;
      RECT 2633.395 1048.035 2633.675 1049.345 ;
      RECT 2629.755 1048.035 2630.035 1049.255 ;
      RECT 2570.675 1048.035 2570.955 1049.155 ;
      RECT 2566.755 1048.035 2567.035 1049.2 ;
      RECT 2562.835 1048.035 2563.115 1048.93 ;
      RECT 2558.915 1048.035 2559.195 1049.155 ;
      RECT 2554.995 1048.035 2555.275 1064.6 ;
      RECT 2507.955 1048.035 2508.235 1049.3 ;
      RECT 2504.315 1048.035 2504.595 1049.265 ;
      RECT 2500.675 1048.035 2500.955 1049.32 ;
      RECT 2497.035 1048.035 2497.315 1049.36 ;
      RECT 2493.395 1048.035 2493.675 1049.345 ;
      RECT 2489.755 1048.035 2490.035 1049.255 ;
      RECT 2430.675 1048.035 2430.955 1049.155 ;
      RECT 2426.755 1048.035 2427.035 1049.2 ;
      RECT 2422.835 1048.035 2423.115 1048.93 ;
      RECT 2418.915 1048.035 2419.195 1049.155 ;
      RECT 2414.995 1048.035 2415.275 1064.6 ;
      RECT 2367.955 1048.035 2368.235 1049.3 ;
      RECT 2364.315 1048.035 2364.595 1049.265 ;
      RECT 2360.675 1048.035 2360.955 1049.32 ;
      RECT 2357.035 1048.035 2357.315 1049.36 ;
      RECT 2353.395 1048.035 2353.675 1049.345 ;
      RECT 2349.755 1048.035 2350.035 1049.255 ;
      RECT 2290.675 1048.035 2290.955 1049.155 ;
      RECT 2286.755 1048.035 2287.035 1049.2 ;
      RECT 2282.835 1048.035 2283.115 1048.93 ;
      RECT 2278.915 1048.035 2279.195 1049.155 ;
      RECT 2274.995 1048.035 2275.275 1064.6 ;
      RECT 2227.955 1048.035 2228.235 1049.3 ;
      RECT 2224.315 1048.035 2224.595 1049.265 ;
      RECT 2220.675 1048.035 2220.955 1049.32 ;
      RECT 2217.035 1048.035 2217.315 1049.36 ;
      RECT 2213.395 1048.035 2213.675 1049.345 ;
      RECT 2209.755 1048.035 2210.035 1049.255 ;
      RECT 2150.675 1048.035 2150.955 1049.155 ;
      RECT 2146.755 1048.035 2147.035 1049.2 ;
      RECT 2142.835 1048.035 2143.115 1048.93 ;
      RECT 2138.915 1048.035 2139.195 1049.155 ;
      RECT 2134.995 1048.035 2135.275 1064.6 ;
      RECT 2087.955 1048.035 2088.235 1049.3 ;
      RECT 2084.315 1048.035 2084.595 1049.265 ;
      RECT 2080.675 1048.035 2080.955 1049.32 ;
      RECT 2077.035 1048.035 2077.315 1049.36 ;
      RECT 2073.395 1048.035 2073.675 1049.345 ;
      RECT 2069.755 1048.035 2070.035 1049.255 ;
      RECT 2010.675 1048.035 2010.955 1049.155 ;
      RECT 2006.755 1048.035 2007.035 1049.2 ;
      RECT 2002.835 1048.035 2003.115 1048.93 ;
      RECT 1998.915 1048.035 1999.195 1049.155 ;
      RECT 1994.995 1048.035 1995.275 1064.6 ;
      RECT 1947.955 1048.035 1948.235 1049.3 ;
      RECT 1944.315 1048.035 1944.595 1049.265 ;
      RECT 1940.675 1048.035 1940.955 1049.32 ;
      RECT 1937.035 1048.035 1937.315 1049.36 ;
      RECT 1933.395 1048.035 1933.675 1049.345 ;
      RECT 1929.755 1048.035 1930.035 1049.255 ;
      RECT 1870.675 1048.035 1870.955 1049.155 ;
      RECT 1866.755 1048.035 1867.035 1049.2 ;
      RECT 1862.835 1048.035 1863.115 1048.93 ;
      RECT 1858.915 1048.035 1859.195 1049.155 ;
      RECT 1854.995 1048.035 1855.275 1064.6 ;
      RECT 1807.955 1048.035 1808.235 1049.3 ;
      RECT 1804.315 1048.035 1804.595 1049.265 ;
      RECT 1800.675 1048.035 1800.955 1049.32 ;
      RECT 1797.035 1048.035 1797.315 1049.36 ;
      RECT 1793.395 1048.035 1793.675 1049.345 ;
      RECT 1789.755 1048.035 1790.035 1049.255 ;
      RECT 1730.675 1048.035 1730.955 1049.155 ;
      RECT 1726.755 1048.035 1727.035 1049.2 ;
      RECT 1722.835 1048.035 1723.115 1048.93 ;
      RECT 1718.915 1048.035 1719.195 1049.155 ;
      RECT 1714.995 1048.035 1715.275 1064.6 ;
      RECT 1667.955 1048.035 1668.235 1049.3 ;
      RECT 1664.315 1048.035 1664.595 1049.265 ;
      RECT 1660.675 1048.035 1660.955 1049.32 ;
      RECT 1657.035 1048.035 1657.315 1049.36 ;
      RECT 1653.395 1048.035 1653.675 1049.345 ;
      RECT 1649.755 1048.035 1650.035 1049.255 ;
      RECT 1590.675 1048.035 1590.955 1049.155 ;
      RECT 1586.755 1048.035 1587.035 1049.2 ;
      RECT 1582.835 1048.035 1583.115 1048.93 ;
      RECT 1578.915 1048.035 1579.195 1049.155 ;
      RECT 1574.995 1048.035 1575.275 1064.6 ;
      RECT 1527.955 1048.035 1528.235 1049.3 ;
      RECT 1524.315 1048.035 1524.595 1049.265 ;
      RECT 1520.675 1048.035 1520.955 1049.32 ;
      RECT 1517.035 1048.035 1517.315 1049.36 ;
      RECT 1513.395 1048.035 1513.675 1049.345 ;
      RECT 1509.755 1048.035 1510.035 1049.255 ;
      RECT 1450.675 1048.035 1450.955 1049.155 ;
      RECT 1446.755 1048.035 1447.035 1049.2 ;
      RECT 1442.835 1048.035 1443.115 1048.93 ;
      RECT 1438.915 1048.035 1439.195 1049.155 ;
      RECT 1434.995 1048.035 1435.275 1064.6 ;
      RECT 1387.955 1048.035 1388.235 1049.3 ;
      RECT 1384.315 1048.035 1384.595 1049.265 ;
      RECT 1380.675 1048.035 1380.955 1049.32 ;
      RECT 1377.035 1048.035 1377.315 1049.36 ;
      RECT 1373.395 1048.035 1373.675 1049.345 ;
      RECT 1369.755 1048.035 1370.035 1049.255 ;
      RECT 1310.675 1048.035 1310.955 1049.155 ;
      RECT 1306.755 1048.035 1307.035 1049.2 ;
      RECT 1302.835 1048.035 1303.115 1048.93 ;
      RECT 1298.915 1048.035 1299.195 1049.155 ;
      RECT 1294.995 1048.035 1295.275 1064.6 ;
      RECT 1247.955 1048.035 1248.235 1049.3 ;
      RECT 1244.315 1048.035 1244.595 1049.265 ;
      RECT 1240.675 1048.035 1240.955 1049.32 ;
      RECT 1237.035 1048.035 1237.315 1049.36 ;
      RECT 1233.395 1048.035 1233.675 1049.345 ;
      RECT 1229.755 1048.035 1230.035 1049.255 ;
      RECT 1170.675 1048.035 1170.955 1049.155 ;
      RECT 1166.755 1048.035 1167.035 1049.2 ;
      RECT 1162.835 1048.035 1163.115 1048.93 ;
      RECT 1158.915 1048.035 1159.195 1049.155 ;
      RECT 1154.995 1048.035 1155.275 1064.6 ;
      RECT 929.89 9258.575 1013.435 9259.995 ;
      RECT 913.47 9297.09 1013.435 9298.51 ;
      RECT 897.05 9330.58 1013.435 9332 ;
      RECT 880.63 9369.09 1013.435 9370.51 ;
      RECT 864.21 9402.575 1013.435 9403.995 ;
      RECT 847.79 9441.09 1013.435 9442.51 ;
      RECT 990 9497.56 1010 9527.56 ;
      RECT 990 9529.56 1010 9559.56 ;
      RECT 990 9617.56 1010 9647.56 ;
      RECT 990 9649.56 1010 9679.56 ;
      RECT 990 9737.56 1010 9767.56 ;
      RECT 990 9769.56 1010 9799.56 ;
      RECT 990 9857.56 1010 9887.56 ;
      RECT 990 9889.56 1010 9919.56 ;
      RECT 1007.765 1048.035 1008.045 1111.38 ;
      RECT 1007.205 1048.035 1007.485 1111.38 ;
      RECT 1006.645 1048.035 1006.925 1111.38 ;
      RECT 1006.085 1048.035 1006.365 1111.38 ;
      RECT 1005.525 1048.035 1005.805 1111.38 ;
      RECT 1004.965 1048.035 1005.245 1111.38 ;
      RECT 1004.405 1048.035 1004.685 1111.38 ;
      RECT 1003.845 1048.035 1004.125 1111.38 ;
      RECT 971.03 1116.59 1001.84 1117.79 ;
      RECT 954.83 1118.99 1001.84 1120.19 ;
      RECT 938.63 1121.39 1001.84 1122.59 ;
      RECT 922.43 1123.79 1001.84 1124.99 ;
      RECT 922.43 1126.185 1001.84 1127.385 ;
    LAYER M2 SPACING 0.28 ;
      RECT 13630.255 1047.855 19161.9 10000 ;
      RECT 19156.575 1046.435 19161.9 10000 ;
      RECT 19028.655 1046.435 19151.535 10000 ;
      RECT 19025.015 1046.435 19027.535 10000 ;
      RECT 19021.375 1046.435 19023.895 10000 ;
      RECT 19017.735 1046.435 19020.255 10000 ;
      RECT 19014.095 1046.435 19016.615 10000 ;
      RECT 19010.455 1046.435 19012.975 10000 ;
      RECT 18951.375 1046.435 19009.335 10000 ;
      RECT 18947.455 1046.435 18950.255 10000 ;
      RECT 18943.535 1046.435 18946.335 10000 ;
      RECT 18939.615 1046.435 18942.415 10000 ;
      RECT 18935.695 1046.435 18938.495 10000 ;
      RECT 18888.655 1046.435 18934.575 10000 ;
      RECT 18885.015 1046.435 18887.535 10000 ;
      RECT 18881.375 1046.435 18883.895 10000 ;
      RECT 18877.735 1046.435 18880.255 10000 ;
      RECT 18874.095 1046.435 18876.615 10000 ;
      RECT 18870.455 1046.435 18872.975 10000 ;
      RECT 18811.375 1046.435 18869.335 10000 ;
      RECT 18807.455 1046.435 18810.255 10000 ;
      RECT 18803.535 1046.435 18806.335 10000 ;
      RECT 18799.615 1046.435 18802.415 10000 ;
      RECT 18795.695 1046.435 18798.495 10000 ;
      RECT 18748.655 1046.435 18794.575 10000 ;
      RECT 18745.015 1046.435 18747.535 10000 ;
      RECT 18741.375 1046.435 18743.895 10000 ;
      RECT 18737.735 1046.435 18740.255 10000 ;
      RECT 18734.095 1046.435 18736.615 10000 ;
      RECT 18730.455 1046.435 18732.975 10000 ;
      RECT 18671.375 1046.435 18729.335 10000 ;
      RECT 18667.455 1046.435 18670.255 10000 ;
      RECT 18663.535 1046.435 18666.335 10000 ;
      RECT 18659.615 1046.435 18662.415 10000 ;
      RECT 18655.695 1046.435 18658.495 10000 ;
      RECT 18608.655 1046.435 18654.575 10000 ;
      RECT 18605.015 1046.435 18607.535 10000 ;
      RECT 18601.375 1046.435 18603.895 10000 ;
      RECT 18597.735 1046.435 18600.255 10000 ;
      RECT 18594.095 1046.435 18596.615 10000 ;
      RECT 18590.455 1046.435 18592.975 10000 ;
      RECT 18531.375 1046.435 18589.335 10000 ;
      RECT 18527.455 1046.435 18530.255 10000 ;
      RECT 18523.535 1046.435 18526.335 10000 ;
      RECT 18519.615 1046.435 18522.415 10000 ;
      RECT 18515.695 1046.435 18518.495 10000 ;
      RECT 18468.655 1046.435 18514.575 10000 ;
      RECT 18465.015 1046.435 18467.535 10000 ;
      RECT 18461.375 1046.435 18463.895 10000 ;
      RECT 18457.735 1046.435 18460.255 10000 ;
      RECT 18454.095 1046.435 18456.615 10000 ;
      RECT 18450.455 1046.435 18452.975 10000 ;
      RECT 18391.375 1046.435 18449.335 10000 ;
      RECT 18387.455 1046.435 18390.255 10000 ;
      RECT 18383.535 1046.435 18386.335 10000 ;
      RECT 18379.615 1046.435 18382.415 10000 ;
      RECT 18375.695 1046.435 18378.495 10000 ;
      RECT 18328.655 1046.435 18374.575 10000 ;
      RECT 18325.015 1046.435 18327.535 10000 ;
      RECT 18321.375 1046.435 18323.895 10000 ;
      RECT 18317.735 1046.435 18320.255 10000 ;
      RECT 18314.095 1046.435 18316.615 10000 ;
      RECT 18310.455 1046.435 18312.975 10000 ;
      RECT 18251.375 1046.435 18309.335 10000 ;
      RECT 18247.455 1046.435 18250.255 10000 ;
      RECT 18243.535 1046.435 18246.335 10000 ;
      RECT 18239.615 1046.435 18242.415 10000 ;
      RECT 18235.695 1046.435 18238.495 10000 ;
      RECT 18188.655 1046.435 18234.575 10000 ;
      RECT 18185.015 1046.435 18187.535 10000 ;
      RECT 18181.375 1046.435 18183.895 10000 ;
      RECT 18177.735 1046.435 18180.255 10000 ;
      RECT 18174.095 1046.435 18176.615 10000 ;
      RECT 18170.455 1046.435 18172.975 10000 ;
      RECT 18111.375 1046.435 18169.335 10000 ;
      RECT 18107.455 1046.435 18110.255 10000 ;
      RECT 18103.535 1046.435 18106.335 10000 ;
      RECT 18099.615 1046.435 18102.415 10000 ;
      RECT 18095.695 1046.435 18098.495 10000 ;
      RECT 18048.655 1046.435 18094.575 10000 ;
      RECT 18045.015 1046.435 18047.535 10000 ;
      RECT 18041.375 1046.435 18043.895 10000 ;
      RECT 18037.735 1046.435 18040.255 10000 ;
      RECT 18034.095 1046.435 18036.615 10000 ;
      RECT 18030.455 1046.435 18032.975 10000 ;
      RECT 17971.375 1046.435 18029.335 10000 ;
      RECT 17967.455 1046.435 17970.255 10000 ;
      RECT 17963.535 1046.435 17966.335 10000 ;
      RECT 17959.615 1046.435 17962.415 10000 ;
      RECT 17955.695 1046.435 17958.495 10000 ;
      RECT 17908.655 1046.435 17954.575 10000 ;
      RECT 17905.015 1046.435 17907.535 10000 ;
      RECT 17901.375 1046.435 17903.895 10000 ;
      RECT 17897.735 1046.435 17900.255 10000 ;
      RECT 17894.095 1046.435 17896.615 10000 ;
      RECT 17890.455 1046.435 17892.975 10000 ;
      RECT 17831.375 1046.435 17889.335 10000 ;
      RECT 17827.455 1046.435 17830.255 10000 ;
      RECT 17823.535 1046.435 17826.335 10000 ;
      RECT 17819.615 1046.435 17822.415 10000 ;
      RECT 17815.695 1046.435 17818.495 10000 ;
      RECT 17768.655 1046.435 17814.575 10000 ;
      RECT 17765.015 1046.435 17767.535 10000 ;
      RECT 17761.375 1046.435 17763.895 10000 ;
      RECT 17757.735 1046.435 17760.255 10000 ;
      RECT 17754.095 1046.435 17756.615 10000 ;
      RECT 17750.455 1046.435 17752.975 10000 ;
      RECT 17691.375 1046.435 17749.335 10000 ;
      RECT 17687.455 1046.435 17690.255 10000 ;
      RECT 17683.535 1046.435 17686.335 10000 ;
      RECT 17679.615 1046.435 17682.415 10000 ;
      RECT 17675.695 1046.435 17678.495 10000 ;
      RECT 17628.655 1046.435 17674.575 10000 ;
      RECT 17625.015 1046.435 17627.535 10000 ;
      RECT 17621.375 1046.435 17623.895 10000 ;
      RECT 17617.735 1046.435 17620.255 10000 ;
      RECT 17614.095 1046.435 17616.615 10000 ;
      RECT 17610.455 1046.435 17612.975 10000 ;
      RECT 17551.375 1046.435 17609.335 10000 ;
      RECT 17547.455 1046.435 17550.255 10000 ;
      RECT 17543.535 1046.435 17546.335 10000 ;
      RECT 17539.615 1046.435 17542.415 10000 ;
      RECT 17535.695 1046.435 17538.495 10000 ;
      RECT 17488.655 1046.435 17534.575 10000 ;
      RECT 17485.015 1046.435 17487.535 10000 ;
      RECT 17481.375 1046.435 17483.895 10000 ;
      RECT 17477.735 1046.435 17480.255 10000 ;
      RECT 17474.095 1046.435 17476.615 10000 ;
      RECT 17470.455 1046.435 17472.975 10000 ;
      RECT 17411.375 1046.435 17469.335 10000 ;
      RECT 17407.455 1046.435 17410.255 10000 ;
      RECT 17403.535 1046.435 17406.335 10000 ;
      RECT 17399.615 1046.435 17402.415 10000 ;
      RECT 17395.695 1046.435 17398.495 10000 ;
      RECT 17348.655 1046.435 17394.575 10000 ;
      RECT 17345.015 1046.435 17347.535 10000 ;
      RECT 17341.375 1046.435 17343.895 10000 ;
      RECT 17337.735 1046.435 17340.255 10000 ;
      RECT 17334.095 1046.435 17336.615 10000 ;
      RECT 17330.455 1046.435 17332.975 10000 ;
      RECT 17271.375 1046.435 17329.335 10000 ;
      RECT 17267.455 1046.435 17270.255 10000 ;
      RECT 17263.535 1046.435 17266.335 10000 ;
      RECT 17259.615 1046.435 17262.415 10000 ;
      RECT 17255.695 1046.435 17258.495 10000 ;
      RECT 17208.655 1046.435 17254.575 10000 ;
      RECT 17205.015 1046.435 17207.535 10000 ;
      RECT 17201.375 1046.435 17203.895 10000 ;
      RECT 17197.735 1046.435 17200.255 10000 ;
      RECT 17194.095 1046.435 17196.615 10000 ;
      RECT 17190.455 1046.435 17192.975 10000 ;
      RECT 17131.375 1046.435 17189.335 10000 ;
      RECT 17127.455 1046.435 17130.255 10000 ;
      RECT 17123.535 1046.435 17126.335 10000 ;
      RECT 17119.615 1046.435 17122.415 10000 ;
      RECT 17115.695 1046.435 17118.495 10000 ;
      RECT 17068.655 1046.435 17114.575 10000 ;
      RECT 17065.015 1046.435 17067.535 10000 ;
      RECT 17061.375 1046.435 17063.895 10000 ;
      RECT 17057.735 1046.435 17060.255 10000 ;
      RECT 17054.095 1046.435 17056.615 10000 ;
      RECT 17050.455 1046.435 17052.975 10000 ;
      RECT 16991.375 1046.435 17049.335 10000 ;
      RECT 16987.455 1046.435 16990.255 10000 ;
      RECT 16983.535 1046.435 16986.335 10000 ;
      RECT 16979.615 1046.435 16982.415 10000 ;
      RECT 16975.695 1046.435 16978.495 10000 ;
      RECT 16928.655 1046.435 16974.575 10000 ;
      RECT 16925.015 1046.435 16927.535 10000 ;
      RECT 16921.375 1046.435 16923.895 10000 ;
      RECT 16917.735 1046.435 16920.255 10000 ;
      RECT 16914.095 1046.435 16916.615 10000 ;
      RECT 16910.455 1046.435 16912.975 10000 ;
      RECT 16851.375 1046.435 16909.335 10000 ;
      RECT 16847.455 1046.435 16850.255 10000 ;
      RECT 16843.535 1046.435 16846.335 10000 ;
      RECT 16839.615 1046.435 16842.415 10000 ;
      RECT 16835.695 1046.435 16838.495 10000 ;
      RECT 16788.655 1046.435 16834.575 10000 ;
      RECT 16785.015 1046.435 16787.535 10000 ;
      RECT 16781.375 1046.435 16783.895 10000 ;
      RECT 16777.735 1046.435 16780.255 10000 ;
      RECT 16774.095 1046.435 16776.615 10000 ;
      RECT 16770.455 1046.435 16772.975 10000 ;
      RECT 16711.375 1046.435 16769.335 10000 ;
      RECT 16707.455 1046.435 16710.255 10000 ;
      RECT 16703.535 1046.435 16706.335 10000 ;
      RECT 16699.615 1046.435 16702.415 10000 ;
      RECT 16695.695 1046.435 16698.495 10000 ;
      RECT 16648.655 1046.435 16694.575 10000 ;
      RECT 16645.015 1046.435 16647.535 10000 ;
      RECT 16641.375 1046.435 16643.895 10000 ;
      RECT 16637.735 1046.435 16640.255 10000 ;
      RECT 16634.095 1046.435 16636.615 10000 ;
      RECT 16630.455 1046.435 16632.975 10000 ;
      RECT 16571.375 1046.435 16629.335 10000 ;
      RECT 16567.455 1046.435 16570.255 10000 ;
      RECT 16563.535 1046.435 16566.335 10000 ;
      RECT 16559.615 1046.435 16562.415 10000 ;
      RECT 16555.695 1046.435 16558.495 10000 ;
      RECT 16508.655 1046.435 16554.575 10000 ;
      RECT 16505.015 1046.435 16507.535 10000 ;
      RECT 16501.375 1046.435 16503.895 10000 ;
      RECT 16497.735 1046.435 16500.255 10000 ;
      RECT 16494.095 1046.435 16496.615 10000 ;
      RECT 16490.455 1046.435 16492.975 10000 ;
      RECT 16431.375 1046.435 16489.335 10000 ;
      RECT 16427.455 1046.435 16430.255 10000 ;
      RECT 16423.535 1046.435 16426.335 10000 ;
      RECT 16419.615 1046.435 16422.415 10000 ;
      RECT 16415.695 1046.435 16418.495 10000 ;
      RECT 16368.655 1046.435 16414.575 10000 ;
      RECT 16365.015 1046.435 16367.535 10000 ;
      RECT 16361.375 1046.435 16363.895 10000 ;
      RECT 16357.735 1046.435 16360.255 10000 ;
      RECT 16354.095 1046.435 16356.615 10000 ;
      RECT 16350.455 1046.435 16352.975 10000 ;
      RECT 16291.375 1046.435 16349.335 10000 ;
      RECT 16287.455 1046.435 16290.255 10000 ;
      RECT 16283.535 1046.435 16286.335 10000 ;
      RECT 16279.615 1046.435 16282.415 10000 ;
      RECT 16275.695 1046.435 16278.495 10000 ;
      RECT 16228.655 1046.435 16274.575 10000 ;
      RECT 16225.015 1046.435 16227.535 10000 ;
      RECT 16221.375 1046.435 16223.895 10000 ;
      RECT 16217.735 1046.435 16220.255 10000 ;
      RECT 16214.095 1046.435 16216.615 10000 ;
      RECT 16210.455 1046.435 16212.975 10000 ;
      RECT 16151.375 1046.435 16209.335 10000 ;
      RECT 16147.455 1046.435 16150.255 10000 ;
      RECT 16143.535 1046.435 16146.335 10000 ;
      RECT 16139.615 1046.435 16142.415 10000 ;
      RECT 16135.695 1046.435 16138.495 10000 ;
      RECT 16088.655 1046.435 16134.575 10000 ;
      RECT 16085.015 1046.435 16087.535 10000 ;
      RECT 16081.375 1046.435 16083.895 10000 ;
      RECT 16077.735 1046.435 16080.255 10000 ;
      RECT 16074.095 1046.435 16076.615 10000 ;
      RECT 16070.455 1046.435 16072.975 10000 ;
      RECT 16011.375 1046.435 16069.335 10000 ;
      RECT 16007.455 1046.435 16010.255 10000 ;
      RECT 16003.535 1046.435 16006.335 10000 ;
      RECT 15999.615 1046.435 16002.415 10000 ;
      RECT 15995.695 1046.435 15998.495 10000 ;
      RECT 15948.655 1046.435 15994.575 10000 ;
      RECT 15945.015 1046.435 15947.535 10000 ;
      RECT 15941.375 1046.435 15943.895 10000 ;
      RECT 15937.735 1046.435 15940.255 10000 ;
      RECT 15934.095 1046.435 15936.615 10000 ;
      RECT 15930.455 1046.435 15932.975 10000 ;
      RECT 15871.375 1046.435 15929.335 10000 ;
      RECT 15867.455 1046.435 15870.255 10000 ;
      RECT 15863.535 1046.435 15866.335 10000 ;
      RECT 15859.615 1046.435 15862.415 10000 ;
      RECT 15855.695 1046.435 15858.495 10000 ;
      RECT 15808.655 1046.435 15854.575 10000 ;
      RECT 15805.015 1046.435 15807.535 10000 ;
      RECT 15801.375 1046.435 15803.895 10000 ;
      RECT 15797.735 1046.435 15800.255 10000 ;
      RECT 15794.095 1046.435 15796.615 10000 ;
      RECT 15790.455 1046.435 15792.975 10000 ;
      RECT 15731.375 1046.435 15789.335 10000 ;
      RECT 15727.455 1046.435 15730.255 10000 ;
      RECT 15723.535 1046.435 15726.335 10000 ;
      RECT 15719.615 1046.435 15722.415 10000 ;
      RECT 15715.695 1046.435 15718.495 10000 ;
      RECT 15668.655 1046.435 15714.575 10000 ;
      RECT 15665.015 1046.435 15667.535 10000 ;
      RECT 15661.375 1046.435 15663.895 10000 ;
      RECT 15657.735 1046.435 15660.255 10000 ;
      RECT 15654.095 1046.435 15656.615 10000 ;
      RECT 15650.455 1046.435 15652.975 10000 ;
      RECT 15591.375 1046.435 15649.335 10000 ;
      RECT 15587.455 1046.435 15590.255 10000 ;
      RECT 15583.535 1046.435 15586.335 10000 ;
      RECT 15579.615 1046.435 15582.415 10000 ;
      RECT 15575.695 1046.435 15578.495 10000 ;
      RECT 15528.655 1046.435 15574.575 10000 ;
      RECT 15525.015 1046.435 15527.535 10000 ;
      RECT 15521.375 1046.435 15523.895 10000 ;
      RECT 15517.735 1046.435 15520.255 10000 ;
      RECT 15514.095 1046.435 15516.615 10000 ;
      RECT 15510.455 1046.435 15512.975 10000 ;
      RECT 15451.375 1046.435 15509.335 10000 ;
      RECT 15447.455 1046.435 15450.255 10000 ;
      RECT 15443.535 1046.435 15446.335 10000 ;
      RECT 15439.615 1046.435 15442.415 10000 ;
      RECT 15435.695 1046.435 15438.495 10000 ;
      RECT 15388.655 1046.435 15434.575 10000 ;
      RECT 15385.015 1046.435 15387.535 10000 ;
      RECT 15381.375 1046.435 15383.895 10000 ;
      RECT 15377.735 1046.435 15380.255 10000 ;
      RECT 15374.095 1046.435 15376.615 10000 ;
      RECT 15370.455 1046.435 15372.975 10000 ;
      RECT 15311.375 1046.435 15369.335 10000 ;
      RECT 15307.455 1046.435 15310.255 10000 ;
      RECT 15303.535 1046.435 15306.335 10000 ;
      RECT 15299.615 1046.435 15302.415 10000 ;
      RECT 15295.695 1046.435 15298.495 10000 ;
      RECT 15248.655 1046.435 15294.575 10000 ;
      RECT 15245.015 1046.435 15247.535 10000 ;
      RECT 15241.375 1046.435 15243.895 10000 ;
      RECT 15237.735 1046.435 15240.255 10000 ;
      RECT 15234.095 1046.435 15236.615 10000 ;
      RECT 15230.455 1046.435 15232.975 10000 ;
      RECT 15171.375 1046.435 15229.335 10000 ;
      RECT 15167.455 1046.435 15170.255 10000 ;
      RECT 15163.535 1046.435 15166.335 10000 ;
      RECT 15159.615 1046.435 15162.415 10000 ;
      RECT 15155.695 1046.435 15158.495 10000 ;
      RECT 15108.655 1046.435 15154.575 10000 ;
      RECT 15105.015 1046.435 15107.535 10000 ;
      RECT 15101.375 1046.435 15103.895 10000 ;
      RECT 15097.735 1046.435 15100.255 10000 ;
      RECT 15094.095 1046.435 15096.615 10000 ;
      RECT 15090.455 1046.435 15092.975 10000 ;
      RECT 15031.375 1046.435 15089.335 10000 ;
      RECT 15027.455 1046.435 15030.255 10000 ;
      RECT 15023.535 1046.435 15026.335 10000 ;
      RECT 15019.615 1046.435 15022.415 10000 ;
      RECT 15015.695 1046.435 15018.495 10000 ;
      RECT 14968.655 1046.435 15014.575 10000 ;
      RECT 14965.015 1046.435 14967.535 10000 ;
      RECT 14961.375 1046.435 14963.895 10000 ;
      RECT 14957.735 1046.435 14960.255 10000 ;
      RECT 14954.095 1046.435 14956.615 10000 ;
      RECT 14950.455 1046.435 14952.975 10000 ;
      RECT 14891.375 1046.435 14949.335 10000 ;
      RECT 14887.455 1046.435 14890.255 10000 ;
      RECT 14883.535 1046.435 14886.335 10000 ;
      RECT 14879.615 1046.435 14882.415 10000 ;
      RECT 14875.695 1046.435 14878.495 10000 ;
      RECT 14828.655 1046.435 14874.575 10000 ;
      RECT 14825.015 1046.435 14827.535 10000 ;
      RECT 14821.375 1046.435 14823.895 10000 ;
      RECT 14817.735 1046.435 14820.255 10000 ;
      RECT 14814.095 1046.435 14816.615 10000 ;
      RECT 14810.455 1046.435 14812.975 10000 ;
      RECT 14751.375 1046.435 14809.335 10000 ;
      RECT 14747.455 1046.435 14750.255 10000 ;
      RECT 14743.535 1046.435 14746.335 10000 ;
      RECT 14739.615 1046.435 14742.415 10000 ;
      RECT 14735.695 1046.435 14738.495 10000 ;
      RECT 14688.655 1046.435 14734.575 10000 ;
      RECT 14685.015 1046.435 14687.535 10000 ;
      RECT 14681.375 1046.435 14683.895 10000 ;
      RECT 14677.735 1046.435 14680.255 10000 ;
      RECT 14674.095 1046.435 14676.615 10000 ;
      RECT 14670.455 1046.435 14672.975 10000 ;
      RECT 14611.375 1046.435 14669.335 10000 ;
      RECT 14607.455 1046.435 14610.255 10000 ;
      RECT 14603.535 1046.435 14606.335 10000 ;
      RECT 14599.615 1046.435 14602.415 10000 ;
      RECT 14595.695 1046.435 14598.495 10000 ;
      RECT 14548.655 1046.435 14594.575 10000 ;
      RECT 14545.015 1046.435 14547.535 10000 ;
      RECT 14541.375 1046.435 14543.895 10000 ;
      RECT 14537.735 1046.435 14540.255 10000 ;
      RECT 14534.095 1046.435 14536.615 10000 ;
      RECT 14530.455 1046.435 14532.975 10000 ;
      RECT 14471.375 1046.435 14529.335 10000 ;
      RECT 14467.455 1046.435 14470.255 10000 ;
      RECT 14463.535 1046.435 14466.335 10000 ;
      RECT 14459.615 1046.435 14462.415 10000 ;
      RECT 14455.695 1046.435 14458.495 10000 ;
      RECT 14408.655 1046.435 14454.575 10000 ;
      RECT 14405.015 1046.435 14407.535 10000 ;
      RECT 14401.375 1046.435 14403.895 10000 ;
      RECT 14397.735 1046.435 14400.255 10000 ;
      RECT 14394.095 1046.435 14396.615 10000 ;
      RECT 14390.455 1046.435 14392.975 10000 ;
      RECT 14331.375 1046.435 14389.335 10000 ;
      RECT 14327.455 1046.435 14330.255 10000 ;
      RECT 14323.535 1046.435 14326.335 10000 ;
      RECT 14319.615 1046.435 14322.415 10000 ;
      RECT 14315.695 1046.435 14318.495 10000 ;
      RECT 14268.655 1046.435 14314.575 10000 ;
      RECT 14265.015 1046.435 14267.535 10000 ;
      RECT 14261.375 1046.435 14263.895 10000 ;
      RECT 14257.735 1046.435 14260.255 10000 ;
      RECT 14254.095 1046.435 14256.615 10000 ;
      RECT 14250.455 1046.435 14252.975 10000 ;
      RECT 14191.375 1046.435 14249.335 10000 ;
      RECT 14187.455 1046.435 14190.255 10000 ;
      RECT 14183.535 1046.435 14186.335 10000 ;
      RECT 14179.615 1046.435 14182.415 10000 ;
      RECT 14175.695 1046.435 14178.495 10000 ;
      RECT 14128.655 1046.435 14174.575 10000 ;
      RECT 14125.015 1046.435 14127.535 10000 ;
      RECT 14121.375 1046.435 14123.895 10000 ;
      RECT 14117.735 1046.435 14120.255 10000 ;
      RECT 14114.095 1046.435 14116.615 10000 ;
      RECT 14110.455 1046.435 14112.975 10000 ;
      RECT 14051.375 1046.435 14109.335 10000 ;
      RECT 14047.455 1046.435 14050.255 10000 ;
      RECT 14043.535 1046.435 14046.335 10000 ;
      RECT 14039.615 1046.435 14042.415 10000 ;
      RECT 14035.695 1046.435 14038.495 10000 ;
      RECT 13988.655 1046.435 14034.575 10000 ;
      RECT 13985.015 1046.435 13987.535 10000 ;
      RECT 13981.375 1046.435 13983.895 10000 ;
      RECT 13977.735 1046.435 13980.255 10000 ;
      RECT 13974.095 1046.435 13976.615 10000 ;
      RECT 13970.455 1046.435 13972.975 10000 ;
      RECT 13911.375 1046.435 13969.335 10000 ;
      RECT 13907.455 1046.435 13910.255 10000 ;
      RECT 13903.535 1046.435 13906.335 10000 ;
      RECT 13899.615 1046.435 13902.415 10000 ;
      RECT 13895.695 1046.435 13898.495 10000 ;
      RECT 13848.655 1046.435 13894.575 10000 ;
      RECT 13845.015 1046.435 13847.535 10000 ;
      RECT 13841.375 1046.435 13843.895 10000 ;
      RECT 13837.735 1046.435 13840.255 10000 ;
      RECT 13834.095 1046.435 13836.615 10000 ;
      RECT 13830.455 1046.435 13832.975 10000 ;
      RECT 13771.375 1046.435 13829.335 10000 ;
      RECT 13767.455 1046.435 13770.255 10000 ;
      RECT 13763.535 1046.435 13766.335 10000 ;
      RECT 13759.615 1046.435 13762.415 10000 ;
      RECT 13755.695 1046.435 13758.495 10000 ;
      RECT 13708.655 1046.435 13754.575 10000 ;
      RECT 13705.015 1046.435 13707.535 10000 ;
      RECT 13701.375 1046.435 13703.895 10000 ;
      RECT 13697.735 1046.435 13700.255 10000 ;
      RECT 13694.095 1046.435 13696.615 10000 ;
      RECT 13690.455 1046.435 13692.975 10000 ;
      RECT 13631.375 1046.435 13689.335 10000 ;
      RECT 998.1 1047.855 13630.255 10000 ;
      RECT 13627.455 1046.435 13630.255 10000 ;
      RECT 13623.535 1046.435 13626.335 10000 ;
      RECT 13619.615 1046.435 13622.415 10000 ;
      RECT 13615.695 1046.435 13618.495 10000 ;
      RECT 13568.655 1046.435 13614.575 10000 ;
      RECT 13565.015 1046.435 13567.535 10000 ;
      RECT 13561.375 1046.435 13563.895 10000 ;
      RECT 13557.735 1046.435 13560.255 10000 ;
      RECT 13554.095 1046.435 13556.615 10000 ;
      RECT 13550.455 1046.435 13552.975 10000 ;
      RECT 13491.375 1046.435 13549.335 10000 ;
      RECT 13487.455 1046.435 13490.255 10000 ;
      RECT 13483.535 1046.435 13486.335 10000 ;
      RECT 13479.615 1046.435 13482.415 10000 ;
      RECT 13475.695 1046.435 13478.495 10000 ;
      RECT 13428.655 1046.435 13474.575 10000 ;
      RECT 13425.015 1046.435 13427.535 10000 ;
      RECT 13421.375 1046.435 13423.895 10000 ;
      RECT 13417.735 1046.435 13420.255 10000 ;
      RECT 13414.095 1046.435 13416.615 10000 ;
      RECT 13410.455 1046.435 13412.975 10000 ;
      RECT 13351.375 1046.435 13409.335 10000 ;
      RECT 13347.455 1046.435 13350.255 10000 ;
      RECT 13343.535 1046.435 13346.335 10000 ;
      RECT 13339.615 1046.435 13342.415 10000 ;
      RECT 13335.695 1046.435 13338.495 10000 ;
      RECT 13288.655 1046.435 13334.575 10000 ;
      RECT 13285.015 1046.435 13287.535 10000 ;
      RECT 13281.375 1046.435 13283.895 10000 ;
      RECT 13277.735 1046.435 13280.255 10000 ;
      RECT 13274.095 1046.435 13276.615 10000 ;
      RECT 13270.455 1046.435 13272.975 10000 ;
      RECT 13211.375 1046.435 13269.335 10000 ;
      RECT 13207.455 1046.435 13210.255 10000 ;
      RECT 13203.535 1046.435 13206.335 10000 ;
      RECT 13199.615 1046.435 13202.415 10000 ;
      RECT 13195.695 1046.435 13198.495 10000 ;
      RECT 13148.655 1046.435 13194.575 10000 ;
      RECT 13145.015 1046.435 13147.535 10000 ;
      RECT 13141.375 1046.435 13143.895 10000 ;
      RECT 13137.735 1046.435 13140.255 10000 ;
      RECT 13134.095 1046.435 13136.615 10000 ;
      RECT 13130.455 1046.435 13132.975 10000 ;
      RECT 13071.375 1046.435 13129.335 10000 ;
      RECT 13067.455 1046.435 13070.255 10000 ;
      RECT 13063.535 1046.435 13066.335 10000 ;
      RECT 13059.615 1046.435 13062.415 10000 ;
      RECT 13055.695 1046.435 13058.495 10000 ;
      RECT 13008.655 1046.435 13054.575 10000 ;
      RECT 13005.015 1046.435 13007.535 10000 ;
      RECT 13001.375 1046.435 13003.895 10000 ;
      RECT 12997.735 1046.435 13000.255 10000 ;
      RECT 12994.095 1046.435 12996.615 10000 ;
      RECT 12990.455 1046.435 12992.975 10000 ;
      RECT 12931.375 1046.435 12989.335 10000 ;
      RECT 12927.455 1046.435 12930.255 10000 ;
      RECT 12923.535 1046.435 12926.335 10000 ;
      RECT 12919.615 1046.435 12922.415 10000 ;
      RECT 12915.695 1046.435 12918.495 10000 ;
      RECT 12868.655 1046.435 12914.575 10000 ;
      RECT 12865.015 1046.435 12867.535 10000 ;
      RECT 12861.375 1046.435 12863.895 10000 ;
      RECT 12857.735 1046.435 12860.255 10000 ;
      RECT 12854.095 1046.435 12856.615 10000 ;
      RECT 12850.455 1046.435 12852.975 10000 ;
      RECT 12791.375 1046.435 12849.335 10000 ;
      RECT 12787.455 1046.435 12790.255 10000 ;
      RECT 12783.535 1046.435 12786.335 10000 ;
      RECT 12779.615 1046.435 12782.415 10000 ;
      RECT 12775.695 1046.435 12778.495 10000 ;
      RECT 12728.655 1046.435 12774.575 10000 ;
      RECT 12725.015 1046.435 12727.535 10000 ;
      RECT 12721.375 1046.435 12723.895 10000 ;
      RECT 12717.735 1046.435 12720.255 10000 ;
      RECT 12714.095 1046.435 12716.615 10000 ;
      RECT 12710.455 1046.435 12712.975 10000 ;
      RECT 12651.375 1046.435 12709.335 10000 ;
      RECT 12647.455 1046.435 12650.255 10000 ;
      RECT 12643.535 1046.435 12646.335 10000 ;
      RECT 12639.615 1046.435 12642.415 10000 ;
      RECT 12635.695 1046.435 12638.495 10000 ;
      RECT 12588.655 1046.435 12634.575 10000 ;
      RECT 12585.015 1046.435 12587.535 10000 ;
      RECT 12581.375 1046.435 12583.895 10000 ;
      RECT 12577.735 1046.435 12580.255 10000 ;
      RECT 12574.095 1046.435 12576.615 10000 ;
      RECT 12570.455 1046.435 12572.975 10000 ;
      RECT 12511.375 1046.435 12569.335 10000 ;
      RECT 12507.455 1046.435 12510.255 10000 ;
      RECT 12503.535 1046.435 12506.335 10000 ;
      RECT 12499.615 1046.435 12502.415 10000 ;
      RECT 12495.695 1046.435 12498.495 10000 ;
      RECT 12448.655 1046.435 12494.575 10000 ;
      RECT 12445.015 1046.435 12447.535 10000 ;
      RECT 12441.375 1046.435 12443.895 10000 ;
      RECT 12437.735 1046.435 12440.255 10000 ;
      RECT 12434.095 1046.435 12436.615 10000 ;
      RECT 12430.455 1046.435 12432.975 10000 ;
      RECT 12371.375 1046.435 12429.335 10000 ;
      RECT 12367.455 1046.435 12370.255 10000 ;
      RECT 12363.535 1046.435 12366.335 10000 ;
      RECT 12359.615 1046.435 12362.415 10000 ;
      RECT 12355.695 1046.435 12358.495 10000 ;
      RECT 12308.655 1046.435 12354.575 10000 ;
      RECT 12305.015 1046.435 12307.535 10000 ;
      RECT 12301.375 1046.435 12303.895 10000 ;
      RECT 12297.735 1046.435 12300.255 10000 ;
      RECT 12294.095 1046.435 12296.615 10000 ;
      RECT 12290.455 1046.435 12292.975 10000 ;
      RECT 12231.375 1046.435 12289.335 10000 ;
      RECT 12227.455 1046.435 12230.255 10000 ;
      RECT 12223.535 1046.435 12226.335 10000 ;
      RECT 12219.615 1046.435 12222.415 10000 ;
      RECT 12215.695 1046.435 12218.495 10000 ;
      RECT 12168.655 1046.435 12214.575 10000 ;
      RECT 12165.015 1046.435 12167.535 10000 ;
      RECT 12161.375 1046.435 12163.895 10000 ;
      RECT 12157.735 1046.435 12160.255 10000 ;
      RECT 12154.095 1046.435 12156.615 10000 ;
      RECT 12150.455 1046.435 12152.975 10000 ;
      RECT 12091.375 1046.435 12149.335 10000 ;
      RECT 12087.455 1046.435 12090.255 10000 ;
      RECT 12083.535 1046.435 12086.335 10000 ;
      RECT 12079.615 1046.435 12082.415 10000 ;
      RECT 12075.695 1046.435 12078.495 10000 ;
      RECT 12028.655 1046.435 12074.575 10000 ;
      RECT 12025.015 1046.435 12027.535 10000 ;
      RECT 12021.375 1046.435 12023.895 10000 ;
      RECT 12017.735 1046.435 12020.255 10000 ;
      RECT 12014.095 1046.435 12016.615 10000 ;
      RECT 12010.455 1046.435 12012.975 10000 ;
      RECT 11951.375 1046.435 12009.335 10000 ;
      RECT 11947.455 1046.435 11950.255 10000 ;
      RECT 11943.535 1046.435 11946.335 10000 ;
      RECT 11939.615 1046.435 11942.415 10000 ;
      RECT 11935.695 1046.435 11938.495 10000 ;
      RECT 11888.655 1046.435 11934.575 10000 ;
      RECT 11885.015 1046.435 11887.535 10000 ;
      RECT 11881.375 1046.435 11883.895 10000 ;
      RECT 11877.735 1046.435 11880.255 10000 ;
      RECT 11874.095 1046.435 11876.615 10000 ;
      RECT 11870.455 1046.435 11872.975 10000 ;
      RECT 11811.375 1046.435 11869.335 10000 ;
      RECT 11807.455 1046.435 11810.255 10000 ;
      RECT 11803.535 1046.435 11806.335 10000 ;
      RECT 11799.615 1046.435 11802.415 10000 ;
      RECT 11795.695 1046.435 11798.495 10000 ;
      RECT 11748.655 1046.435 11794.575 10000 ;
      RECT 11745.015 1046.435 11747.535 10000 ;
      RECT 11741.375 1046.435 11743.895 10000 ;
      RECT 11737.735 1046.435 11740.255 10000 ;
      RECT 11734.095 1046.435 11736.615 10000 ;
      RECT 11730.455 1046.435 11732.975 10000 ;
      RECT 11671.375 1046.435 11729.335 10000 ;
      RECT 11667.455 1046.435 11670.255 10000 ;
      RECT 11663.535 1046.435 11666.335 10000 ;
      RECT 11659.615 1046.435 11662.415 10000 ;
      RECT 11655.695 1046.435 11658.495 10000 ;
      RECT 11608.655 1046.435 11654.575 10000 ;
      RECT 11605.015 1046.435 11607.535 10000 ;
      RECT 11601.375 1046.435 11603.895 10000 ;
      RECT 11597.735 1046.435 11600.255 10000 ;
      RECT 11594.095 1046.435 11596.615 10000 ;
      RECT 11590.455 1046.435 11592.975 10000 ;
      RECT 11531.375 1046.435 11589.335 10000 ;
      RECT 11527.455 1046.435 11530.255 10000 ;
      RECT 11523.535 1046.435 11526.335 10000 ;
      RECT 11519.615 1046.435 11522.415 10000 ;
      RECT 11515.695 1046.435 11518.495 10000 ;
      RECT 11468.655 1046.435 11514.575 10000 ;
      RECT 11465.015 1046.435 11467.535 10000 ;
      RECT 11461.375 1046.435 11463.895 10000 ;
      RECT 11457.735 1046.435 11460.255 10000 ;
      RECT 11454.095 1046.435 11456.615 10000 ;
      RECT 11450.455 1046.435 11452.975 10000 ;
      RECT 11391.375 1046.435 11449.335 10000 ;
      RECT 11387.455 1046.435 11390.255 10000 ;
      RECT 11383.535 1046.435 11386.335 10000 ;
      RECT 11379.615 1046.435 11382.415 10000 ;
      RECT 11375.695 1046.435 11378.495 10000 ;
      RECT 11328.655 1046.435 11374.575 10000 ;
      RECT 11325.015 1046.435 11327.535 10000 ;
      RECT 11321.375 1046.435 11323.895 10000 ;
      RECT 11317.735 1046.435 11320.255 10000 ;
      RECT 11314.095 1046.435 11316.615 10000 ;
      RECT 11310.455 1046.435 11312.975 10000 ;
      RECT 11251.375 1046.435 11309.335 10000 ;
      RECT 11247.455 1046.435 11250.255 10000 ;
      RECT 11243.535 1046.435 11246.335 10000 ;
      RECT 11239.615 1046.435 11242.415 10000 ;
      RECT 11235.695 1046.435 11238.495 10000 ;
      RECT 11188.655 1046.435 11234.575 10000 ;
      RECT 11185.015 1046.435 11187.535 10000 ;
      RECT 11181.375 1046.435 11183.895 10000 ;
      RECT 11177.735 1046.435 11180.255 10000 ;
      RECT 11174.095 1046.435 11176.615 10000 ;
      RECT 11170.455 1046.435 11172.975 10000 ;
      RECT 11111.375 1046.435 11169.335 10000 ;
      RECT 11107.455 1046.435 11110.255 10000 ;
      RECT 11103.535 1046.435 11106.335 10000 ;
      RECT 11099.615 1046.435 11102.415 10000 ;
      RECT 11095.695 1046.435 11098.495 10000 ;
      RECT 11048.655 1046.435 11094.575 10000 ;
      RECT 11045.015 1046.435 11047.535 10000 ;
      RECT 11041.375 1046.435 11043.895 10000 ;
      RECT 11037.735 1046.435 11040.255 10000 ;
      RECT 11034.095 1046.435 11036.615 10000 ;
      RECT 11030.455 1046.435 11032.975 10000 ;
      RECT 10971.375 1046.435 11029.335 10000 ;
      RECT 10967.455 1046.435 10970.255 10000 ;
      RECT 10963.535 1046.435 10966.335 10000 ;
      RECT 10959.615 1046.435 10962.415 10000 ;
      RECT 10955.695 1046.435 10958.495 10000 ;
      RECT 10908.655 1046.435 10954.575 10000 ;
      RECT 10905.015 1046.435 10907.535 10000 ;
      RECT 10901.375 1046.435 10903.895 10000 ;
      RECT 10897.735 1046.435 10900.255 10000 ;
      RECT 10894.095 1046.435 10896.615 10000 ;
      RECT 10890.455 1046.435 10892.975 10000 ;
      RECT 10831.375 1046.435 10889.335 10000 ;
      RECT 10827.455 1046.435 10830.255 10000 ;
      RECT 10823.535 1046.435 10826.335 10000 ;
      RECT 10819.615 1046.435 10822.415 10000 ;
      RECT 10815.695 1046.435 10818.495 10000 ;
      RECT 10768.655 1046.435 10814.575 10000 ;
      RECT 10765.015 1046.435 10767.535 10000 ;
      RECT 10761.375 1046.435 10763.895 10000 ;
      RECT 10757.735 1046.435 10760.255 10000 ;
      RECT 10754.095 1046.435 10756.615 10000 ;
      RECT 10750.455 1046.435 10752.975 10000 ;
      RECT 10691.375 1046.435 10749.335 10000 ;
      RECT 10687.455 1046.435 10690.255 10000 ;
      RECT 10683.535 1046.435 10686.335 10000 ;
      RECT 10679.615 1046.435 10682.415 10000 ;
      RECT 10675.695 1046.435 10678.495 10000 ;
      RECT 10628.655 1046.435 10674.575 10000 ;
      RECT 10625.015 1046.435 10627.535 10000 ;
      RECT 10621.375 1046.435 10623.895 10000 ;
      RECT 10617.735 1046.435 10620.255 10000 ;
      RECT 10614.095 1046.435 10616.615 10000 ;
      RECT 10610.455 1046.435 10612.975 10000 ;
      RECT 10551.375 1046.435 10609.335 10000 ;
      RECT 10547.455 1046.435 10550.255 10000 ;
      RECT 10543.535 1046.435 10546.335 10000 ;
      RECT 10539.615 1046.435 10542.415 10000 ;
      RECT 10535.695 1046.435 10538.495 10000 ;
      RECT 10488.655 1046.435 10534.575 10000 ;
      RECT 10485.015 1046.435 10487.535 10000 ;
      RECT 10481.375 1046.435 10483.895 10000 ;
      RECT 10477.735 1046.435 10480.255 10000 ;
      RECT 10474.095 1046.435 10476.615 10000 ;
      RECT 10470.455 1046.435 10472.975 10000 ;
      RECT 10411.375 1046.435 10469.335 10000 ;
      RECT 10407.455 1046.435 10410.255 10000 ;
      RECT 10403.535 1046.435 10406.335 10000 ;
      RECT 10399.615 1046.435 10402.415 10000 ;
      RECT 10395.695 1046.435 10398.495 10000 ;
      RECT 10348.655 1046.435 10394.575 10000 ;
      RECT 10345.015 1046.435 10347.535 10000 ;
      RECT 10341.375 1046.435 10343.895 10000 ;
      RECT 10337.735 1046.435 10340.255 10000 ;
      RECT 10334.095 1046.435 10336.615 10000 ;
      RECT 10330.455 1046.435 10332.975 10000 ;
      RECT 10271.375 1046.435 10329.335 10000 ;
      RECT 10267.455 1046.435 10270.255 10000 ;
      RECT 10263.535 1046.435 10266.335 10000 ;
      RECT 10259.615 1046.435 10262.415 10000 ;
      RECT 10255.695 1046.435 10258.495 10000 ;
      RECT 10208.655 1046.435 10254.575 10000 ;
      RECT 10205.015 1046.435 10207.535 10000 ;
      RECT 10201.375 1046.435 10203.895 10000 ;
      RECT 10197.735 1046.435 10200.255 10000 ;
      RECT 10194.095 1046.435 10196.615 10000 ;
      RECT 10190.455 1046.435 10192.975 10000 ;
      RECT 10131.375 1046.435 10189.335 10000 ;
      RECT 10127.455 1046.435 10130.255 10000 ;
      RECT 10123.535 1046.435 10126.335 10000 ;
      RECT 10119.615 1046.435 10122.415 10000 ;
      RECT 10115.695 1046.435 10118.495 10000 ;
      RECT 10102.375 1047.71 10114.575 10000 ;
      RECT 10104.055 1046.435 10114.575 10000 ;
      RECT 10100.695 1046.435 10100.975 10000 ;
      RECT 10099.015 1046.435 10099.295 10000 ;
      RECT 10097.335 1046.435 10097.615 10000 ;
      RECT 10095.655 1046.435 10095.935 10000 ;
      RECT 10093.975 1046.435 10094.255 10000 ;
      RECT 10092.295 1046.435 10092.575 10000 ;
      RECT 10090.615 1046.435 10090.895 10000 ;
      RECT 10088.935 1046.435 10089.215 10000 ;
      RECT 10087.255 1046.435 10087.535 10000 ;
      RECT 10085.575 1046.435 10085.855 10000 ;
      RECT 10083.895 1046.435 10084.175 10000 ;
      RECT 10082.215 1046.435 10082.495 10000 ;
      RECT 10080.535 1046.435 10080.815 10000 ;
      RECT 10068.655 1046.435 10079.135 10000 ;
      RECT 10065.015 1046.435 10067.535 10000 ;
      RECT 10061.375 1046.435 10063.895 10000 ;
      RECT 10057.735 1046.435 10060.255 10000 ;
      RECT 10054.095 1046.435 10056.615 10000 ;
      RECT 10050.455 1046.435 10052.975 10000 ;
      RECT 9991.375 1046.435 10049.335 10000 ;
      RECT 9987.455 1046.435 9990.255 10000 ;
      RECT 9983.535 1046.435 9986.335 10000 ;
      RECT 9979.615 1046.435 9982.415 10000 ;
      RECT 9975.695 1046.435 9978.495 10000 ;
      RECT 9928.655 1046.435 9974.575 10000 ;
      RECT 9925.015 1046.435 9927.535 10000 ;
      RECT 9921.375 1046.435 9923.895 10000 ;
      RECT 9917.735 1046.435 9920.255 10000 ;
      RECT 9914.095 1046.435 9916.615 10000 ;
      RECT 9910.455 1046.435 9912.975 10000 ;
      RECT 9851.375 1046.435 9909.335 10000 ;
      RECT 9847.455 1046.435 9850.255 10000 ;
      RECT 9843.535 1046.435 9846.335 10000 ;
      RECT 9839.615 1046.435 9842.415 10000 ;
      RECT 9835.695 1046.435 9838.495 10000 ;
      RECT 9788.655 1046.435 9834.575 10000 ;
      RECT 9785.015 1046.435 9787.535 10000 ;
      RECT 9781.375 1046.435 9783.895 10000 ;
      RECT 9777.735 1046.435 9780.255 10000 ;
      RECT 9774.095 1046.435 9776.615 10000 ;
      RECT 9770.455 1046.435 9772.975 10000 ;
      RECT 9711.375 1046.435 9769.335 10000 ;
      RECT 9707.455 1046.435 9710.255 10000 ;
      RECT 9703.535 1046.435 9706.335 10000 ;
      RECT 9699.615 1046.435 9702.415 10000 ;
      RECT 9695.695 1046.435 9698.495 10000 ;
      RECT 9648.655 1046.435 9694.575 10000 ;
      RECT 9645.015 1046.435 9647.535 10000 ;
      RECT 9641.375 1046.435 9643.895 10000 ;
      RECT 9637.735 1046.435 9640.255 10000 ;
      RECT 9634.095 1046.435 9636.615 10000 ;
      RECT 9630.455 1046.435 9632.975 10000 ;
      RECT 9571.375 1046.435 9629.335 10000 ;
      RECT 9567.455 1046.435 9570.255 10000 ;
      RECT 9563.535 1046.435 9566.335 10000 ;
      RECT 9559.615 1046.435 9562.415 10000 ;
      RECT 9555.695 1046.435 9558.495 10000 ;
      RECT 9508.655 1046.435 9554.575 10000 ;
      RECT 9505.015 1046.435 9507.535 10000 ;
      RECT 9501.375 1046.435 9503.895 10000 ;
      RECT 9497.735 1046.435 9500.255 10000 ;
      RECT 9494.095 1046.435 9496.615 10000 ;
      RECT 9490.455 1046.435 9492.975 10000 ;
      RECT 9431.375 1046.435 9489.335 10000 ;
      RECT 9427.455 1046.435 9430.255 10000 ;
      RECT 9423.535 1046.435 9426.335 10000 ;
      RECT 9419.615 1046.435 9422.415 10000 ;
      RECT 9415.695 1046.435 9418.495 10000 ;
      RECT 9368.655 1046.435 9414.575 10000 ;
      RECT 9365.015 1046.435 9367.535 10000 ;
      RECT 9361.375 1046.435 9363.895 10000 ;
      RECT 9357.735 1046.435 9360.255 10000 ;
      RECT 9354.095 1046.435 9356.615 10000 ;
      RECT 9350.455 1046.435 9352.975 10000 ;
      RECT 9291.375 1046.435 9349.335 10000 ;
      RECT 9287.455 1046.435 9290.255 10000 ;
      RECT 9283.535 1046.435 9286.335 10000 ;
      RECT 9279.615 1046.435 9282.415 10000 ;
      RECT 9275.695 1046.435 9278.495 10000 ;
      RECT 9228.655 1046.435 9274.575 10000 ;
      RECT 9225.015 1046.435 9227.535 10000 ;
      RECT 9221.375 1046.435 9223.895 10000 ;
      RECT 9217.735 1046.435 9220.255 10000 ;
      RECT 9214.095 1046.435 9216.615 10000 ;
      RECT 9210.455 1046.435 9212.975 10000 ;
      RECT 9151.375 1046.435 9209.335 10000 ;
      RECT 9147.455 1046.435 9150.255 10000 ;
      RECT 9143.535 1046.435 9146.335 10000 ;
      RECT 9139.615 1046.435 9142.415 10000 ;
      RECT 9135.695 1046.435 9138.495 10000 ;
      RECT 9088.655 1046.435 9134.575 10000 ;
      RECT 9085.015 1046.435 9087.535 10000 ;
      RECT 9081.375 1046.435 9083.895 10000 ;
      RECT 9077.735 1046.435 9080.255 10000 ;
      RECT 9074.095 1046.435 9076.615 10000 ;
      RECT 9070.455 1046.435 9072.975 10000 ;
      RECT 9011.375 1046.435 9069.335 10000 ;
      RECT 9007.455 1046.435 9010.255 10000 ;
      RECT 9003.535 1046.435 9006.335 10000 ;
      RECT 8999.615 1046.435 9002.415 10000 ;
      RECT 8995.695 1046.435 8998.495 10000 ;
      RECT 8948.655 1046.435 8994.575 10000 ;
      RECT 8945.015 1046.435 8947.535 10000 ;
      RECT 8941.375 1046.435 8943.895 10000 ;
      RECT 8937.735 1046.435 8940.255 10000 ;
      RECT 8934.095 1046.435 8936.615 10000 ;
      RECT 8930.455 1046.435 8932.975 10000 ;
      RECT 8871.375 1046.435 8929.335 10000 ;
      RECT 8867.455 1046.435 8870.255 10000 ;
      RECT 8863.535 1046.435 8866.335 10000 ;
      RECT 8859.615 1046.435 8862.415 10000 ;
      RECT 8855.695 1046.435 8858.495 10000 ;
      RECT 8808.655 1046.435 8854.575 10000 ;
      RECT 8805.015 1046.435 8807.535 10000 ;
      RECT 8801.375 1046.435 8803.895 10000 ;
      RECT 8797.735 1046.435 8800.255 10000 ;
      RECT 8794.095 1046.435 8796.615 10000 ;
      RECT 8790.455 1046.435 8792.975 10000 ;
      RECT 8731.375 1046.435 8789.335 10000 ;
      RECT 8727.455 1046.435 8730.255 10000 ;
      RECT 8723.535 1046.435 8726.335 10000 ;
      RECT 8719.615 1046.435 8722.415 10000 ;
      RECT 8715.695 1046.435 8718.495 10000 ;
      RECT 8668.655 1046.435 8714.575 10000 ;
      RECT 8665.015 1046.435 8667.535 10000 ;
      RECT 8661.375 1046.435 8663.895 10000 ;
      RECT 8657.735 1046.435 8660.255 10000 ;
      RECT 8654.095 1046.435 8656.615 10000 ;
      RECT 8650.455 1046.435 8652.975 10000 ;
      RECT 8591.375 1046.435 8649.335 10000 ;
      RECT 8587.455 1046.435 8590.255 10000 ;
      RECT 8583.535 1046.435 8586.335 10000 ;
      RECT 8579.615 1046.435 8582.415 10000 ;
      RECT 8575.695 1046.435 8578.495 10000 ;
      RECT 8528.655 1046.435 8574.575 10000 ;
      RECT 8525.015 1046.435 8527.535 10000 ;
      RECT 8521.375 1046.435 8523.895 10000 ;
      RECT 8517.735 1046.435 8520.255 10000 ;
      RECT 8514.095 1046.435 8516.615 10000 ;
      RECT 8510.455 1046.435 8512.975 10000 ;
      RECT 8451.375 1046.435 8509.335 10000 ;
      RECT 8447.455 1046.435 8450.255 10000 ;
      RECT 8443.535 1046.435 8446.335 10000 ;
      RECT 8439.615 1046.435 8442.415 10000 ;
      RECT 8435.695 1046.435 8438.495 10000 ;
      RECT 8388.655 1046.435 8434.575 10000 ;
      RECT 8385.015 1046.435 8387.535 10000 ;
      RECT 8381.375 1046.435 8383.895 10000 ;
      RECT 8377.735 1046.435 8380.255 10000 ;
      RECT 8374.095 1046.435 8376.615 10000 ;
      RECT 8370.455 1046.435 8372.975 10000 ;
      RECT 8311.375 1046.435 8369.335 10000 ;
      RECT 8307.455 1046.435 8310.255 10000 ;
      RECT 8303.535 1046.435 8306.335 10000 ;
      RECT 8299.615 1046.435 8302.415 10000 ;
      RECT 8295.695 1046.435 8298.495 10000 ;
      RECT 8248.655 1046.435 8294.575 10000 ;
      RECT 8245.015 1046.435 8247.535 10000 ;
      RECT 8241.375 1046.435 8243.895 10000 ;
      RECT 8237.735 1046.435 8240.255 10000 ;
      RECT 8234.095 1046.435 8236.615 10000 ;
      RECT 8230.455 1046.435 8232.975 10000 ;
      RECT 8171.375 1046.435 8229.335 10000 ;
      RECT 8167.455 1046.435 8170.255 10000 ;
      RECT 8163.535 1046.435 8166.335 10000 ;
      RECT 8159.615 1046.435 8162.415 10000 ;
      RECT 8155.695 1046.435 8158.495 10000 ;
      RECT 8108.655 1046.435 8154.575 10000 ;
      RECT 8105.015 1046.435 8107.535 10000 ;
      RECT 8101.375 1046.435 8103.895 10000 ;
      RECT 8097.735 1046.435 8100.255 10000 ;
      RECT 8094.095 1046.435 8096.615 10000 ;
      RECT 8090.455 1046.435 8092.975 10000 ;
      RECT 8031.375 1046.435 8089.335 10000 ;
      RECT 8027.455 1046.435 8030.255 10000 ;
      RECT 8023.535 1046.435 8026.335 10000 ;
      RECT 8019.615 1046.435 8022.415 10000 ;
      RECT 8015.695 1046.435 8018.495 10000 ;
      RECT 7968.655 1046.435 8014.575 10000 ;
      RECT 7965.015 1046.435 7967.535 10000 ;
      RECT 7961.375 1046.435 7963.895 10000 ;
      RECT 7957.735 1046.435 7960.255 10000 ;
      RECT 7954.095 1046.435 7956.615 10000 ;
      RECT 7950.455 1046.435 7952.975 10000 ;
      RECT 7891.375 1046.435 7949.335 10000 ;
      RECT 7887.455 1046.435 7890.255 10000 ;
      RECT 7883.535 1046.435 7886.335 10000 ;
      RECT 7879.615 1046.435 7882.415 10000 ;
      RECT 7875.695 1046.435 7878.495 10000 ;
      RECT 7828.655 1046.435 7874.575 10000 ;
      RECT 7825.015 1046.435 7827.535 10000 ;
      RECT 7821.375 1046.435 7823.895 10000 ;
      RECT 7817.735 1046.435 7820.255 10000 ;
      RECT 7814.095 1046.435 7816.615 10000 ;
      RECT 7810.455 1046.435 7812.975 10000 ;
      RECT 7751.375 1046.435 7809.335 10000 ;
      RECT 7747.455 1046.435 7750.255 10000 ;
      RECT 7743.535 1046.435 7746.335 10000 ;
      RECT 7739.615 1046.435 7742.415 10000 ;
      RECT 7735.695 1046.435 7738.495 10000 ;
      RECT 7688.655 1046.435 7734.575 10000 ;
      RECT 7685.015 1046.435 7687.535 10000 ;
      RECT 7681.375 1046.435 7683.895 10000 ;
      RECT 7677.735 1046.435 7680.255 10000 ;
      RECT 7674.095 1046.435 7676.615 10000 ;
      RECT 7670.455 1046.435 7672.975 10000 ;
      RECT 7611.375 1046.435 7669.335 10000 ;
      RECT 7607.455 1046.435 7610.255 10000 ;
      RECT 7603.535 1046.435 7606.335 10000 ;
      RECT 7599.615 1046.435 7602.415 10000 ;
      RECT 7595.695 1046.435 7598.495 10000 ;
      RECT 7548.655 1046.435 7594.575 10000 ;
      RECT 7545.015 1046.435 7547.535 10000 ;
      RECT 7541.375 1046.435 7543.895 10000 ;
      RECT 7537.735 1046.435 7540.255 10000 ;
      RECT 7534.095 1046.435 7536.615 10000 ;
      RECT 7530.455 1046.435 7532.975 10000 ;
      RECT 7471.375 1046.435 7529.335 10000 ;
      RECT 7467.455 1046.435 7470.255 10000 ;
      RECT 7463.535 1046.435 7466.335 10000 ;
      RECT 7459.615 1046.435 7462.415 10000 ;
      RECT 7455.695 1046.435 7458.495 10000 ;
      RECT 7408.655 1046.435 7454.575 10000 ;
      RECT 7405.015 1046.435 7407.535 10000 ;
      RECT 7401.375 1046.435 7403.895 10000 ;
      RECT 7397.735 1046.435 7400.255 10000 ;
      RECT 7394.095 1046.435 7396.615 10000 ;
      RECT 7390.455 1046.435 7392.975 10000 ;
      RECT 7331.375 1046.435 7389.335 10000 ;
      RECT 7327.455 1046.435 7330.255 10000 ;
      RECT 7323.535 1046.435 7326.335 10000 ;
      RECT 7319.615 1046.435 7322.415 10000 ;
      RECT 7315.695 1046.435 7318.495 10000 ;
      RECT 7268.655 1046.435 7314.575 10000 ;
      RECT 7265.015 1046.435 7267.535 10000 ;
      RECT 7261.375 1046.435 7263.895 10000 ;
      RECT 7257.735 1046.435 7260.255 10000 ;
      RECT 7254.095 1046.435 7256.615 10000 ;
      RECT 7250.455 1046.435 7252.975 10000 ;
      RECT 7191.375 1046.435 7249.335 10000 ;
      RECT 7187.455 1046.435 7190.255 10000 ;
      RECT 7183.535 1046.435 7186.335 10000 ;
      RECT 7179.615 1046.435 7182.415 10000 ;
      RECT 7175.695 1046.435 7178.495 10000 ;
      RECT 7128.655 1046.435 7174.575 10000 ;
      RECT 7125.015 1046.435 7127.535 10000 ;
      RECT 7121.375 1046.435 7123.895 10000 ;
      RECT 7117.735 1046.435 7120.255 10000 ;
      RECT 7114.095 1046.435 7116.615 10000 ;
      RECT 7110.455 1046.435 7112.975 10000 ;
      RECT 7051.375 1046.435 7109.335 10000 ;
      RECT 7047.455 1046.435 7050.255 10000 ;
      RECT 7043.535 1046.435 7046.335 10000 ;
      RECT 7039.615 1046.435 7042.415 10000 ;
      RECT 7035.695 1046.435 7038.495 10000 ;
      RECT 6988.655 1046.435 7034.575 10000 ;
      RECT 6985.015 1046.435 6987.535 10000 ;
      RECT 6981.375 1046.435 6983.895 10000 ;
      RECT 6977.735 1046.435 6980.255 10000 ;
      RECT 6974.095 1046.435 6976.615 10000 ;
      RECT 6970.455 1046.435 6972.975 10000 ;
      RECT 6911.375 1046.435 6969.335 10000 ;
      RECT 6907.455 1046.435 6910.255 10000 ;
      RECT 6903.535 1046.435 6906.335 10000 ;
      RECT 6899.615 1046.435 6902.415 10000 ;
      RECT 6895.695 1046.435 6898.495 10000 ;
      RECT 6848.655 1046.435 6894.575 10000 ;
      RECT 6845.015 1046.435 6847.535 10000 ;
      RECT 6841.375 1046.435 6843.895 10000 ;
      RECT 6837.735 1046.435 6840.255 10000 ;
      RECT 6834.095 1046.435 6836.615 10000 ;
      RECT 6830.455 1046.435 6832.975 10000 ;
      RECT 6771.375 1046.435 6829.335 10000 ;
      RECT 6767.455 1046.435 6770.255 10000 ;
      RECT 6763.535 1046.435 6766.335 10000 ;
      RECT 6759.615 1046.435 6762.415 10000 ;
      RECT 6755.695 1046.435 6758.495 10000 ;
      RECT 6708.655 1046.435 6754.575 10000 ;
      RECT 6705.015 1046.435 6707.535 10000 ;
      RECT 6701.375 1046.435 6703.895 10000 ;
      RECT 6697.735 1046.435 6700.255 10000 ;
      RECT 6694.095 1046.435 6696.615 10000 ;
      RECT 6690.455 1046.435 6692.975 10000 ;
      RECT 6631.375 1046.435 6689.335 10000 ;
      RECT 6627.455 1046.435 6630.255 10000 ;
      RECT 6623.535 1046.435 6626.335 10000 ;
      RECT 6619.615 1046.435 6622.415 10000 ;
      RECT 6615.695 1046.435 6618.495 10000 ;
      RECT 6568.655 1046.435 6614.575 10000 ;
      RECT 6565.015 1046.435 6567.535 10000 ;
      RECT 6561.375 1046.435 6563.895 10000 ;
      RECT 6557.735 1046.435 6560.255 10000 ;
      RECT 6554.095 1046.435 6556.615 10000 ;
      RECT 6550.455 1046.435 6552.975 10000 ;
      RECT 6491.375 1046.435 6549.335 10000 ;
      RECT 6487.455 1046.435 6490.255 10000 ;
      RECT 6483.535 1046.435 6486.335 10000 ;
      RECT 6479.615 1046.435 6482.415 10000 ;
      RECT 6475.695 1046.435 6478.495 10000 ;
      RECT 6428.655 1046.435 6474.575 10000 ;
      RECT 6425.015 1046.435 6427.535 10000 ;
      RECT 6421.375 1046.435 6423.895 10000 ;
      RECT 6417.735 1046.435 6420.255 10000 ;
      RECT 6414.095 1046.435 6416.615 10000 ;
      RECT 6410.455 1046.435 6412.975 10000 ;
      RECT 6351.375 1046.435 6409.335 10000 ;
      RECT 6347.455 1046.435 6350.255 10000 ;
      RECT 6343.535 1046.435 6346.335 10000 ;
      RECT 6339.615 1046.435 6342.415 10000 ;
      RECT 6335.695 1046.435 6338.495 10000 ;
      RECT 6288.655 1046.435 6334.575 10000 ;
      RECT 6285.015 1046.435 6287.535 10000 ;
      RECT 6281.375 1046.435 6283.895 10000 ;
      RECT 6277.735 1046.435 6280.255 10000 ;
      RECT 6274.095 1046.435 6276.615 10000 ;
      RECT 6270.455 1046.435 6272.975 10000 ;
      RECT 6211.375 1046.435 6269.335 10000 ;
      RECT 6207.455 1046.435 6210.255 10000 ;
      RECT 6203.535 1046.435 6206.335 10000 ;
      RECT 6199.615 1046.435 6202.415 10000 ;
      RECT 6195.695 1046.435 6198.495 10000 ;
      RECT 6148.655 1046.435 6194.575 10000 ;
      RECT 6145.015 1046.435 6147.535 10000 ;
      RECT 6141.375 1046.435 6143.895 10000 ;
      RECT 6137.735 1046.435 6140.255 10000 ;
      RECT 6134.095 1046.435 6136.615 10000 ;
      RECT 6130.455 1046.435 6132.975 10000 ;
      RECT 6071.375 1046.435 6129.335 10000 ;
      RECT 6067.455 1046.435 6070.255 10000 ;
      RECT 6063.535 1046.435 6066.335 10000 ;
      RECT 6059.615 1046.435 6062.415 10000 ;
      RECT 6055.695 1046.435 6058.495 10000 ;
      RECT 6008.655 1046.435 6054.575 10000 ;
      RECT 6005.015 1046.435 6007.535 10000 ;
      RECT 6001.375 1046.435 6003.895 10000 ;
      RECT 5997.735 1046.435 6000.255 10000 ;
      RECT 5994.095 1046.435 5996.615 10000 ;
      RECT 5990.455 1046.435 5992.975 10000 ;
      RECT 5931.375 1046.435 5989.335 10000 ;
      RECT 5927.455 1046.435 5930.255 10000 ;
      RECT 5923.535 1046.435 5926.335 10000 ;
      RECT 5919.615 1046.435 5922.415 10000 ;
      RECT 5915.695 1046.435 5918.495 10000 ;
      RECT 5868.655 1046.435 5914.575 10000 ;
      RECT 5865.015 1046.435 5867.535 10000 ;
      RECT 5861.375 1046.435 5863.895 10000 ;
      RECT 5857.735 1046.435 5860.255 10000 ;
      RECT 5854.095 1046.435 5856.615 10000 ;
      RECT 5850.455 1046.435 5852.975 10000 ;
      RECT 5791.375 1046.435 5849.335 10000 ;
      RECT 5787.455 1046.435 5790.255 10000 ;
      RECT 5783.535 1046.435 5786.335 10000 ;
      RECT 5779.615 1046.435 5782.415 10000 ;
      RECT 5775.695 1046.435 5778.495 10000 ;
      RECT 5728.655 1046.435 5774.575 10000 ;
      RECT 5725.015 1046.435 5727.535 10000 ;
      RECT 5721.375 1046.435 5723.895 10000 ;
      RECT 5717.735 1046.435 5720.255 10000 ;
      RECT 5714.095 1046.435 5716.615 10000 ;
      RECT 5710.455 1046.435 5712.975 10000 ;
      RECT 5651.375 1046.435 5709.335 10000 ;
      RECT 5647.455 1046.435 5650.255 10000 ;
      RECT 5643.535 1046.435 5646.335 10000 ;
      RECT 5639.615 1046.435 5642.415 10000 ;
      RECT 5635.695 1046.435 5638.495 10000 ;
      RECT 5588.655 1046.435 5634.575 10000 ;
      RECT 5585.015 1046.435 5587.535 10000 ;
      RECT 5581.375 1046.435 5583.895 10000 ;
      RECT 5577.735 1046.435 5580.255 10000 ;
      RECT 5574.095 1046.435 5576.615 10000 ;
      RECT 5570.455 1046.435 5572.975 10000 ;
      RECT 5511.375 1046.435 5569.335 10000 ;
      RECT 5507.455 1046.435 5510.255 10000 ;
      RECT 5503.535 1046.435 5506.335 10000 ;
      RECT 5499.615 1046.435 5502.415 10000 ;
      RECT 5495.695 1046.435 5498.495 10000 ;
      RECT 5448.655 1046.435 5494.575 10000 ;
      RECT 5445.015 1046.435 5447.535 10000 ;
      RECT 5441.375 1046.435 5443.895 10000 ;
      RECT 5437.735 1046.435 5440.255 10000 ;
      RECT 5434.095 1046.435 5436.615 10000 ;
      RECT 5430.455 1046.435 5432.975 10000 ;
      RECT 5371.375 1046.435 5429.335 10000 ;
      RECT 5367.455 1046.435 5370.255 10000 ;
      RECT 5363.535 1046.435 5366.335 10000 ;
      RECT 5359.615 1046.435 5362.415 10000 ;
      RECT 5355.695 1046.435 5358.495 10000 ;
      RECT 5308.655 1046.435 5354.575 10000 ;
      RECT 5305.015 1046.435 5307.535 10000 ;
      RECT 5301.375 1046.435 5303.895 10000 ;
      RECT 5297.735 1046.435 5300.255 10000 ;
      RECT 5294.095 1046.435 5296.615 10000 ;
      RECT 5290.455 1046.435 5292.975 10000 ;
      RECT 5231.375 1046.435 5289.335 10000 ;
      RECT 5227.455 1046.435 5230.255 10000 ;
      RECT 5223.535 1046.435 5226.335 10000 ;
      RECT 5219.615 1046.435 5222.415 10000 ;
      RECT 5215.695 1046.435 5218.495 10000 ;
      RECT 5168.655 1046.435 5214.575 10000 ;
      RECT 5165.015 1046.435 5167.535 10000 ;
      RECT 5161.375 1046.435 5163.895 10000 ;
      RECT 5157.735 1046.435 5160.255 10000 ;
      RECT 5154.095 1046.435 5156.615 10000 ;
      RECT 5150.455 1046.435 5152.975 10000 ;
      RECT 5091.375 1046.435 5149.335 10000 ;
      RECT 5087.455 1046.435 5090.255 10000 ;
      RECT 5083.535 1046.435 5086.335 10000 ;
      RECT 5079.615 1046.435 5082.415 10000 ;
      RECT 5075.695 1046.435 5078.495 10000 ;
      RECT 5028.655 1046.435 5074.575 10000 ;
      RECT 5025.015 1046.435 5027.535 10000 ;
      RECT 5021.375 1046.435 5023.895 10000 ;
      RECT 5017.735 1046.435 5020.255 10000 ;
      RECT 5014.095 1046.435 5016.615 10000 ;
      RECT 5010.455 1046.435 5012.975 10000 ;
      RECT 4951.375 1046.435 5009.335 10000 ;
      RECT 4947.455 1046.435 4950.255 10000 ;
      RECT 4943.535 1046.435 4946.335 10000 ;
      RECT 4939.615 1046.435 4942.415 10000 ;
      RECT 4935.695 1046.435 4938.495 10000 ;
      RECT 4888.655 1046.435 4934.575 10000 ;
      RECT 4885.015 1046.435 4887.535 10000 ;
      RECT 4881.375 1046.435 4883.895 10000 ;
      RECT 4877.735 1046.435 4880.255 10000 ;
      RECT 4874.095 1046.435 4876.615 10000 ;
      RECT 4870.455 1046.435 4872.975 10000 ;
      RECT 4811.375 1046.435 4869.335 10000 ;
      RECT 4807.455 1046.435 4810.255 10000 ;
      RECT 4803.535 1046.435 4806.335 10000 ;
      RECT 4799.615 1046.435 4802.415 10000 ;
      RECT 4795.695 1046.435 4798.495 10000 ;
      RECT 4748.655 1046.435 4794.575 10000 ;
      RECT 4745.015 1046.435 4747.535 10000 ;
      RECT 4741.375 1046.435 4743.895 10000 ;
      RECT 4737.735 1046.435 4740.255 10000 ;
      RECT 4734.095 1046.435 4736.615 10000 ;
      RECT 4730.455 1046.435 4732.975 10000 ;
      RECT 4671.375 1046.435 4729.335 10000 ;
      RECT 4667.455 1046.435 4670.255 10000 ;
      RECT 4663.535 1046.435 4666.335 10000 ;
      RECT 4659.615 1046.435 4662.415 10000 ;
      RECT 4655.695 1046.435 4658.495 10000 ;
      RECT 4608.655 1046.435 4654.575 10000 ;
      RECT 4605.015 1046.435 4607.535 10000 ;
      RECT 4601.375 1046.435 4603.895 10000 ;
      RECT 4597.735 1046.435 4600.255 10000 ;
      RECT 4594.095 1046.435 4596.615 10000 ;
      RECT 4590.455 1046.435 4592.975 10000 ;
      RECT 4531.375 1046.435 4589.335 10000 ;
      RECT 4527.455 1046.435 4530.255 10000 ;
      RECT 4523.535 1046.435 4526.335 10000 ;
      RECT 4519.615 1046.435 4522.415 10000 ;
      RECT 4515.695 1046.435 4518.495 10000 ;
      RECT 4468.655 1046.435 4514.575 10000 ;
      RECT 4465.015 1046.435 4467.535 10000 ;
      RECT 4461.375 1046.435 4463.895 10000 ;
      RECT 4457.735 1046.435 4460.255 10000 ;
      RECT 4454.095 1046.435 4456.615 10000 ;
      RECT 4450.455 1046.435 4452.975 10000 ;
      RECT 4391.375 1046.435 4449.335 10000 ;
      RECT 4387.455 1046.435 4390.255 10000 ;
      RECT 4383.535 1046.435 4386.335 10000 ;
      RECT 4379.615 1046.435 4382.415 10000 ;
      RECT 4375.695 1046.435 4378.495 10000 ;
      RECT 4328.655 1046.435 4374.575 10000 ;
      RECT 4325.015 1046.435 4327.535 10000 ;
      RECT 4321.375 1046.435 4323.895 10000 ;
      RECT 4317.735 1046.435 4320.255 10000 ;
      RECT 4314.095 1046.435 4316.615 10000 ;
      RECT 4310.455 1046.435 4312.975 10000 ;
      RECT 4251.375 1046.435 4309.335 10000 ;
      RECT 4247.455 1046.435 4250.255 10000 ;
      RECT 4243.535 1046.435 4246.335 10000 ;
      RECT 4239.615 1046.435 4242.415 10000 ;
      RECT 4235.695 1046.435 4238.495 10000 ;
      RECT 4188.655 1046.435 4234.575 10000 ;
      RECT 4185.015 1046.435 4187.535 10000 ;
      RECT 4181.375 1046.435 4183.895 10000 ;
      RECT 4177.735 1046.435 4180.255 10000 ;
      RECT 4174.095 1046.435 4176.615 10000 ;
      RECT 4170.455 1046.435 4172.975 10000 ;
      RECT 4111.375 1046.435 4169.335 10000 ;
      RECT 4107.455 1046.435 4110.255 10000 ;
      RECT 4103.535 1046.435 4106.335 10000 ;
      RECT 4099.615 1046.435 4102.415 10000 ;
      RECT 4095.695 1046.435 4098.495 10000 ;
      RECT 4048.655 1046.435 4094.575 10000 ;
      RECT 4045.015 1046.435 4047.535 10000 ;
      RECT 4041.375 1046.435 4043.895 10000 ;
      RECT 4037.735 1046.435 4040.255 10000 ;
      RECT 4034.095 1046.435 4036.615 10000 ;
      RECT 4030.455 1046.435 4032.975 10000 ;
      RECT 3971.375 1046.435 4029.335 10000 ;
      RECT 3967.455 1046.435 3970.255 10000 ;
      RECT 3963.535 1046.435 3966.335 10000 ;
      RECT 3959.615 1046.435 3962.415 10000 ;
      RECT 3955.695 1046.435 3958.495 10000 ;
      RECT 3908.655 1046.435 3954.575 10000 ;
      RECT 3905.015 1046.435 3907.535 10000 ;
      RECT 3901.375 1046.435 3903.895 10000 ;
      RECT 3897.735 1046.435 3900.255 10000 ;
      RECT 3894.095 1046.435 3896.615 10000 ;
      RECT 3890.455 1046.435 3892.975 10000 ;
      RECT 3831.375 1046.435 3889.335 10000 ;
      RECT 3827.455 1046.435 3830.255 10000 ;
      RECT 3823.535 1046.435 3826.335 10000 ;
      RECT 3819.615 1046.435 3822.415 10000 ;
      RECT 3815.695 1046.435 3818.495 10000 ;
      RECT 3768.655 1046.435 3814.575 10000 ;
      RECT 3765.015 1046.435 3767.535 10000 ;
      RECT 3761.375 1046.435 3763.895 10000 ;
      RECT 3757.735 1046.435 3760.255 10000 ;
      RECT 3754.095 1046.435 3756.615 10000 ;
      RECT 3750.455 1046.435 3752.975 10000 ;
      RECT 3691.375 1046.435 3749.335 10000 ;
      RECT 3687.455 1046.435 3690.255 10000 ;
      RECT 3683.535 1046.435 3686.335 10000 ;
      RECT 3679.615 1046.435 3682.415 10000 ;
      RECT 3675.695 1046.435 3678.495 10000 ;
      RECT 3628.655 1046.435 3674.575 10000 ;
      RECT 3625.015 1046.435 3627.535 10000 ;
      RECT 3621.375 1046.435 3623.895 10000 ;
      RECT 3617.735 1046.435 3620.255 10000 ;
      RECT 3614.095 1046.435 3616.615 10000 ;
      RECT 3610.455 1046.435 3612.975 10000 ;
      RECT 3551.375 1046.435 3609.335 10000 ;
      RECT 3547.455 1046.435 3550.255 10000 ;
      RECT 3543.535 1046.435 3546.335 10000 ;
      RECT 3539.615 1046.435 3542.415 10000 ;
      RECT 3535.695 1046.435 3538.495 10000 ;
      RECT 3488.655 1046.435 3534.575 10000 ;
      RECT 3485.015 1046.435 3487.535 10000 ;
      RECT 3481.375 1046.435 3483.895 10000 ;
      RECT 3477.735 1046.435 3480.255 10000 ;
      RECT 3474.095 1046.435 3476.615 10000 ;
      RECT 3470.455 1046.435 3472.975 10000 ;
      RECT 3411.375 1046.435 3469.335 10000 ;
      RECT 3407.455 1046.435 3410.255 10000 ;
      RECT 3403.535 1046.435 3406.335 10000 ;
      RECT 3399.615 1046.435 3402.415 10000 ;
      RECT 3395.695 1046.435 3398.495 10000 ;
      RECT 3348.655 1046.435 3394.575 10000 ;
      RECT 3345.015 1046.435 3347.535 10000 ;
      RECT 3341.375 1046.435 3343.895 10000 ;
      RECT 3337.735 1046.435 3340.255 10000 ;
      RECT 3334.095 1046.435 3336.615 10000 ;
      RECT 3330.455 1046.435 3332.975 10000 ;
      RECT 3271.375 1046.435 3329.335 10000 ;
      RECT 3267.455 1046.435 3270.255 10000 ;
      RECT 3263.535 1046.435 3266.335 10000 ;
      RECT 3259.615 1046.435 3262.415 10000 ;
      RECT 3255.695 1046.435 3258.495 10000 ;
      RECT 3208.655 1046.435 3254.575 10000 ;
      RECT 3205.015 1046.435 3207.535 10000 ;
      RECT 3201.375 1046.435 3203.895 10000 ;
      RECT 3197.735 1046.435 3200.255 10000 ;
      RECT 3194.095 1046.435 3196.615 10000 ;
      RECT 3190.455 1046.435 3192.975 10000 ;
      RECT 3131.375 1046.435 3189.335 10000 ;
      RECT 3127.455 1046.435 3130.255 10000 ;
      RECT 3123.535 1046.435 3126.335 10000 ;
      RECT 3119.615 1046.435 3122.415 10000 ;
      RECT 3115.695 1046.435 3118.495 10000 ;
      RECT 3068.655 1046.435 3114.575 10000 ;
      RECT 3065.015 1046.435 3067.535 10000 ;
      RECT 3061.375 1046.435 3063.895 10000 ;
      RECT 3057.735 1046.435 3060.255 10000 ;
      RECT 3054.095 1046.435 3056.615 10000 ;
      RECT 3050.455 1046.435 3052.975 10000 ;
      RECT 2991.375 1046.435 3049.335 10000 ;
      RECT 2987.455 1046.435 2990.255 10000 ;
      RECT 2983.535 1046.435 2986.335 10000 ;
      RECT 2979.615 1046.435 2982.415 10000 ;
      RECT 2975.695 1046.435 2978.495 10000 ;
      RECT 2928.655 1046.435 2974.575 10000 ;
      RECT 2925.015 1046.435 2927.535 10000 ;
      RECT 2921.375 1046.435 2923.895 10000 ;
      RECT 2917.735 1046.435 2920.255 10000 ;
      RECT 2914.095 1046.435 2916.615 10000 ;
      RECT 2910.455 1046.435 2912.975 10000 ;
      RECT 2851.375 1046.435 2909.335 10000 ;
      RECT 2847.455 1046.435 2850.255 10000 ;
      RECT 2843.535 1046.435 2846.335 10000 ;
      RECT 2839.615 1046.435 2842.415 10000 ;
      RECT 2835.695 1046.435 2838.495 10000 ;
      RECT 2788.655 1046.435 2834.575 10000 ;
      RECT 2785.015 1046.435 2787.535 10000 ;
      RECT 2781.375 1046.435 2783.895 10000 ;
      RECT 2777.735 1046.435 2780.255 10000 ;
      RECT 2774.095 1046.435 2776.615 10000 ;
      RECT 2770.455 1046.435 2772.975 10000 ;
      RECT 2711.375 1046.435 2769.335 10000 ;
      RECT 2707.455 1046.435 2710.255 10000 ;
      RECT 2703.535 1046.435 2706.335 10000 ;
      RECT 2699.615 1046.435 2702.415 10000 ;
      RECT 2695.695 1046.435 2698.495 10000 ;
      RECT 2648.655 1046.435 2694.575 10000 ;
      RECT 2645.015 1046.435 2647.535 10000 ;
      RECT 2641.375 1046.435 2643.895 10000 ;
      RECT 2637.735 1046.435 2640.255 10000 ;
      RECT 2634.095 1046.435 2636.615 10000 ;
      RECT 2630.455 1046.435 2632.975 10000 ;
      RECT 2571.375 1046.435 2629.335 10000 ;
      RECT 2567.455 1046.435 2570.255 10000 ;
      RECT 2563.535 1046.435 2566.335 10000 ;
      RECT 2559.615 1046.435 2562.415 10000 ;
      RECT 2555.695 1046.435 2558.495 10000 ;
      RECT 2508.655 1046.435 2554.575 10000 ;
      RECT 2505.015 1046.435 2507.535 10000 ;
      RECT 2501.375 1046.435 2503.895 10000 ;
      RECT 2497.735 1046.435 2500.255 10000 ;
      RECT 2494.095 1046.435 2496.615 10000 ;
      RECT 2490.455 1046.435 2492.975 10000 ;
      RECT 2431.375 1046.435 2489.335 10000 ;
      RECT 2427.455 1046.435 2430.255 10000 ;
      RECT 2423.535 1046.435 2426.335 10000 ;
      RECT 2419.615 1046.435 2422.415 10000 ;
      RECT 2415.695 1046.435 2418.495 10000 ;
      RECT 2368.655 1046.435 2414.575 10000 ;
      RECT 2365.015 1046.435 2367.535 10000 ;
      RECT 2361.375 1046.435 2363.895 10000 ;
      RECT 2357.735 1046.435 2360.255 10000 ;
      RECT 2354.095 1046.435 2356.615 10000 ;
      RECT 2350.455 1046.435 2352.975 10000 ;
      RECT 2291.375 1046.435 2349.335 10000 ;
      RECT 2287.455 1046.435 2290.255 10000 ;
      RECT 2283.535 1046.435 2286.335 10000 ;
      RECT 2279.615 1046.435 2282.415 10000 ;
      RECT 2275.695 1046.435 2278.495 10000 ;
      RECT 2228.655 1046.435 2274.575 10000 ;
      RECT 2225.015 1046.435 2227.535 10000 ;
      RECT 2221.375 1046.435 2223.895 10000 ;
      RECT 2217.735 1046.435 2220.255 10000 ;
      RECT 2214.095 1046.435 2216.615 10000 ;
      RECT 2210.455 1046.435 2212.975 10000 ;
      RECT 2151.375 1046.435 2209.335 10000 ;
      RECT 2147.455 1046.435 2150.255 10000 ;
      RECT 2143.535 1046.435 2146.335 10000 ;
      RECT 2139.615 1046.435 2142.415 10000 ;
      RECT 2135.695 1046.435 2138.495 10000 ;
      RECT 2088.655 1046.435 2134.575 10000 ;
      RECT 2085.015 1046.435 2087.535 10000 ;
      RECT 2081.375 1046.435 2083.895 10000 ;
      RECT 2077.735 1046.435 2080.255 10000 ;
      RECT 2074.095 1046.435 2076.615 10000 ;
      RECT 2070.455 1046.435 2072.975 10000 ;
      RECT 2011.375 1046.435 2069.335 10000 ;
      RECT 2007.455 1046.435 2010.255 10000 ;
      RECT 2003.535 1046.435 2006.335 10000 ;
      RECT 1999.615 1046.435 2002.415 10000 ;
      RECT 1995.695 1046.435 1998.495 10000 ;
      RECT 1948.655 1046.435 1994.575 10000 ;
      RECT 1945.015 1046.435 1947.535 10000 ;
      RECT 1941.375 1046.435 1943.895 10000 ;
      RECT 1937.735 1046.435 1940.255 10000 ;
      RECT 1934.095 1046.435 1936.615 10000 ;
      RECT 1930.455 1046.435 1932.975 10000 ;
      RECT 1871.375 1046.435 1929.335 10000 ;
      RECT 1867.455 1046.435 1870.255 10000 ;
      RECT 1863.535 1046.435 1866.335 10000 ;
      RECT 1859.615 1046.435 1862.415 10000 ;
      RECT 1855.695 1046.435 1858.495 10000 ;
      RECT 1808.655 1046.435 1854.575 10000 ;
      RECT 1805.015 1046.435 1807.535 10000 ;
      RECT 1801.375 1046.435 1803.895 10000 ;
      RECT 1797.735 1046.435 1800.255 10000 ;
      RECT 1794.095 1046.435 1796.615 10000 ;
      RECT 1790.455 1046.435 1792.975 10000 ;
      RECT 1731.375 1046.435 1789.335 10000 ;
      RECT 1727.455 1046.435 1730.255 10000 ;
      RECT 1723.535 1046.435 1726.335 10000 ;
      RECT 1719.615 1046.435 1722.415 10000 ;
      RECT 1715.695 1046.435 1718.495 10000 ;
      RECT 1668.655 1046.435 1714.575 10000 ;
      RECT 1665.015 1046.435 1667.535 10000 ;
      RECT 1661.375 1046.435 1663.895 10000 ;
      RECT 1657.735 1046.435 1660.255 10000 ;
      RECT 1654.095 1046.435 1656.615 10000 ;
      RECT 1650.455 1046.435 1652.975 10000 ;
      RECT 1591.375 1046.435 1649.335 10000 ;
      RECT 1587.455 1046.435 1590.255 10000 ;
      RECT 1583.535 1046.435 1586.335 10000 ;
      RECT 1579.615 1046.435 1582.415 10000 ;
      RECT 1575.695 1046.435 1578.495 10000 ;
      RECT 1528.655 1046.435 1574.575 10000 ;
      RECT 1525.015 1046.435 1527.535 10000 ;
      RECT 1521.375 1046.435 1523.895 10000 ;
      RECT 1517.735 1046.435 1520.255 10000 ;
      RECT 1514.095 1046.435 1516.615 10000 ;
      RECT 1510.455 1046.435 1512.975 10000 ;
      RECT 1451.375 1046.435 1509.335 10000 ;
      RECT 1447.455 1046.435 1450.255 10000 ;
      RECT 1443.535 1046.435 1446.335 10000 ;
      RECT 1439.615 1046.435 1442.415 10000 ;
      RECT 1435.695 1046.435 1438.495 10000 ;
      RECT 1388.655 1046.435 1434.575 10000 ;
      RECT 1385.015 1046.435 1387.535 10000 ;
      RECT 1381.375 1046.435 1383.895 10000 ;
      RECT 1377.735 1046.435 1380.255 10000 ;
      RECT 1374.095 1046.435 1376.615 10000 ;
      RECT 1370.455 1046.435 1372.975 10000 ;
      RECT 1311.375 1046.435 1369.335 10000 ;
      RECT 1307.455 1046.435 1310.255 10000 ;
      RECT 1303.535 1046.435 1306.335 10000 ;
      RECT 1299.615 1046.435 1302.415 10000 ;
      RECT 1295.695 1046.435 1298.495 10000 ;
      RECT 1248.655 1046.435 1294.575 10000 ;
      RECT 1245.015 1046.435 1247.535 10000 ;
      RECT 1241.375 1046.435 1243.895 10000 ;
      RECT 1237.735 1046.435 1240.255 10000 ;
      RECT 1234.095 1046.435 1236.615 10000 ;
      RECT 1230.455 1046.435 1232.975 10000 ;
      RECT 1171.375 1046.435 1229.335 10000 ;
      RECT 1167.455 1046.435 1170.255 10000 ;
      RECT 1163.535 1046.435 1166.335 10000 ;
      RECT 1159.615 1046.435 1162.415 10000 ;
      RECT 1155.695 1046.435 1158.495 10000 ;
      RECT 1008.465 1046.435 1154.575 10000 ;
      RECT 998.1 1046.435 1003.425 10000 ;
      RECT 10102.375 1046.435 10102.655 10000 ;
    LAYER M3 ;
      RECT 0.5 9996.5 20199.5 9999.5 ;
      RECT 20196.5 0.5 20199.5 9999.5 ;
      RECT 0.5 0.5 3.5 9999.5 ;
      RECT 0.5 0.5 20199.5 3.5 ;
      RECT 4.1 9990 20195.9 9995.9 ;
      RECT 20190 4.1 20195.9 9995.9 ;
      RECT 4.1 4.1 10 9995.9 ;
      RECT 4.1 4.1 20195.9 10 ;
      RECT 19150 9497.56 19170 9527.56 ;
      RECT 19150 9529.56 19170 9559.56 ;
      RECT 19150 9617.56 19170 9647.56 ;
      RECT 19150 9649.56 19170 9679.56 ;
      RECT 19150 9737.56 19170 9767.56 ;
      RECT 19150 9769.56 19170 9799.56 ;
      RECT 19150 9857.56 19170 9887.56 ;
      RECT 19150 9889.56 19170 9919.56 ;
      RECT 19158.16 1119.19 19167.9 1119.99 ;
      RECT 19158.16 1121.59 19167.9 1122.39 ;
      RECT 19158.16 1123.99 19167.9 1124.79 ;
      RECT 19158.16 1126.39 19167.9 1127.19 ;
      RECT 19158.16 1364.42 19167.75 1365.49 ;
      RECT 19158.16 1367.4 19167.75 1368.47 ;
      RECT 19146.82 9258.62 19161.76 9259.94 ;
      RECT 19146.82 9297.14 19161.76 9298.46 ;
      RECT 19146.82 9330.63 19161.76 9331.95 ;
      RECT 19146.82 9369.135 19161.76 9370.455 ;
      RECT 19146.82 9402.63 19161.76 9403.95 ;
      RECT 19146.82 9441.145 19161.76 9442.465 ;
      RECT 19014.355 1046.935 19039.355 1189.16 ;
      RECT 18988.355 1046.935 19012.355 1189.16 ;
      RECT 18937.745 1046.935 18961.745 1118.84 ;
      RECT 18924.745 1046.935 18935.745 1118.84 ;
      RECT 18874.355 1046.935 18899.355 1189.16 ;
      RECT 18848.355 1046.935 18872.355 1189.16 ;
      RECT 18797.745 1046.935 18821.745 1118.84 ;
      RECT 18784.745 1046.935 18795.745 1118.84 ;
      RECT 18734.355 1046.935 18759.355 1189.16 ;
      RECT 18708.355 1046.935 18732.355 1189.16 ;
      RECT 18657.745 1046.935 18681.745 1118.84 ;
      RECT 18644.745 1046.935 18655.745 1118.84 ;
      RECT 18594.355 1046.935 18619.355 1189.16 ;
      RECT 18568.355 1046.935 18592.355 1189.16 ;
      RECT 18517.745 1046.935 18541.745 1118.84 ;
      RECT 18504.745 1046.935 18515.745 1118.84 ;
      RECT 18454.355 1046.935 18479.355 1189.16 ;
      RECT 18428.355 1046.935 18452.355 1189.16 ;
      RECT 18377.745 1046.935 18401.745 1118.84 ;
      RECT 18364.745 1046.935 18375.745 1118.84 ;
      RECT 18314.355 1046.935 18339.355 1189.16 ;
      RECT 18288.355 1046.935 18312.355 1189.16 ;
      RECT 18237.745 1046.935 18261.745 1118.84 ;
      RECT 18224.745 1046.935 18235.745 1118.84 ;
      RECT 18174.355 1046.935 18199.355 1189.16 ;
      RECT 18148.355 1046.935 18172.355 1189.16 ;
      RECT 18097.745 1046.935 18121.745 1118.84 ;
      RECT 18084.745 1046.935 18095.745 1118.84 ;
      RECT 18034.355 1046.935 18059.355 1189.16 ;
      RECT 18008.355 1046.935 18032.355 1189.16 ;
      RECT 17957.745 1046.935 17981.745 1118.84 ;
      RECT 17944.745 1046.935 17955.745 1118.84 ;
      RECT 17894.355 1046.935 17919.355 1189.16 ;
      RECT 17868.355 1046.935 17892.355 1189.16 ;
      RECT 17817.745 1046.935 17841.745 1118.84 ;
      RECT 17804.745 1046.935 17815.745 1118.84 ;
      RECT 17754.355 1046.935 17779.355 1189.16 ;
      RECT 17728.355 1046.935 17752.355 1189.16 ;
      RECT 17677.745 1046.935 17701.745 1118.84 ;
      RECT 17664.745 1046.935 17675.745 1118.84 ;
      RECT 17614.355 1046.935 17639.355 1189.16 ;
      RECT 17588.355 1046.935 17612.355 1189.16 ;
      RECT 17537.745 1046.935 17561.745 1118.84 ;
      RECT 17524.745 1046.935 17535.745 1118.84 ;
      RECT 17474.355 1046.935 17499.355 1189.16 ;
      RECT 17448.355 1046.935 17472.355 1189.16 ;
      RECT 17397.745 1046.935 17421.745 1118.84 ;
      RECT 17384.745 1046.935 17395.745 1118.84 ;
      RECT 17334.355 1046.935 17359.355 1189.16 ;
      RECT 17308.355 1046.935 17332.355 1189.16 ;
      RECT 17257.745 1046.935 17281.745 1118.84 ;
      RECT 17244.745 1046.935 17255.745 1118.84 ;
      RECT 17194.355 1046.935 17219.355 1189.16 ;
      RECT 17168.355 1046.935 17192.355 1189.16 ;
      RECT 17117.745 1046.935 17141.745 1118.84 ;
      RECT 17104.745 1046.935 17115.745 1118.84 ;
      RECT 17054.355 1046.935 17079.355 1189.16 ;
      RECT 17028.355 1046.935 17052.355 1189.16 ;
      RECT 16977.745 1046.935 17001.745 1118.84 ;
      RECT 16964.745 1046.935 16975.745 1118.84 ;
      RECT 16914.355 1046.935 16939.355 1189.16 ;
      RECT 16888.355 1046.935 16912.355 1189.16 ;
      RECT 16837.745 1046.935 16861.745 1118.84 ;
      RECT 16824.745 1046.935 16835.745 1118.84 ;
      RECT 16774.355 1046.935 16799.355 1189.16 ;
      RECT 16748.355 1046.935 16772.355 1189.16 ;
      RECT 16697.745 1046.935 16721.745 1118.84 ;
      RECT 16684.745 1046.935 16695.745 1118.84 ;
      RECT 16634.355 1046.935 16659.355 1189.16 ;
      RECT 16608.355 1046.935 16632.355 1189.16 ;
      RECT 16557.745 1046.935 16581.745 1118.84 ;
      RECT 16544.745 1046.935 16555.745 1118.84 ;
      RECT 16494.355 1046.935 16519.355 1189.16 ;
      RECT 16468.355 1046.935 16492.355 1189.16 ;
      RECT 16417.745 1046.935 16441.745 1118.84 ;
      RECT 16404.745 1046.935 16415.745 1118.84 ;
      RECT 16354.355 1046.935 16379.355 1189.16 ;
      RECT 16328.355 1046.935 16352.355 1189.16 ;
      RECT 16277.745 1046.935 16301.745 1118.84 ;
      RECT 16264.745 1046.935 16275.745 1118.84 ;
      RECT 16214.355 1046.935 16239.355 1189.16 ;
      RECT 16188.355 1046.935 16212.355 1189.16 ;
      RECT 16137.745 1046.935 16161.745 1118.84 ;
      RECT 16124.745 1046.935 16135.745 1118.84 ;
      RECT 16074.355 1046.935 16099.355 1189.16 ;
      RECT 16048.355 1046.935 16072.355 1189.16 ;
      RECT 15997.745 1046.935 16021.745 1118.84 ;
      RECT 15984.745 1046.935 15995.745 1118.84 ;
      RECT 15934.355 1046.935 15959.355 1189.16 ;
      RECT 15908.355 1046.935 15932.355 1189.16 ;
      RECT 15857.745 1046.935 15881.745 1118.84 ;
      RECT 15844.745 1046.935 15855.745 1118.84 ;
      RECT 15794.355 1046.935 15819.355 1189.16 ;
      RECT 15768.355 1046.935 15792.355 1189.16 ;
      RECT 15717.745 1046.935 15741.745 1118.84 ;
      RECT 15704.745 1046.935 15715.745 1118.84 ;
      RECT 15654.355 1046.935 15679.355 1189.16 ;
      RECT 15628.355 1046.935 15652.355 1189.16 ;
      RECT 15577.745 1046.935 15601.745 1118.84 ;
      RECT 15564.745 1046.935 15575.745 1118.84 ;
      RECT 15514.355 1046.935 15539.355 1189.16 ;
      RECT 15488.355 1046.935 15512.355 1189.16 ;
      RECT 15437.745 1046.935 15461.745 1118.84 ;
      RECT 15424.745 1046.935 15435.745 1118.84 ;
      RECT 15374.355 1046.935 15399.355 1189.16 ;
      RECT 15348.355 1046.935 15372.355 1189.16 ;
      RECT 15297.745 1046.935 15321.745 1118.84 ;
      RECT 15284.745 1046.935 15295.745 1118.84 ;
      RECT 15234.355 1046.935 15259.355 1189.16 ;
      RECT 15208.355 1046.935 15232.355 1189.16 ;
      RECT 15157.745 1046.935 15181.745 1118.84 ;
      RECT 15144.745 1046.935 15155.745 1118.84 ;
      RECT 15094.355 1046.935 15119.355 1189.16 ;
      RECT 15068.355 1046.935 15092.355 1189.16 ;
      RECT 15017.745 1046.935 15041.745 1118.84 ;
      RECT 15004.745 1046.935 15015.745 1118.84 ;
      RECT 14954.355 1046.935 14979.355 1189.16 ;
      RECT 14928.355 1046.935 14952.355 1189.16 ;
      RECT 14877.745 1046.935 14901.745 1118.84 ;
      RECT 14864.745 1046.935 14875.745 1118.84 ;
      RECT 14814.355 1046.935 14839.355 1189.16 ;
      RECT 14788.355 1046.935 14812.355 1189.16 ;
      RECT 14737.745 1046.935 14761.745 1118.84 ;
      RECT 14724.745 1046.935 14735.745 1118.84 ;
      RECT 14674.355 1046.935 14699.355 1189.16 ;
      RECT 14648.355 1046.935 14672.355 1189.16 ;
      RECT 14597.745 1046.935 14621.745 1118.84 ;
      RECT 14584.745 1046.935 14595.745 1118.84 ;
      RECT 14534.355 1046.935 14559.355 1189.16 ;
      RECT 14508.355 1046.935 14532.355 1189.16 ;
      RECT 14457.745 1046.935 14481.745 1118.84 ;
      RECT 14444.745 1046.935 14455.745 1118.84 ;
      RECT 14394.355 1046.935 14419.355 1189.16 ;
      RECT 14368.355 1046.935 14392.355 1189.16 ;
      RECT 14317.745 1046.935 14341.745 1118.84 ;
      RECT 14304.745 1046.935 14315.745 1118.84 ;
      RECT 14254.355 1046.935 14279.355 1189.16 ;
      RECT 14228.355 1046.935 14252.355 1189.16 ;
      RECT 14177.745 1046.935 14201.745 1118.84 ;
      RECT 14164.745 1046.935 14175.745 1118.84 ;
      RECT 14114.355 1046.935 14139.355 1189.16 ;
      RECT 14088.355 1046.935 14112.355 1189.16 ;
      RECT 14037.745 1046.935 14061.745 1118.84 ;
      RECT 14024.745 1046.935 14035.745 1118.84 ;
      RECT 13974.355 1046.935 13999.355 1189.16 ;
      RECT 13948.355 1046.935 13972.355 1189.16 ;
      RECT 13897.745 1046.935 13921.745 1118.84 ;
      RECT 13884.745 1046.935 13895.745 1118.84 ;
      RECT 13834.355 1046.935 13859.355 1189.16 ;
      RECT 13808.355 1046.935 13832.355 1189.16 ;
      RECT 13757.745 1046.935 13781.745 1118.84 ;
      RECT 13744.745 1046.935 13755.745 1118.84 ;
      RECT 13694.355 1046.935 13719.355 1189.16 ;
      RECT 13668.355 1046.935 13692.355 1189.16 ;
      RECT 13617.745 1046.935 13641.745 1118.84 ;
      RECT 13604.745 1046.935 13615.745 1118.84 ;
      RECT 13554.355 1046.935 13579.355 1189.16 ;
      RECT 13528.355 1046.935 13552.355 1189.16 ;
      RECT 13477.745 1046.935 13501.745 1118.84 ;
      RECT 13464.745 1046.935 13475.745 1118.84 ;
      RECT 13414.355 1046.935 13439.355 1189.16 ;
      RECT 13388.355 1046.935 13412.355 1189.16 ;
      RECT 13337.745 1046.935 13361.745 1118.84 ;
      RECT 13324.745 1046.935 13335.745 1118.84 ;
      RECT 13274.355 1046.935 13299.355 1189.16 ;
      RECT 13248.355 1046.935 13272.355 1189.16 ;
      RECT 13197.745 1046.935 13221.745 1118.84 ;
      RECT 13184.745 1046.935 13195.745 1118.84 ;
      RECT 13134.355 1046.935 13159.355 1189.16 ;
      RECT 13108.355 1046.935 13132.355 1189.16 ;
      RECT 13057.745 1046.935 13081.745 1118.84 ;
      RECT 13044.745 1046.935 13055.745 1118.84 ;
      RECT 12994.355 1046.935 13019.355 1189.16 ;
      RECT 12968.355 1046.935 12992.355 1189.16 ;
      RECT 12917.745 1046.935 12941.745 1118.84 ;
      RECT 12904.745 1046.935 12915.745 1118.84 ;
      RECT 12854.355 1046.935 12879.355 1189.16 ;
      RECT 12828.355 1046.935 12852.355 1189.16 ;
      RECT 12777.745 1046.935 12801.745 1118.84 ;
      RECT 12764.745 1046.935 12775.745 1118.84 ;
      RECT 12714.355 1046.935 12739.355 1189.16 ;
      RECT 12688.355 1046.935 12712.355 1189.16 ;
      RECT 12637.745 1046.935 12661.745 1118.84 ;
      RECT 12624.745 1046.935 12635.745 1118.84 ;
      RECT 12574.355 1046.935 12599.355 1189.16 ;
      RECT 12548.355 1046.935 12572.355 1189.16 ;
      RECT 12497.745 1046.935 12521.745 1118.84 ;
      RECT 12484.745 1046.935 12495.745 1118.84 ;
      RECT 12434.355 1046.935 12459.355 1189.16 ;
      RECT 12408.355 1046.935 12432.355 1189.16 ;
      RECT 12357.745 1046.935 12381.745 1118.84 ;
      RECT 12344.745 1046.935 12355.745 1118.84 ;
      RECT 12294.355 1046.935 12319.355 1189.16 ;
      RECT 12268.355 1046.935 12292.355 1189.16 ;
      RECT 12217.745 1046.935 12241.745 1118.84 ;
      RECT 12204.745 1046.935 12215.745 1118.84 ;
      RECT 12154.355 1046.935 12179.355 1189.16 ;
      RECT 12128.355 1046.935 12152.355 1189.16 ;
      RECT 12077.745 1046.935 12101.745 1118.84 ;
      RECT 12064.745 1046.935 12075.745 1118.84 ;
      RECT 12014.355 1046.935 12039.355 1189.16 ;
      RECT 11988.355 1046.935 12012.355 1189.16 ;
      RECT 11937.745 1046.935 11961.745 1118.84 ;
      RECT 11924.745 1046.935 11935.745 1118.84 ;
      RECT 11874.355 1046.935 11899.355 1189.16 ;
      RECT 11848.355 1046.935 11872.355 1189.16 ;
      RECT 11797.745 1046.935 11821.745 1118.84 ;
      RECT 11784.745 1046.935 11795.745 1118.84 ;
      RECT 11734.355 1046.935 11759.355 1189.16 ;
      RECT 11708.355 1046.935 11732.355 1189.16 ;
      RECT 11657.745 1046.935 11681.745 1118.84 ;
      RECT 11644.745 1046.935 11655.745 1118.84 ;
      RECT 11594.355 1046.935 11619.355 1189.16 ;
      RECT 11568.355 1046.935 11592.355 1189.16 ;
      RECT 11517.745 1046.935 11541.745 1118.84 ;
      RECT 11504.745 1046.935 11515.745 1118.84 ;
      RECT 11454.355 1046.935 11479.355 1189.16 ;
      RECT 11428.355 1046.935 11452.355 1189.16 ;
      RECT 11377.745 1046.935 11401.745 1118.84 ;
      RECT 11364.745 1046.935 11375.745 1118.84 ;
      RECT 11314.355 1046.935 11339.355 1189.16 ;
      RECT 11288.355 1046.935 11312.355 1189.16 ;
      RECT 11237.745 1046.935 11261.745 1118.84 ;
      RECT 11224.745 1046.935 11235.745 1118.84 ;
      RECT 11174.355 1046.935 11199.355 1189.16 ;
      RECT 11148.355 1046.935 11172.355 1189.16 ;
      RECT 11097.745 1046.935 11121.745 1118.84 ;
      RECT 11084.745 1046.935 11095.745 1118.84 ;
      RECT 11034.355 1046.935 11059.355 1189.16 ;
      RECT 11008.355 1046.935 11032.355 1189.16 ;
      RECT 10957.745 1046.935 10981.745 1118.84 ;
      RECT 10944.745 1046.935 10955.745 1118.84 ;
      RECT 10894.355 1046.935 10919.355 1189.16 ;
      RECT 10868.355 1046.935 10892.355 1189.16 ;
      RECT 10817.745 1046.935 10841.745 1118.84 ;
      RECT 10804.745 1046.935 10815.745 1118.84 ;
      RECT 10754.355 1046.935 10779.355 1189.16 ;
      RECT 10728.355 1046.935 10752.355 1189.16 ;
      RECT 10677.745 1046.935 10701.745 1118.84 ;
      RECT 10664.745 1046.935 10675.745 1118.84 ;
      RECT 10614.355 1046.935 10639.355 1189.16 ;
      RECT 10588.355 1046.935 10612.355 1189.16 ;
      RECT 10537.745 1046.935 10561.745 1118.84 ;
      RECT 10524.745 1046.935 10535.745 1118.84 ;
      RECT 10474.355 1046.935 10499.355 1189.16 ;
      RECT 10448.355 1046.935 10472.355 1189.16 ;
      RECT 10397.745 1046.935 10421.745 1118.84 ;
      RECT 10384.745 1046.935 10395.745 1118.84 ;
      RECT 10334.355 1046.935 10359.355 1189.16 ;
      RECT 10308.355 1046.935 10332.355 1189.16 ;
      RECT 10257.745 1046.935 10281.745 1118.84 ;
      RECT 10244.745 1046.935 10255.745 1118.84 ;
      RECT 10194.355 1046.935 10219.355 1189.16 ;
      RECT 10168.355 1046.935 10192.355 1189.16 ;
      RECT 10117.745 1046.935 10141.745 1118.84 ;
      RECT 10104.745 1046.935 10115.745 1118.84 ;
      RECT 10091.745 1046.935 10102.745 1156.96 ;
      RECT 10054.355 1046.935 10079.355 1189.16 ;
      RECT 10028.355 1046.935 10052.355 1189.16 ;
      RECT 9977.745 1046.935 10001.745 1118.84 ;
      RECT 9964.745 1046.935 9975.745 1118.84 ;
      RECT 9914.355 1046.935 9939.355 1189.16 ;
      RECT 9888.355 1046.935 9912.355 1189.16 ;
      RECT 9837.745 1046.935 9861.745 1118.84 ;
      RECT 9824.745 1046.935 9835.745 1118.84 ;
      RECT 9774.355 1046.935 9799.355 1189.16 ;
      RECT 9748.355 1046.935 9772.355 1189.16 ;
      RECT 9697.745 1046.935 9721.745 1118.84 ;
      RECT 9684.745 1046.935 9695.745 1118.84 ;
      RECT 9634.355 1046.935 9659.355 1189.16 ;
      RECT 9608.355 1046.935 9632.355 1189.16 ;
      RECT 9557.745 1046.935 9581.745 1118.84 ;
      RECT 9544.745 1046.935 9555.745 1118.84 ;
      RECT 9494.355 1046.935 9519.355 1189.16 ;
      RECT 9468.355 1046.935 9492.355 1189.16 ;
      RECT 9417.745 1046.935 9441.745 1118.84 ;
      RECT 9404.745 1046.935 9415.745 1118.84 ;
      RECT 9354.355 1046.935 9379.355 1189.16 ;
      RECT 9328.355 1046.935 9352.355 1189.16 ;
      RECT 9277.745 1046.935 9301.745 1118.84 ;
      RECT 9264.745 1046.935 9275.745 1118.84 ;
      RECT 9214.355 1046.935 9239.355 1189.16 ;
      RECT 9188.355 1046.935 9212.355 1189.16 ;
      RECT 9137.745 1046.935 9161.745 1118.84 ;
      RECT 9124.745 1046.935 9135.745 1118.84 ;
      RECT 9074.355 1046.935 9099.355 1189.16 ;
      RECT 9048.355 1046.935 9072.355 1189.16 ;
      RECT 8997.745 1046.935 9021.745 1118.84 ;
      RECT 8984.745 1046.935 8995.745 1118.84 ;
      RECT 8934.355 1046.935 8959.355 1189.16 ;
      RECT 8908.355 1046.935 8932.355 1189.16 ;
      RECT 8857.745 1046.935 8881.745 1118.84 ;
      RECT 8844.745 1046.935 8855.745 1118.84 ;
      RECT 8794.355 1046.935 8819.355 1189.16 ;
      RECT 8768.355 1046.935 8792.355 1189.16 ;
      RECT 8717.745 1046.935 8741.745 1118.84 ;
      RECT 8704.745 1046.935 8715.745 1118.84 ;
      RECT 8654.355 1046.935 8679.355 1189.16 ;
      RECT 8628.355 1046.935 8652.355 1189.16 ;
      RECT 8577.745 1046.935 8601.745 1118.84 ;
      RECT 8564.745 1046.935 8575.745 1118.84 ;
      RECT 8514.355 1046.935 8539.355 1189.16 ;
      RECT 8488.355 1046.935 8512.355 1189.16 ;
      RECT 8437.745 1046.935 8461.745 1118.84 ;
      RECT 8424.745 1046.935 8435.745 1118.84 ;
      RECT 8374.355 1046.935 8399.355 1189.16 ;
      RECT 8348.355 1046.935 8372.355 1189.16 ;
      RECT 8297.745 1046.935 8321.745 1118.84 ;
      RECT 8284.745 1046.935 8295.745 1118.84 ;
      RECT 8234.355 1046.935 8259.355 1189.16 ;
      RECT 8208.355 1046.935 8232.355 1189.16 ;
      RECT 8157.745 1046.935 8181.745 1118.84 ;
      RECT 8144.745 1046.935 8155.745 1118.84 ;
      RECT 8094.355 1046.935 8119.355 1189.16 ;
      RECT 8068.355 1046.935 8092.355 1189.16 ;
      RECT 8017.745 1046.935 8041.745 1118.84 ;
      RECT 8004.745 1046.935 8015.745 1118.84 ;
      RECT 7954.355 1046.935 7979.355 1189.16 ;
      RECT 7928.355 1046.935 7952.355 1189.16 ;
      RECT 7877.745 1046.935 7901.745 1118.84 ;
      RECT 7864.745 1046.935 7875.745 1118.84 ;
      RECT 7814.355 1046.935 7839.355 1189.16 ;
      RECT 7788.355 1046.935 7812.355 1189.16 ;
      RECT 7737.745 1046.935 7761.745 1118.84 ;
      RECT 7724.745 1046.935 7735.745 1118.84 ;
      RECT 7674.355 1046.935 7699.355 1189.16 ;
      RECT 7648.355 1046.935 7672.355 1189.16 ;
      RECT 7597.745 1046.935 7621.745 1118.84 ;
      RECT 7584.745 1046.935 7595.745 1118.84 ;
      RECT 7534.355 1046.935 7559.355 1189.16 ;
      RECT 7508.355 1046.935 7532.355 1189.16 ;
      RECT 7457.745 1046.935 7481.745 1118.84 ;
      RECT 7444.745 1046.935 7455.745 1118.84 ;
      RECT 7394.355 1046.935 7419.355 1189.16 ;
      RECT 7368.355 1046.935 7392.355 1189.16 ;
      RECT 7317.745 1046.935 7341.745 1118.84 ;
      RECT 7304.745 1046.935 7315.745 1118.84 ;
      RECT 7254.355 1046.935 7279.355 1189.16 ;
      RECT 7228.355 1046.935 7252.355 1189.16 ;
      RECT 7177.745 1046.935 7201.745 1118.84 ;
      RECT 7164.745 1046.935 7175.745 1118.84 ;
      RECT 7114.355 1046.935 7139.355 1189.16 ;
      RECT 7088.355 1046.935 7112.355 1189.16 ;
      RECT 7037.745 1046.935 7061.745 1118.84 ;
      RECT 7024.745 1046.935 7035.745 1118.84 ;
      RECT 6974.355 1046.935 6999.355 1189.16 ;
      RECT 6948.355 1046.935 6972.355 1189.16 ;
      RECT 6897.745 1046.935 6921.745 1118.84 ;
      RECT 6884.745 1046.935 6895.745 1118.84 ;
      RECT 6834.355 1046.935 6859.355 1189.16 ;
      RECT 6808.355 1046.935 6832.355 1189.16 ;
      RECT 6757.745 1046.935 6781.745 1118.84 ;
      RECT 6744.745 1046.935 6755.745 1118.84 ;
      RECT 6694.355 1046.935 6719.355 1189.16 ;
      RECT 6668.355 1046.935 6692.355 1189.16 ;
      RECT 6617.745 1046.935 6641.745 1118.84 ;
      RECT 6604.745 1046.935 6615.745 1118.84 ;
      RECT 6554.355 1046.935 6579.355 1189.16 ;
      RECT 6528.355 1046.935 6552.355 1189.16 ;
      RECT 6477.745 1046.935 6501.745 1118.84 ;
      RECT 6464.745 1046.935 6475.745 1118.84 ;
      RECT 6414.355 1046.935 6439.355 1189.16 ;
      RECT 6388.355 1046.935 6412.355 1189.16 ;
      RECT 6337.745 1046.935 6361.745 1118.84 ;
      RECT 6324.745 1046.935 6335.745 1118.84 ;
      RECT 6274.355 1046.935 6299.355 1189.16 ;
      RECT 6248.355 1046.935 6272.355 1189.16 ;
      RECT 6197.745 1046.935 6221.745 1118.84 ;
      RECT 6184.745 1046.935 6195.745 1118.84 ;
      RECT 6134.355 1046.935 6159.355 1189.16 ;
      RECT 6108.355 1046.935 6132.355 1189.16 ;
      RECT 6057.745 1046.935 6081.745 1118.84 ;
      RECT 6044.745 1046.935 6055.745 1118.84 ;
      RECT 5994.355 1046.935 6019.355 1189.16 ;
      RECT 5968.355 1046.935 5992.355 1189.16 ;
      RECT 5917.745 1046.935 5941.745 1118.84 ;
      RECT 5904.745 1046.935 5915.745 1118.84 ;
      RECT 5854.355 1046.935 5879.355 1189.16 ;
      RECT 5828.355 1046.935 5852.355 1189.16 ;
      RECT 5777.745 1046.935 5801.745 1118.84 ;
      RECT 5764.745 1046.935 5775.745 1118.84 ;
      RECT 5714.355 1046.935 5739.355 1189.16 ;
      RECT 5688.355 1046.935 5712.355 1189.16 ;
      RECT 5637.745 1046.935 5661.745 1118.84 ;
      RECT 5624.745 1046.935 5635.745 1118.84 ;
      RECT 5574.355 1046.935 5599.355 1189.16 ;
      RECT 5548.355 1046.935 5572.355 1189.16 ;
      RECT 5497.745 1046.935 5521.745 1118.84 ;
      RECT 5484.745 1046.935 5495.745 1118.84 ;
      RECT 5434.355 1046.935 5459.355 1189.16 ;
      RECT 5408.355 1046.935 5432.355 1189.16 ;
      RECT 5357.745 1046.935 5381.745 1118.84 ;
      RECT 5344.745 1046.935 5355.745 1118.84 ;
      RECT 5294.355 1046.935 5319.355 1189.16 ;
      RECT 5268.355 1046.935 5292.355 1189.16 ;
      RECT 5217.745 1046.935 5241.745 1118.84 ;
      RECT 5204.745 1046.935 5215.745 1118.84 ;
      RECT 5154.355 1046.935 5179.355 1189.16 ;
      RECT 5128.355 1046.935 5152.355 1189.16 ;
      RECT 5077.745 1046.935 5101.745 1118.84 ;
      RECT 5064.745 1046.935 5075.745 1118.84 ;
      RECT 5014.355 1046.935 5039.355 1189.16 ;
      RECT 4988.355 1046.935 5012.355 1189.16 ;
      RECT 4937.745 1046.935 4961.745 1118.84 ;
      RECT 4924.745 1046.935 4935.745 1118.84 ;
      RECT 4874.355 1046.935 4899.355 1189.16 ;
      RECT 4848.355 1046.935 4872.355 1189.16 ;
      RECT 4797.745 1046.935 4821.745 1118.84 ;
      RECT 4784.745 1046.935 4795.745 1118.84 ;
      RECT 4734.355 1046.935 4759.355 1189.16 ;
      RECT 4708.355 1046.935 4732.355 1189.16 ;
      RECT 4657.745 1046.935 4681.745 1118.84 ;
      RECT 4644.745 1046.935 4655.745 1118.84 ;
      RECT 4594.355 1046.935 4619.355 1189.16 ;
      RECT 4568.355 1046.935 4592.355 1189.16 ;
      RECT 4517.745 1046.935 4541.745 1118.84 ;
      RECT 4504.745 1046.935 4515.745 1118.84 ;
      RECT 4454.355 1046.935 4479.355 1189.16 ;
      RECT 4428.355 1046.935 4452.355 1189.16 ;
      RECT 4377.745 1046.935 4401.745 1118.84 ;
      RECT 4364.745 1046.935 4375.745 1118.84 ;
      RECT 4314.355 1046.935 4339.355 1189.16 ;
      RECT 4288.355 1046.935 4312.355 1189.16 ;
      RECT 4237.745 1046.935 4261.745 1118.84 ;
      RECT 4224.745 1046.935 4235.745 1118.84 ;
      RECT 4174.355 1046.935 4199.355 1189.16 ;
      RECT 4148.355 1046.935 4172.355 1189.16 ;
      RECT 4097.745 1046.935 4121.745 1118.84 ;
      RECT 4084.745 1046.935 4095.745 1118.84 ;
      RECT 4034.355 1046.935 4059.355 1189.16 ;
      RECT 4008.355 1046.935 4032.355 1189.16 ;
      RECT 3957.745 1046.935 3981.745 1118.84 ;
      RECT 3944.745 1046.935 3955.745 1118.84 ;
      RECT 3894.355 1046.935 3919.355 1189.16 ;
      RECT 3868.355 1046.935 3892.355 1189.16 ;
      RECT 3817.745 1046.935 3841.745 1118.84 ;
      RECT 3804.745 1046.935 3815.745 1118.84 ;
      RECT 3754.355 1046.935 3779.355 1189.16 ;
      RECT 3728.355 1046.935 3752.355 1189.16 ;
      RECT 3677.745 1046.935 3701.745 1118.84 ;
      RECT 3664.745 1046.935 3675.745 1118.84 ;
      RECT 3614.355 1046.935 3639.355 1189.16 ;
      RECT 3588.355 1046.935 3612.355 1189.16 ;
      RECT 3537.745 1046.935 3561.745 1118.84 ;
      RECT 3524.745 1046.935 3535.745 1118.84 ;
      RECT 3474.355 1046.935 3499.355 1189.16 ;
      RECT 3448.355 1046.935 3472.355 1189.16 ;
      RECT 3397.745 1046.935 3421.745 1118.84 ;
      RECT 3384.745 1046.935 3395.745 1118.84 ;
      RECT 3334.355 1046.935 3359.355 1189.16 ;
      RECT 3308.355 1046.935 3332.355 1189.16 ;
      RECT 3257.745 1046.935 3281.745 1118.84 ;
      RECT 3244.745 1046.935 3255.745 1118.84 ;
      RECT 3194.355 1046.935 3219.355 1189.16 ;
      RECT 3168.355 1046.935 3192.355 1189.16 ;
      RECT 3117.745 1046.935 3141.745 1118.84 ;
      RECT 3104.745 1046.935 3115.745 1118.84 ;
      RECT 3054.355 1046.935 3079.355 1189.16 ;
      RECT 3028.355 1046.935 3052.355 1189.16 ;
      RECT 2977.745 1046.935 3001.745 1118.84 ;
      RECT 2964.745 1046.935 2975.745 1118.84 ;
      RECT 2914.355 1046.935 2939.355 1189.16 ;
      RECT 2888.355 1046.935 2912.355 1189.16 ;
      RECT 2837.745 1046.935 2861.745 1118.84 ;
      RECT 2824.745 1046.935 2835.745 1118.84 ;
      RECT 2774.355 1046.935 2799.355 1189.16 ;
      RECT 2748.355 1046.935 2772.355 1189.16 ;
      RECT 2697.745 1046.935 2721.745 1118.84 ;
      RECT 2684.745 1046.935 2695.745 1118.84 ;
      RECT 2634.355 1046.935 2659.355 1189.16 ;
      RECT 2608.355 1046.935 2632.355 1189.16 ;
      RECT 2557.745 1046.935 2581.745 1118.84 ;
      RECT 2544.745 1046.935 2555.745 1118.84 ;
      RECT 2494.355 1046.935 2519.355 1189.16 ;
      RECT 2468.355 1046.935 2492.355 1189.16 ;
      RECT 2417.745 1046.935 2441.745 1118.84 ;
      RECT 2404.745 1046.935 2415.745 1118.84 ;
      RECT 2354.355 1046.935 2379.355 1189.16 ;
      RECT 2328.355 1046.935 2352.355 1189.16 ;
      RECT 2277.745 1046.935 2301.745 1118.84 ;
      RECT 2264.745 1046.935 2275.745 1118.84 ;
      RECT 2214.355 1046.935 2239.355 1189.16 ;
      RECT 2188.355 1046.935 2212.355 1189.16 ;
      RECT 2137.745 1046.935 2161.745 1118.84 ;
      RECT 2124.745 1046.935 2135.745 1118.84 ;
      RECT 2074.355 1046.935 2099.355 1189.16 ;
      RECT 2048.355 1046.935 2072.355 1189.16 ;
      RECT 1997.745 1046.935 2021.745 1118.84 ;
      RECT 1984.745 1046.935 1995.745 1118.84 ;
      RECT 1934.355 1046.935 1959.355 1189.16 ;
      RECT 1908.355 1046.935 1932.355 1189.16 ;
      RECT 1857.745 1046.935 1881.745 1118.84 ;
      RECT 1844.745 1046.935 1855.745 1118.84 ;
      RECT 1794.355 1046.935 1819.355 1189.16 ;
      RECT 1768.355 1046.935 1792.355 1189.16 ;
      RECT 1717.745 1046.935 1741.745 1118.84 ;
      RECT 1704.745 1046.935 1715.745 1118.84 ;
      RECT 1654.355 1046.935 1679.355 1189.16 ;
      RECT 1628.355 1046.935 1652.355 1189.16 ;
      RECT 1577.745 1046.935 1601.745 1118.84 ;
      RECT 1564.745 1046.935 1575.745 1118.84 ;
      RECT 1514.355 1046.935 1539.355 1189.16 ;
      RECT 1488.355 1046.935 1512.355 1189.16 ;
      RECT 1437.745 1046.935 1461.745 1118.84 ;
      RECT 1424.745 1046.935 1435.745 1118.84 ;
      RECT 1374.355 1046.935 1399.355 1189.16 ;
      RECT 1348.355 1046.935 1372.355 1189.16 ;
      RECT 1297.745 1046.935 1321.745 1118.84 ;
      RECT 1284.745 1046.935 1295.745 1118.84 ;
      RECT 1234.355 1046.935 1259.355 1189.16 ;
      RECT 1208.355 1046.935 1232.355 1189.16 ;
      RECT 1157.745 1046.935 1181.745 1118.84 ;
      RECT 1144.745 1046.935 1155.745 1118.84 ;
      RECT 998.24 9258.62 1013.18 9259.94 ;
      RECT 998.24 9297.14 1013.18 9298.46 ;
      RECT 998.24 9330.63 1013.18 9331.95 ;
      RECT 998.24 9369.135 1013.18 9370.455 ;
      RECT 998.24 9402.63 1013.18 9403.95 ;
      RECT 998.24 9441.145 1013.18 9442.465 ;
      RECT 990 9497.56 1010 9527.56 ;
      RECT 990 9529.56 1010 9559.56 ;
      RECT 990 9617.56 1010 9647.56 ;
      RECT 990 9649.56 1010 9679.56 ;
      RECT 990 9737.56 1010 9767.56 ;
      RECT 990 9769.56 1010 9799.56 ;
      RECT 990 9857.56 1010 9887.56 ;
      RECT 990 9889.56 1010 9919.56 ;
      RECT 992.1 1116.79 1001.84 1117.59 ;
      RECT 992.1 1119.19 1001.84 1119.99 ;
      RECT 992.1 1121.59 1001.84 1122.39 ;
      RECT 992.1 1123.99 1001.84 1124.79 ;
      RECT 992.1 1126.39 1001.84 1127.19 ;
    LAYER M3 SPACING 0.28 ;
      RECT 13623.535 1047.855 19161.9 10000 ;
      RECT 19156.575 1046.435 19161.9 10000 ;
      RECT 19014.095 1046.935 19151.535 10000 ;
      RECT 19028.655 1046.435 19151.535 10000 ;
      RECT 18874.095 1046.935 19012.975 10000 ;
      RECT 19010.455 1046.435 19012.975 10000 ;
      RECT 18734.095 1046.935 18872.975 10000 ;
      RECT 18870.455 1046.435 18872.975 10000 ;
      RECT 18594.095 1046.935 18732.975 10000 ;
      RECT 18730.455 1046.435 18732.975 10000 ;
      RECT 18454.095 1046.935 18592.975 10000 ;
      RECT 18590.455 1046.435 18592.975 10000 ;
      RECT 18314.095 1046.935 18452.975 10000 ;
      RECT 18450.455 1046.435 18452.975 10000 ;
      RECT 18174.095 1046.935 18312.975 10000 ;
      RECT 18310.455 1046.435 18312.975 10000 ;
      RECT 18034.095 1046.935 18172.975 10000 ;
      RECT 18170.455 1046.435 18172.975 10000 ;
      RECT 17894.095 1046.935 18032.975 10000 ;
      RECT 18030.455 1046.435 18032.975 10000 ;
      RECT 17754.095 1046.935 17892.975 10000 ;
      RECT 17890.455 1046.435 17892.975 10000 ;
      RECT 17614.095 1046.935 17752.975 10000 ;
      RECT 17750.455 1046.435 17752.975 10000 ;
      RECT 17474.095 1046.935 17612.975 10000 ;
      RECT 17610.455 1046.435 17612.975 10000 ;
      RECT 17334.095 1046.935 17472.975 10000 ;
      RECT 17470.455 1046.435 17472.975 10000 ;
      RECT 17194.095 1046.935 17332.975 10000 ;
      RECT 17330.455 1046.435 17332.975 10000 ;
      RECT 17054.095 1046.935 17192.975 10000 ;
      RECT 17190.455 1046.435 17192.975 10000 ;
      RECT 16914.095 1046.935 17052.975 10000 ;
      RECT 17050.455 1046.435 17052.975 10000 ;
      RECT 16774.095 1046.935 16912.975 10000 ;
      RECT 16910.455 1046.435 16912.975 10000 ;
      RECT 16634.095 1046.935 16772.975 10000 ;
      RECT 16770.455 1046.435 16772.975 10000 ;
      RECT 16494.095 1046.935 16632.975 10000 ;
      RECT 16630.455 1046.435 16632.975 10000 ;
      RECT 16354.095 1046.935 16492.975 10000 ;
      RECT 16490.455 1046.435 16492.975 10000 ;
      RECT 16214.095 1046.935 16352.975 10000 ;
      RECT 16350.455 1046.435 16352.975 10000 ;
      RECT 16074.095 1046.935 16212.975 10000 ;
      RECT 16210.455 1046.435 16212.975 10000 ;
      RECT 15934.095 1046.935 16072.975 10000 ;
      RECT 16070.455 1046.435 16072.975 10000 ;
      RECT 15794.095 1046.935 15932.975 10000 ;
      RECT 15930.455 1046.435 15932.975 10000 ;
      RECT 15654.095 1046.935 15792.975 10000 ;
      RECT 15790.455 1046.435 15792.975 10000 ;
      RECT 15514.095 1046.935 15652.975 10000 ;
      RECT 15650.455 1046.435 15652.975 10000 ;
      RECT 15374.095 1046.935 15512.975 10000 ;
      RECT 15510.455 1046.435 15512.975 10000 ;
      RECT 15234.095 1046.935 15372.975 10000 ;
      RECT 15370.455 1046.435 15372.975 10000 ;
      RECT 15094.095 1046.935 15232.975 10000 ;
      RECT 15230.455 1046.435 15232.975 10000 ;
      RECT 14954.095 1046.935 15092.975 10000 ;
      RECT 15090.455 1046.435 15092.975 10000 ;
      RECT 14814.095 1046.935 14952.975 10000 ;
      RECT 14950.455 1046.435 14952.975 10000 ;
      RECT 14674.095 1046.935 14812.975 10000 ;
      RECT 14810.455 1046.435 14812.975 10000 ;
      RECT 14534.095 1046.935 14672.975 10000 ;
      RECT 14670.455 1046.435 14672.975 10000 ;
      RECT 14394.095 1046.935 14532.975 10000 ;
      RECT 14530.455 1046.435 14532.975 10000 ;
      RECT 14254.095 1046.935 14392.975 10000 ;
      RECT 14390.455 1046.435 14392.975 10000 ;
      RECT 14114.095 1046.935 14252.975 10000 ;
      RECT 14250.455 1046.435 14252.975 10000 ;
      RECT 13974.095 1046.935 14112.975 10000 ;
      RECT 14110.455 1046.435 14112.975 10000 ;
      RECT 13834.095 1046.935 13972.975 10000 ;
      RECT 13970.455 1046.435 13972.975 10000 ;
      RECT 13694.095 1046.935 13832.975 10000 ;
      RECT 13830.455 1046.435 13832.975 10000 ;
      RECT 13623.535 1046.935 13692.975 10000 ;
      RECT 13690.455 1046.435 13692.975 10000 ;
      RECT 19025.015 1046.435 19027.535 10000 ;
      RECT 19021.375 1046.435 19023.895 10000 ;
      RECT 19017.735 1046.435 19020.255 10000 ;
      RECT 19014.095 1046.435 19016.615 10000 ;
      RECT 18951.375 1046.435 19009.335 10000 ;
      RECT 18947.455 1046.435 18950.255 10000 ;
      RECT 18943.535 1046.435 18946.335 10000 ;
      RECT 18939.615 1046.435 18942.415 10000 ;
      RECT 18935.695 1046.435 18938.495 10000 ;
      RECT 18888.655 1046.435 18934.575 10000 ;
      RECT 18885.015 1046.435 18887.535 10000 ;
      RECT 18881.375 1046.435 18883.895 10000 ;
      RECT 18877.735 1046.435 18880.255 10000 ;
      RECT 18874.095 1046.435 18876.615 10000 ;
      RECT 18811.375 1046.435 18869.335 10000 ;
      RECT 18807.455 1046.435 18810.255 10000 ;
      RECT 18803.535 1046.435 18806.335 10000 ;
      RECT 18799.615 1046.435 18802.415 10000 ;
      RECT 18795.695 1046.435 18798.495 10000 ;
      RECT 18748.655 1046.435 18794.575 10000 ;
      RECT 18745.015 1046.435 18747.535 10000 ;
      RECT 18741.375 1046.435 18743.895 10000 ;
      RECT 18737.735 1046.435 18740.255 10000 ;
      RECT 18734.095 1046.435 18736.615 10000 ;
      RECT 18671.375 1046.435 18729.335 10000 ;
      RECT 18667.455 1046.435 18670.255 10000 ;
      RECT 18663.535 1046.435 18666.335 10000 ;
      RECT 18659.615 1046.435 18662.415 10000 ;
      RECT 18655.695 1046.435 18658.495 10000 ;
      RECT 18608.655 1046.435 18654.575 10000 ;
      RECT 18605.015 1046.435 18607.535 10000 ;
      RECT 18601.375 1046.435 18603.895 10000 ;
      RECT 18597.735 1046.435 18600.255 10000 ;
      RECT 18594.095 1046.435 18596.615 10000 ;
      RECT 18531.375 1046.435 18589.335 10000 ;
      RECT 18527.455 1046.435 18530.255 10000 ;
      RECT 18523.535 1046.435 18526.335 10000 ;
      RECT 18519.615 1046.435 18522.415 10000 ;
      RECT 18515.695 1046.435 18518.495 10000 ;
      RECT 18468.655 1046.435 18514.575 10000 ;
      RECT 18465.015 1046.435 18467.535 10000 ;
      RECT 18461.375 1046.435 18463.895 10000 ;
      RECT 18457.735 1046.435 18460.255 10000 ;
      RECT 18454.095 1046.435 18456.615 10000 ;
      RECT 18391.375 1046.435 18449.335 10000 ;
      RECT 18387.455 1046.435 18390.255 10000 ;
      RECT 18383.535 1046.435 18386.335 10000 ;
      RECT 18379.615 1046.435 18382.415 10000 ;
      RECT 18375.695 1046.435 18378.495 10000 ;
      RECT 18328.655 1046.435 18374.575 10000 ;
      RECT 18325.015 1046.435 18327.535 10000 ;
      RECT 18321.375 1046.435 18323.895 10000 ;
      RECT 18317.735 1046.435 18320.255 10000 ;
      RECT 18314.095 1046.435 18316.615 10000 ;
      RECT 18251.375 1046.435 18309.335 10000 ;
      RECT 18247.455 1046.435 18250.255 10000 ;
      RECT 18243.535 1046.435 18246.335 10000 ;
      RECT 18239.615 1046.435 18242.415 10000 ;
      RECT 18235.695 1046.435 18238.495 10000 ;
      RECT 18188.655 1046.435 18234.575 10000 ;
      RECT 18185.015 1046.435 18187.535 10000 ;
      RECT 18181.375 1046.435 18183.895 10000 ;
      RECT 18177.735 1046.435 18180.255 10000 ;
      RECT 18174.095 1046.435 18176.615 10000 ;
      RECT 18111.375 1046.435 18169.335 10000 ;
      RECT 18107.455 1046.435 18110.255 10000 ;
      RECT 18103.535 1046.435 18106.335 10000 ;
      RECT 18099.615 1046.435 18102.415 10000 ;
      RECT 18095.695 1046.435 18098.495 10000 ;
      RECT 18048.655 1046.435 18094.575 10000 ;
      RECT 18045.015 1046.435 18047.535 10000 ;
      RECT 18041.375 1046.435 18043.895 10000 ;
      RECT 18037.735 1046.435 18040.255 10000 ;
      RECT 18034.095 1046.435 18036.615 10000 ;
      RECT 17971.375 1046.435 18029.335 10000 ;
      RECT 17967.455 1046.435 17970.255 10000 ;
      RECT 17963.535 1046.435 17966.335 10000 ;
      RECT 17959.615 1046.435 17962.415 10000 ;
      RECT 17955.695 1046.435 17958.495 10000 ;
      RECT 17908.655 1046.435 17954.575 10000 ;
      RECT 17905.015 1046.435 17907.535 10000 ;
      RECT 17901.375 1046.435 17903.895 10000 ;
      RECT 17897.735 1046.435 17900.255 10000 ;
      RECT 17894.095 1046.435 17896.615 10000 ;
      RECT 17831.375 1046.435 17889.335 10000 ;
      RECT 17827.455 1046.435 17830.255 10000 ;
      RECT 17823.535 1046.435 17826.335 10000 ;
      RECT 17819.615 1046.435 17822.415 10000 ;
      RECT 17815.695 1046.435 17818.495 10000 ;
      RECT 17768.655 1046.435 17814.575 10000 ;
      RECT 17765.015 1046.435 17767.535 10000 ;
      RECT 17761.375 1046.435 17763.895 10000 ;
      RECT 17757.735 1046.435 17760.255 10000 ;
      RECT 17754.095 1046.435 17756.615 10000 ;
      RECT 17691.375 1046.435 17749.335 10000 ;
      RECT 17687.455 1046.435 17690.255 10000 ;
      RECT 17683.535 1046.435 17686.335 10000 ;
      RECT 17679.615 1046.435 17682.415 10000 ;
      RECT 17675.695 1046.435 17678.495 10000 ;
      RECT 17628.655 1046.435 17674.575 10000 ;
      RECT 17625.015 1046.435 17627.535 10000 ;
      RECT 17621.375 1046.435 17623.895 10000 ;
      RECT 17617.735 1046.435 17620.255 10000 ;
      RECT 17614.095 1046.435 17616.615 10000 ;
      RECT 17551.375 1046.435 17609.335 10000 ;
      RECT 17547.455 1046.435 17550.255 10000 ;
      RECT 17543.535 1046.435 17546.335 10000 ;
      RECT 17539.615 1046.435 17542.415 10000 ;
      RECT 17535.695 1046.435 17538.495 10000 ;
      RECT 17488.655 1046.435 17534.575 10000 ;
      RECT 17485.015 1046.435 17487.535 10000 ;
      RECT 17481.375 1046.435 17483.895 10000 ;
      RECT 17477.735 1046.435 17480.255 10000 ;
      RECT 17474.095 1046.435 17476.615 10000 ;
      RECT 17411.375 1046.435 17469.335 10000 ;
      RECT 17407.455 1046.435 17410.255 10000 ;
      RECT 17403.535 1046.435 17406.335 10000 ;
      RECT 17399.615 1046.435 17402.415 10000 ;
      RECT 17395.695 1046.435 17398.495 10000 ;
      RECT 17348.655 1046.435 17394.575 10000 ;
      RECT 17345.015 1046.435 17347.535 10000 ;
      RECT 17341.375 1046.435 17343.895 10000 ;
      RECT 17337.735 1046.435 17340.255 10000 ;
      RECT 17334.095 1046.435 17336.615 10000 ;
      RECT 17271.375 1046.435 17329.335 10000 ;
      RECT 17267.455 1046.435 17270.255 10000 ;
      RECT 17263.535 1046.435 17266.335 10000 ;
      RECT 17259.615 1046.435 17262.415 10000 ;
      RECT 17255.695 1046.435 17258.495 10000 ;
      RECT 17208.655 1046.435 17254.575 10000 ;
      RECT 17205.015 1046.435 17207.535 10000 ;
      RECT 17201.375 1046.435 17203.895 10000 ;
      RECT 17197.735 1046.435 17200.255 10000 ;
      RECT 17194.095 1046.435 17196.615 10000 ;
      RECT 17131.375 1046.435 17189.335 10000 ;
      RECT 17127.455 1046.435 17130.255 10000 ;
      RECT 17123.535 1046.435 17126.335 10000 ;
      RECT 17119.615 1046.435 17122.415 10000 ;
      RECT 17115.695 1046.435 17118.495 10000 ;
      RECT 17068.655 1046.435 17114.575 10000 ;
      RECT 17065.015 1046.435 17067.535 10000 ;
      RECT 17061.375 1046.435 17063.895 10000 ;
      RECT 17057.735 1046.435 17060.255 10000 ;
      RECT 17054.095 1046.435 17056.615 10000 ;
      RECT 16991.375 1046.435 17049.335 10000 ;
      RECT 16987.455 1046.435 16990.255 10000 ;
      RECT 16983.535 1046.435 16986.335 10000 ;
      RECT 16979.615 1046.435 16982.415 10000 ;
      RECT 16975.695 1046.435 16978.495 10000 ;
      RECT 16928.655 1046.435 16974.575 10000 ;
      RECT 16925.015 1046.435 16927.535 10000 ;
      RECT 16921.375 1046.435 16923.895 10000 ;
      RECT 16917.735 1046.435 16920.255 10000 ;
      RECT 16914.095 1046.435 16916.615 10000 ;
      RECT 16851.375 1046.435 16909.335 10000 ;
      RECT 16847.455 1046.435 16850.255 10000 ;
      RECT 16843.535 1046.435 16846.335 10000 ;
      RECT 16839.615 1046.435 16842.415 10000 ;
      RECT 16835.695 1046.435 16838.495 10000 ;
      RECT 16788.655 1046.435 16834.575 10000 ;
      RECT 16785.015 1046.435 16787.535 10000 ;
      RECT 16781.375 1046.435 16783.895 10000 ;
      RECT 16777.735 1046.435 16780.255 10000 ;
      RECT 16774.095 1046.435 16776.615 10000 ;
      RECT 16711.375 1046.435 16769.335 10000 ;
      RECT 16707.455 1046.435 16710.255 10000 ;
      RECT 16703.535 1046.435 16706.335 10000 ;
      RECT 16699.615 1046.435 16702.415 10000 ;
      RECT 16695.695 1046.435 16698.495 10000 ;
      RECT 16648.655 1046.435 16694.575 10000 ;
      RECT 16645.015 1046.435 16647.535 10000 ;
      RECT 16641.375 1046.435 16643.895 10000 ;
      RECT 16637.735 1046.435 16640.255 10000 ;
      RECT 16634.095 1046.435 16636.615 10000 ;
      RECT 16571.375 1046.435 16629.335 10000 ;
      RECT 16567.455 1046.435 16570.255 10000 ;
      RECT 16563.535 1046.435 16566.335 10000 ;
      RECT 16559.615 1046.435 16562.415 10000 ;
      RECT 16555.695 1046.435 16558.495 10000 ;
      RECT 16508.655 1046.435 16554.575 10000 ;
      RECT 16505.015 1046.435 16507.535 10000 ;
      RECT 16501.375 1046.435 16503.895 10000 ;
      RECT 16497.735 1046.435 16500.255 10000 ;
      RECT 16494.095 1046.435 16496.615 10000 ;
      RECT 16431.375 1046.435 16489.335 10000 ;
      RECT 16427.455 1046.435 16430.255 10000 ;
      RECT 16423.535 1046.435 16426.335 10000 ;
      RECT 16419.615 1046.435 16422.415 10000 ;
      RECT 16415.695 1046.435 16418.495 10000 ;
      RECT 16368.655 1046.435 16414.575 10000 ;
      RECT 16365.015 1046.435 16367.535 10000 ;
      RECT 16361.375 1046.435 16363.895 10000 ;
      RECT 16357.735 1046.435 16360.255 10000 ;
      RECT 16354.095 1046.435 16356.615 10000 ;
      RECT 16291.375 1046.435 16349.335 10000 ;
      RECT 16287.455 1046.435 16290.255 10000 ;
      RECT 16283.535 1046.435 16286.335 10000 ;
      RECT 16279.615 1046.435 16282.415 10000 ;
      RECT 16275.695 1046.435 16278.495 10000 ;
      RECT 16228.655 1046.435 16274.575 10000 ;
      RECT 16225.015 1046.435 16227.535 10000 ;
      RECT 16221.375 1046.435 16223.895 10000 ;
      RECT 16217.735 1046.435 16220.255 10000 ;
      RECT 16214.095 1046.435 16216.615 10000 ;
      RECT 16151.375 1046.435 16209.335 10000 ;
      RECT 16147.455 1046.435 16150.255 10000 ;
      RECT 16143.535 1046.435 16146.335 10000 ;
      RECT 16139.615 1046.435 16142.415 10000 ;
      RECT 16135.695 1046.435 16138.495 10000 ;
      RECT 16088.655 1046.435 16134.575 10000 ;
      RECT 16085.015 1046.435 16087.535 10000 ;
      RECT 16081.375 1046.435 16083.895 10000 ;
      RECT 16077.735 1046.435 16080.255 10000 ;
      RECT 16074.095 1046.435 16076.615 10000 ;
      RECT 16011.375 1046.435 16069.335 10000 ;
      RECT 16007.455 1046.435 16010.255 10000 ;
      RECT 16003.535 1046.435 16006.335 10000 ;
      RECT 15999.615 1046.435 16002.415 10000 ;
      RECT 15995.695 1046.435 15998.495 10000 ;
      RECT 15948.655 1046.435 15994.575 10000 ;
      RECT 15945.015 1046.435 15947.535 10000 ;
      RECT 15941.375 1046.435 15943.895 10000 ;
      RECT 15937.735 1046.435 15940.255 10000 ;
      RECT 15934.095 1046.435 15936.615 10000 ;
      RECT 15871.375 1046.435 15929.335 10000 ;
      RECT 15867.455 1046.435 15870.255 10000 ;
      RECT 15863.535 1046.435 15866.335 10000 ;
      RECT 15859.615 1046.435 15862.415 10000 ;
      RECT 15855.695 1046.435 15858.495 10000 ;
      RECT 15808.655 1046.435 15854.575 10000 ;
      RECT 15805.015 1046.435 15807.535 10000 ;
      RECT 15801.375 1046.435 15803.895 10000 ;
      RECT 15797.735 1046.435 15800.255 10000 ;
      RECT 15794.095 1046.435 15796.615 10000 ;
      RECT 15731.375 1046.435 15789.335 10000 ;
      RECT 15727.455 1046.435 15730.255 10000 ;
      RECT 15723.535 1046.435 15726.335 10000 ;
      RECT 15719.615 1046.435 15722.415 10000 ;
      RECT 15715.695 1046.435 15718.495 10000 ;
      RECT 15668.655 1046.435 15714.575 10000 ;
      RECT 15665.015 1046.435 15667.535 10000 ;
      RECT 15661.375 1046.435 15663.895 10000 ;
      RECT 15657.735 1046.435 15660.255 10000 ;
      RECT 15654.095 1046.435 15656.615 10000 ;
      RECT 15591.375 1046.435 15649.335 10000 ;
      RECT 15587.455 1046.435 15590.255 10000 ;
      RECT 15583.535 1046.435 15586.335 10000 ;
      RECT 15579.615 1046.435 15582.415 10000 ;
      RECT 15575.695 1046.435 15578.495 10000 ;
      RECT 15528.655 1046.435 15574.575 10000 ;
      RECT 15525.015 1046.435 15527.535 10000 ;
      RECT 15521.375 1046.435 15523.895 10000 ;
      RECT 15517.735 1046.435 15520.255 10000 ;
      RECT 15514.095 1046.435 15516.615 10000 ;
      RECT 15451.375 1046.435 15509.335 10000 ;
      RECT 15447.455 1046.435 15450.255 10000 ;
      RECT 15443.535 1046.435 15446.335 10000 ;
      RECT 15439.615 1046.435 15442.415 10000 ;
      RECT 15435.695 1046.435 15438.495 10000 ;
      RECT 15388.655 1046.435 15434.575 10000 ;
      RECT 15385.015 1046.435 15387.535 10000 ;
      RECT 15381.375 1046.435 15383.895 10000 ;
      RECT 15377.735 1046.435 15380.255 10000 ;
      RECT 15374.095 1046.435 15376.615 10000 ;
      RECT 15311.375 1046.435 15369.335 10000 ;
      RECT 15307.455 1046.435 15310.255 10000 ;
      RECT 15303.535 1046.435 15306.335 10000 ;
      RECT 15299.615 1046.435 15302.415 10000 ;
      RECT 15295.695 1046.435 15298.495 10000 ;
      RECT 15248.655 1046.435 15294.575 10000 ;
      RECT 15245.015 1046.435 15247.535 10000 ;
      RECT 15241.375 1046.435 15243.895 10000 ;
      RECT 15237.735 1046.435 15240.255 10000 ;
      RECT 15234.095 1046.435 15236.615 10000 ;
      RECT 15171.375 1046.435 15229.335 10000 ;
      RECT 15167.455 1046.435 15170.255 10000 ;
      RECT 15163.535 1046.435 15166.335 10000 ;
      RECT 15159.615 1046.435 15162.415 10000 ;
      RECT 15155.695 1046.435 15158.495 10000 ;
      RECT 15108.655 1046.435 15154.575 10000 ;
      RECT 15105.015 1046.435 15107.535 10000 ;
      RECT 15101.375 1046.435 15103.895 10000 ;
      RECT 15097.735 1046.435 15100.255 10000 ;
      RECT 15094.095 1046.435 15096.615 10000 ;
      RECT 15031.375 1046.435 15089.335 10000 ;
      RECT 15027.455 1046.435 15030.255 10000 ;
      RECT 15023.535 1046.435 15026.335 10000 ;
      RECT 15019.615 1046.435 15022.415 10000 ;
      RECT 15015.695 1046.435 15018.495 10000 ;
      RECT 14968.655 1046.435 15014.575 10000 ;
      RECT 14965.015 1046.435 14967.535 10000 ;
      RECT 14961.375 1046.435 14963.895 10000 ;
      RECT 14957.735 1046.435 14960.255 10000 ;
      RECT 14954.095 1046.435 14956.615 10000 ;
      RECT 14891.375 1046.435 14949.335 10000 ;
      RECT 14887.455 1046.435 14890.255 10000 ;
      RECT 14883.535 1046.435 14886.335 10000 ;
      RECT 14879.615 1046.435 14882.415 10000 ;
      RECT 14875.695 1046.435 14878.495 10000 ;
      RECT 14828.655 1046.435 14874.575 10000 ;
      RECT 14825.015 1046.435 14827.535 10000 ;
      RECT 14821.375 1046.435 14823.895 10000 ;
      RECT 14817.735 1046.435 14820.255 10000 ;
      RECT 14814.095 1046.435 14816.615 10000 ;
      RECT 14751.375 1046.435 14809.335 10000 ;
      RECT 14747.455 1046.435 14750.255 10000 ;
      RECT 14743.535 1046.435 14746.335 10000 ;
      RECT 14739.615 1046.435 14742.415 10000 ;
      RECT 14735.695 1046.435 14738.495 10000 ;
      RECT 14688.655 1046.435 14734.575 10000 ;
      RECT 14685.015 1046.435 14687.535 10000 ;
      RECT 14681.375 1046.435 14683.895 10000 ;
      RECT 14677.735 1046.435 14680.255 10000 ;
      RECT 14674.095 1046.435 14676.615 10000 ;
      RECT 14611.375 1046.435 14669.335 10000 ;
      RECT 14607.455 1046.435 14610.255 10000 ;
      RECT 14603.535 1046.435 14606.335 10000 ;
      RECT 14599.615 1046.435 14602.415 10000 ;
      RECT 14595.695 1046.435 14598.495 10000 ;
      RECT 14548.655 1046.435 14594.575 10000 ;
      RECT 14545.015 1046.435 14547.535 10000 ;
      RECT 14541.375 1046.435 14543.895 10000 ;
      RECT 14537.735 1046.435 14540.255 10000 ;
      RECT 14534.095 1046.435 14536.615 10000 ;
      RECT 14471.375 1046.435 14529.335 10000 ;
      RECT 14467.455 1046.435 14470.255 10000 ;
      RECT 14463.535 1046.435 14466.335 10000 ;
      RECT 14459.615 1046.435 14462.415 10000 ;
      RECT 14455.695 1046.435 14458.495 10000 ;
      RECT 14408.655 1046.435 14454.575 10000 ;
      RECT 14405.015 1046.435 14407.535 10000 ;
      RECT 14401.375 1046.435 14403.895 10000 ;
      RECT 14397.735 1046.435 14400.255 10000 ;
      RECT 14394.095 1046.435 14396.615 10000 ;
      RECT 14331.375 1046.435 14389.335 10000 ;
      RECT 14327.455 1046.435 14330.255 10000 ;
      RECT 14323.535 1046.435 14326.335 10000 ;
      RECT 14319.615 1046.435 14322.415 10000 ;
      RECT 14315.695 1046.435 14318.495 10000 ;
      RECT 14268.655 1046.435 14314.575 10000 ;
      RECT 14265.015 1046.435 14267.535 10000 ;
      RECT 14261.375 1046.435 14263.895 10000 ;
      RECT 14257.735 1046.435 14260.255 10000 ;
      RECT 14254.095 1046.435 14256.615 10000 ;
      RECT 14191.375 1046.435 14249.335 10000 ;
      RECT 14187.455 1046.435 14190.255 10000 ;
      RECT 14183.535 1046.435 14186.335 10000 ;
      RECT 14179.615 1046.435 14182.415 10000 ;
      RECT 14175.695 1046.435 14178.495 10000 ;
      RECT 14128.655 1046.435 14174.575 10000 ;
      RECT 14125.015 1046.435 14127.535 10000 ;
      RECT 14121.375 1046.435 14123.895 10000 ;
      RECT 14117.735 1046.435 14120.255 10000 ;
      RECT 14114.095 1046.435 14116.615 10000 ;
      RECT 14051.375 1046.435 14109.335 10000 ;
      RECT 14047.455 1046.435 14050.255 10000 ;
      RECT 14043.535 1046.435 14046.335 10000 ;
      RECT 14039.615 1046.435 14042.415 10000 ;
      RECT 14035.695 1046.435 14038.495 10000 ;
      RECT 13988.655 1046.435 14034.575 10000 ;
      RECT 13985.015 1046.435 13987.535 10000 ;
      RECT 13981.375 1046.435 13983.895 10000 ;
      RECT 13977.735 1046.435 13980.255 10000 ;
      RECT 13974.095 1046.435 13976.615 10000 ;
      RECT 13911.375 1046.435 13969.335 10000 ;
      RECT 13907.455 1046.435 13910.255 10000 ;
      RECT 13903.535 1046.435 13906.335 10000 ;
      RECT 13899.615 1046.435 13902.415 10000 ;
      RECT 13895.695 1046.435 13898.495 10000 ;
      RECT 13848.655 1046.435 13894.575 10000 ;
      RECT 13845.015 1046.435 13847.535 10000 ;
      RECT 13841.375 1046.435 13843.895 10000 ;
      RECT 13837.735 1046.435 13840.255 10000 ;
      RECT 13834.095 1046.435 13836.615 10000 ;
      RECT 13771.375 1046.435 13829.335 10000 ;
      RECT 13767.455 1046.435 13770.255 10000 ;
      RECT 13763.535 1046.435 13766.335 10000 ;
      RECT 13759.615 1046.435 13762.415 10000 ;
      RECT 13755.695 1046.435 13758.495 10000 ;
      RECT 13708.655 1046.435 13754.575 10000 ;
      RECT 13705.015 1046.435 13707.535 10000 ;
      RECT 13701.375 1046.435 13703.895 10000 ;
      RECT 13697.735 1046.435 13700.255 10000 ;
      RECT 13694.095 1046.435 13696.615 10000 ;
      RECT 13631.375 1046.435 13689.335 10000 ;
      RECT 13627.455 1046.435 13630.255 10000 ;
      RECT 13623.535 1046.435 13626.335 10000 ;
      RECT 998.1 1047.855 13623.535 10000 ;
      RECT 13554.095 1046.935 13623.535 10000 ;
      RECT 13414.095 1046.935 13552.975 10000 ;
      RECT 13550.455 1046.435 13552.975 10000 ;
      RECT 13274.095 1046.935 13412.975 10000 ;
      RECT 13410.455 1046.435 13412.975 10000 ;
      RECT 13134.095 1046.935 13272.975 10000 ;
      RECT 13270.455 1046.435 13272.975 10000 ;
      RECT 12994.095 1046.935 13132.975 10000 ;
      RECT 13130.455 1046.435 13132.975 10000 ;
      RECT 12854.095 1046.935 12992.975 10000 ;
      RECT 12990.455 1046.435 12992.975 10000 ;
      RECT 12714.095 1046.935 12852.975 10000 ;
      RECT 12850.455 1046.435 12852.975 10000 ;
      RECT 12574.095 1046.935 12712.975 10000 ;
      RECT 12710.455 1046.435 12712.975 10000 ;
      RECT 12434.095 1046.935 12572.975 10000 ;
      RECT 12570.455 1046.435 12572.975 10000 ;
      RECT 12294.095 1046.935 12432.975 10000 ;
      RECT 12430.455 1046.435 12432.975 10000 ;
      RECT 12154.095 1046.935 12292.975 10000 ;
      RECT 12290.455 1046.435 12292.975 10000 ;
      RECT 12014.095 1046.935 12152.975 10000 ;
      RECT 12150.455 1046.435 12152.975 10000 ;
      RECT 11874.095 1046.935 12012.975 10000 ;
      RECT 12010.455 1046.435 12012.975 10000 ;
      RECT 11734.095 1046.935 11872.975 10000 ;
      RECT 11870.455 1046.435 11872.975 10000 ;
      RECT 11594.095 1046.935 11732.975 10000 ;
      RECT 11730.455 1046.435 11732.975 10000 ;
      RECT 11454.095 1046.935 11592.975 10000 ;
      RECT 11590.455 1046.435 11592.975 10000 ;
      RECT 11314.095 1046.935 11452.975 10000 ;
      RECT 11450.455 1046.435 11452.975 10000 ;
      RECT 11174.095 1046.935 11312.975 10000 ;
      RECT 11310.455 1046.435 11312.975 10000 ;
      RECT 11034.095 1046.935 11172.975 10000 ;
      RECT 11170.455 1046.435 11172.975 10000 ;
      RECT 10894.095 1046.935 11032.975 10000 ;
      RECT 11030.455 1046.435 11032.975 10000 ;
      RECT 10754.095 1046.935 10892.975 10000 ;
      RECT 10890.455 1046.435 10892.975 10000 ;
      RECT 10614.095 1046.935 10752.975 10000 ;
      RECT 10750.455 1046.435 10752.975 10000 ;
      RECT 10474.095 1046.935 10612.975 10000 ;
      RECT 10610.455 1046.435 10612.975 10000 ;
      RECT 10334.095 1046.935 10472.975 10000 ;
      RECT 10470.455 1046.435 10472.975 10000 ;
      RECT 10194.095 1046.935 10332.975 10000 ;
      RECT 10330.455 1046.435 10332.975 10000 ;
      RECT 10091.745 1047.71 10192.975 10000 ;
      RECT 10190.455 1046.435 10192.975 10000 ;
      RECT 10090.615 1046.435 10090.895 10000 ;
      RECT 10088.935 1046.435 10089.215 10000 ;
      RECT 10087.255 1046.435 10087.535 10000 ;
      RECT 10085.575 1046.435 10085.855 10000 ;
      RECT 10083.895 1046.435 10084.175 10000 ;
      RECT 10082.215 1046.435 10082.495 10000 ;
      RECT 10080.535 1046.435 10080.815 10000 ;
      RECT 10054.095 1046.935 10079.355 10000 ;
      RECT 9914.095 1046.935 10052.975 10000 ;
      RECT 10050.455 1046.435 10052.975 10000 ;
      RECT 9774.095 1046.935 9912.975 10000 ;
      RECT 9910.455 1046.435 9912.975 10000 ;
      RECT 9634.095 1046.935 9772.975 10000 ;
      RECT 9770.455 1046.435 9772.975 10000 ;
      RECT 9494.095 1046.935 9632.975 10000 ;
      RECT 9630.455 1046.435 9632.975 10000 ;
      RECT 9354.095 1046.935 9492.975 10000 ;
      RECT 9490.455 1046.435 9492.975 10000 ;
      RECT 9214.095 1046.935 9352.975 10000 ;
      RECT 9350.455 1046.435 9352.975 10000 ;
      RECT 9074.095 1046.935 9212.975 10000 ;
      RECT 9210.455 1046.435 9212.975 10000 ;
      RECT 8934.095 1046.935 9072.975 10000 ;
      RECT 9070.455 1046.435 9072.975 10000 ;
      RECT 8794.095 1046.935 8932.975 10000 ;
      RECT 8930.455 1046.435 8932.975 10000 ;
      RECT 8654.095 1046.935 8792.975 10000 ;
      RECT 8790.455 1046.435 8792.975 10000 ;
      RECT 8514.095 1046.935 8652.975 10000 ;
      RECT 8650.455 1046.435 8652.975 10000 ;
      RECT 8374.095 1046.935 8512.975 10000 ;
      RECT 8510.455 1046.435 8512.975 10000 ;
      RECT 8234.095 1046.935 8372.975 10000 ;
      RECT 8370.455 1046.435 8372.975 10000 ;
      RECT 8094.095 1046.935 8232.975 10000 ;
      RECT 8230.455 1046.435 8232.975 10000 ;
      RECT 7954.095 1046.935 8092.975 10000 ;
      RECT 8090.455 1046.435 8092.975 10000 ;
      RECT 7814.095 1046.935 7952.975 10000 ;
      RECT 7950.455 1046.435 7952.975 10000 ;
      RECT 7674.095 1046.935 7812.975 10000 ;
      RECT 7810.455 1046.435 7812.975 10000 ;
      RECT 7534.095 1046.935 7672.975 10000 ;
      RECT 7670.455 1046.435 7672.975 10000 ;
      RECT 7394.095 1046.935 7532.975 10000 ;
      RECT 7530.455 1046.435 7532.975 10000 ;
      RECT 7254.095 1046.935 7392.975 10000 ;
      RECT 7390.455 1046.435 7392.975 10000 ;
      RECT 7114.095 1046.935 7252.975 10000 ;
      RECT 7250.455 1046.435 7252.975 10000 ;
      RECT 6974.095 1046.935 7112.975 10000 ;
      RECT 7110.455 1046.435 7112.975 10000 ;
      RECT 6834.095 1046.935 6972.975 10000 ;
      RECT 6970.455 1046.435 6972.975 10000 ;
      RECT 6694.095 1046.935 6832.975 10000 ;
      RECT 6830.455 1046.435 6832.975 10000 ;
      RECT 6554.095 1046.935 6692.975 10000 ;
      RECT 6690.455 1046.435 6692.975 10000 ;
      RECT 6414.095 1046.935 6552.975 10000 ;
      RECT 6550.455 1046.435 6552.975 10000 ;
      RECT 6274.095 1046.935 6412.975 10000 ;
      RECT 6410.455 1046.435 6412.975 10000 ;
      RECT 6134.095 1046.935 6272.975 10000 ;
      RECT 6270.455 1046.435 6272.975 10000 ;
      RECT 5994.095 1046.935 6132.975 10000 ;
      RECT 6130.455 1046.435 6132.975 10000 ;
      RECT 5854.095 1046.935 5992.975 10000 ;
      RECT 5990.455 1046.435 5992.975 10000 ;
      RECT 5714.095 1046.935 5852.975 10000 ;
      RECT 5850.455 1046.435 5852.975 10000 ;
      RECT 5574.095 1046.935 5712.975 10000 ;
      RECT 5710.455 1046.435 5712.975 10000 ;
      RECT 5434.095 1046.935 5572.975 10000 ;
      RECT 5570.455 1046.435 5572.975 10000 ;
      RECT 5294.095 1046.935 5432.975 10000 ;
      RECT 5430.455 1046.435 5432.975 10000 ;
      RECT 5154.095 1046.935 5292.975 10000 ;
      RECT 5290.455 1046.435 5292.975 10000 ;
      RECT 5014.095 1046.935 5152.975 10000 ;
      RECT 5150.455 1046.435 5152.975 10000 ;
      RECT 4874.095 1046.935 5012.975 10000 ;
      RECT 5010.455 1046.435 5012.975 10000 ;
      RECT 4734.095 1046.935 4872.975 10000 ;
      RECT 4870.455 1046.435 4872.975 10000 ;
      RECT 4594.095 1046.935 4732.975 10000 ;
      RECT 4730.455 1046.435 4732.975 10000 ;
      RECT 4454.095 1046.935 4592.975 10000 ;
      RECT 4590.455 1046.435 4592.975 10000 ;
      RECT 4314.095 1046.935 4452.975 10000 ;
      RECT 4450.455 1046.435 4452.975 10000 ;
      RECT 4174.095 1046.935 4312.975 10000 ;
      RECT 4310.455 1046.435 4312.975 10000 ;
      RECT 4034.095 1046.935 4172.975 10000 ;
      RECT 4170.455 1046.435 4172.975 10000 ;
      RECT 3894.095 1046.935 4032.975 10000 ;
      RECT 4030.455 1046.435 4032.975 10000 ;
      RECT 3754.095 1046.935 3892.975 10000 ;
      RECT 3890.455 1046.435 3892.975 10000 ;
      RECT 3614.095 1046.935 3752.975 10000 ;
      RECT 3750.455 1046.435 3752.975 10000 ;
      RECT 3474.095 1046.935 3612.975 10000 ;
      RECT 3610.455 1046.435 3612.975 10000 ;
      RECT 3334.095 1046.935 3472.975 10000 ;
      RECT 3470.455 1046.435 3472.975 10000 ;
      RECT 3194.095 1046.935 3332.975 10000 ;
      RECT 3330.455 1046.435 3332.975 10000 ;
      RECT 3054.095 1046.935 3192.975 10000 ;
      RECT 3190.455 1046.435 3192.975 10000 ;
      RECT 2914.095 1046.935 3052.975 10000 ;
      RECT 3050.455 1046.435 3052.975 10000 ;
      RECT 2774.095 1046.935 2912.975 10000 ;
      RECT 2910.455 1046.435 2912.975 10000 ;
      RECT 2634.095 1046.935 2772.975 10000 ;
      RECT 2770.455 1046.435 2772.975 10000 ;
      RECT 2494.095 1046.935 2632.975 10000 ;
      RECT 2630.455 1046.435 2632.975 10000 ;
      RECT 2354.095 1046.935 2492.975 10000 ;
      RECT 2490.455 1046.435 2492.975 10000 ;
      RECT 2214.095 1046.935 2352.975 10000 ;
      RECT 2350.455 1046.435 2352.975 10000 ;
      RECT 2074.095 1046.935 2212.975 10000 ;
      RECT 2210.455 1046.435 2212.975 10000 ;
      RECT 1934.095 1046.935 2072.975 10000 ;
      RECT 2070.455 1046.435 2072.975 10000 ;
      RECT 1794.095 1046.935 1932.975 10000 ;
      RECT 1930.455 1046.435 1932.975 10000 ;
      RECT 1654.095 1046.935 1792.975 10000 ;
      RECT 1790.455 1046.435 1792.975 10000 ;
      RECT 1514.095 1046.935 1652.975 10000 ;
      RECT 1650.455 1046.435 1652.975 10000 ;
      RECT 1374.095 1046.935 1512.975 10000 ;
      RECT 1510.455 1046.435 1512.975 10000 ;
      RECT 1234.095 1046.935 1372.975 10000 ;
      RECT 1370.455 1046.435 1372.975 10000 ;
      RECT 1008.465 1046.935 1232.975 10000 ;
      RECT 1230.455 1046.435 1232.975 10000 ;
      RECT 998.1 1046.435 1003.425 10000 ;
      RECT 10104.055 1046.935 10192.975 10000 ;
      RECT 10091.745 1046.935 10102.745 10000 ;
      RECT 13619.615 1046.435 13622.415 10000 ;
      RECT 13615.695 1046.435 13618.495 10000 ;
      RECT 13568.655 1046.435 13614.575 10000 ;
      RECT 13565.015 1046.435 13567.535 10000 ;
      RECT 13561.375 1046.435 13563.895 10000 ;
      RECT 13557.735 1046.435 13560.255 10000 ;
      RECT 13554.095 1046.435 13556.615 10000 ;
      RECT 13491.375 1046.435 13549.335 10000 ;
      RECT 13487.455 1046.435 13490.255 10000 ;
      RECT 13483.535 1046.435 13486.335 10000 ;
      RECT 13479.615 1046.435 13482.415 10000 ;
      RECT 13475.695 1046.435 13478.495 10000 ;
      RECT 13428.655 1046.435 13474.575 10000 ;
      RECT 13425.015 1046.435 13427.535 10000 ;
      RECT 13421.375 1046.435 13423.895 10000 ;
      RECT 13417.735 1046.435 13420.255 10000 ;
      RECT 13414.095 1046.435 13416.615 10000 ;
      RECT 13351.375 1046.435 13409.335 10000 ;
      RECT 13347.455 1046.435 13350.255 10000 ;
      RECT 13343.535 1046.435 13346.335 10000 ;
      RECT 13339.615 1046.435 13342.415 10000 ;
      RECT 13335.695 1046.435 13338.495 10000 ;
      RECT 13288.655 1046.435 13334.575 10000 ;
      RECT 13285.015 1046.435 13287.535 10000 ;
      RECT 13281.375 1046.435 13283.895 10000 ;
      RECT 13277.735 1046.435 13280.255 10000 ;
      RECT 13274.095 1046.435 13276.615 10000 ;
      RECT 13211.375 1046.435 13269.335 10000 ;
      RECT 13207.455 1046.435 13210.255 10000 ;
      RECT 13203.535 1046.435 13206.335 10000 ;
      RECT 13199.615 1046.435 13202.415 10000 ;
      RECT 13195.695 1046.435 13198.495 10000 ;
      RECT 13148.655 1046.435 13194.575 10000 ;
      RECT 13145.015 1046.435 13147.535 10000 ;
      RECT 13141.375 1046.435 13143.895 10000 ;
      RECT 13137.735 1046.435 13140.255 10000 ;
      RECT 13134.095 1046.435 13136.615 10000 ;
      RECT 13071.375 1046.435 13129.335 10000 ;
      RECT 13067.455 1046.435 13070.255 10000 ;
      RECT 13063.535 1046.435 13066.335 10000 ;
      RECT 13059.615 1046.435 13062.415 10000 ;
      RECT 13055.695 1046.435 13058.495 10000 ;
      RECT 13008.655 1046.435 13054.575 10000 ;
      RECT 13005.015 1046.435 13007.535 10000 ;
      RECT 13001.375 1046.435 13003.895 10000 ;
      RECT 12997.735 1046.435 13000.255 10000 ;
      RECT 12994.095 1046.435 12996.615 10000 ;
      RECT 12931.375 1046.435 12989.335 10000 ;
      RECT 12927.455 1046.435 12930.255 10000 ;
      RECT 12923.535 1046.435 12926.335 10000 ;
      RECT 12919.615 1046.435 12922.415 10000 ;
      RECT 12915.695 1046.435 12918.495 10000 ;
      RECT 12868.655 1046.435 12914.575 10000 ;
      RECT 12865.015 1046.435 12867.535 10000 ;
      RECT 12861.375 1046.435 12863.895 10000 ;
      RECT 12857.735 1046.435 12860.255 10000 ;
      RECT 12854.095 1046.435 12856.615 10000 ;
      RECT 12791.375 1046.435 12849.335 10000 ;
      RECT 12787.455 1046.435 12790.255 10000 ;
      RECT 12783.535 1046.435 12786.335 10000 ;
      RECT 12779.615 1046.435 12782.415 10000 ;
      RECT 12775.695 1046.435 12778.495 10000 ;
      RECT 12728.655 1046.435 12774.575 10000 ;
      RECT 12725.015 1046.435 12727.535 10000 ;
      RECT 12721.375 1046.435 12723.895 10000 ;
      RECT 12717.735 1046.435 12720.255 10000 ;
      RECT 12714.095 1046.435 12716.615 10000 ;
      RECT 12651.375 1046.435 12709.335 10000 ;
      RECT 12647.455 1046.435 12650.255 10000 ;
      RECT 12643.535 1046.435 12646.335 10000 ;
      RECT 12639.615 1046.435 12642.415 10000 ;
      RECT 12635.695 1046.435 12638.495 10000 ;
      RECT 12588.655 1046.435 12634.575 10000 ;
      RECT 12585.015 1046.435 12587.535 10000 ;
      RECT 12581.375 1046.435 12583.895 10000 ;
      RECT 12577.735 1046.435 12580.255 10000 ;
      RECT 12574.095 1046.435 12576.615 10000 ;
      RECT 12511.375 1046.435 12569.335 10000 ;
      RECT 12507.455 1046.435 12510.255 10000 ;
      RECT 12503.535 1046.435 12506.335 10000 ;
      RECT 12499.615 1046.435 12502.415 10000 ;
      RECT 12495.695 1046.435 12498.495 10000 ;
      RECT 12448.655 1046.435 12494.575 10000 ;
      RECT 12445.015 1046.435 12447.535 10000 ;
      RECT 12441.375 1046.435 12443.895 10000 ;
      RECT 12437.735 1046.435 12440.255 10000 ;
      RECT 12434.095 1046.435 12436.615 10000 ;
      RECT 12371.375 1046.435 12429.335 10000 ;
      RECT 12367.455 1046.435 12370.255 10000 ;
      RECT 12363.535 1046.435 12366.335 10000 ;
      RECT 12359.615 1046.435 12362.415 10000 ;
      RECT 12355.695 1046.435 12358.495 10000 ;
      RECT 12308.655 1046.435 12354.575 10000 ;
      RECT 12305.015 1046.435 12307.535 10000 ;
      RECT 12301.375 1046.435 12303.895 10000 ;
      RECT 12297.735 1046.435 12300.255 10000 ;
      RECT 12294.095 1046.435 12296.615 10000 ;
      RECT 12231.375 1046.435 12289.335 10000 ;
      RECT 12227.455 1046.435 12230.255 10000 ;
      RECT 12223.535 1046.435 12226.335 10000 ;
      RECT 12219.615 1046.435 12222.415 10000 ;
      RECT 12215.695 1046.435 12218.495 10000 ;
      RECT 12168.655 1046.435 12214.575 10000 ;
      RECT 12165.015 1046.435 12167.535 10000 ;
      RECT 12161.375 1046.435 12163.895 10000 ;
      RECT 12157.735 1046.435 12160.255 10000 ;
      RECT 12154.095 1046.435 12156.615 10000 ;
      RECT 12091.375 1046.435 12149.335 10000 ;
      RECT 12087.455 1046.435 12090.255 10000 ;
      RECT 12083.535 1046.435 12086.335 10000 ;
      RECT 12079.615 1046.435 12082.415 10000 ;
      RECT 12075.695 1046.435 12078.495 10000 ;
      RECT 12028.655 1046.435 12074.575 10000 ;
      RECT 12025.015 1046.435 12027.535 10000 ;
      RECT 12021.375 1046.435 12023.895 10000 ;
      RECT 12017.735 1046.435 12020.255 10000 ;
      RECT 12014.095 1046.435 12016.615 10000 ;
      RECT 11951.375 1046.435 12009.335 10000 ;
      RECT 11947.455 1046.435 11950.255 10000 ;
      RECT 11943.535 1046.435 11946.335 10000 ;
      RECT 11939.615 1046.435 11942.415 10000 ;
      RECT 11935.695 1046.435 11938.495 10000 ;
      RECT 11888.655 1046.435 11934.575 10000 ;
      RECT 11885.015 1046.435 11887.535 10000 ;
      RECT 11881.375 1046.435 11883.895 10000 ;
      RECT 11877.735 1046.435 11880.255 10000 ;
      RECT 11874.095 1046.435 11876.615 10000 ;
      RECT 11811.375 1046.435 11869.335 10000 ;
      RECT 11807.455 1046.435 11810.255 10000 ;
      RECT 11803.535 1046.435 11806.335 10000 ;
      RECT 11799.615 1046.435 11802.415 10000 ;
      RECT 11795.695 1046.435 11798.495 10000 ;
      RECT 11748.655 1046.435 11794.575 10000 ;
      RECT 11745.015 1046.435 11747.535 10000 ;
      RECT 11741.375 1046.435 11743.895 10000 ;
      RECT 11737.735 1046.435 11740.255 10000 ;
      RECT 11734.095 1046.435 11736.615 10000 ;
      RECT 11671.375 1046.435 11729.335 10000 ;
      RECT 11667.455 1046.435 11670.255 10000 ;
      RECT 11663.535 1046.435 11666.335 10000 ;
      RECT 11659.615 1046.435 11662.415 10000 ;
      RECT 11655.695 1046.435 11658.495 10000 ;
      RECT 11608.655 1046.435 11654.575 10000 ;
      RECT 11605.015 1046.435 11607.535 10000 ;
      RECT 11601.375 1046.435 11603.895 10000 ;
      RECT 11597.735 1046.435 11600.255 10000 ;
      RECT 11594.095 1046.435 11596.615 10000 ;
      RECT 11531.375 1046.435 11589.335 10000 ;
      RECT 11527.455 1046.435 11530.255 10000 ;
      RECT 11523.535 1046.435 11526.335 10000 ;
      RECT 11519.615 1046.435 11522.415 10000 ;
      RECT 11515.695 1046.435 11518.495 10000 ;
      RECT 11468.655 1046.435 11514.575 10000 ;
      RECT 11465.015 1046.435 11467.535 10000 ;
      RECT 11461.375 1046.435 11463.895 10000 ;
      RECT 11457.735 1046.435 11460.255 10000 ;
      RECT 11454.095 1046.435 11456.615 10000 ;
      RECT 11391.375 1046.435 11449.335 10000 ;
      RECT 11387.455 1046.435 11390.255 10000 ;
      RECT 11383.535 1046.435 11386.335 10000 ;
      RECT 11379.615 1046.435 11382.415 10000 ;
      RECT 11375.695 1046.435 11378.495 10000 ;
      RECT 11328.655 1046.435 11374.575 10000 ;
      RECT 11325.015 1046.435 11327.535 10000 ;
      RECT 11321.375 1046.435 11323.895 10000 ;
      RECT 11317.735 1046.435 11320.255 10000 ;
      RECT 11314.095 1046.435 11316.615 10000 ;
      RECT 11251.375 1046.435 11309.335 10000 ;
      RECT 11247.455 1046.435 11250.255 10000 ;
      RECT 11243.535 1046.435 11246.335 10000 ;
      RECT 11239.615 1046.435 11242.415 10000 ;
      RECT 11235.695 1046.435 11238.495 10000 ;
      RECT 11188.655 1046.435 11234.575 10000 ;
      RECT 11185.015 1046.435 11187.535 10000 ;
      RECT 11181.375 1046.435 11183.895 10000 ;
      RECT 11177.735 1046.435 11180.255 10000 ;
      RECT 11174.095 1046.435 11176.615 10000 ;
      RECT 11111.375 1046.435 11169.335 10000 ;
      RECT 11107.455 1046.435 11110.255 10000 ;
      RECT 11103.535 1046.435 11106.335 10000 ;
      RECT 11099.615 1046.435 11102.415 10000 ;
      RECT 11095.695 1046.435 11098.495 10000 ;
      RECT 11048.655 1046.435 11094.575 10000 ;
      RECT 11045.015 1046.435 11047.535 10000 ;
      RECT 11041.375 1046.435 11043.895 10000 ;
      RECT 11037.735 1046.435 11040.255 10000 ;
      RECT 11034.095 1046.435 11036.615 10000 ;
      RECT 10971.375 1046.435 11029.335 10000 ;
      RECT 10967.455 1046.435 10970.255 10000 ;
      RECT 10963.535 1046.435 10966.335 10000 ;
      RECT 10959.615 1046.435 10962.415 10000 ;
      RECT 10955.695 1046.435 10958.495 10000 ;
      RECT 10908.655 1046.435 10954.575 10000 ;
      RECT 10905.015 1046.435 10907.535 10000 ;
      RECT 10901.375 1046.435 10903.895 10000 ;
      RECT 10897.735 1046.435 10900.255 10000 ;
      RECT 10894.095 1046.435 10896.615 10000 ;
      RECT 10831.375 1046.435 10889.335 10000 ;
      RECT 10827.455 1046.435 10830.255 10000 ;
      RECT 10823.535 1046.435 10826.335 10000 ;
      RECT 10819.615 1046.435 10822.415 10000 ;
      RECT 10815.695 1046.435 10818.495 10000 ;
      RECT 10768.655 1046.435 10814.575 10000 ;
      RECT 10765.015 1046.435 10767.535 10000 ;
      RECT 10761.375 1046.435 10763.895 10000 ;
      RECT 10757.735 1046.435 10760.255 10000 ;
      RECT 10754.095 1046.435 10756.615 10000 ;
      RECT 10691.375 1046.435 10749.335 10000 ;
      RECT 10687.455 1046.435 10690.255 10000 ;
      RECT 10683.535 1046.435 10686.335 10000 ;
      RECT 10679.615 1046.435 10682.415 10000 ;
      RECT 10675.695 1046.435 10678.495 10000 ;
      RECT 10628.655 1046.435 10674.575 10000 ;
      RECT 10625.015 1046.435 10627.535 10000 ;
      RECT 10621.375 1046.435 10623.895 10000 ;
      RECT 10617.735 1046.435 10620.255 10000 ;
      RECT 10614.095 1046.435 10616.615 10000 ;
      RECT 10551.375 1046.435 10609.335 10000 ;
      RECT 10547.455 1046.435 10550.255 10000 ;
      RECT 10543.535 1046.435 10546.335 10000 ;
      RECT 10539.615 1046.435 10542.415 10000 ;
      RECT 10535.695 1046.435 10538.495 10000 ;
      RECT 10488.655 1046.435 10534.575 10000 ;
      RECT 10485.015 1046.435 10487.535 10000 ;
      RECT 10481.375 1046.435 10483.895 10000 ;
      RECT 10477.735 1046.435 10480.255 10000 ;
      RECT 10474.095 1046.435 10476.615 10000 ;
      RECT 10411.375 1046.435 10469.335 10000 ;
      RECT 10407.455 1046.435 10410.255 10000 ;
      RECT 10403.535 1046.435 10406.335 10000 ;
      RECT 10399.615 1046.435 10402.415 10000 ;
      RECT 10395.695 1046.435 10398.495 10000 ;
      RECT 10348.655 1046.435 10394.575 10000 ;
      RECT 10345.015 1046.435 10347.535 10000 ;
      RECT 10341.375 1046.435 10343.895 10000 ;
      RECT 10337.735 1046.435 10340.255 10000 ;
      RECT 10334.095 1046.435 10336.615 10000 ;
      RECT 10271.375 1046.435 10329.335 10000 ;
      RECT 10267.455 1046.435 10270.255 10000 ;
      RECT 10263.535 1046.435 10266.335 10000 ;
      RECT 10259.615 1046.435 10262.415 10000 ;
      RECT 10255.695 1046.435 10258.495 10000 ;
      RECT 10208.655 1046.435 10254.575 10000 ;
      RECT 10205.015 1046.435 10207.535 10000 ;
      RECT 10201.375 1046.435 10203.895 10000 ;
      RECT 10197.735 1046.435 10200.255 10000 ;
      RECT 10194.095 1046.435 10196.615 10000 ;
      RECT 10131.375 1046.435 10189.335 10000 ;
      RECT 10127.455 1046.435 10130.255 10000 ;
      RECT 10123.535 1046.435 10126.335 10000 ;
      RECT 10119.615 1046.435 10122.415 10000 ;
      RECT 10115.695 1046.435 10118.495 10000 ;
      RECT 10104.055 1046.435 10114.575 10000 ;
      RECT 10102.375 1046.435 10102.655 10000 ;
      RECT 10100.695 1046.435 10100.975 10000 ;
      RECT 10099.015 1046.435 10099.295 10000 ;
      RECT 10097.335 1046.435 10097.615 10000 ;
      RECT 10095.655 1046.435 10095.935 10000 ;
      RECT 10093.975 1046.435 10094.255 10000 ;
      RECT 10092.295 1046.435 10092.575 10000 ;
      RECT 10068.655 1046.435 10079.135 10000 ;
      RECT 10065.015 1046.435 10067.535 10000 ;
      RECT 10061.375 1046.435 10063.895 10000 ;
      RECT 10057.735 1046.435 10060.255 10000 ;
      RECT 10054.095 1046.435 10056.615 10000 ;
      RECT 9991.375 1046.435 10049.335 10000 ;
      RECT 9987.455 1046.435 9990.255 10000 ;
      RECT 9983.535 1046.435 9986.335 10000 ;
      RECT 9979.615 1046.435 9982.415 10000 ;
      RECT 9975.695 1046.435 9978.495 10000 ;
      RECT 9928.655 1046.435 9974.575 10000 ;
      RECT 9925.015 1046.435 9927.535 10000 ;
      RECT 9921.375 1046.435 9923.895 10000 ;
      RECT 9917.735 1046.435 9920.255 10000 ;
      RECT 9914.095 1046.435 9916.615 10000 ;
      RECT 9851.375 1046.435 9909.335 10000 ;
      RECT 9847.455 1046.435 9850.255 10000 ;
      RECT 9843.535 1046.435 9846.335 10000 ;
      RECT 9839.615 1046.435 9842.415 10000 ;
      RECT 9835.695 1046.435 9838.495 10000 ;
      RECT 9788.655 1046.435 9834.575 10000 ;
      RECT 9785.015 1046.435 9787.535 10000 ;
      RECT 9781.375 1046.435 9783.895 10000 ;
      RECT 9777.735 1046.435 9780.255 10000 ;
      RECT 9774.095 1046.435 9776.615 10000 ;
      RECT 9711.375 1046.435 9769.335 10000 ;
      RECT 9707.455 1046.435 9710.255 10000 ;
      RECT 9703.535 1046.435 9706.335 10000 ;
      RECT 9699.615 1046.435 9702.415 10000 ;
      RECT 9695.695 1046.435 9698.495 10000 ;
      RECT 9648.655 1046.435 9694.575 10000 ;
      RECT 9645.015 1046.435 9647.535 10000 ;
      RECT 9641.375 1046.435 9643.895 10000 ;
      RECT 9637.735 1046.435 9640.255 10000 ;
      RECT 9634.095 1046.435 9636.615 10000 ;
      RECT 9571.375 1046.435 9629.335 10000 ;
      RECT 9567.455 1046.435 9570.255 10000 ;
      RECT 9563.535 1046.435 9566.335 10000 ;
      RECT 9559.615 1046.435 9562.415 10000 ;
      RECT 9555.695 1046.435 9558.495 10000 ;
      RECT 9508.655 1046.435 9554.575 10000 ;
      RECT 9505.015 1046.435 9507.535 10000 ;
      RECT 9501.375 1046.435 9503.895 10000 ;
      RECT 9497.735 1046.435 9500.255 10000 ;
      RECT 9494.095 1046.435 9496.615 10000 ;
      RECT 9431.375 1046.435 9489.335 10000 ;
      RECT 9427.455 1046.435 9430.255 10000 ;
      RECT 9423.535 1046.435 9426.335 10000 ;
      RECT 9419.615 1046.435 9422.415 10000 ;
      RECT 9415.695 1046.435 9418.495 10000 ;
      RECT 9368.655 1046.435 9414.575 10000 ;
      RECT 9365.015 1046.435 9367.535 10000 ;
      RECT 9361.375 1046.435 9363.895 10000 ;
      RECT 9357.735 1046.435 9360.255 10000 ;
      RECT 9354.095 1046.435 9356.615 10000 ;
      RECT 9291.375 1046.435 9349.335 10000 ;
      RECT 9287.455 1046.435 9290.255 10000 ;
      RECT 9283.535 1046.435 9286.335 10000 ;
      RECT 9279.615 1046.435 9282.415 10000 ;
      RECT 9275.695 1046.435 9278.495 10000 ;
      RECT 9228.655 1046.435 9274.575 10000 ;
      RECT 9225.015 1046.435 9227.535 10000 ;
      RECT 9221.375 1046.435 9223.895 10000 ;
      RECT 9217.735 1046.435 9220.255 10000 ;
      RECT 9214.095 1046.435 9216.615 10000 ;
      RECT 9151.375 1046.435 9209.335 10000 ;
      RECT 9147.455 1046.435 9150.255 10000 ;
      RECT 9143.535 1046.435 9146.335 10000 ;
      RECT 9139.615 1046.435 9142.415 10000 ;
      RECT 9135.695 1046.435 9138.495 10000 ;
      RECT 9088.655 1046.435 9134.575 10000 ;
      RECT 9085.015 1046.435 9087.535 10000 ;
      RECT 9081.375 1046.435 9083.895 10000 ;
      RECT 9077.735 1046.435 9080.255 10000 ;
      RECT 9074.095 1046.435 9076.615 10000 ;
      RECT 9011.375 1046.435 9069.335 10000 ;
      RECT 9007.455 1046.435 9010.255 10000 ;
      RECT 9003.535 1046.435 9006.335 10000 ;
      RECT 8999.615 1046.435 9002.415 10000 ;
      RECT 8995.695 1046.435 8998.495 10000 ;
      RECT 8948.655 1046.435 8994.575 10000 ;
      RECT 8945.015 1046.435 8947.535 10000 ;
      RECT 8941.375 1046.435 8943.895 10000 ;
      RECT 8937.735 1046.435 8940.255 10000 ;
      RECT 8934.095 1046.435 8936.615 10000 ;
      RECT 8871.375 1046.435 8929.335 10000 ;
      RECT 8867.455 1046.435 8870.255 10000 ;
      RECT 8863.535 1046.435 8866.335 10000 ;
      RECT 8859.615 1046.435 8862.415 10000 ;
      RECT 8855.695 1046.435 8858.495 10000 ;
      RECT 8808.655 1046.435 8854.575 10000 ;
      RECT 8805.015 1046.435 8807.535 10000 ;
      RECT 8801.375 1046.435 8803.895 10000 ;
      RECT 8797.735 1046.435 8800.255 10000 ;
      RECT 8794.095 1046.435 8796.615 10000 ;
      RECT 8731.375 1046.435 8789.335 10000 ;
      RECT 8727.455 1046.435 8730.255 10000 ;
      RECT 8723.535 1046.435 8726.335 10000 ;
      RECT 8719.615 1046.435 8722.415 10000 ;
      RECT 8715.695 1046.435 8718.495 10000 ;
      RECT 8668.655 1046.435 8714.575 10000 ;
      RECT 8665.015 1046.435 8667.535 10000 ;
      RECT 8661.375 1046.435 8663.895 10000 ;
      RECT 8657.735 1046.435 8660.255 10000 ;
      RECT 8654.095 1046.435 8656.615 10000 ;
      RECT 8591.375 1046.435 8649.335 10000 ;
      RECT 8587.455 1046.435 8590.255 10000 ;
      RECT 8583.535 1046.435 8586.335 10000 ;
      RECT 8579.615 1046.435 8582.415 10000 ;
      RECT 8575.695 1046.435 8578.495 10000 ;
      RECT 8528.655 1046.435 8574.575 10000 ;
      RECT 8525.015 1046.435 8527.535 10000 ;
      RECT 8521.375 1046.435 8523.895 10000 ;
      RECT 8517.735 1046.435 8520.255 10000 ;
      RECT 8514.095 1046.435 8516.615 10000 ;
      RECT 8451.375 1046.435 8509.335 10000 ;
      RECT 8447.455 1046.435 8450.255 10000 ;
      RECT 8443.535 1046.435 8446.335 10000 ;
      RECT 8439.615 1046.435 8442.415 10000 ;
      RECT 8435.695 1046.435 8438.495 10000 ;
      RECT 8388.655 1046.435 8434.575 10000 ;
      RECT 8385.015 1046.435 8387.535 10000 ;
      RECT 8381.375 1046.435 8383.895 10000 ;
      RECT 8377.735 1046.435 8380.255 10000 ;
      RECT 8374.095 1046.435 8376.615 10000 ;
      RECT 8311.375 1046.435 8369.335 10000 ;
      RECT 8307.455 1046.435 8310.255 10000 ;
      RECT 8303.535 1046.435 8306.335 10000 ;
      RECT 8299.615 1046.435 8302.415 10000 ;
      RECT 8295.695 1046.435 8298.495 10000 ;
      RECT 8248.655 1046.435 8294.575 10000 ;
      RECT 8245.015 1046.435 8247.535 10000 ;
      RECT 8241.375 1046.435 8243.895 10000 ;
      RECT 8237.735 1046.435 8240.255 10000 ;
      RECT 8234.095 1046.435 8236.615 10000 ;
      RECT 8171.375 1046.435 8229.335 10000 ;
      RECT 8167.455 1046.435 8170.255 10000 ;
      RECT 8163.535 1046.435 8166.335 10000 ;
      RECT 8159.615 1046.435 8162.415 10000 ;
      RECT 8155.695 1046.435 8158.495 10000 ;
      RECT 8108.655 1046.435 8154.575 10000 ;
      RECT 8105.015 1046.435 8107.535 10000 ;
      RECT 8101.375 1046.435 8103.895 10000 ;
      RECT 8097.735 1046.435 8100.255 10000 ;
      RECT 8094.095 1046.435 8096.615 10000 ;
      RECT 8031.375 1046.435 8089.335 10000 ;
      RECT 8027.455 1046.435 8030.255 10000 ;
      RECT 8023.535 1046.435 8026.335 10000 ;
      RECT 8019.615 1046.435 8022.415 10000 ;
      RECT 8015.695 1046.435 8018.495 10000 ;
      RECT 7968.655 1046.435 8014.575 10000 ;
      RECT 7965.015 1046.435 7967.535 10000 ;
      RECT 7961.375 1046.435 7963.895 10000 ;
      RECT 7957.735 1046.435 7960.255 10000 ;
      RECT 7954.095 1046.435 7956.615 10000 ;
      RECT 7891.375 1046.435 7949.335 10000 ;
      RECT 7887.455 1046.435 7890.255 10000 ;
      RECT 7883.535 1046.435 7886.335 10000 ;
      RECT 7879.615 1046.435 7882.415 10000 ;
      RECT 7875.695 1046.435 7878.495 10000 ;
      RECT 7828.655 1046.435 7874.575 10000 ;
      RECT 7825.015 1046.435 7827.535 10000 ;
      RECT 7821.375 1046.435 7823.895 10000 ;
      RECT 7817.735 1046.435 7820.255 10000 ;
      RECT 7814.095 1046.435 7816.615 10000 ;
      RECT 7751.375 1046.435 7809.335 10000 ;
      RECT 7747.455 1046.435 7750.255 10000 ;
      RECT 7743.535 1046.435 7746.335 10000 ;
      RECT 7739.615 1046.435 7742.415 10000 ;
      RECT 7735.695 1046.435 7738.495 10000 ;
      RECT 7688.655 1046.435 7734.575 10000 ;
      RECT 7685.015 1046.435 7687.535 10000 ;
      RECT 7681.375 1046.435 7683.895 10000 ;
      RECT 7677.735 1046.435 7680.255 10000 ;
      RECT 7674.095 1046.435 7676.615 10000 ;
      RECT 7611.375 1046.435 7669.335 10000 ;
      RECT 7607.455 1046.435 7610.255 10000 ;
      RECT 7603.535 1046.435 7606.335 10000 ;
      RECT 7599.615 1046.435 7602.415 10000 ;
      RECT 7595.695 1046.435 7598.495 10000 ;
      RECT 7548.655 1046.435 7594.575 10000 ;
      RECT 7545.015 1046.435 7547.535 10000 ;
      RECT 7541.375 1046.435 7543.895 10000 ;
      RECT 7537.735 1046.435 7540.255 10000 ;
      RECT 7534.095 1046.435 7536.615 10000 ;
      RECT 7471.375 1046.435 7529.335 10000 ;
      RECT 7467.455 1046.435 7470.255 10000 ;
      RECT 7463.535 1046.435 7466.335 10000 ;
      RECT 7459.615 1046.435 7462.415 10000 ;
      RECT 7455.695 1046.435 7458.495 10000 ;
      RECT 7408.655 1046.435 7454.575 10000 ;
      RECT 7405.015 1046.435 7407.535 10000 ;
      RECT 7401.375 1046.435 7403.895 10000 ;
      RECT 7397.735 1046.435 7400.255 10000 ;
      RECT 7394.095 1046.435 7396.615 10000 ;
      RECT 7331.375 1046.435 7389.335 10000 ;
      RECT 7327.455 1046.435 7330.255 10000 ;
      RECT 7323.535 1046.435 7326.335 10000 ;
      RECT 7319.615 1046.435 7322.415 10000 ;
      RECT 7315.695 1046.435 7318.495 10000 ;
      RECT 7268.655 1046.435 7314.575 10000 ;
      RECT 7265.015 1046.435 7267.535 10000 ;
      RECT 7261.375 1046.435 7263.895 10000 ;
      RECT 7257.735 1046.435 7260.255 10000 ;
      RECT 7254.095 1046.435 7256.615 10000 ;
      RECT 7191.375 1046.435 7249.335 10000 ;
      RECT 7187.455 1046.435 7190.255 10000 ;
      RECT 7183.535 1046.435 7186.335 10000 ;
      RECT 7179.615 1046.435 7182.415 10000 ;
      RECT 7175.695 1046.435 7178.495 10000 ;
      RECT 7128.655 1046.435 7174.575 10000 ;
      RECT 7125.015 1046.435 7127.535 10000 ;
      RECT 7121.375 1046.435 7123.895 10000 ;
      RECT 7117.735 1046.435 7120.255 10000 ;
      RECT 7114.095 1046.435 7116.615 10000 ;
      RECT 7051.375 1046.435 7109.335 10000 ;
      RECT 7047.455 1046.435 7050.255 10000 ;
      RECT 7043.535 1046.435 7046.335 10000 ;
      RECT 7039.615 1046.435 7042.415 10000 ;
      RECT 7035.695 1046.435 7038.495 10000 ;
      RECT 6988.655 1046.435 7034.575 10000 ;
      RECT 6985.015 1046.435 6987.535 10000 ;
      RECT 6981.375 1046.435 6983.895 10000 ;
      RECT 6977.735 1046.435 6980.255 10000 ;
      RECT 6974.095 1046.435 6976.615 10000 ;
      RECT 6911.375 1046.435 6969.335 10000 ;
      RECT 6907.455 1046.435 6910.255 10000 ;
      RECT 6903.535 1046.435 6906.335 10000 ;
      RECT 6899.615 1046.435 6902.415 10000 ;
      RECT 6895.695 1046.435 6898.495 10000 ;
      RECT 6848.655 1046.435 6894.575 10000 ;
      RECT 6845.015 1046.435 6847.535 10000 ;
      RECT 6841.375 1046.435 6843.895 10000 ;
      RECT 6837.735 1046.435 6840.255 10000 ;
      RECT 6834.095 1046.435 6836.615 10000 ;
      RECT 6771.375 1046.435 6829.335 10000 ;
      RECT 6767.455 1046.435 6770.255 10000 ;
      RECT 6763.535 1046.435 6766.335 10000 ;
      RECT 6759.615 1046.435 6762.415 10000 ;
      RECT 6755.695 1046.435 6758.495 10000 ;
      RECT 6708.655 1046.435 6754.575 10000 ;
      RECT 6705.015 1046.435 6707.535 10000 ;
      RECT 6701.375 1046.435 6703.895 10000 ;
      RECT 6697.735 1046.435 6700.255 10000 ;
      RECT 6694.095 1046.435 6696.615 10000 ;
      RECT 6631.375 1046.435 6689.335 10000 ;
      RECT 6627.455 1046.435 6630.255 10000 ;
      RECT 6623.535 1046.435 6626.335 10000 ;
      RECT 6619.615 1046.435 6622.415 10000 ;
      RECT 6615.695 1046.435 6618.495 10000 ;
      RECT 6568.655 1046.435 6614.575 10000 ;
      RECT 6565.015 1046.435 6567.535 10000 ;
      RECT 6561.375 1046.435 6563.895 10000 ;
      RECT 6557.735 1046.435 6560.255 10000 ;
      RECT 6554.095 1046.435 6556.615 10000 ;
      RECT 6491.375 1046.435 6549.335 10000 ;
      RECT 6487.455 1046.435 6490.255 10000 ;
      RECT 6483.535 1046.435 6486.335 10000 ;
      RECT 6479.615 1046.435 6482.415 10000 ;
      RECT 6475.695 1046.435 6478.495 10000 ;
      RECT 6428.655 1046.435 6474.575 10000 ;
      RECT 6425.015 1046.435 6427.535 10000 ;
      RECT 6421.375 1046.435 6423.895 10000 ;
      RECT 6417.735 1046.435 6420.255 10000 ;
      RECT 6414.095 1046.435 6416.615 10000 ;
      RECT 6351.375 1046.435 6409.335 10000 ;
      RECT 6347.455 1046.435 6350.255 10000 ;
      RECT 6343.535 1046.435 6346.335 10000 ;
      RECT 6339.615 1046.435 6342.415 10000 ;
      RECT 6335.695 1046.435 6338.495 10000 ;
      RECT 6288.655 1046.435 6334.575 10000 ;
      RECT 6285.015 1046.435 6287.535 10000 ;
      RECT 6281.375 1046.435 6283.895 10000 ;
      RECT 6277.735 1046.435 6280.255 10000 ;
      RECT 6274.095 1046.435 6276.615 10000 ;
      RECT 6211.375 1046.435 6269.335 10000 ;
      RECT 6207.455 1046.435 6210.255 10000 ;
      RECT 6203.535 1046.435 6206.335 10000 ;
      RECT 6199.615 1046.435 6202.415 10000 ;
      RECT 6195.695 1046.435 6198.495 10000 ;
      RECT 6148.655 1046.435 6194.575 10000 ;
      RECT 6145.015 1046.435 6147.535 10000 ;
      RECT 6141.375 1046.435 6143.895 10000 ;
      RECT 6137.735 1046.435 6140.255 10000 ;
      RECT 6134.095 1046.435 6136.615 10000 ;
      RECT 6071.375 1046.435 6129.335 10000 ;
      RECT 6067.455 1046.435 6070.255 10000 ;
      RECT 6063.535 1046.435 6066.335 10000 ;
      RECT 6059.615 1046.435 6062.415 10000 ;
      RECT 6055.695 1046.435 6058.495 10000 ;
      RECT 6008.655 1046.435 6054.575 10000 ;
      RECT 6005.015 1046.435 6007.535 10000 ;
      RECT 6001.375 1046.435 6003.895 10000 ;
      RECT 5997.735 1046.435 6000.255 10000 ;
      RECT 5994.095 1046.435 5996.615 10000 ;
      RECT 5931.375 1046.435 5989.335 10000 ;
      RECT 5927.455 1046.435 5930.255 10000 ;
      RECT 5923.535 1046.435 5926.335 10000 ;
      RECT 5919.615 1046.435 5922.415 10000 ;
      RECT 5915.695 1046.435 5918.495 10000 ;
      RECT 5868.655 1046.435 5914.575 10000 ;
      RECT 5865.015 1046.435 5867.535 10000 ;
      RECT 5861.375 1046.435 5863.895 10000 ;
      RECT 5857.735 1046.435 5860.255 10000 ;
      RECT 5854.095 1046.435 5856.615 10000 ;
      RECT 5791.375 1046.435 5849.335 10000 ;
      RECT 5787.455 1046.435 5790.255 10000 ;
      RECT 5783.535 1046.435 5786.335 10000 ;
      RECT 5779.615 1046.435 5782.415 10000 ;
      RECT 5775.695 1046.435 5778.495 10000 ;
      RECT 5728.655 1046.435 5774.575 10000 ;
      RECT 5725.015 1046.435 5727.535 10000 ;
      RECT 5721.375 1046.435 5723.895 10000 ;
      RECT 5717.735 1046.435 5720.255 10000 ;
      RECT 5714.095 1046.435 5716.615 10000 ;
      RECT 5651.375 1046.435 5709.335 10000 ;
      RECT 5647.455 1046.435 5650.255 10000 ;
      RECT 5643.535 1046.435 5646.335 10000 ;
      RECT 5639.615 1046.435 5642.415 10000 ;
      RECT 5635.695 1046.435 5638.495 10000 ;
      RECT 5588.655 1046.435 5634.575 10000 ;
      RECT 5585.015 1046.435 5587.535 10000 ;
      RECT 5581.375 1046.435 5583.895 10000 ;
      RECT 5577.735 1046.435 5580.255 10000 ;
      RECT 5574.095 1046.435 5576.615 10000 ;
      RECT 5511.375 1046.435 5569.335 10000 ;
      RECT 5507.455 1046.435 5510.255 10000 ;
      RECT 5503.535 1046.435 5506.335 10000 ;
      RECT 5499.615 1046.435 5502.415 10000 ;
      RECT 5495.695 1046.435 5498.495 10000 ;
      RECT 5448.655 1046.435 5494.575 10000 ;
      RECT 5445.015 1046.435 5447.535 10000 ;
      RECT 5441.375 1046.435 5443.895 10000 ;
      RECT 5437.735 1046.435 5440.255 10000 ;
      RECT 5434.095 1046.435 5436.615 10000 ;
      RECT 5371.375 1046.435 5429.335 10000 ;
      RECT 5367.455 1046.435 5370.255 10000 ;
      RECT 5363.535 1046.435 5366.335 10000 ;
      RECT 5359.615 1046.435 5362.415 10000 ;
      RECT 5355.695 1046.435 5358.495 10000 ;
      RECT 5308.655 1046.435 5354.575 10000 ;
      RECT 5305.015 1046.435 5307.535 10000 ;
      RECT 5301.375 1046.435 5303.895 10000 ;
      RECT 5297.735 1046.435 5300.255 10000 ;
      RECT 5294.095 1046.435 5296.615 10000 ;
      RECT 5231.375 1046.435 5289.335 10000 ;
      RECT 5227.455 1046.435 5230.255 10000 ;
      RECT 5223.535 1046.435 5226.335 10000 ;
      RECT 5219.615 1046.435 5222.415 10000 ;
      RECT 5215.695 1046.435 5218.495 10000 ;
      RECT 5168.655 1046.435 5214.575 10000 ;
      RECT 5165.015 1046.435 5167.535 10000 ;
      RECT 5161.375 1046.435 5163.895 10000 ;
      RECT 5157.735 1046.435 5160.255 10000 ;
      RECT 5154.095 1046.435 5156.615 10000 ;
      RECT 5091.375 1046.435 5149.335 10000 ;
      RECT 5087.455 1046.435 5090.255 10000 ;
      RECT 5083.535 1046.435 5086.335 10000 ;
      RECT 5079.615 1046.435 5082.415 10000 ;
      RECT 5075.695 1046.435 5078.495 10000 ;
      RECT 5028.655 1046.435 5074.575 10000 ;
      RECT 5025.015 1046.435 5027.535 10000 ;
      RECT 5021.375 1046.435 5023.895 10000 ;
      RECT 5017.735 1046.435 5020.255 10000 ;
      RECT 5014.095 1046.435 5016.615 10000 ;
      RECT 4951.375 1046.435 5009.335 10000 ;
      RECT 4947.455 1046.435 4950.255 10000 ;
      RECT 4943.535 1046.435 4946.335 10000 ;
      RECT 4939.615 1046.435 4942.415 10000 ;
      RECT 4935.695 1046.435 4938.495 10000 ;
      RECT 4888.655 1046.435 4934.575 10000 ;
      RECT 4885.015 1046.435 4887.535 10000 ;
      RECT 4881.375 1046.435 4883.895 10000 ;
      RECT 4877.735 1046.435 4880.255 10000 ;
      RECT 4874.095 1046.435 4876.615 10000 ;
      RECT 4811.375 1046.435 4869.335 10000 ;
      RECT 4807.455 1046.435 4810.255 10000 ;
      RECT 4803.535 1046.435 4806.335 10000 ;
      RECT 4799.615 1046.435 4802.415 10000 ;
      RECT 4795.695 1046.435 4798.495 10000 ;
      RECT 4748.655 1046.435 4794.575 10000 ;
      RECT 4745.015 1046.435 4747.535 10000 ;
      RECT 4741.375 1046.435 4743.895 10000 ;
      RECT 4737.735 1046.435 4740.255 10000 ;
      RECT 4734.095 1046.435 4736.615 10000 ;
      RECT 4671.375 1046.435 4729.335 10000 ;
      RECT 4667.455 1046.435 4670.255 10000 ;
      RECT 4663.535 1046.435 4666.335 10000 ;
      RECT 4659.615 1046.435 4662.415 10000 ;
      RECT 4655.695 1046.435 4658.495 10000 ;
      RECT 4608.655 1046.435 4654.575 10000 ;
      RECT 4605.015 1046.435 4607.535 10000 ;
      RECT 4601.375 1046.435 4603.895 10000 ;
      RECT 4597.735 1046.435 4600.255 10000 ;
      RECT 4594.095 1046.435 4596.615 10000 ;
      RECT 4531.375 1046.435 4589.335 10000 ;
      RECT 4527.455 1046.435 4530.255 10000 ;
      RECT 4523.535 1046.435 4526.335 10000 ;
      RECT 4519.615 1046.435 4522.415 10000 ;
      RECT 4515.695 1046.435 4518.495 10000 ;
      RECT 4468.655 1046.435 4514.575 10000 ;
      RECT 4465.015 1046.435 4467.535 10000 ;
      RECT 4461.375 1046.435 4463.895 10000 ;
      RECT 4457.735 1046.435 4460.255 10000 ;
      RECT 4454.095 1046.435 4456.615 10000 ;
      RECT 4391.375 1046.435 4449.335 10000 ;
      RECT 4387.455 1046.435 4390.255 10000 ;
      RECT 4383.535 1046.435 4386.335 10000 ;
      RECT 4379.615 1046.435 4382.415 10000 ;
      RECT 4375.695 1046.435 4378.495 10000 ;
      RECT 4328.655 1046.435 4374.575 10000 ;
      RECT 4325.015 1046.435 4327.535 10000 ;
      RECT 4321.375 1046.435 4323.895 10000 ;
      RECT 4317.735 1046.435 4320.255 10000 ;
      RECT 4314.095 1046.435 4316.615 10000 ;
      RECT 4251.375 1046.435 4309.335 10000 ;
      RECT 4247.455 1046.435 4250.255 10000 ;
      RECT 4243.535 1046.435 4246.335 10000 ;
      RECT 4239.615 1046.435 4242.415 10000 ;
      RECT 4235.695 1046.435 4238.495 10000 ;
      RECT 4188.655 1046.435 4234.575 10000 ;
      RECT 4185.015 1046.435 4187.535 10000 ;
      RECT 4181.375 1046.435 4183.895 10000 ;
      RECT 4177.735 1046.435 4180.255 10000 ;
      RECT 4174.095 1046.435 4176.615 10000 ;
      RECT 4111.375 1046.435 4169.335 10000 ;
      RECT 4107.455 1046.435 4110.255 10000 ;
      RECT 4103.535 1046.435 4106.335 10000 ;
      RECT 4099.615 1046.435 4102.415 10000 ;
      RECT 4095.695 1046.435 4098.495 10000 ;
      RECT 4048.655 1046.435 4094.575 10000 ;
      RECT 4045.015 1046.435 4047.535 10000 ;
      RECT 4041.375 1046.435 4043.895 10000 ;
      RECT 4037.735 1046.435 4040.255 10000 ;
      RECT 4034.095 1046.435 4036.615 10000 ;
      RECT 3971.375 1046.435 4029.335 10000 ;
      RECT 3967.455 1046.435 3970.255 10000 ;
      RECT 3963.535 1046.435 3966.335 10000 ;
      RECT 3959.615 1046.435 3962.415 10000 ;
      RECT 3955.695 1046.435 3958.495 10000 ;
      RECT 3908.655 1046.435 3954.575 10000 ;
      RECT 3905.015 1046.435 3907.535 10000 ;
      RECT 3901.375 1046.435 3903.895 10000 ;
      RECT 3897.735 1046.435 3900.255 10000 ;
      RECT 3894.095 1046.435 3896.615 10000 ;
      RECT 3831.375 1046.435 3889.335 10000 ;
      RECT 3827.455 1046.435 3830.255 10000 ;
      RECT 3823.535 1046.435 3826.335 10000 ;
      RECT 3819.615 1046.435 3822.415 10000 ;
      RECT 3815.695 1046.435 3818.495 10000 ;
      RECT 3768.655 1046.435 3814.575 10000 ;
      RECT 3765.015 1046.435 3767.535 10000 ;
      RECT 3761.375 1046.435 3763.895 10000 ;
      RECT 3757.735 1046.435 3760.255 10000 ;
      RECT 3754.095 1046.435 3756.615 10000 ;
      RECT 3691.375 1046.435 3749.335 10000 ;
      RECT 3687.455 1046.435 3690.255 10000 ;
      RECT 3683.535 1046.435 3686.335 10000 ;
      RECT 3679.615 1046.435 3682.415 10000 ;
      RECT 3675.695 1046.435 3678.495 10000 ;
      RECT 3628.655 1046.435 3674.575 10000 ;
      RECT 3625.015 1046.435 3627.535 10000 ;
      RECT 3621.375 1046.435 3623.895 10000 ;
      RECT 3617.735 1046.435 3620.255 10000 ;
      RECT 3614.095 1046.435 3616.615 10000 ;
      RECT 3551.375 1046.435 3609.335 10000 ;
      RECT 3547.455 1046.435 3550.255 10000 ;
      RECT 3543.535 1046.435 3546.335 10000 ;
      RECT 3539.615 1046.435 3542.415 10000 ;
      RECT 3535.695 1046.435 3538.495 10000 ;
      RECT 3488.655 1046.435 3534.575 10000 ;
      RECT 3485.015 1046.435 3487.535 10000 ;
      RECT 3481.375 1046.435 3483.895 10000 ;
      RECT 3477.735 1046.435 3480.255 10000 ;
      RECT 3474.095 1046.435 3476.615 10000 ;
      RECT 3411.375 1046.435 3469.335 10000 ;
      RECT 3407.455 1046.435 3410.255 10000 ;
      RECT 3403.535 1046.435 3406.335 10000 ;
      RECT 3399.615 1046.435 3402.415 10000 ;
      RECT 3395.695 1046.435 3398.495 10000 ;
      RECT 3348.655 1046.435 3394.575 10000 ;
      RECT 3345.015 1046.435 3347.535 10000 ;
      RECT 3341.375 1046.435 3343.895 10000 ;
      RECT 3337.735 1046.435 3340.255 10000 ;
      RECT 3334.095 1046.435 3336.615 10000 ;
      RECT 3271.375 1046.435 3329.335 10000 ;
      RECT 3267.455 1046.435 3270.255 10000 ;
      RECT 3263.535 1046.435 3266.335 10000 ;
      RECT 3259.615 1046.435 3262.415 10000 ;
      RECT 3255.695 1046.435 3258.495 10000 ;
      RECT 3208.655 1046.435 3254.575 10000 ;
      RECT 3205.015 1046.435 3207.535 10000 ;
      RECT 3201.375 1046.435 3203.895 10000 ;
      RECT 3197.735 1046.435 3200.255 10000 ;
      RECT 3194.095 1046.435 3196.615 10000 ;
      RECT 3131.375 1046.435 3189.335 10000 ;
      RECT 3127.455 1046.435 3130.255 10000 ;
      RECT 3123.535 1046.435 3126.335 10000 ;
      RECT 3119.615 1046.435 3122.415 10000 ;
      RECT 3115.695 1046.435 3118.495 10000 ;
      RECT 3068.655 1046.435 3114.575 10000 ;
      RECT 3065.015 1046.435 3067.535 10000 ;
      RECT 3061.375 1046.435 3063.895 10000 ;
      RECT 3057.735 1046.435 3060.255 10000 ;
      RECT 3054.095 1046.435 3056.615 10000 ;
      RECT 2991.375 1046.435 3049.335 10000 ;
      RECT 2987.455 1046.435 2990.255 10000 ;
      RECT 2983.535 1046.435 2986.335 10000 ;
      RECT 2979.615 1046.435 2982.415 10000 ;
      RECT 2975.695 1046.435 2978.495 10000 ;
      RECT 2928.655 1046.435 2974.575 10000 ;
      RECT 2925.015 1046.435 2927.535 10000 ;
      RECT 2921.375 1046.435 2923.895 10000 ;
      RECT 2917.735 1046.435 2920.255 10000 ;
      RECT 2914.095 1046.435 2916.615 10000 ;
      RECT 2851.375 1046.435 2909.335 10000 ;
      RECT 2847.455 1046.435 2850.255 10000 ;
      RECT 2843.535 1046.435 2846.335 10000 ;
      RECT 2839.615 1046.435 2842.415 10000 ;
      RECT 2835.695 1046.435 2838.495 10000 ;
      RECT 2788.655 1046.435 2834.575 10000 ;
      RECT 2785.015 1046.435 2787.535 10000 ;
      RECT 2781.375 1046.435 2783.895 10000 ;
      RECT 2777.735 1046.435 2780.255 10000 ;
      RECT 2774.095 1046.435 2776.615 10000 ;
      RECT 2711.375 1046.435 2769.335 10000 ;
      RECT 2707.455 1046.435 2710.255 10000 ;
      RECT 2703.535 1046.435 2706.335 10000 ;
      RECT 2699.615 1046.435 2702.415 10000 ;
      RECT 2695.695 1046.435 2698.495 10000 ;
      RECT 2648.655 1046.435 2694.575 10000 ;
      RECT 2645.015 1046.435 2647.535 10000 ;
      RECT 2641.375 1046.435 2643.895 10000 ;
      RECT 2637.735 1046.435 2640.255 10000 ;
      RECT 2634.095 1046.435 2636.615 10000 ;
      RECT 2571.375 1046.435 2629.335 10000 ;
      RECT 2567.455 1046.435 2570.255 10000 ;
      RECT 2563.535 1046.435 2566.335 10000 ;
      RECT 2559.615 1046.435 2562.415 10000 ;
      RECT 2555.695 1046.435 2558.495 10000 ;
      RECT 2508.655 1046.435 2554.575 10000 ;
      RECT 2505.015 1046.435 2507.535 10000 ;
      RECT 2501.375 1046.435 2503.895 10000 ;
      RECT 2497.735 1046.435 2500.255 10000 ;
      RECT 2494.095 1046.435 2496.615 10000 ;
      RECT 2431.375 1046.435 2489.335 10000 ;
      RECT 2427.455 1046.435 2430.255 10000 ;
      RECT 2423.535 1046.435 2426.335 10000 ;
      RECT 2419.615 1046.435 2422.415 10000 ;
      RECT 2415.695 1046.435 2418.495 10000 ;
      RECT 2368.655 1046.435 2414.575 10000 ;
      RECT 2365.015 1046.435 2367.535 10000 ;
      RECT 2361.375 1046.435 2363.895 10000 ;
      RECT 2357.735 1046.435 2360.255 10000 ;
      RECT 2354.095 1046.435 2356.615 10000 ;
      RECT 2291.375 1046.435 2349.335 10000 ;
      RECT 2287.455 1046.435 2290.255 10000 ;
      RECT 2283.535 1046.435 2286.335 10000 ;
      RECT 2279.615 1046.435 2282.415 10000 ;
      RECT 2275.695 1046.435 2278.495 10000 ;
      RECT 2228.655 1046.435 2274.575 10000 ;
      RECT 2225.015 1046.435 2227.535 10000 ;
      RECT 2221.375 1046.435 2223.895 10000 ;
      RECT 2217.735 1046.435 2220.255 10000 ;
      RECT 2214.095 1046.435 2216.615 10000 ;
      RECT 2151.375 1046.435 2209.335 10000 ;
      RECT 2147.455 1046.435 2150.255 10000 ;
      RECT 2143.535 1046.435 2146.335 10000 ;
      RECT 2139.615 1046.435 2142.415 10000 ;
      RECT 2135.695 1046.435 2138.495 10000 ;
      RECT 2088.655 1046.435 2134.575 10000 ;
      RECT 2085.015 1046.435 2087.535 10000 ;
      RECT 2081.375 1046.435 2083.895 10000 ;
      RECT 2077.735 1046.435 2080.255 10000 ;
      RECT 2074.095 1046.435 2076.615 10000 ;
      RECT 2011.375 1046.435 2069.335 10000 ;
      RECT 2007.455 1046.435 2010.255 10000 ;
      RECT 2003.535 1046.435 2006.335 10000 ;
      RECT 1999.615 1046.435 2002.415 10000 ;
      RECT 1995.695 1046.435 1998.495 10000 ;
      RECT 1948.655 1046.435 1994.575 10000 ;
      RECT 1945.015 1046.435 1947.535 10000 ;
      RECT 1941.375 1046.435 1943.895 10000 ;
      RECT 1937.735 1046.435 1940.255 10000 ;
      RECT 1934.095 1046.435 1936.615 10000 ;
      RECT 1871.375 1046.435 1929.335 10000 ;
      RECT 1867.455 1046.435 1870.255 10000 ;
      RECT 1863.535 1046.435 1866.335 10000 ;
      RECT 1859.615 1046.435 1862.415 10000 ;
      RECT 1855.695 1046.435 1858.495 10000 ;
      RECT 1808.655 1046.435 1854.575 10000 ;
      RECT 1805.015 1046.435 1807.535 10000 ;
      RECT 1801.375 1046.435 1803.895 10000 ;
      RECT 1797.735 1046.435 1800.255 10000 ;
      RECT 1794.095 1046.435 1796.615 10000 ;
      RECT 1731.375 1046.435 1789.335 10000 ;
      RECT 1727.455 1046.435 1730.255 10000 ;
      RECT 1723.535 1046.435 1726.335 10000 ;
      RECT 1719.615 1046.435 1722.415 10000 ;
      RECT 1715.695 1046.435 1718.495 10000 ;
      RECT 1668.655 1046.435 1714.575 10000 ;
      RECT 1665.015 1046.435 1667.535 10000 ;
      RECT 1661.375 1046.435 1663.895 10000 ;
      RECT 1657.735 1046.435 1660.255 10000 ;
      RECT 1654.095 1046.435 1656.615 10000 ;
      RECT 1591.375 1046.435 1649.335 10000 ;
      RECT 1587.455 1046.435 1590.255 10000 ;
      RECT 1583.535 1046.435 1586.335 10000 ;
      RECT 1579.615 1046.435 1582.415 10000 ;
      RECT 1575.695 1046.435 1578.495 10000 ;
      RECT 1528.655 1046.435 1574.575 10000 ;
      RECT 1525.015 1046.435 1527.535 10000 ;
      RECT 1521.375 1046.435 1523.895 10000 ;
      RECT 1517.735 1046.435 1520.255 10000 ;
      RECT 1514.095 1046.435 1516.615 10000 ;
      RECT 1451.375 1046.435 1509.335 10000 ;
      RECT 1447.455 1046.435 1450.255 10000 ;
      RECT 1443.535 1046.435 1446.335 10000 ;
      RECT 1439.615 1046.435 1442.415 10000 ;
      RECT 1435.695 1046.435 1438.495 10000 ;
      RECT 1388.655 1046.435 1434.575 10000 ;
      RECT 1385.015 1046.435 1387.535 10000 ;
      RECT 1381.375 1046.435 1383.895 10000 ;
      RECT 1377.735 1046.435 1380.255 10000 ;
      RECT 1374.095 1046.435 1376.615 10000 ;
      RECT 1311.375 1046.435 1369.335 10000 ;
      RECT 1307.455 1046.435 1310.255 10000 ;
      RECT 1303.535 1046.435 1306.335 10000 ;
      RECT 1299.615 1046.435 1302.415 10000 ;
      RECT 1295.695 1046.435 1298.495 10000 ;
      RECT 1248.655 1046.435 1294.575 10000 ;
      RECT 1245.015 1046.435 1247.535 10000 ;
      RECT 1241.375 1046.435 1243.895 10000 ;
      RECT 1237.735 1046.435 1240.255 10000 ;
      RECT 1234.095 1046.435 1236.615 10000 ;
      RECT 1171.375 1046.435 1229.335 10000 ;
      RECT 1167.455 1046.435 1170.255 10000 ;
      RECT 1163.535 1046.435 1166.335 10000 ;
      RECT 1159.615 1046.435 1162.415 10000 ;
      RECT 1155.695 1046.435 1158.495 10000 ;
      RECT 1008.465 1046.435 1154.575 10000 ;
    LAYER M4 ;
      RECT 4.1 9990 20195.9 9995.9 ;
      RECT 20190 4.1 20195.9 9995.9 ;
      RECT 4.1 4.1 10 9995.9 ;
      RECT 4.1 4.1 20195.9 10 ;
      RECT 19160.9 9258.575 19161.9 9259.995 ;
      RECT 19146.82 9258.62 19161.9 9259.94 ;
      RECT 19160.9 9297.09 19161.9 9298.51 ;
      RECT 19146.82 9297.14 19161.9 9298.46 ;
      RECT 19160.9 9330.575 19161.9 9331.995 ;
      RECT 19146.82 9330.63 19161.9 9331.95 ;
      RECT 19160.9 9369.09 19161.9 9370.51 ;
      RECT 19146.82 9369.135 19161.9 9370.455 ;
      RECT 19160.9 9402.575 19161.9 9403.995 ;
      RECT 19146.82 9402.63 19161.9 9403.95 ;
      RECT 19160.9 9441.09 19161.9 9442.51 ;
      RECT 19146.82 9441.145 19161.9 9442.465 ;
      RECT 998.1 9258.575 999.1 9259.995 ;
      RECT 998.1 9258.62 1013.18 9259.94 ;
      RECT 998.1 9297.09 999.1 9298.51 ;
      RECT 998.1 9297.14 1013.18 9298.46 ;
      RECT 998.1 9330.575 999.1 9331.995 ;
      RECT 998.1 9330.63 1013.18 9331.95 ;
      RECT 998.1 9369.09 999.1 9370.51 ;
      RECT 998.1 9369.135 1013.18 9370.455 ;
      RECT 998.1 9402.575 999.1 9403.995 ;
      RECT 998.1 9402.63 1013.18 9403.95 ;
      RECT 998.1 9441.09 999.1 9442.51 ;
      RECT 998.1 9441.145 1013.18 9442.465 ;
      RECT 19150 9497.56 19170 9527.56 ;
      RECT 19150 9529.56 19170 9559.56 ;
      RECT 19150 9617.56 19170 9647.56 ;
      RECT 19150 9649.56 19170 9679.56 ;
      RECT 19150 9737.56 19170 9767.56 ;
      RECT 19150 9769.56 19170 9799.56 ;
      RECT 19150 9857.56 19170 9887.56 ;
      RECT 19150 9889.56 19170 9919.56 ;
      RECT 19158.16 1055.685 19167.9 1056.485 ;
      RECT 19158.16 1088.01 19167.9 1088.81 ;
      RECT 19158.16 1119.19 19167.9 1119.99 ;
      RECT 19158.16 1121.59 19167.9 1122.39 ;
      RECT 19158.16 1123.99 19167.9 1124.79 ;
      RECT 19158.16 1126.39 19167.9 1127.19 ;
      RECT 19158.16 1364.42 19167.75 1365.49 ;
      RECT 19158.16 1367.4 19167.75 1368.47 ;
      RECT 19032.505 1048.035 19032.785 1177.59 ;
      RECT 19031.945 1048.035 19032.225 1201.16 ;
      RECT 19031.385 1046.935 19031.665 1201.4 ;
      RECT 19030.825 1048.035 19031.105 1201.64 ;
      RECT 19030.265 1046.935 19030.545 1201.885 ;
      RECT 19029.705 1048.035 19029.985 1202.125 ;
      RECT 19029.145 1046.935 19029.425 1202.365 ;
      RECT 19028.585 1048.035 19028.865 1202.605 ;
      RECT 19028.025 1048.035 19028.305 1202.845 ;
      RECT 19027.465 1048.035 19027.745 1188.465 ;
      RECT 19026.905 1048.035 19027.185 1188.225 ;
      RECT 19026.345 1048.035 19026.625 1187.985 ;
      RECT 19025.785 1048.035 19026.065 1187.745 ;
      RECT 19025.225 1048.035 19025.505 1187.505 ;
      RECT 19024.665 1048.035 19024.945 1187.265 ;
      RECT 19024.105 1048.035 19024.385 1187.025 ;
      RECT 19023.545 1048.035 19023.825 1186.785 ;
      RECT 19022.985 1048.035 19023.265 1186.545 ;
      RECT 19022.425 1048.035 19022.705 1186.305 ;
      RECT 19021.865 1046.935 19022.145 1186.065 ;
      RECT 19021.305 1048.035 19021.585 1185.825 ;
      RECT 19020.745 1046.935 19021.025 1185.585 ;
      RECT 19020.185 1048.035 19020.465 1185.345 ;
      RECT 19006.185 1046.935 19006.465 1191.465 ;
      RECT 19005.625 1048.035 19005.905 1191.225 ;
      RECT 19005.065 1048.035 19005.345 1190.985 ;
      RECT 19004.505 1048.035 19004.785 1190.745 ;
      RECT 19003.945 1048.035 19004.225 1190.505 ;
      RECT 19003.385 1048.035 19003.665 1190.265 ;
      RECT 19002.825 1048.035 19003.105 1190.025 ;
      RECT 19002.265 1048.035 19002.545 1189.785 ;
      RECT 19001.705 1048.035 19001.985 1189.545 ;
      RECT 19001.145 1046.935 19001.425 1189.305 ;
      RECT 19000.585 1048.035 19000.865 1189.065 ;
      RECT 19000.025 1046.935 19000.305 1188.825 ;
      RECT 18999.465 1048.035 18999.745 1188.585 ;
      RECT 18998.905 1048.035 18999.185 1188.345 ;
      RECT 18998.345 1048.035 18998.625 1188.105 ;
      RECT 18997.785 1048.035 18998.065 1187.865 ;
      RECT 18997.225 1048.035 18997.505 1187.625 ;
      RECT 18996.665 1048.035 18996.945 1187.385 ;
      RECT 18996.105 1048.035 18996.385 1187.145 ;
      RECT 18995.545 1048.035 18995.825 1186.905 ;
      RECT 18994.985 1048.035 18995.265 1186.665 ;
      RECT 18994.425 1048.035 18994.705 1186.425 ;
      RECT 18993.865 1048.035 18994.145 1186.185 ;
      RECT 18954.665 1048.035 18954.945 1193.09 ;
      RECT 18954.105 1048.035 18954.385 1193.33 ;
      RECT 18953.545 1048.035 18953.825 1193.57 ;
      RECT 18952.985 1046.935 18953.265 1193.81 ;
      RECT 18952.425 1048.035 18952.705 1194.05 ;
      RECT 18951.865 1046.935 18952.145 1194.29 ;
      RECT 18951.305 1048.035 18951.585 1194.53 ;
      RECT 18950.745 1048.035 18951.025 1194.77 ;
      RECT 18950.185 1048.035 18950.465 1195.01 ;
      RECT 18949.625 1046.935 18949.905 1195.25 ;
      RECT 18949.065 1048.035 18949.345 1195.49 ;
      RECT 18948.505 1046.935 18948.785 1195.73 ;
      RECT 18947.945 1048.035 18948.225 1195.97 ;
      RECT 18947.385 1046.935 18947.665 1196.21 ;
      RECT 18946.825 1048.035 18947.105 1196.45 ;
      RECT 18946.265 1048.035 18946.545 1196.69 ;
      RECT 18945.705 1048.035 18945.985 1196.69 ;
      RECT 18945.145 1048.035 18945.425 1196.45 ;
      RECT 18944.585 1048.035 18944.865 1196.21 ;
      RECT 18944.025 1048.035 18944.305 1195.97 ;
      RECT 18943.465 1048.035 18943.745 1195.73 ;
      RECT 18942.905 1048.035 18943.185 1195.49 ;
      RECT 18942.345 1048.035 18942.625 1195.25 ;
      RECT 18941.785 1048.035 18942.065 1195.01 ;
      RECT 18941.225 1048.035 18941.505 1194.77 ;
      RECT 18932.265 1048.035 18932.545 1194.285 ;
      RECT 18931.705 1046.935 18931.985 1194.045 ;
      RECT 18931.145 1048.035 18931.425 1193.805 ;
      RECT 18930.585 1046.935 18930.865 1193.565 ;
      RECT 18930.025 1048.035 18930.305 1193.325 ;
      RECT 18929.465 1046.935 18929.745 1193.085 ;
      RECT 18928.905 1048.035 18929.185 1192.845 ;
      RECT 18928.345 1048.035 18928.625 1192.605 ;
      RECT 18927.785 1048.035 18928.065 1192.365 ;
      RECT 18927.225 1048.035 18927.505 1192.125 ;
      RECT 18926.665 1048.035 18926.945 1191.885 ;
      RECT 18926.105 1048.035 18926.385 1191.645 ;
      RECT 18925.545 1048.035 18925.825 1191.405 ;
      RECT 18924.985 1048.035 18925.265 1191.165 ;
      RECT 18922.465 1046.935 18922.745 1192.885 ;
      RECT 18921.905 1048.035 18922.185 1192.645 ;
      RECT 18921.345 1046.935 18921.625 1192.405 ;
      RECT 18920.785 1048.035 18921.065 1192.165 ;
      RECT 18920.225 1048.035 18920.505 1191.925 ;
      RECT 18919.665 1048.035 18919.945 1191.685 ;
      RECT 18919.105 1048.035 18919.385 1191.445 ;
      RECT 18918.545 1048.035 18918.825 1191.205 ;
      RECT 18892.505 1048.035 18892.785 1188.855 ;
      RECT 18891.945 1048.035 18892.225 1189.095 ;
      RECT 18891.385 1048.035 18891.665 1189.335 ;
      RECT 18890.825 1048.035 18891.105 1189.58 ;
      RECT 18890.265 1048.035 18890.545 1189.82 ;
      RECT 18889.705 1048.035 18889.985 1190.06 ;
      RECT 18889.145 1048.035 18889.425 1190.06 ;
      RECT 18888.585 1048.035 18888.865 1189.82 ;
      RECT 18888.025 1048.035 18888.305 1189.58 ;
      RECT 18887.465 1046.935 18887.745 1189.34 ;
      RECT 18886.905 1048.035 18887.185 1189.1 ;
      RECT 18886.345 1046.935 18886.625 1188.86 ;
      RECT 18885.785 1048.035 18886.065 1188.62 ;
      RECT 18885.225 1048.035 18885.505 1188.38 ;
      RECT 18884.665 1048.035 18884.945 1188.14 ;
      RECT 18884.105 1046.935 18884.385 1187.9 ;
      RECT 18883.545 1048.035 18883.825 1187.66 ;
      RECT 18882.985 1046.935 18883.265 1187.42 ;
      RECT 18882.425 1048.035 18882.705 1187.18 ;
      RECT 18881.865 1046.935 18882.145 1186.94 ;
      RECT 18881.305 1048.035 18881.585 1186.7 ;
      RECT 18880.745 1048.035 18881.025 1186.46 ;
      RECT 18880.185 1048.035 18880.465 1186.22 ;
      RECT 18879.625 1048.035 18879.905 1185.98 ;
      RECT 18866.185 1048.035 18866.465 1191.78 ;
      RECT 18865.625 1048.035 18865.905 1191.54 ;
      RECT 18865.065 1048.035 18865.345 1191.3 ;
      RECT 18864.505 1048.035 18864.785 1191.06 ;
      RECT 18863.945 1048.035 18864.225 1190.82 ;
      RECT 18863.385 1048.035 18863.665 1190.58 ;
      RECT 18862.825 1048.035 18863.105 1190.34 ;
      RECT 18862.265 1048.035 18862.545 1190.1 ;
      RECT 18861.705 1046.935 18861.985 1189.86 ;
      RECT 18861.145 1048.035 18861.425 1189.62 ;
      RECT 18860.585 1046.935 18860.865 1189.3 ;
      RECT 18860.025 1048.035 18860.305 1189.14 ;
      RECT 18859.465 1046.935 18859.745 1188.9 ;
      RECT 18858.905 1048.035 18859.185 1188.66 ;
      RECT 18858.345 1048.035 18858.625 1188.42 ;
      RECT 18857.785 1048.035 18858.065 1188.18 ;
      RECT 18857.225 1048.035 18857.505 1187.94 ;
      RECT 18856.665 1048.035 18856.945 1187.7 ;
      RECT 18856.105 1048.035 18856.385 1187.46 ;
      RECT 18855.545 1048.035 18855.825 1187.22 ;
      RECT 18854.985 1048.035 18855.265 1186.98 ;
      RECT 18854.425 1046.935 18854.705 1186.74 ;
      RECT 18853.865 1048.035 18854.145 1186.5 ;
      RECT 18853.305 1046.935 18853.585 1186.26 ;
      RECT 18814.105 1048.035 18814.385 1191.87 ;
      RECT 18813.545 1048.035 18813.825 1192.11 ;
      RECT 18812.985 1048.035 18813.265 1192.35 ;
      RECT 18812.425 1048.035 18812.705 1192.59 ;
      RECT 18811.865 1048.035 18812.145 1192.83 ;
      RECT 18811.305 1048.035 18811.585 1193.07 ;
      RECT 18810.745 1048.035 18811.025 1193.31 ;
      RECT 18810.185 1048.035 18810.465 1193.55 ;
      RECT 18809.625 1048.035 18809.905 1193.79 ;
      RECT 18809.065 1048.035 18809.345 1194.03 ;
      RECT 18808.505 1048.035 18808.785 1194.27 ;
      RECT 18807.945 1048.035 18808.225 1194.51 ;
      RECT 18807.385 1048.035 18807.665 1194.75 ;
      RECT 18806.825 1048.035 18807.105 1194.75 ;
      RECT 18806.265 1046.935 18806.545 1194.51 ;
      RECT 18805.705 1048.035 18805.985 1194.27 ;
      RECT 18805.145 1046.935 18805.425 1194.03 ;
      RECT 18804.585 1048.035 18804.865 1193.79 ;
      RECT 18804.025 1048.035 18804.305 1193.55 ;
      RECT 18803.465 1048.035 18803.745 1193.31 ;
      RECT 18802.905 1046.935 18803.185 1193.045 ;
      RECT 18802.345 1048.035 18802.625 1192.805 ;
      RECT 18801.785 1046.935 18802.065 1192.565 ;
      RECT 18801.225 1048.035 18801.505 1192.325 ;
      RECT 18792.265 1046.935 18792.545 1186.16 ;
      RECT 18791.705 1048.035 18791.985 1186.4 ;
      RECT 18791.145 1048.035 18791.425 1186.64 ;
      RECT 18790.585 1048.035 18790.865 1186.64 ;
      RECT 18790.025 1048.035 18790.305 1186.4 ;
      RECT 18789.465 1048.035 18789.745 1186.16 ;
      RECT 18788.905 1048.035 18789.185 1185.92 ;
      RECT 18788.345 1048.035 18788.625 1185.68 ;
      RECT 18787.785 1048.035 18788.065 1185.44 ;
      RECT 18787.225 1048.035 18787.505 1185.2 ;
      RECT 18786.665 1048.035 18786.945 1184.96 ;
      RECT 18786.105 1048.035 18786.385 1184.72 ;
      RECT 18785.545 1048.035 18785.825 1184.48 ;
      RECT 18784.985 1046.935 18785.265 1184.24 ;
      RECT 18782.465 1048.035 18782.745 1185.96 ;
      RECT 18781.905 1046.935 18782.185 1185.72 ;
      RECT 18781.345 1048.035 18781.625 1185.48 ;
      RECT 18780.785 1046.935 18781.065 1185.24 ;
      RECT 18780.225 1048.035 18780.505 1185 ;
      RECT 18779.665 1048.035 18779.945 1184.76 ;
      RECT 18779.105 1048.035 18779.385 1184.52 ;
      RECT 18753.065 1048.035 18753.345 1187.305 ;
      RECT 18752.505 1048.035 18752.785 1187.545 ;
      RECT 18751.945 1048.035 18752.225 1187.785 ;
      RECT 18751.385 1048.035 18751.665 1188.025 ;
      RECT 18750.825 1048.035 18751.105 1188.265 ;
      RECT 18750.265 1046.935 18750.545 1188.505 ;
      RECT 18749.705 1048.035 18749.985 1188.745 ;
      RECT 18749.145 1046.935 18749.425 1188.985 ;
      RECT 18748.585 1048.035 18748.865 1189.225 ;
      RECT 18748.025 1048.035 18748.305 1189.465 ;
      RECT 18747.465 1048.035 18747.745 1189.705 ;
      RECT 18746.905 1048.035 18747.185 1189.945 ;
      RECT 18746.345 1048.035 18746.625 1190.185 ;
      RECT 18745.785 1048.035 18746.065 1190.425 ;
      RECT 18745.225 1048.035 18745.505 1190.665 ;
      RECT 18744.665 1048.035 18744.945 1190.665 ;
      RECT 18744.105 1048.035 18744.385 1190.425 ;
      RECT 18743.545 1048.035 18743.825 1190.185 ;
      RECT 18742.985 1048.035 18743.265 1189.945 ;
      RECT 18742.425 1048.035 18742.705 1189.7 ;
      RECT 18741.865 1048.035 18742.145 1189.46 ;
      RECT 18741.305 1048.035 18741.585 1189.22 ;
      RECT 18740.745 1046.935 18741.025 1188.98 ;
      RECT 18740.185 1048.035 18740.465 1188.74 ;
      RECT 18726.745 1046.935 18727.025 1186.22 ;
      RECT 18726.185 1048.035 18726.465 1185.98 ;
      RECT 18725.625 1048.035 18725.905 1185.74 ;
      RECT 18725.065 1048.035 18725.345 1185.5 ;
      RECT 18724.505 1046.935 18724.785 1185.26 ;
      RECT 18723.945 1048.035 18724.225 1185.02 ;
      RECT 18723.385 1046.935 18723.665 1184.78 ;
      RECT 18722.825 1048.035 18723.105 1184.54 ;
      RECT 18722.265 1046.935 18722.545 1184.3 ;
      RECT 18721.705 1048.035 18721.985 1184.06 ;
      RECT 18721.145 1048.035 18721.425 1183.82 ;
      RECT 18720.585 1048.035 18720.865 1183.58 ;
      RECT 18720.025 1048.035 18720.305 1183.34 ;
      RECT 18719.465 1048.035 18719.745 1183.1 ;
      RECT 18718.905 1048.035 18719.185 1182.86 ;
      RECT 18718.345 1048.035 18718.625 1182.62 ;
      RECT 18717.785 1048.035 18718.065 1182.38 ;
      RECT 18717.225 1048.035 18717.505 1182.14 ;
      RECT 18716.665 1048.035 18716.945 1181.9 ;
      RECT 18716.105 1048.035 18716.385 1181.66 ;
      RECT 18715.545 1048.035 18715.825 1181.42 ;
      RECT 18714.985 1046.935 18715.265 1181.18 ;
      RECT 18714.425 1048.035 18714.705 1180.94 ;
      RECT 18713.865 1046.935 18714.145 1180.7 ;
      RECT 18674.105 1048.035 18674.385 1191.17 ;
      RECT 18673.545 1046.935 18673.825 1191.41 ;
      RECT 18672.985 1048.035 18673.265 1191.65 ;
      RECT 18672.425 1048.035 18672.705 1191.89 ;
      RECT 18671.865 1048.035 18672.145 1192.13 ;
      RECT 18671.305 1048.035 18671.585 1192.37 ;
      RECT 18670.745 1048.035 18671.025 1192.61 ;
      RECT 18670.185 1048.035 18670.465 1192.855 ;
      RECT 18669.625 1048.035 18669.905 1193.095 ;
      RECT 18669.065 1048.035 18669.345 1193.335 ;
      RECT 18668.505 1046.935 18668.785 1193.575 ;
      RECT 18667.945 1048.035 18668.225 1193.815 ;
      RECT 18667.385 1046.935 18667.665 1194.055 ;
      RECT 18666.825 1048.035 18667.105 1194.295 ;
      RECT 18666.265 1048.035 18666.545 1194.535 ;
      RECT 18665.705 1048.035 18665.985 1194.775 ;
      RECT 18665.145 1048.035 18665.425 1195.015 ;
      RECT 18664.585 1048.035 18664.865 1195.255 ;
      RECT 18664.025 1048.035 18664.305 1195.495 ;
      RECT 18663.465 1048.035 18663.745 1195.735 ;
      RECT 18662.905 1048.035 18663.185 1195.975 ;
      RECT 18662.345 1048.035 18662.625 1196.215 ;
      RECT 18661.785 1048.035 18662.065 1196.455 ;
      RECT 18661.225 1048.035 18661.505 1196.695 ;
      RECT 18652.265 1048.035 18652.545 1192.28 ;
      RECT 18651.705 1048.035 18651.985 1192.04 ;
      RECT 18651.145 1048.035 18651.425 1191.8 ;
      RECT 18650.585 1046.935 18650.865 1191.56 ;
      RECT 18650.025 1048.035 18650.305 1191.32 ;
      RECT 18649.465 1046.935 18649.745 1191.08 ;
      RECT 18648.905 1048.035 18649.185 1190.84 ;
      RECT 18648.345 1048.035 18648.625 1190.6 ;
      RECT 18647.785 1048.035 18648.065 1190.36 ;
      RECT 18647.225 1046.935 18647.505 1190.12 ;
      RECT 18646.665 1048.035 18646.945 1189.88 ;
      RECT 18646.105 1046.935 18646.385 1189.64 ;
      RECT 18645.545 1048.035 18645.825 1189.4 ;
      RECT 18644.985 1046.935 18645.265 1189.16 ;
      RECT 18642.465 1048.035 18642.745 1181.56 ;
      RECT 18641.905 1048.035 18642.185 1181.32 ;
      RECT 18641.345 1048.035 18641.625 1181.08 ;
      RECT 18640.785 1048.035 18641.065 1180.84 ;
      RECT 18640.225 1048.035 18640.505 1180.6 ;
      RECT 18639.665 1048.035 18639.945 1180.36 ;
      RECT 18639.105 1048.035 18639.385 1180.12 ;
      RECT 18613.065 1048.035 18613.345 1193.995 ;
      RECT 18612.505 1048.035 18612.785 1194.235 ;
      RECT 18611.945 1048.035 18612.225 1194.475 ;
      RECT 18611.385 1048.035 18611.665 1194.715 ;
      RECT 18610.825 1048.035 18611.105 1194.955 ;
      RECT 18610.265 1046.935 18610.545 1194.955 ;
      RECT 18609.705 1048.035 18609.985 1194.715 ;
      RECT 18609.145 1046.935 18609.425 1194.47 ;
      RECT 18608.585 1048.035 18608.865 1194.23 ;
      RECT 18608.025 1046.935 18608.305 1193.99 ;
      RECT 18607.465 1048.035 18607.745 1193.75 ;
      RECT 18606.905 1048.035 18607.185 1193.51 ;
      RECT 18606.345 1048.035 18606.625 1193.27 ;
      RECT 18605.785 1048.035 18606.065 1193.03 ;
      RECT 18605.225 1048.035 18605.505 1192.79 ;
      RECT 18604.665 1048.035 18604.945 1192.55 ;
      RECT 18604.105 1048.035 18604.385 1192.31 ;
      RECT 18603.545 1048.035 18603.825 1192.07 ;
      RECT 18602.985 1046.935 18603.265 1191.83 ;
      RECT 18602.425 1048.035 18602.705 1191.59 ;
      RECT 18601.865 1046.935 18602.145 1191.35 ;
      RECT 18601.305 1048.035 18601.585 1191.11 ;
      RECT 18600.745 1048.035 18601.025 1190.87 ;
      RECT 18600.185 1048.035 18600.465 1190.63 ;
      RECT 18586.745 1048.035 18587.025 1194.03 ;
      RECT 18586.185 1048.035 18586.465 1194.27 ;
      RECT 18585.625 1048.035 18585.905 1194.515 ;
      RECT 18585.065 1048.035 18585.345 1194.755 ;
      RECT 18584.505 1048.035 18584.785 1194.995 ;
      RECT 18583.945 1048.035 18584.225 1194.995 ;
      RECT 18583.385 1048.035 18583.665 1194.755 ;
      RECT 18582.825 1048.035 18583.105 1194.515 ;
      RECT 18582.265 1048.035 18582.545 1187.5 ;
      RECT 18581.705 1048.035 18581.985 1187.26 ;
      RECT 18581.145 1048.035 18581.425 1187.02 ;
      RECT 18580.585 1046.935 18580.865 1186.78 ;
      RECT 18580.025 1048.035 18580.305 1186.54 ;
      RECT 18579.465 1046.935 18579.745 1186.3 ;
      RECT 18578.905 1048.035 18579.185 1186.06 ;
      RECT 18578.345 1048.035 18578.625 1185.82 ;
      RECT 18577.785 1048.035 18578.065 1185.58 ;
      RECT 18577.225 1046.935 18577.505 1185.34 ;
      RECT 18576.665 1048.035 18576.945 1185.1 ;
      RECT 18576.105 1046.935 18576.385 1184.86 ;
      RECT 18575.545 1048.035 18575.825 1184.62 ;
      RECT 18574.985 1046.935 18575.265 1184.38 ;
      RECT 18574.425 1048.035 18574.705 1184.14 ;
      RECT 18573.865 1048.035 18574.145 1183.9 ;
      RECT 18533.545 1048.035 18533.825 1192.795 ;
      RECT 18532.985 1048.035 18533.265 1193.035 ;
      RECT 18532.425 1048.035 18532.705 1193.28 ;
      RECT 18531.865 1048.035 18532.145 1193.52 ;
      RECT 18531.305 1048.035 18531.585 1193.76 ;
      RECT 18530.745 1048.035 18531.025 1194 ;
      RECT 18530.185 1048.035 18530.465 1194.24 ;
      RECT 18529.625 1048.035 18529.905 1194.48 ;
      RECT 18529.065 1048.035 18529.345 1194.72 ;
      RECT 18528.505 1048.035 18528.785 1194.96 ;
      RECT 18527.945 1046.935 18528.225 1195.2 ;
      RECT 18527.385 1048.035 18527.665 1195.44 ;
      RECT 18526.825 1046.935 18527.105 1195.68 ;
      RECT 18526.265 1048.035 18526.545 1195.92 ;
      RECT 18525.705 1046.935 18525.985 1196.16 ;
      RECT 18525.145 1048.035 18525.425 1196.16 ;
      RECT 18524.585 1048.035 18524.865 1195.92 ;
      RECT 18524.025 1048.035 18524.305 1195.68 ;
      RECT 18523.465 1048.035 18523.745 1195.44 ;
      RECT 18522.905 1048.035 18523.185 1195.2 ;
      RECT 18522.345 1048.035 18522.625 1194.96 ;
      RECT 18521.785 1048.035 18522.065 1194.72 ;
      RECT 18521.225 1048.035 18521.505 1194.48 ;
      RECT 18512.265 1046.935 18512.545 1194.51 ;
      RECT 18511.705 1048.035 18511.985 1194.75 ;
      RECT 18511.145 1046.935 18511.425 1194.99 ;
      RECT 18510.585 1048.035 18510.865 1195.205 ;
      RECT 18510.025 1048.035 18510.305 1194.78 ;
      RECT 18509.465 1048.035 18509.745 1194.54 ;
      RECT 18508.905 1048.035 18509.185 1194.3 ;
      RECT 18508.345 1048.035 18508.625 1194.06 ;
      RECT 18507.785 1048.035 18508.065 1193.82 ;
      RECT 18507.225 1048.035 18507.505 1193.58 ;
      RECT 18506.665 1048.035 18506.945 1193.34 ;
      RECT 18506.105 1048.035 18506.385 1193.1 ;
      RECT 18505.545 1048.035 18505.825 1192.86 ;
      RECT 18504.985 1048.035 18505.265 1192.62 ;
      RECT 18502.465 1048.035 18502.745 1191.795 ;
      RECT 18501.905 1048.035 18502.185 1191.555 ;
      RECT 18501.345 1048.035 18501.625 1191.315 ;
      RECT 18500.785 1046.935 18501.065 1191.075 ;
      RECT 18500.225 1048.035 18500.505 1190.835 ;
      RECT 18499.665 1046.935 18499.945 1190.595 ;
      RECT 18499.105 1048.035 18499.385 1190.355 ;
      RECT 18498.545 1048.035 18498.825 1190.115 ;
      RECT 18471.945 1048.035 18472.225 1201.16 ;
      RECT 18471.385 1046.935 18471.665 1201.4 ;
      RECT 18470.825 1048.035 18471.105 1201.64 ;
      RECT 18470.265 1046.935 18470.545 1201.885 ;
      RECT 18469.705 1048.035 18469.985 1202.125 ;
      RECT 18469.145 1046.935 18469.425 1202.365 ;
      RECT 18468.585 1048.035 18468.865 1202.605 ;
      RECT 18468.025 1048.035 18468.305 1202.845 ;
      RECT 18467.465 1048.035 18467.745 1188.465 ;
      RECT 18466.905 1048.035 18467.185 1188.225 ;
      RECT 18466.345 1048.035 18466.625 1187.985 ;
      RECT 18465.785 1048.035 18466.065 1187.745 ;
      RECT 18465.225 1048.035 18465.505 1187.505 ;
      RECT 18464.665 1048.035 18464.945 1187.265 ;
      RECT 18464.105 1048.035 18464.385 1187.025 ;
      RECT 18463.545 1048.035 18463.825 1186.785 ;
      RECT 18462.985 1048.035 18463.265 1186.545 ;
      RECT 18462.425 1048.035 18462.705 1186.305 ;
      RECT 18461.865 1046.935 18462.145 1186.065 ;
      RECT 18461.305 1048.035 18461.585 1185.825 ;
      RECT 18460.745 1046.935 18461.025 1185.585 ;
      RECT 18460.185 1048.035 18460.465 1185.345 ;
      RECT 18446.185 1046.935 18446.465 1191.465 ;
      RECT 18445.625 1048.035 18445.905 1191.225 ;
      RECT 18445.065 1048.035 18445.345 1190.985 ;
      RECT 18444.505 1048.035 18444.785 1190.745 ;
      RECT 18443.945 1048.035 18444.225 1190.505 ;
      RECT 18443.385 1048.035 18443.665 1190.265 ;
      RECT 18442.825 1048.035 18443.105 1190.025 ;
      RECT 18442.265 1048.035 18442.545 1189.785 ;
      RECT 18441.705 1048.035 18441.985 1189.545 ;
      RECT 18441.145 1046.935 18441.425 1189.305 ;
      RECT 18440.585 1048.035 18440.865 1189.065 ;
      RECT 18440.025 1046.935 18440.305 1188.825 ;
      RECT 18439.465 1048.035 18439.745 1188.585 ;
      RECT 18438.905 1048.035 18439.185 1188.345 ;
      RECT 18438.345 1048.035 18438.625 1188.105 ;
      RECT 18437.785 1048.035 18438.065 1187.865 ;
      RECT 18437.225 1048.035 18437.505 1187.625 ;
      RECT 18436.665 1048.035 18436.945 1187.385 ;
      RECT 18436.105 1048.035 18436.385 1187.145 ;
      RECT 18435.545 1048.035 18435.825 1186.905 ;
      RECT 18434.985 1048.035 18435.265 1186.665 ;
      RECT 18434.425 1048.035 18434.705 1186.425 ;
      RECT 18433.865 1048.035 18434.145 1186.185 ;
      RECT 18394.665 1048.035 18394.945 1193.09 ;
      RECT 18394.105 1048.035 18394.385 1193.33 ;
      RECT 18393.545 1048.035 18393.825 1193.57 ;
      RECT 18392.985 1046.935 18393.265 1193.81 ;
      RECT 18392.425 1048.035 18392.705 1194.05 ;
      RECT 18391.865 1046.935 18392.145 1194.29 ;
      RECT 18391.305 1048.035 18391.585 1194.53 ;
      RECT 18390.745 1048.035 18391.025 1194.77 ;
      RECT 18390.185 1048.035 18390.465 1195.01 ;
      RECT 18389.625 1046.935 18389.905 1195.25 ;
      RECT 18389.065 1048.035 18389.345 1195.49 ;
      RECT 18388.505 1046.935 18388.785 1195.73 ;
      RECT 18387.945 1048.035 18388.225 1195.97 ;
      RECT 18387.385 1046.935 18387.665 1196.21 ;
      RECT 18386.825 1048.035 18387.105 1196.45 ;
      RECT 18386.265 1048.035 18386.545 1196.69 ;
      RECT 18385.705 1048.035 18385.985 1196.69 ;
      RECT 18385.145 1048.035 18385.425 1196.45 ;
      RECT 18384.585 1048.035 18384.865 1196.21 ;
      RECT 18384.025 1048.035 18384.305 1195.97 ;
      RECT 18383.465 1048.035 18383.745 1195.73 ;
      RECT 18382.905 1048.035 18383.185 1195.49 ;
      RECT 18382.345 1048.035 18382.625 1195.25 ;
      RECT 18381.785 1048.035 18382.065 1195.01 ;
      RECT 18381.225 1048.035 18381.505 1194.77 ;
      RECT 18372.265 1048.035 18372.545 1194.285 ;
      RECT 18371.705 1046.935 18371.985 1194.045 ;
      RECT 18371.145 1048.035 18371.425 1193.805 ;
      RECT 18370.585 1046.935 18370.865 1193.565 ;
      RECT 18370.025 1048.035 18370.305 1193.325 ;
      RECT 18369.465 1046.935 18369.745 1193.085 ;
      RECT 18368.905 1048.035 18369.185 1192.845 ;
      RECT 18368.345 1048.035 18368.625 1192.605 ;
      RECT 18367.785 1048.035 18368.065 1192.365 ;
      RECT 18367.225 1048.035 18367.505 1192.125 ;
      RECT 18366.665 1048.035 18366.945 1191.885 ;
      RECT 18366.105 1048.035 18366.385 1191.645 ;
      RECT 18365.545 1048.035 18365.825 1191.405 ;
      RECT 18364.985 1048.035 18365.265 1191.165 ;
      RECT 18362.465 1046.935 18362.745 1192.885 ;
      RECT 18361.905 1048.035 18362.185 1192.645 ;
      RECT 18361.345 1046.935 18361.625 1192.405 ;
      RECT 18360.785 1048.035 18361.065 1192.165 ;
      RECT 18360.225 1048.035 18360.505 1191.925 ;
      RECT 18359.665 1048.035 18359.945 1191.685 ;
      RECT 18359.105 1048.035 18359.385 1191.445 ;
      RECT 18358.545 1048.035 18358.825 1191.205 ;
      RECT 18332.505 1048.035 18332.785 1188.855 ;
      RECT 18331.945 1048.035 18332.225 1189.095 ;
      RECT 18331.385 1048.035 18331.665 1189.335 ;
      RECT 18330.825 1048.035 18331.105 1189.58 ;
      RECT 18330.265 1048.035 18330.545 1189.82 ;
      RECT 18329.705 1048.035 18329.985 1190.06 ;
      RECT 18329.145 1048.035 18329.425 1190.06 ;
      RECT 18328.585 1048.035 18328.865 1189.82 ;
      RECT 18328.025 1048.035 18328.305 1189.58 ;
      RECT 18327.465 1046.935 18327.745 1189.34 ;
      RECT 18326.905 1048.035 18327.185 1189.1 ;
      RECT 18326.345 1046.935 18326.625 1188.86 ;
      RECT 18325.785 1048.035 18326.065 1188.62 ;
      RECT 18325.225 1048.035 18325.505 1188.38 ;
      RECT 18324.665 1048.035 18324.945 1188.14 ;
      RECT 18324.105 1046.935 18324.385 1187.9 ;
      RECT 18323.545 1048.035 18323.825 1187.66 ;
      RECT 18322.985 1046.935 18323.265 1187.42 ;
      RECT 18322.425 1048.035 18322.705 1187.18 ;
      RECT 18321.865 1046.935 18322.145 1186.94 ;
      RECT 18321.305 1048.035 18321.585 1186.7 ;
      RECT 18320.745 1048.035 18321.025 1186.46 ;
      RECT 18320.185 1048.035 18320.465 1186.22 ;
      RECT 18319.625 1048.035 18319.905 1185.98 ;
      RECT 18306.185 1048.035 18306.465 1191.78 ;
      RECT 18305.625 1048.035 18305.905 1191.54 ;
      RECT 18305.065 1048.035 18305.345 1191.3 ;
      RECT 18304.505 1048.035 18304.785 1191.06 ;
      RECT 18303.945 1048.035 18304.225 1190.82 ;
      RECT 18303.385 1048.035 18303.665 1190.58 ;
      RECT 18302.825 1048.035 18303.105 1190.34 ;
      RECT 18302.265 1048.035 18302.545 1190.1 ;
      RECT 18301.705 1046.935 18301.985 1189.86 ;
      RECT 18301.145 1048.035 18301.425 1189.62 ;
      RECT 18300.585 1046.935 18300.865 1189.3 ;
      RECT 18300.025 1048.035 18300.305 1189.14 ;
      RECT 18299.465 1046.935 18299.745 1188.9 ;
      RECT 18298.905 1048.035 18299.185 1188.66 ;
      RECT 18298.345 1048.035 18298.625 1188.42 ;
      RECT 18297.785 1048.035 18298.065 1188.18 ;
      RECT 18297.225 1048.035 18297.505 1187.94 ;
      RECT 18296.665 1048.035 18296.945 1187.7 ;
      RECT 18296.105 1048.035 18296.385 1187.46 ;
      RECT 18295.545 1048.035 18295.825 1187.22 ;
      RECT 18294.985 1048.035 18295.265 1186.98 ;
      RECT 18294.425 1046.935 18294.705 1186.74 ;
      RECT 18293.865 1048.035 18294.145 1186.5 ;
      RECT 18293.305 1046.935 18293.585 1186.26 ;
      RECT 18254.105 1048.035 18254.385 1191.87 ;
      RECT 18253.545 1048.035 18253.825 1192.11 ;
      RECT 18252.985 1048.035 18253.265 1192.35 ;
      RECT 18252.425 1048.035 18252.705 1192.59 ;
      RECT 18251.865 1048.035 18252.145 1192.83 ;
      RECT 18251.305 1048.035 18251.585 1193.07 ;
      RECT 18250.745 1048.035 18251.025 1193.31 ;
      RECT 18250.185 1048.035 18250.465 1193.55 ;
      RECT 18249.625 1048.035 18249.905 1193.79 ;
      RECT 18249.065 1048.035 18249.345 1194.03 ;
      RECT 18248.505 1048.035 18248.785 1194.27 ;
      RECT 18247.945 1048.035 18248.225 1194.51 ;
      RECT 18247.385 1048.035 18247.665 1194.75 ;
      RECT 18246.825 1048.035 18247.105 1194.75 ;
      RECT 18246.265 1046.935 18246.545 1194.51 ;
      RECT 18245.705 1048.035 18245.985 1194.27 ;
      RECT 18245.145 1046.935 18245.425 1194.03 ;
      RECT 18244.585 1048.035 18244.865 1193.79 ;
      RECT 18244.025 1048.035 18244.305 1193.55 ;
      RECT 18243.465 1048.035 18243.745 1193.31 ;
      RECT 18242.905 1046.935 18243.185 1193.045 ;
      RECT 18242.345 1048.035 18242.625 1192.805 ;
      RECT 18241.785 1046.935 18242.065 1192.565 ;
      RECT 18241.225 1048.035 18241.505 1192.325 ;
      RECT 18232.265 1046.935 18232.545 1186.16 ;
      RECT 18231.705 1048.035 18231.985 1186.4 ;
      RECT 18231.145 1048.035 18231.425 1186.64 ;
      RECT 18230.585 1048.035 18230.865 1186.64 ;
      RECT 18230.025 1048.035 18230.305 1186.4 ;
      RECT 18229.465 1048.035 18229.745 1186.16 ;
      RECT 18228.905 1048.035 18229.185 1185.92 ;
      RECT 18228.345 1048.035 18228.625 1185.68 ;
      RECT 18227.785 1048.035 18228.065 1185.44 ;
      RECT 18227.225 1048.035 18227.505 1185.2 ;
      RECT 18226.665 1048.035 18226.945 1184.96 ;
      RECT 18226.105 1048.035 18226.385 1184.72 ;
      RECT 18225.545 1048.035 18225.825 1184.48 ;
      RECT 18224.985 1046.935 18225.265 1184.24 ;
      RECT 18222.465 1048.035 18222.745 1185.96 ;
      RECT 18221.905 1046.935 18222.185 1185.72 ;
      RECT 18221.345 1048.035 18221.625 1185.48 ;
      RECT 18220.785 1046.935 18221.065 1185.24 ;
      RECT 18220.225 1048.035 18220.505 1185 ;
      RECT 18219.665 1048.035 18219.945 1184.76 ;
      RECT 18219.105 1048.035 18219.385 1184.52 ;
      RECT 18193.065 1048.035 18193.345 1187.305 ;
      RECT 18192.505 1048.035 18192.785 1187.545 ;
      RECT 18191.945 1048.035 18192.225 1187.785 ;
      RECT 18191.385 1048.035 18191.665 1188.025 ;
      RECT 18190.825 1048.035 18191.105 1188.265 ;
      RECT 18190.265 1046.935 18190.545 1188.505 ;
      RECT 18189.705 1048.035 18189.985 1188.745 ;
      RECT 18189.145 1046.935 18189.425 1188.985 ;
      RECT 18188.585 1048.035 18188.865 1189.225 ;
      RECT 18188.025 1048.035 18188.305 1189.465 ;
      RECT 18187.465 1048.035 18187.745 1189.705 ;
      RECT 18186.905 1048.035 18187.185 1189.945 ;
      RECT 18186.345 1048.035 18186.625 1190.185 ;
      RECT 18185.785 1048.035 18186.065 1190.425 ;
      RECT 18185.225 1048.035 18185.505 1190.665 ;
      RECT 18184.665 1048.035 18184.945 1190.665 ;
      RECT 18184.105 1048.035 18184.385 1190.425 ;
      RECT 18183.545 1048.035 18183.825 1190.185 ;
      RECT 18182.985 1048.035 18183.265 1189.945 ;
      RECT 18182.425 1048.035 18182.705 1189.7 ;
      RECT 18181.865 1048.035 18182.145 1189.46 ;
      RECT 18181.305 1048.035 18181.585 1189.22 ;
      RECT 18180.745 1046.935 18181.025 1188.98 ;
      RECT 18180.185 1048.035 18180.465 1188.74 ;
      RECT 18166.745 1046.935 18167.025 1186.22 ;
      RECT 18166.185 1048.035 18166.465 1185.98 ;
      RECT 18165.625 1048.035 18165.905 1185.74 ;
      RECT 18165.065 1048.035 18165.345 1185.5 ;
      RECT 18164.505 1046.935 18164.785 1185.26 ;
      RECT 18163.945 1048.035 18164.225 1185.02 ;
      RECT 18163.385 1046.935 18163.665 1184.78 ;
      RECT 18162.825 1048.035 18163.105 1184.54 ;
      RECT 18162.265 1046.935 18162.545 1184.3 ;
      RECT 18161.705 1048.035 18161.985 1184.06 ;
      RECT 18161.145 1048.035 18161.425 1183.82 ;
      RECT 18160.585 1048.035 18160.865 1183.58 ;
      RECT 18160.025 1048.035 18160.305 1183.34 ;
      RECT 18159.465 1048.035 18159.745 1183.1 ;
      RECT 18158.905 1048.035 18159.185 1182.86 ;
      RECT 18158.345 1048.035 18158.625 1182.62 ;
      RECT 18157.785 1048.035 18158.065 1182.38 ;
      RECT 18157.225 1048.035 18157.505 1182.14 ;
      RECT 18156.665 1048.035 18156.945 1181.9 ;
      RECT 18156.105 1048.035 18156.385 1181.66 ;
      RECT 18155.545 1048.035 18155.825 1181.42 ;
      RECT 18154.985 1046.935 18155.265 1181.18 ;
      RECT 18154.425 1048.035 18154.705 1180.94 ;
      RECT 18153.865 1046.935 18154.145 1180.7 ;
      RECT 18114.105 1048.035 18114.385 1191.17 ;
      RECT 18113.545 1046.935 18113.825 1191.41 ;
      RECT 18112.985 1048.035 18113.265 1191.65 ;
      RECT 18112.425 1048.035 18112.705 1191.89 ;
      RECT 18111.865 1048.035 18112.145 1192.13 ;
      RECT 18111.305 1048.035 18111.585 1192.37 ;
      RECT 18110.745 1048.035 18111.025 1192.61 ;
      RECT 18110.185 1048.035 18110.465 1192.855 ;
      RECT 18109.625 1048.035 18109.905 1193.095 ;
      RECT 18109.065 1048.035 18109.345 1193.335 ;
      RECT 18108.505 1046.935 18108.785 1193.575 ;
      RECT 18107.945 1048.035 18108.225 1193.815 ;
      RECT 18107.385 1046.935 18107.665 1194.055 ;
      RECT 18106.825 1048.035 18107.105 1194.295 ;
      RECT 18106.265 1048.035 18106.545 1194.535 ;
      RECT 18105.705 1048.035 18105.985 1194.775 ;
      RECT 18105.145 1048.035 18105.425 1195.015 ;
      RECT 18104.585 1048.035 18104.865 1195.255 ;
      RECT 18104.025 1048.035 18104.305 1195.495 ;
      RECT 18103.465 1048.035 18103.745 1195.735 ;
      RECT 18102.905 1048.035 18103.185 1195.975 ;
      RECT 18102.345 1048.035 18102.625 1196.215 ;
      RECT 18101.785 1048.035 18102.065 1196.455 ;
      RECT 18101.225 1048.035 18101.505 1196.695 ;
      RECT 18092.265 1048.035 18092.545 1192.28 ;
      RECT 18091.705 1048.035 18091.985 1192.04 ;
      RECT 18091.145 1048.035 18091.425 1191.8 ;
      RECT 18090.585 1046.935 18090.865 1191.56 ;
      RECT 18090.025 1048.035 18090.305 1191.32 ;
      RECT 18089.465 1046.935 18089.745 1191.08 ;
      RECT 18088.905 1048.035 18089.185 1190.84 ;
      RECT 18088.345 1048.035 18088.625 1190.6 ;
      RECT 18087.785 1048.035 18088.065 1190.36 ;
      RECT 18087.225 1046.935 18087.505 1190.12 ;
      RECT 18086.665 1048.035 18086.945 1189.88 ;
      RECT 18086.105 1046.935 18086.385 1189.64 ;
      RECT 18085.545 1048.035 18085.825 1189.4 ;
      RECT 18084.985 1046.935 18085.265 1189.16 ;
      RECT 18082.465 1048.035 18082.745 1181.56 ;
      RECT 18081.905 1048.035 18082.185 1181.32 ;
      RECT 18081.345 1048.035 18081.625 1181.08 ;
      RECT 18080.785 1048.035 18081.065 1180.84 ;
      RECT 18080.225 1048.035 18080.505 1180.6 ;
      RECT 18079.665 1048.035 18079.945 1180.36 ;
      RECT 18079.105 1048.035 18079.385 1180.12 ;
      RECT 18053.065 1048.035 18053.345 1193.995 ;
      RECT 18052.505 1048.035 18052.785 1194.235 ;
      RECT 18051.945 1048.035 18052.225 1194.475 ;
      RECT 18051.385 1048.035 18051.665 1194.715 ;
      RECT 18050.825 1048.035 18051.105 1194.955 ;
      RECT 18050.265 1046.935 18050.545 1194.955 ;
      RECT 18049.705 1048.035 18049.985 1194.715 ;
      RECT 18049.145 1046.935 18049.425 1194.47 ;
      RECT 18048.585 1048.035 18048.865 1194.23 ;
      RECT 18048.025 1046.935 18048.305 1193.99 ;
      RECT 18047.465 1048.035 18047.745 1193.75 ;
      RECT 18046.905 1048.035 18047.185 1193.51 ;
      RECT 18046.345 1048.035 18046.625 1193.27 ;
      RECT 18045.785 1048.035 18046.065 1193.03 ;
      RECT 18045.225 1048.035 18045.505 1192.79 ;
      RECT 18044.665 1048.035 18044.945 1192.55 ;
      RECT 18044.105 1048.035 18044.385 1192.31 ;
      RECT 18043.545 1048.035 18043.825 1192.07 ;
      RECT 18042.985 1046.935 18043.265 1191.83 ;
      RECT 18042.425 1048.035 18042.705 1191.59 ;
      RECT 18041.865 1046.935 18042.145 1191.35 ;
      RECT 18041.305 1048.035 18041.585 1191.11 ;
      RECT 18040.745 1048.035 18041.025 1190.87 ;
      RECT 18040.185 1048.035 18040.465 1190.63 ;
      RECT 18026.745 1048.035 18027.025 1194.03 ;
      RECT 18026.185 1048.035 18026.465 1194.27 ;
      RECT 18025.625 1048.035 18025.905 1194.515 ;
      RECT 18025.065 1048.035 18025.345 1194.755 ;
      RECT 18024.505 1048.035 18024.785 1194.995 ;
      RECT 18023.945 1048.035 18024.225 1194.995 ;
      RECT 18023.385 1048.035 18023.665 1194.755 ;
      RECT 18022.825 1048.035 18023.105 1194.515 ;
      RECT 18022.265 1048.035 18022.545 1187.5 ;
      RECT 18021.705 1048.035 18021.985 1187.26 ;
      RECT 18021.145 1048.035 18021.425 1187.02 ;
      RECT 18020.585 1046.935 18020.865 1186.78 ;
      RECT 18020.025 1048.035 18020.305 1186.54 ;
      RECT 18019.465 1046.935 18019.745 1186.3 ;
      RECT 18018.905 1048.035 18019.185 1186.06 ;
      RECT 18018.345 1048.035 18018.625 1185.82 ;
      RECT 18017.785 1048.035 18018.065 1185.58 ;
      RECT 18017.225 1046.935 18017.505 1185.34 ;
      RECT 18016.665 1048.035 18016.945 1185.1 ;
      RECT 18016.105 1046.935 18016.385 1184.86 ;
      RECT 18015.545 1048.035 18015.825 1184.62 ;
      RECT 18014.985 1046.935 18015.265 1184.38 ;
      RECT 18014.425 1048.035 18014.705 1184.14 ;
      RECT 18013.865 1048.035 18014.145 1183.9 ;
      RECT 17973.545 1048.035 17973.825 1192.795 ;
      RECT 17972.985 1048.035 17973.265 1193.035 ;
      RECT 17972.425 1048.035 17972.705 1193.28 ;
      RECT 17971.865 1048.035 17972.145 1193.52 ;
      RECT 17971.305 1048.035 17971.585 1193.76 ;
      RECT 17970.745 1048.035 17971.025 1194 ;
      RECT 17970.185 1048.035 17970.465 1194.24 ;
      RECT 17969.625 1048.035 17969.905 1194.48 ;
      RECT 17969.065 1048.035 17969.345 1194.72 ;
      RECT 17968.505 1048.035 17968.785 1194.96 ;
      RECT 17967.945 1046.935 17968.225 1195.2 ;
      RECT 17967.385 1048.035 17967.665 1195.44 ;
      RECT 17966.825 1046.935 17967.105 1195.68 ;
      RECT 17966.265 1048.035 17966.545 1195.92 ;
      RECT 17965.705 1046.935 17965.985 1196.16 ;
      RECT 17965.145 1048.035 17965.425 1196.16 ;
      RECT 17964.585 1048.035 17964.865 1195.92 ;
      RECT 17964.025 1048.035 17964.305 1195.68 ;
      RECT 17963.465 1048.035 17963.745 1195.44 ;
      RECT 17962.905 1048.035 17963.185 1195.2 ;
      RECT 17962.345 1048.035 17962.625 1194.96 ;
      RECT 17961.785 1048.035 17962.065 1194.72 ;
      RECT 17961.225 1048.035 17961.505 1194.48 ;
      RECT 17952.265 1046.935 17952.545 1194.51 ;
      RECT 17951.705 1048.035 17951.985 1194.75 ;
      RECT 17951.145 1046.935 17951.425 1194.99 ;
      RECT 17950.585 1048.035 17950.865 1195.205 ;
      RECT 17950.025 1048.035 17950.305 1194.78 ;
      RECT 17949.465 1048.035 17949.745 1194.54 ;
      RECT 17948.905 1048.035 17949.185 1194.3 ;
      RECT 17948.345 1048.035 17948.625 1194.06 ;
      RECT 17947.785 1048.035 17948.065 1193.82 ;
      RECT 17947.225 1048.035 17947.505 1193.58 ;
      RECT 17946.665 1048.035 17946.945 1193.34 ;
      RECT 17946.105 1048.035 17946.385 1193.1 ;
      RECT 17945.545 1048.035 17945.825 1192.86 ;
      RECT 17944.985 1048.035 17945.265 1192.62 ;
      RECT 17942.465 1048.035 17942.745 1191.795 ;
      RECT 17941.905 1048.035 17942.185 1191.555 ;
      RECT 17941.345 1048.035 17941.625 1191.315 ;
      RECT 17940.785 1046.935 17941.065 1191.075 ;
      RECT 17940.225 1048.035 17940.505 1190.835 ;
      RECT 17939.665 1046.935 17939.945 1190.595 ;
      RECT 17939.105 1048.035 17939.385 1190.355 ;
      RECT 17938.545 1048.035 17938.825 1190.115 ;
      RECT 17911.945 1048.035 17912.225 1201.16 ;
      RECT 17911.385 1046.935 17911.665 1201.4 ;
      RECT 17910.825 1048.035 17911.105 1201.64 ;
      RECT 17910.265 1046.935 17910.545 1201.885 ;
      RECT 17909.705 1048.035 17909.985 1202.125 ;
      RECT 17909.145 1046.935 17909.425 1202.365 ;
      RECT 17908.585 1048.035 17908.865 1202.605 ;
      RECT 17908.025 1048.035 17908.305 1202.845 ;
      RECT 17907.465 1048.035 17907.745 1188.465 ;
      RECT 17906.905 1048.035 17907.185 1188.225 ;
      RECT 17906.345 1048.035 17906.625 1187.985 ;
      RECT 17905.785 1048.035 17906.065 1187.745 ;
      RECT 17905.225 1048.035 17905.505 1187.505 ;
      RECT 17904.665 1048.035 17904.945 1187.265 ;
      RECT 17904.105 1048.035 17904.385 1187.025 ;
      RECT 17903.545 1048.035 17903.825 1186.785 ;
      RECT 17902.985 1048.035 17903.265 1186.545 ;
      RECT 17902.425 1048.035 17902.705 1186.305 ;
      RECT 17901.865 1046.935 17902.145 1186.065 ;
      RECT 17901.305 1048.035 17901.585 1185.825 ;
      RECT 17900.745 1046.935 17901.025 1185.585 ;
      RECT 17900.185 1048.035 17900.465 1185.345 ;
      RECT 17886.185 1046.935 17886.465 1191.465 ;
      RECT 17885.625 1048.035 17885.905 1191.225 ;
      RECT 17885.065 1048.035 17885.345 1190.985 ;
      RECT 17884.505 1048.035 17884.785 1190.745 ;
      RECT 17883.945 1048.035 17884.225 1190.505 ;
      RECT 17883.385 1048.035 17883.665 1190.265 ;
      RECT 17882.825 1048.035 17883.105 1190.025 ;
      RECT 17882.265 1048.035 17882.545 1189.785 ;
      RECT 17881.705 1048.035 17881.985 1189.545 ;
      RECT 17881.145 1046.935 17881.425 1189.305 ;
      RECT 17880.585 1048.035 17880.865 1189.065 ;
      RECT 17880.025 1046.935 17880.305 1188.825 ;
      RECT 17879.465 1048.035 17879.745 1188.585 ;
      RECT 17878.905 1048.035 17879.185 1188.345 ;
      RECT 17878.345 1048.035 17878.625 1188.105 ;
      RECT 17877.785 1048.035 17878.065 1187.865 ;
      RECT 17877.225 1048.035 17877.505 1187.625 ;
      RECT 17876.665 1048.035 17876.945 1187.385 ;
      RECT 17876.105 1048.035 17876.385 1187.145 ;
      RECT 17875.545 1048.035 17875.825 1186.905 ;
      RECT 17874.985 1048.035 17875.265 1186.665 ;
      RECT 17874.425 1048.035 17874.705 1186.425 ;
      RECT 17873.865 1048.035 17874.145 1186.185 ;
      RECT 17834.665 1048.035 17834.945 1193.09 ;
      RECT 17834.105 1048.035 17834.385 1193.33 ;
      RECT 17833.545 1048.035 17833.825 1193.57 ;
      RECT 17832.985 1046.935 17833.265 1193.81 ;
      RECT 17832.425 1048.035 17832.705 1194.05 ;
      RECT 17831.865 1046.935 17832.145 1194.29 ;
      RECT 17831.305 1048.035 17831.585 1194.53 ;
      RECT 17830.745 1048.035 17831.025 1194.77 ;
      RECT 17830.185 1048.035 17830.465 1195.01 ;
      RECT 17829.625 1046.935 17829.905 1195.25 ;
      RECT 17829.065 1048.035 17829.345 1195.49 ;
      RECT 17828.505 1046.935 17828.785 1195.73 ;
      RECT 17827.945 1048.035 17828.225 1195.97 ;
      RECT 17827.385 1046.935 17827.665 1196.21 ;
      RECT 17826.825 1048.035 17827.105 1196.45 ;
      RECT 17826.265 1048.035 17826.545 1196.69 ;
      RECT 17825.705 1048.035 17825.985 1196.69 ;
      RECT 17825.145 1048.035 17825.425 1196.45 ;
      RECT 17824.585 1048.035 17824.865 1196.21 ;
      RECT 17824.025 1048.035 17824.305 1195.97 ;
      RECT 17823.465 1048.035 17823.745 1195.73 ;
      RECT 17822.905 1048.035 17823.185 1195.49 ;
      RECT 17822.345 1048.035 17822.625 1195.25 ;
      RECT 17821.785 1048.035 17822.065 1195.01 ;
      RECT 17821.225 1048.035 17821.505 1194.77 ;
      RECT 17812.265 1048.035 17812.545 1194.285 ;
      RECT 17811.705 1046.935 17811.985 1194.045 ;
      RECT 17811.145 1048.035 17811.425 1193.805 ;
      RECT 17810.585 1046.935 17810.865 1193.565 ;
      RECT 17810.025 1048.035 17810.305 1193.325 ;
      RECT 17809.465 1046.935 17809.745 1193.085 ;
      RECT 17808.905 1048.035 17809.185 1192.845 ;
      RECT 17808.345 1048.035 17808.625 1192.605 ;
      RECT 17807.785 1048.035 17808.065 1192.365 ;
      RECT 17807.225 1048.035 17807.505 1192.125 ;
      RECT 17806.665 1048.035 17806.945 1191.885 ;
      RECT 17806.105 1048.035 17806.385 1191.645 ;
      RECT 17805.545 1048.035 17805.825 1191.405 ;
      RECT 17804.985 1048.035 17805.265 1191.165 ;
      RECT 17802.465 1046.935 17802.745 1192.885 ;
      RECT 17801.905 1048.035 17802.185 1192.645 ;
      RECT 17801.345 1046.935 17801.625 1192.405 ;
      RECT 17800.785 1048.035 17801.065 1192.165 ;
      RECT 17800.225 1048.035 17800.505 1191.925 ;
      RECT 17799.665 1048.035 17799.945 1191.685 ;
      RECT 17799.105 1048.035 17799.385 1191.445 ;
      RECT 17798.545 1048.035 17798.825 1191.205 ;
      RECT 17772.505 1048.035 17772.785 1188.855 ;
      RECT 17771.945 1048.035 17772.225 1189.095 ;
      RECT 17771.385 1048.035 17771.665 1189.335 ;
      RECT 17770.825 1048.035 17771.105 1189.58 ;
      RECT 17770.265 1048.035 17770.545 1189.82 ;
      RECT 17769.705 1048.035 17769.985 1190.06 ;
      RECT 17769.145 1048.035 17769.425 1190.06 ;
      RECT 17768.585 1048.035 17768.865 1189.82 ;
      RECT 17768.025 1048.035 17768.305 1189.58 ;
      RECT 17767.465 1046.935 17767.745 1189.34 ;
      RECT 17766.905 1048.035 17767.185 1189.1 ;
      RECT 17766.345 1046.935 17766.625 1188.86 ;
      RECT 17765.785 1048.035 17766.065 1188.62 ;
      RECT 17765.225 1048.035 17765.505 1188.38 ;
      RECT 17764.665 1048.035 17764.945 1188.14 ;
      RECT 17764.105 1046.935 17764.385 1187.9 ;
      RECT 17763.545 1048.035 17763.825 1187.66 ;
      RECT 17762.985 1046.935 17763.265 1187.42 ;
      RECT 17762.425 1048.035 17762.705 1187.18 ;
      RECT 17761.865 1046.935 17762.145 1186.94 ;
      RECT 17761.305 1048.035 17761.585 1186.7 ;
      RECT 17760.745 1048.035 17761.025 1186.46 ;
      RECT 17760.185 1048.035 17760.465 1186.22 ;
      RECT 17759.625 1048.035 17759.905 1185.98 ;
      RECT 17746.185 1048.035 17746.465 1191.78 ;
      RECT 17745.625 1048.035 17745.905 1191.54 ;
      RECT 17745.065 1048.035 17745.345 1191.3 ;
      RECT 17744.505 1048.035 17744.785 1191.06 ;
      RECT 17743.945 1048.035 17744.225 1190.82 ;
      RECT 17743.385 1048.035 17743.665 1190.58 ;
      RECT 17742.825 1048.035 17743.105 1190.34 ;
      RECT 17742.265 1048.035 17742.545 1190.1 ;
      RECT 17741.705 1046.935 17741.985 1189.86 ;
      RECT 17741.145 1048.035 17741.425 1189.62 ;
      RECT 17740.585 1046.935 17740.865 1189.3 ;
      RECT 17740.025 1048.035 17740.305 1189.14 ;
      RECT 17739.465 1046.935 17739.745 1188.9 ;
      RECT 17738.905 1048.035 17739.185 1188.66 ;
      RECT 17738.345 1048.035 17738.625 1188.42 ;
      RECT 17737.785 1048.035 17738.065 1188.18 ;
      RECT 17737.225 1048.035 17737.505 1187.94 ;
      RECT 17736.665 1048.035 17736.945 1187.7 ;
      RECT 17736.105 1048.035 17736.385 1187.46 ;
      RECT 17735.545 1048.035 17735.825 1187.22 ;
      RECT 17734.985 1048.035 17735.265 1186.98 ;
      RECT 17734.425 1046.935 17734.705 1186.74 ;
      RECT 17733.865 1048.035 17734.145 1186.5 ;
      RECT 17733.305 1046.935 17733.585 1186.26 ;
      RECT 17694.105 1048.035 17694.385 1191.87 ;
      RECT 17693.545 1048.035 17693.825 1192.11 ;
      RECT 17692.985 1048.035 17693.265 1192.35 ;
      RECT 17692.425 1048.035 17692.705 1192.59 ;
      RECT 17691.865 1048.035 17692.145 1192.83 ;
      RECT 17691.305 1048.035 17691.585 1193.07 ;
      RECT 17690.745 1048.035 17691.025 1193.31 ;
      RECT 17690.185 1048.035 17690.465 1193.55 ;
      RECT 17689.625 1048.035 17689.905 1193.79 ;
      RECT 17689.065 1048.035 17689.345 1194.03 ;
      RECT 17688.505 1048.035 17688.785 1194.27 ;
      RECT 17687.945 1048.035 17688.225 1194.51 ;
      RECT 17687.385 1048.035 17687.665 1194.75 ;
      RECT 17686.825 1048.035 17687.105 1194.75 ;
      RECT 17686.265 1046.935 17686.545 1194.51 ;
      RECT 17685.705 1048.035 17685.985 1194.27 ;
      RECT 17685.145 1046.935 17685.425 1194.03 ;
      RECT 17684.585 1048.035 17684.865 1193.79 ;
      RECT 17684.025 1048.035 17684.305 1193.55 ;
      RECT 17683.465 1048.035 17683.745 1193.31 ;
      RECT 17682.905 1046.935 17683.185 1193.045 ;
      RECT 17682.345 1048.035 17682.625 1192.805 ;
      RECT 17681.785 1046.935 17682.065 1192.565 ;
      RECT 17681.225 1048.035 17681.505 1192.325 ;
      RECT 17672.265 1046.935 17672.545 1186.16 ;
      RECT 17671.705 1048.035 17671.985 1186.4 ;
      RECT 17671.145 1048.035 17671.425 1186.64 ;
      RECT 17670.585 1048.035 17670.865 1186.64 ;
      RECT 17670.025 1048.035 17670.305 1186.4 ;
      RECT 17669.465 1048.035 17669.745 1186.16 ;
      RECT 17668.905 1048.035 17669.185 1185.92 ;
      RECT 17668.345 1048.035 17668.625 1185.68 ;
      RECT 17667.785 1048.035 17668.065 1185.44 ;
      RECT 17667.225 1048.035 17667.505 1185.2 ;
      RECT 17666.665 1048.035 17666.945 1184.96 ;
      RECT 17666.105 1048.035 17666.385 1184.72 ;
      RECT 17665.545 1048.035 17665.825 1184.48 ;
      RECT 17664.985 1046.935 17665.265 1184.24 ;
      RECT 17662.465 1048.035 17662.745 1185.96 ;
      RECT 17661.905 1046.935 17662.185 1185.72 ;
      RECT 17661.345 1048.035 17661.625 1185.48 ;
      RECT 17660.785 1046.935 17661.065 1185.24 ;
      RECT 17660.225 1048.035 17660.505 1185 ;
      RECT 17659.665 1048.035 17659.945 1184.76 ;
      RECT 17659.105 1048.035 17659.385 1184.52 ;
      RECT 17633.065 1048.035 17633.345 1187.305 ;
      RECT 17632.505 1048.035 17632.785 1187.545 ;
      RECT 17631.945 1048.035 17632.225 1187.785 ;
      RECT 17631.385 1048.035 17631.665 1188.025 ;
      RECT 17630.825 1048.035 17631.105 1188.265 ;
      RECT 17630.265 1046.935 17630.545 1188.505 ;
      RECT 17629.705 1048.035 17629.985 1188.745 ;
      RECT 17629.145 1046.935 17629.425 1188.985 ;
      RECT 17628.585 1048.035 17628.865 1189.225 ;
      RECT 17628.025 1048.035 17628.305 1189.465 ;
      RECT 17627.465 1048.035 17627.745 1189.705 ;
      RECT 17626.905 1048.035 17627.185 1189.945 ;
      RECT 17626.345 1048.035 17626.625 1190.185 ;
      RECT 17625.785 1048.035 17626.065 1190.425 ;
      RECT 17625.225 1048.035 17625.505 1190.665 ;
      RECT 17624.665 1048.035 17624.945 1190.665 ;
      RECT 17624.105 1048.035 17624.385 1190.425 ;
      RECT 17623.545 1048.035 17623.825 1190.185 ;
      RECT 17622.985 1048.035 17623.265 1189.945 ;
      RECT 17622.425 1048.035 17622.705 1189.7 ;
      RECT 17621.865 1048.035 17622.145 1189.46 ;
      RECT 17621.305 1048.035 17621.585 1189.22 ;
      RECT 17620.745 1046.935 17621.025 1188.98 ;
      RECT 17620.185 1048.035 17620.465 1188.74 ;
      RECT 17606.745 1046.935 17607.025 1186.22 ;
      RECT 17606.185 1048.035 17606.465 1185.98 ;
      RECT 17605.625 1048.035 17605.905 1185.74 ;
      RECT 17605.065 1048.035 17605.345 1185.5 ;
      RECT 17604.505 1046.935 17604.785 1185.26 ;
      RECT 17603.945 1048.035 17604.225 1185.02 ;
      RECT 17603.385 1046.935 17603.665 1184.78 ;
      RECT 17602.825 1048.035 17603.105 1184.54 ;
      RECT 17602.265 1046.935 17602.545 1184.3 ;
      RECT 17601.705 1048.035 17601.985 1184.06 ;
      RECT 17601.145 1048.035 17601.425 1183.82 ;
      RECT 17600.585 1048.035 17600.865 1183.58 ;
      RECT 17600.025 1048.035 17600.305 1183.34 ;
      RECT 17599.465 1048.035 17599.745 1183.1 ;
      RECT 17598.905 1048.035 17599.185 1182.86 ;
      RECT 17598.345 1048.035 17598.625 1182.62 ;
      RECT 17597.785 1048.035 17598.065 1182.38 ;
      RECT 17597.225 1048.035 17597.505 1182.14 ;
      RECT 17596.665 1048.035 17596.945 1181.9 ;
      RECT 17596.105 1048.035 17596.385 1181.66 ;
      RECT 17595.545 1048.035 17595.825 1181.42 ;
      RECT 17594.985 1046.935 17595.265 1181.18 ;
      RECT 17594.425 1048.035 17594.705 1180.94 ;
      RECT 17593.865 1046.935 17594.145 1180.7 ;
      RECT 17554.105 1048.035 17554.385 1191.17 ;
      RECT 17553.545 1046.935 17553.825 1191.41 ;
      RECT 17552.985 1048.035 17553.265 1191.65 ;
      RECT 17552.425 1048.035 17552.705 1191.89 ;
      RECT 17551.865 1048.035 17552.145 1192.13 ;
      RECT 17551.305 1048.035 17551.585 1192.37 ;
      RECT 17550.745 1048.035 17551.025 1192.61 ;
      RECT 17550.185 1048.035 17550.465 1192.855 ;
      RECT 17549.625 1048.035 17549.905 1193.095 ;
      RECT 17549.065 1048.035 17549.345 1193.335 ;
      RECT 17548.505 1046.935 17548.785 1193.575 ;
      RECT 17547.945 1048.035 17548.225 1193.815 ;
      RECT 17547.385 1046.935 17547.665 1194.055 ;
      RECT 17546.825 1048.035 17547.105 1194.295 ;
      RECT 17546.265 1048.035 17546.545 1194.535 ;
      RECT 17545.705 1048.035 17545.985 1194.775 ;
      RECT 17545.145 1048.035 17545.425 1195.015 ;
      RECT 17544.585 1048.035 17544.865 1195.255 ;
      RECT 17544.025 1048.035 17544.305 1195.495 ;
      RECT 17543.465 1048.035 17543.745 1195.735 ;
      RECT 17542.905 1048.035 17543.185 1195.975 ;
      RECT 17542.345 1048.035 17542.625 1196.215 ;
      RECT 17541.785 1048.035 17542.065 1196.455 ;
      RECT 17541.225 1048.035 17541.505 1196.695 ;
      RECT 17532.265 1048.035 17532.545 1192.28 ;
      RECT 17531.705 1048.035 17531.985 1192.04 ;
      RECT 17531.145 1048.035 17531.425 1191.8 ;
      RECT 17530.585 1046.935 17530.865 1191.56 ;
      RECT 17530.025 1048.035 17530.305 1191.32 ;
      RECT 17529.465 1046.935 17529.745 1191.08 ;
      RECT 17528.905 1048.035 17529.185 1190.84 ;
      RECT 17528.345 1048.035 17528.625 1190.6 ;
      RECT 17527.785 1048.035 17528.065 1190.36 ;
      RECT 17527.225 1046.935 17527.505 1190.12 ;
      RECT 17526.665 1048.035 17526.945 1189.88 ;
      RECT 17526.105 1046.935 17526.385 1189.64 ;
      RECT 17525.545 1048.035 17525.825 1189.4 ;
      RECT 17524.985 1046.935 17525.265 1189.16 ;
      RECT 17522.465 1048.035 17522.745 1181.56 ;
      RECT 17521.905 1048.035 17522.185 1181.32 ;
      RECT 17521.345 1048.035 17521.625 1181.08 ;
      RECT 17520.785 1048.035 17521.065 1180.84 ;
      RECT 17520.225 1048.035 17520.505 1180.6 ;
      RECT 17519.665 1048.035 17519.945 1180.36 ;
      RECT 17519.105 1048.035 17519.385 1180.12 ;
      RECT 17493.065 1048.035 17493.345 1193.995 ;
      RECT 17492.505 1048.035 17492.785 1194.235 ;
      RECT 17491.945 1048.035 17492.225 1194.475 ;
      RECT 17491.385 1048.035 17491.665 1194.715 ;
      RECT 17490.825 1048.035 17491.105 1194.955 ;
      RECT 17490.265 1046.935 17490.545 1194.955 ;
      RECT 17489.705 1048.035 17489.985 1194.715 ;
      RECT 17489.145 1046.935 17489.425 1194.47 ;
      RECT 17488.585 1048.035 17488.865 1194.23 ;
      RECT 17488.025 1046.935 17488.305 1193.99 ;
      RECT 17487.465 1048.035 17487.745 1193.75 ;
      RECT 17486.905 1048.035 17487.185 1193.51 ;
      RECT 17486.345 1048.035 17486.625 1193.27 ;
      RECT 17485.785 1048.035 17486.065 1193.03 ;
      RECT 17485.225 1048.035 17485.505 1192.79 ;
      RECT 17484.665 1048.035 17484.945 1192.55 ;
      RECT 17484.105 1048.035 17484.385 1192.31 ;
      RECT 17483.545 1048.035 17483.825 1192.07 ;
      RECT 17482.985 1046.935 17483.265 1191.83 ;
      RECT 17482.425 1048.035 17482.705 1191.59 ;
      RECT 17481.865 1046.935 17482.145 1191.35 ;
      RECT 17481.305 1048.035 17481.585 1191.11 ;
      RECT 17480.745 1048.035 17481.025 1190.87 ;
      RECT 17480.185 1048.035 17480.465 1190.63 ;
      RECT 17466.745 1048.035 17467.025 1194.03 ;
      RECT 17466.185 1048.035 17466.465 1194.27 ;
      RECT 17465.625 1048.035 17465.905 1194.515 ;
      RECT 17465.065 1048.035 17465.345 1194.755 ;
      RECT 17464.505 1048.035 17464.785 1194.995 ;
      RECT 17463.945 1048.035 17464.225 1194.995 ;
      RECT 17463.385 1048.035 17463.665 1194.755 ;
      RECT 17462.825 1048.035 17463.105 1194.515 ;
      RECT 17462.265 1048.035 17462.545 1187.5 ;
      RECT 17461.705 1048.035 17461.985 1187.26 ;
      RECT 17461.145 1048.035 17461.425 1187.02 ;
      RECT 17460.585 1046.935 17460.865 1186.78 ;
      RECT 17460.025 1048.035 17460.305 1186.54 ;
      RECT 17459.465 1046.935 17459.745 1186.3 ;
      RECT 17458.905 1048.035 17459.185 1186.06 ;
      RECT 17458.345 1048.035 17458.625 1185.82 ;
      RECT 17457.785 1048.035 17458.065 1185.58 ;
      RECT 17457.225 1046.935 17457.505 1185.34 ;
      RECT 17456.665 1048.035 17456.945 1185.1 ;
      RECT 17456.105 1046.935 17456.385 1184.86 ;
      RECT 17455.545 1048.035 17455.825 1184.62 ;
      RECT 17454.985 1046.935 17455.265 1184.38 ;
      RECT 17454.425 1048.035 17454.705 1184.14 ;
      RECT 17453.865 1048.035 17454.145 1183.9 ;
      RECT 17413.545 1048.035 17413.825 1192.795 ;
      RECT 17412.985 1048.035 17413.265 1193.035 ;
      RECT 17412.425 1048.035 17412.705 1193.28 ;
      RECT 17411.865 1048.035 17412.145 1193.52 ;
      RECT 17411.305 1048.035 17411.585 1193.76 ;
      RECT 17410.745 1048.035 17411.025 1194 ;
      RECT 17410.185 1048.035 17410.465 1194.24 ;
      RECT 17409.625 1048.035 17409.905 1194.48 ;
      RECT 17409.065 1048.035 17409.345 1194.72 ;
      RECT 17408.505 1048.035 17408.785 1194.96 ;
      RECT 17407.945 1046.935 17408.225 1195.2 ;
      RECT 17407.385 1048.035 17407.665 1195.44 ;
      RECT 17406.825 1046.935 17407.105 1195.68 ;
      RECT 17406.265 1048.035 17406.545 1195.92 ;
      RECT 17405.705 1046.935 17405.985 1196.16 ;
      RECT 17405.145 1048.035 17405.425 1196.16 ;
      RECT 17404.585 1048.035 17404.865 1195.92 ;
      RECT 17404.025 1048.035 17404.305 1195.68 ;
      RECT 17403.465 1048.035 17403.745 1195.44 ;
      RECT 17402.905 1048.035 17403.185 1195.2 ;
      RECT 17402.345 1048.035 17402.625 1194.96 ;
      RECT 17401.785 1048.035 17402.065 1194.72 ;
      RECT 17401.225 1048.035 17401.505 1194.48 ;
      RECT 17392.265 1046.935 17392.545 1194.51 ;
      RECT 17391.705 1048.035 17391.985 1194.75 ;
      RECT 17391.145 1046.935 17391.425 1194.99 ;
      RECT 17390.585 1048.035 17390.865 1195.205 ;
      RECT 17390.025 1048.035 17390.305 1194.78 ;
      RECT 17389.465 1048.035 17389.745 1194.54 ;
      RECT 17388.905 1048.035 17389.185 1194.3 ;
      RECT 17388.345 1048.035 17388.625 1194.06 ;
      RECT 17387.785 1048.035 17388.065 1193.82 ;
      RECT 17387.225 1048.035 17387.505 1193.58 ;
      RECT 17386.665 1048.035 17386.945 1193.34 ;
      RECT 17386.105 1048.035 17386.385 1193.1 ;
      RECT 17385.545 1048.035 17385.825 1192.86 ;
      RECT 17384.985 1048.035 17385.265 1192.62 ;
      RECT 17382.465 1048.035 17382.745 1191.795 ;
      RECT 17381.905 1048.035 17382.185 1191.555 ;
      RECT 17381.345 1048.035 17381.625 1191.315 ;
      RECT 17380.785 1046.935 17381.065 1191.075 ;
      RECT 17380.225 1048.035 17380.505 1190.835 ;
      RECT 17379.665 1046.935 17379.945 1190.595 ;
      RECT 17379.105 1048.035 17379.385 1190.355 ;
      RECT 17378.545 1048.035 17378.825 1190.115 ;
      RECT 17351.945 1048.035 17352.225 1201.16 ;
      RECT 17351.385 1046.935 17351.665 1201.4 ;
      RECT 17350.825 1048.035 17351.105 1201.64 ;
      RECT 17350.265 1046.935 17350.545 1201.885 ;
      RECT 17349.705 1048.035 17349.985 1202.125 ;
      RECT 17349.145 1046.935 17349.425 1202.365 ;
      RECT 17348.585 1048.035 17348.865 1202.605 ;
      RECT 17348.025 1048.035 17348.305 1202.845 ;
      RECT 17347.465 1048.035 17347.745 1188.465 ;
      RECT 17346.905 1048.035 17347.185 1188.225 ;
      RECT 17346.345 1048.035 17346.625 1187.985 ;
      RECT 17345.785 1048.035 17346.065 1187.745 ;
      RECT 17345.225 1048.035 17345.505 1187.505 ;
      RECT 17344.665 1048.035 17344.945 1187.265 ;
      RECT 17344.105 1048.035 17344.385 1187.025 ;
      RECT 17343.545 1048.035 17343.825 1186.785 ;
      RECT 17342.985 1048.035 17343.265 1186.545 ;
      RECT 17342.425 1048.035 17342.705 1186.305 ;
      RECT 17341.865 1046.935 17342.145 1186.065 ;
      RECT 17341.305 1048.035 17341.585 1185.825 ;
      RECT 17340.745 1046.935 17341.025 1185.585 ;
      RECT 17340.185 1048.035 17340.465 1185.345 ;
      RECT 17326.185 1046.935 17326.465 1191.465 ;
      RECT 17325.625 1048.035 17325.905 1191.225 ;
      RECT 17325.065 1048.035 17325.345 1190.985 ;
      RECT 17324.505 1048.035 17324.785 1190.745 ;
      RECT 17323.945 1048.035 17324.225 1190.505 ;
      RECT 17323.385 1048.035 17323.665 1190.265 ;
      RECT 17322.825 1048.035 17323.105 1190.025 ;
      RECT 17322.265 1048.035 17322.545 1189.785 ;
      RECT 17321.705 1048.035 17321.985 1189.545 ;
      RECT 17321.145 1046.935 17321.425 1189.305 ;
      RECT 17320.585 1048.035 17320.865 1189.065 ;
      RECT 17320.025 1046.935 17320.305 1188.825 ;
      RECT 17319.465 1048.035 17319.745 1188.585 ;
      RECT 17318.905 1048.035 17319.185 1188.345 ;
      RECT 17318.345 1048.035 17318.625 1188.105 ;
      RECT 17317.785 1048.035 17318.065 1187.865 ;
      RECT 17317.225 1048.035 17317.505 1187.625 ;
      RECT 17316.665 1048.035 17316.945 1187.385 ;
      RECT 17316.105 1048.035 17316.385 1187.145 ;
      RECT 17315.545 1048.035 17315.825 1186.905 ;
      RECT 17314.985 1048.035 17315.265 1186.665 ;
      RECT 17314.425 1048.035 17314.705 1186.425 ;
      RECT 17313.865 1048.035 17314.145 1186.185 ;
      RECT 17274.665 1048.035 17274.945 1193.09 ;
      RECT 17274.105 1048.035 17274.385 1193.33 ;
      RECT 17273.545 1048.035 17273.825 1193.57 ;
      RECT 17272.985 1046.935 17273.265 1193.81 ;
      RECT 17272.425 1048.035 17272.705 1194.05 ;
      RECT 17271.865 1046.935 17272.145 1194.29 ;
      RECT 17271.305 1048.035 17271.585 1194.53 ;
      RECT 17270.745 1048.035 17271.025 1194.77 ;
      RECT 17270.185 1048.035 17270.465 1195.01 ;
      RECT 17269.625 1046.935 17269.905 1195.25 ;
      RECT 17269.065 1048.035 17269.345 1195.49 ;
      RECT 17268.505 1046.935 17268.785 1195.73 ;
      RECT 17267.945 1048.035 17268.225 1195.97 ;
      RECT 17267.385 1046.935 17267.665 1196.21 ;
      RECT 17266.825 1048.035 17267.105 1196.45 ;
      RECT 17266.265 1048.035 17266.545 1196.69 ;
      RECT 17265.705 1048.035 17265.985 1196.69 ;
      RECT 17265.145 1048.035 17265.425 1196.45 ;
      RECT 17264.585 1048.035 17264.865 1196.21 ;
      RECT 17264.025 1048.035 17264.305 1195.97 ;
      RECT 17263.465 1048.035 17263.745 1195.73 ;
      RECT 17262.905 1048.035 17263.185 1195.49 ;
      RECT 17262.345 1048.035 17262.625 1195.25 ;
      RECT 17261.785 1048.035 17262.065 1195.01 ;
      RECT 17261.225 1048.035 17261.505 1194.77 ;
      RECT 17252.265 1048.035 17252.545 1194.285 ;
      RECT 17251.705 1046.935 17251.985 1194.045 ;
      RECT 17251.145 1048.035 17251.425 1193.805 ;
      RECT 17250.585 1046.935 17250.865 1193.565 ;
      RECT 17250.025 1048.035 17250.305 1193.325 ;
      RECT 17249.465 1046.935 17249.745 1193.085 ;
      RECT 17248.905 1048.035 17249.185 1192.845 ;
      RECT 17248.345 1048.035 17248.625 1192.605 ;
      RECT 17247.785 1048.035 17248.065 1192.365 ;
      RECT 17247.225 1048.035 17247.505 1192.125 ;
      RECT 17246.665 1048.035 17246.945 1191.885 ;
      RECT 17246.105 1048.035 17246.385 1191.645 ;
      RECT 17245.545 1048.035 17245.825 1191.405 ;
      RECT 17244.985 1048.035 17245.265 1191.165 ;
      RECT 17242.465 1046.935 17242.745 1192.885 ;
      RECT 17241.905 1048.035 17242.185 1192.645 ;
      RECT 17241.345 1046.935 17241.625 1192.405 ;
      RECT 17240.785 1048.035 17241.065 1192.165 ;
      RECT 17240.225 1048.035 17240.505 1191.925 ;
      RECT 17239.665 1048.035 17239.945 1191.685 ;
      RECT 17239.105 1048.035 17239.385 1191.445 ;
      RECT 17238.545 1048.035 17238.825 1191.205 ;
      RECT 17212.505 1048.035 17212.785 1188.855 ;
      RECT 17211.945 1048.035 17212.225 1189.095 ;
      RECT 17211.385 1048.035 17211.665 1189.335 ;
      RECT 17210.825 1048.035 17211.105 1189.58 ;
      RECT 17210.265 1048.035 17210.545 1189.82 ;
      RECT 17209.705 1048.035 17209.985 1190.06 ;
      RECT 17209.145 1048.035 17209.425 1190.06 ;
      RECT 17208.585 1048.035 17208.865 1189.82 ;
      RECT 17208.025 1048.035 17208.305 1189.58 ;
      RECT 17207.465 1046.935 17207.745 1189.34 ;
      RECT 17206.905 1048.035 17207.185 1189.1 ;
      RECT 17206.345 1046.935 17206.625 1188.86 ;
      RECT 17205.785 1048.035 17206.065 1188.62 ;
      RECT 17205.225 1048.035 17205.505 1188.38 ;
      RECT 17204.665 1048.035 17204.945 1188.14 ;
      RECT 17204.105 1046.935 17204.385 1187.9 ;
      RECT 17203.545 1048.035 17203.825 1187.66 ;
      RECT 17202.985 1046.935 17203.265 1187.42 ;
      RECT 17202.425 1048.035 17202.705 1187.18 ;
      RECT 17201.865 1046.935 17202.145 1186.94 ;
      RECT 17201.305 1048.035 17201.585 1186.7 ;
      RECT 17200.745 1048.035 17201.025 1186.46 ;
      RECT 17200.185 1048.035 17200.465 1186.22 ;
      RECT 17199.625 1048.035 17199.905 1185.98 ;
      RECT 17186.185 1048.035 17186.465 1191.78 ;
      RECT 17185.625 1048.035 17185.905 1191.54 ;
      RECT 17185.065 1048.035 17185.345 1191.3 ;
      RECT 17184.505 1048.035 17184.785 1191.06 ;
      RECT 17183.945 1048.035 17184.225 1190.82 ;
      RECT 17183.385 1048.035 17183.665 1190.58 ;
      RECT 17182.825 1048.035 17183.105 1190.34 ;
      RECT 17182.265 1048.035 17182.545 1190.1 ;
      RECT 17181.705 1046.935 17181.985 1189.86 ;
      RECT 17181.145 1048.035 17181.425 1189.62 ;
      RECT 17180.585 1046.935 17180.865 1189.3 ;
      RECT 17180.025 1048.035 17180.305 1189.14 ;
      RECT 17179.465 1046.935 17179.745 1188.9 ;
      RECT 17178.905 1048.035 17179.185 1188.66 ;
      RECT 17178.345 1048.035 17178.625 1188.42 ;
      RECT 17177.785 1048.035 17178.065 1188.18 ;
      RECT 17177.225 1048.035 17177.505 1187.94 ;
      RECT 17176.665 1048.035 17176.945 1187.7 ;
      RECT 17176.105 1048.035 17176.385 1187.46 ;
      RECT 17175.545 1048.035 17175.825 1187.22 ;
      RECT 17174.985 1048.035 17175.265 1186.98 ;
      RECT 17174.425 1046.935 17174.705 1186.74 ;
      RECT 17173.865 1048.035 17174.145 1186.5 ;
      RECT 17173.305 1046.935 17173.585 1186.26 ;
      RECT 17134.105 1048.035 17134.385 1191.87 ;
      RECT 17133.545 1048.035 17133.825 1192.11 ;
      RECT 17132.985 1048.035 17133.265 1192.35 ;
      RECT 17132.425 1048.035 17132.705 1192.59 ;
      RECT 17131.865 1048.035 17132.145 1192.83 ;
      RECT 17131.305 1048.035 17131.585 1193.07 ;
      RECT 17130.745 1048.035 17131.025 1193.31 ;
      RECT 17130.185 1048.035 17130.465 1193.55 ;
      RECT 17129.625 1048.035 17129.905 1193.79 ;
      RECT 17129.065 1048.035 17129.345 1194.03 ;
      RECT 17128.505 1048.035 17128.785 1194.27 ;
      RECT 17127.945 1048.035 17128.225 1194.51 ;
      RECT 17127.385 1048.035 17127.665 1194.75 ;
      RECT 17126.825 1048.035 17127.105 1194.75 ;
      RECT 17126.265 1046.935 17126.545 1194.51 ;
      RECT 17125.705 1048.035 17125.985 1194.27 ;
      RECT 17125.145 1046.935 17125.425 1194.03 ;
      RECT 17124.585 1048.035 17124.865 1193.79 ;
      RECT 17124.025 1048.035 17124.305 1193.55 ;
      RECT 17123.465 1048.035 17123.745 1193.31 ;
      RECT 17122.905 1046.935 17123.185 1193.045 ;
      RECT 17122.345 1048.035 17122.625 1192.805 ;
      RECT 17121.785 1046.935 17122.065 1192.565 ;
      RECT 17121.225 1048.035 17121.505 1192.325 ;
      RECT 17112.265 1046.935 17112.545 1186.16 ;
      RECT 17111.705 1048.035 17111.985 1186.4 ;
      RECT 17111.145 1048.035 17111.425 1186.64 ;
      RECT 17110.585 1048.035 17110.865 1186.64 ;
      RECT 17110.025 1048.035 17110.305 1186.4 ;
      RECT 17109.465 1048.035 17109.745 1186.16 ;
      RECT 17108.905 1048.035 17109.185 1185.92 ;
      RECT 17108.345 1048.035 17108.625 1185.68 ;
      RECT 17107.785 1048.035 17108.065 1185.44 ;
      RECT 17107.225 1048.035 17107.505 1185.2 ;
      RECT 17106.665 1048.035 17106.945 1184.96 ;
      RECT 17106.105 1048.035 17106.385 1184.72 ;
      RECT 17105.545 1048.035 17105.825 1184.48 ;
      RECT 17104.985 1046.935 17105.265 1184.24 ;
      RECT 17102.465 1048.035 17102.745 1185.96 ;
      RECT 17101.905 1046.935 17102.185 1185.72 ;
      RECT 17101.345 1048.035 17101.625 1185.48 ;
      RECT 17100.785 1046.935 17101.065 1185.24 ;
      RECT 17100.225 1048.035 17100.505 1185 ;
      RECT 17099.665 1048.035 17099.945 1184.76 ;
      RECT 17099.105 1048.035 17099.385 1184.52 ;
      RECT 17073.065 1048.035 17073.345 1187.305 ;
      RECT 17072.505 1048.035 17072.785 1187.545 ;
      RECT 17071.945 1048.035 17072.225 1187.785 ;
      RECT 17071.385 1048.035 17071.665 1188.025 ;
      RECT 17070.825 1048.035 17071.105 1188.265 ;
      RECT 17070.265 1046.935 17070.545 1188.505 ;
      RECT 17069.705 1048.035 17069.985 1188.745 ;
      RECT 17069.145 1046.935 17069.425 1188.985 ;
      RECT 17068.585 1048.035 17068.865 1189.225 ;
      RECT 17068.025 1048.035 17068.305 1189.465 ;
      RECT 17067.465 1048.035 17067.745 1189.705 ;
      RECT 17066.905 1048.035 17067.185 1189.945 ;
      RECT 17066.345 1048.035 17066.625 1190.185 ;
      RECT 17065.785 1048.035 17066.065 1190.425 ;
      RECT 17065.225 1048.035 17065.505 1190.665 ;
      RECT 17064.665 1048.035 17064.945 1190.665 ;
      RECT 17064.105 1048.035 17064.385 1190.425 ;
      RECT 17063.545 1048.035 17063.825 1190.185 ;
      RECT 17062.985 1048.035 17063.265 1189.945 ;
      RECT 17062.425 1048.035 17062.705 1189.7 ;
      RECT 17061.865 1048.035 17062.145 1189.46 ;
      RECT 17061.305 1048.035 17061.585 1189.22 ;
      RECT 17060.745 1046.935 17061.025 1188.98 ;
      RECT 17060.185 1048.035 17060.465 1188.74 ;
      RECT 17046.745 1046.935 17047.025 1186.22 ;
      RECT 17046.185 1048.035 17046.465 1185.98 ;
      RECT 17045.625 1048.035 17045.905 1185.74 ;
      RECT 17045.065 1048.035 17045.345 1185.5 ;
      RECT 17044.505 1046.935 17044.785 1185.26 ;
      RECT 17043.945 1048.035 17044.225 1185.02 ;
      RECT 17043.385 1046.935 17043.665 1184.78 ;
      RECT 17042.825 1048.035 17043.105 1184.54 ;
      RECT 17042.265 1046.935 17042.545 1184.3 ;
      RECT 17041.705 1048.035 17041.985 1184.06 ;
      RECT 17041.145 1048.035 17041.425 1183.82 ;
      RECT 17040.585 1048.035 17040.865 1183.58 ;
      RECT 17040.025 1048.035 17040.305 1183.34 ;
      RECT 17039.465 1048.035 17039.745 1183.1 ;
      RECT 17038.905 1048.035 17039.185 1182.86 ;
      RECT 17038.345 1048.035 17038.625 1182.62 ;
      RECT 17037.785 1048.035 17038.065 1182.38 ;
      RECT 17037.225 1048.035 17037.505 1182.14 ;
      RECT 17036.665 1048.035 17036.945 1181.9 ;
      RECT 17036.105 1048.035 17036.385 1181.66 ;
      RECT 17035.545 1048.035 17035.825 1181.42 ;
      RECT 17034.985 1046.935 17035.265 1181.18 ;
      RECT 17034.425 1048.035 17034.705 1180.94 ;
      RECT 17033.865 1046.935 17034.145 1180.7 ;
      RECT 16994.105 1048.035 16994.385 1191.17 ;
      RECT 16993.545 1046.935 16993.825 1191.41 ;
      RECT 16992.985 1048.035 16993.265 1191.65 ;
      RECT 16992.425 1048.035 16992.705 1191.89 ;
      RECT 16991.865 1048.035 16992.145 1192.13 ;
      RECT 16991.305 1048.035 16991.585 1192.37 ;
      RECT 16990.745 1048.035 16991.025 1192.61 ;
      RECT 16990.185 1048.035 16990.465 1192.855 ;
      RECT 16989.625 1048.035 16989.905 1193.095 ;
      RECT 16989.065 1048.035 16989.345 1193.335 ;
      RECT 16988.505 1046.935 16988.785 1193.575 ;
      RECT 16987.945 1048.035 16988.225 1193.815 ;
      RECT 16987.385 1046.935 16987.665 1194.055 ;
      RECT 16986.825 1048.035 16987.105 1194.295 ;
      RECT 16986.265 1048.035 16986.545 1194.535 ;
      RECT 16985.705 1048.035 16985.985 1194.775 ;
      RECT 16985.145 1048.035 16985.425 1195.015 ;
      RECT 16984.585 1048.035 16984.865 1195.255 ;
      RECT 16984.025 1048.035 16984.305 1195.495 ;
      RECT 16983.465 1048.035 16983.745 1195.735 ;
      RECT 16982.905 1048.035 16983.185 1195.975 ;
      RECT 16982.345 1048.035 16982.625 1196.215 ;
      RECT 16981.785 1048.035 16982.065 1196.455 ;
      RECT 16981.225 1048.035 16981.505 1196.695 ;
      RECT 16972.265 1048.035 16972.545 1192.28 ;
      RECT 16971.705 1048.035 16971.985 1192.04 ;
      RECT 16971.145 1048.035 16971.425 1191.8 ;
      RECT 16970.585 1046.935 16970.865 1191.56 ;
      RECT 16970.025 1048.035 16970.305 1191.32 ;
      RECT 16969.465 1046.935 16969.745 1191.08 ;
      RECT 16968.905 1048.035 16969.185 1190.84 ;
      RECT 16968.345 1048.035 16968.625 1190.6 ;
      RECT 16967.785 1048.035 16968.065 1190.36 ;
      RECT 16967.225 1046.935 16967.505 1190.12 ;
      RECT 16966.665 1048.035 16966.945 1189.88 ;
      RECT 16966.105 1046.935 16966.385 1189.64 ;
      RECT 16965.545 1048.035 16965.825 1189.4 ;
      RECT 16964.985 1046.935 16965.265 1189.16 ;
      RECT 16962.465 1048.035 16962.745 1181.56 ;
      RECT 16961.905 1048.035 16962.185 1181.32 ;
      RECT 16961.345 1048.035 16961.625 1181.08 ;
      RECT 16960.785 1048.035 16961.065 1180.84 ;
      RECT 16960.225 1048.035 16960.505 1180.6 ;
      RECT 16959.665 1048.035 16959.945 1180.36 ;
      RECT 16959.105 1048.035 16959.385 1180.12 ;
      RECT 16933.065 1048.035 16933.345 1193.995 ;
      RECT 16932.505 1048.035 16932.785 1194.235 ;
      RECT 16931.945 1048.035 16932.225 1194.475 ;
      RECT 16931.385 1048.035 16931.665 1194.715 ;
      RECT 16930.825 1048.035 16931.105 1194.955 ;
      RECT 16930.265 1046.935 16930.545 1194.955 ;
      RECT 16929.705 1048.035 16929.985 1194.715 ;
      RECT 16929.145 1046.935 16929.425 1194.47 ;
      RECT 16928.585 1048.035 16928.865 1194.23 ;
      RECT 16928.025 1046.935 16928.305 1193.99 ;
      RECT 16927.465 1048.035 16927.745 1193.75 ;
      RECT 16926.905 1048.035 16927.185 1193.51 ;
      RECT 16926.345 1048.035 16926.625 1193.27 ;
      RECT 16925.785 1048.035 16926.065 1193.03 ;
      RECT 16925.225 1048.035 16925.505 1192.79 ;
      RECT 16924.665 1048.035 16924.945 1192.55 ;
      RECT 16924.105 1048.035 16924.385 1192.31 ;
      RECT 16923.545 1048.035 16923.825 1192.07 ;
      RECT 16922.985 1046.935 16923.265 1191.83 ;
      RECT 16922.425 1048.035 16922.705 1191.59 ;
      RECT 16921.865 1046.935 16922.145 1191.35 ;
      RECT 16921.305 1048.035 16921.585 1191.11 ;
      RECT 16920.745 1048.035 16921.025 1190.87 ;
      RECT 16920.185 1048.035 16920.465 1190.63 ;
      RECT 16906.745 1048.035 16907.025 1194.03 ;
      RECT 16906.185 1048.035 16906.465 1194.27 ;
      RECT 16905.625 1048.035 16905.905 1194.515 ;
      RECT 16905.065 1048.035 16905.345 1194.755 ;
      RECT 16904.505 1048.035 16904.785 1194.995 ;
      RECT 16903.945 1048.035 16904.225 1194.995 ;
      RECT 16903.385 1048.035 16903.665 1194.755 ;
      RECT 16902.825 1048.035 16903.105 1194.515 ;
      RECT 16902.265 1048.035 16902.545 1187.5 ;
      RECT 16901.705 1048.035 16901.985 1187.26 ;
      RECT 16901.145 1048.035 16901.425 1187.02 ;
      RECT 16900.585 1046.935 16900.865 1186.78 ;
      RECT 16900.025 1048.035 16900.305 1186.54 ;
      RECT 16899.465 1046.935 16899.745 1186.3 ;
      RECT 16898.905 1048.035 16899.185 1186.06 ;
      RECT 16898.345 1048.035 16898.625 1185.82 ;
      RECT 16897.785 1048.035 16898.065 1185.58 ;
      RECT 16897.225 1046.935 16897.505 1185.34 ;
      RECT 16896.665 1048.035 16896.945 1185.1 ;
      RECT 16896.105 1046.935 16896.385 1184.86 ;
      RECT 16895.545 1048.035 16895.825 1184.62 ;
      RECT 16894.985 1046.935 16895.265 1184.38 ;
      RECT 16894.425 1048.035 16894.705 1184.14 ;
      RECT 16893.865 1048.035 16894.145 1183.9 ;
      RECT 16853.545 1048.035 16853.825 1192.795 ;
      RECT 16852.985 1048.035 16853.265 1193.035 ;
      RECT 16852.425 1048.035 16852.705 1193.28 ;
      RECT 16851.865 1048.035 16852.145 1193.52 ;
      RECT 16851.305 1048.035 16851.585 1193.76 ;
      RECT 16850.745 1048.035 16851.025 1194 ;
      RECT 16850.185 1048.035 16850.465 1194.24 ;
      RECT 16849.625 1048.035 16849.905 1194.48 ;
      RECT 16849.065 1048.035 16849.345 1194.72 ;
      RECT 16848.505 1048.035 16848.785 1194.96 ;
      RECT 16847.945 1046.935 16848.225 1195.2 ;
      RECT 16847.385 1048.035 16847.665 1195.44 ;
      RECT 16846.825 1046.935 16847.105 1195.68 ;
      RECT 16846.265 1048.035 16846.545 1195.92 ;
      RECT 16845.705 1046.935 16845.985 1196.16 ;
      RECT 16845.145 1048.035 16845.425 1196.16 ;
      RECT 16844.585 1048.035 16844.865 1195.92 ;
      RECT 16844.025 1048.035 16844.305 1195.68 ;
      RECT 16843.465 1048.035 16843.745 1195.44 ;
      RECT 16842.905 1048.035 16843.185 1195.2 ;
      RECT 16842.345 1048.035 16842.625 1194.96 ;
      RECT 16841.785 1048.035 16842.065 1194.72 ;
      RECT 16841.225 1048.035 16841.505 1194.48 ;
      RECT 16832.265 1046.935 16832.545 1194.51 ;
      RECT 16831.705 1048.035 16831.985 1194.75 ;
      RECT 16831.145 1046.935 16831.425 1194.99 ;
      RECT 16830.585 1048.035 16830.865 1195.205 ;
      RECT 16830.025 1048.035 16830.305 1194.78 ;
      RECT 16829.465 1048.035 16829.745 1194.54 ;
      RECT 16828.905 1048.035 16829.185 1194.3 ;
      RECT 16828.345 1048.035 16828.625 1194.06 ;
      RECT 16827.785 1048.035 16828.065 1193.82 ;
      RECT 16827.225 1048.035 16827.505 1193.58 ;
      RECT 16826.665 1048.035 16826.945 1193.34 ;
      RECT 16826.105 1048.035 16826.385 1193.1 ;
      RECT 16825.545 1048.035 16825.825 1192.86 ;
      RECT 16824.985 1048.035 16825.265 1192.62 ;
      RECT 16822.465 1048.035 16822.745 1191.795 ;
      RECT 16821.905 1048.035 16822.185 1191.555 ;
      RECT 16821.345 1048.035 16821.625 1191.315 ;
      RECT 16820.785 1046.935 16821.065 1191.075 ;
      RECT 16820.225 1048.035 16820.505 1190.835 ;
      RECT 16819.665 1046.935 16819.945 1190.595 ;
      RECT 16819.105 1048.035 16819.385 1190.355 ;
      RECT 16818.545 1048.035 16818.825 1190.115 ;
      RECT 16791.945 1048.035 16792.225 1201.16 ;
      RECT 16791.385 1046.935 16791.665 1201.4 ;
      RECT 16790.825 1048.035 16791.105 1201.64 ;
      RECT 16790.265 1046.935 16790.545 1201.885 ;
      RECT 16789.705 1048.035 16789.985 1202.125 ;
      RECT 16789.145 1046.935 16789.425 1202.365 ;
      RECT 16788.585 1048.035 16788.865 1202.605 ;
      RECT 16788.025 1048.035 16788.305 1202.845 ;
      RECT 16787.465 1048.035 16787.745 1188.465 ;
      RECT 16786.905 1048.035 16787.185 1188.225 ;
      RECT 16786.345 1048.035 16786.625 1187.985 ;
      RECT 16785.785 1048.035 16786.065 1187.745 ;
      RECT 16785.225 1048.035 16785.505 1187.505 ;
      RECT 16784.665 1048.035 16784.945 1187.265 ;
      RECT 16784.105 1048.035 16784.385 1187.025 ;
      RECT 16783.545 1048.035 16783.825 1186.785 ;
      RECT 16782.985 1048.035 16783.265 1186.545 ;
      RECT 16782.425 1048.035 16782.705 1186.305 ;
      RECT 16781.865 1046.935 16782.145 1186.065 ;
      RECT 16781.305 1048.035 16781.585 1185.825 ;
      RECT 16780.745 1046.935 16781.025 1185.585 ;
      RECT 16780.185 1048.035 16780.465 1185.345 ;
      RECT 16766.185 1046.935 16766.465 1191.465 ;
      RECT 16765.625 1048.035 16765.905 1191.225 ;
      RECT 16765.065 1048.035 16765.345 1190.985 ;
      RECT 16764.505 1048.035 16764.785 1190.745 ;
      RECT 16763.945 1048.035 16764.225 1190.505 ;
      RECT 16763.385 1048.035 16763.665 1190.265 ;
      RECT 16762.825 1048.035 16763.105 1190.025 ;
      RECT 16762.265 1048.035 16762.545 1189.785 ;
      RECT 16761.705 1048.035 16761.985 1189.545 ;
      RECT 16761.145 1046.935 16761.425 1189.305 ;
      RECT 16760.585 1048.035 16760.865 1189.065 ;
      RECT 16760.025 1046.935 16760.305 1188.825 ;
      RECT 16759.465 1048.035 16759.745 1188.585 ;
      RECT 16758.905 1048.035 16759.185 1188.345 ;
      RECT 16758.345 1048.035 16758.625 1188.105 ;
      RECT 16757.785 1048.035 16758.065 1187.865 ;
      RECT 16757.225 1048.035 16757.505 1187.625 ;
      RECT 16756.665 1048.035 16756.945 1187.385 ;
      RECT 16756.105 1048.035 16756.385 1187.145 ;
      RECT 16755.545 1048.035 16755.825 1186.905 ;
      RECT 16754.985 1048.035 16755.265 1186.665 ;
      RECT 16754.425 1048.035 16754.705 1186.425 ;
      RECT 16753.865 1048.035 16754.145 1186.185 ;
      RECT 16714.665 1048.035 16714.945 1193.09 ;
      RECT 16714.105 1048.035 16714.385 1193.33 ;
      RECT 16713.545 1048.035 16713.825 1193.57 ;
      RECT 16712.985 1046.935 16713.265 1193.81 ;
      RECT 16712.425 1048.035 16712.705 1194.05 ;
      RECT 16711.865 1046.935 16712.145 1194.29 ;
      RECT 16711.305 1048.035 16711.585 1194.53 ;
      RECT 16710.745 1048.035 16711.025 1194.77 ;
      RECT 16710.185 1048.035 16710.465 1195.01 ;
      RECT 16709.625 1046.935 16709.905 1195.25 ;
      RECT 16709.065 1048.035 16709.345 1195.49 ;
      RECT 16708.505 1046.935 16708.785 1195.73 ;
      RECT 16707.945 1048.035 16708.225 1195.97 ;
      RECT 16707.385 1046.935 16707.665 1196.21 ;
      RECT 16706.825 1048.035 16707.105 1196.45 ;
      RECT 16706.265 1048.035 16706.545 1196.69 ;
      RECT 16705.705 1048.035 16705.985 1196.69 ;
      RECT 16705.145 1048.035 16705.425 1196.45 ;
      RECT 16704.585 1048.035 16704.865 1196.21 ;
      RECT 16704.025 1048.035 16704.305 1195.97 ;
      RECT 16703.465 1048.035 16703.745 1195.73 ;
      RECT 16702.905 1048.035 16703.185 1195.49 ;
      RECT 16702.345 1048.035 16702.625 1195.25 ;
      RECT 16701.785 1048.035 16702.065 1195.01 ;
      RECT 16701.225 1048.035 16701.505 1194.77 ;
      RECT 16692.265 1048.035 16692.545 1194.285 ;
      RECT 16691.705 1046.935 16691.985 1194.045 ;
      RECT 16691.145 1048.035 16691.425 1193.805 ;
      RECT 16690.585 1046.935 16690.865 1193.565 ;
      RECT 16690.025 1048.035 16690.305 1193.325 ;
      RECT 16689.465 1046.935 16689.745 1193.085 ;
      RECT 16688.905 1048.035 16689.185 1192.845 ;
      RECT 16688.345 1048.035 16688.625 1192.605 ;
      RECT 16687.785 1048.035 16688.065 1192.365 ;
      RECT 16687.225 1048.035 16687.505 1192.125 ;
      RECT 16686.665 1048.035 16686.945 1191.885 ;
      RECT 16686.105 1048.035 16686.385 1191.645 ;
      RECT 16685.545 1048.035 16685.825 1191.405 ;
      RECT 16684.985 1048.035 16685.265 1191.165 ;
      RECT 16682.465 1046.935 16682.745 1192.885 ;
      RECT 16681.905 1048.035 16682.185 1192.645 ;
      RECT 16681.345 1046.935 16681.625 1192.405 ;
      RECT 16680.785 1048.035 16681.065 1192.165 ;
      RECT 16680.225 1048.035 16680.505 1191.925 ;
      RECT 16679.665 1048.035 16679.945 1191.685 ;
      RECT 16679.105 1048.035 16679.385 1191.445 ;
      RECT 16678.545 1048.035 16678.825 1191.205 ;
      RECT 16652.505 1048.035 16652.785 1188.855 ;
      RECT 16651.945 1048.035 16652.225 1189.095 ;
      RECT 16651.385 1048.035 16651.665 1189.335 ;
      RECT 16650.825 1048.035 16651.105 1189.58 ;
      RECT 16650.265 1048.035 16650.545 1189.82 ;
      RECT 16649.705 1048.035 16649.985 1190.06 ;
      RECT 16649.145 1048.035 16649.425 1190.06 ;
      RECT 16648.585 1048.035 16648.865 1189.82 ;
      RECT 16648.025 1048.035 16648.305 1189.58 ;
      RECT 16647.465 1046.935 16647.745 1189.34 ;
      RECT 16646.905 1048.035 16647.185 1189.1 ;
      RECT 16646.345 1046.935 16646.625 1188.86 ;
      RECT 16645.785 1048.035 16646.065 1188.62 ;
      RECT 16645.225 1048.035 16645.505 1188.38 ;
      RECT 16644.665 1048.035 16644.945 1188.14 ;
      RECT 16644.105 1046.935 16644.385 1187.9 ;
      RECT 16643.545 1048.035 16643.825 1187.66 ;
      RECT 16642.985 1046.935 16643.265 1187.42 ;
      RECT 16642.425 1048.035 16642.705 1187.18 ;
      RECT 16641.865 1046.935 16642.145 1186.94 ;
      RECT 16641.305 1048.035 16641.585 1186.7 ;
      RECT 16640.745 1048.035 16641.025 1186.46 ;
      RECT 16640.185 1048.035 16640.465 1186.22 ;
      RECT 16639.625 1048.035 16639.905 1185.98 ;
      RECT 16626.185 1048.035 16626.465 1191.78 ;
      RECT 16625.625 1048.035 16625.905 1191.54 ;
      RECT 16625.065 1048.035 16625.345 1191.3 ;
      RECT 16624.505 1048.035 16624.785 1191.06 ;
      RECT 16623.945 1048.035 16624.225 1190.82 ;
      RECT 16623.385 1048.035 16623.665 1190.58 ;
      RECT 16622.825 1048.035 16623.105 1190.34 ;
      RECT 16622.265 1048.035 16622.545 1190.1 ;
      RECT 16621.705 1046.935 16621.985 1189.86 ;
      RECT 16621.145 1048.035 16621.425 1189.62 ;
      RECT 16620.585 1046.935 16620.865 1189.3 ;
      RECT 16620.025 1048.035 16620.305 1189.14 ;
      RECT 16619.465 1046.935 16619.745 1188.9 ;
      RECT 16618.905 1048.035 16619.185 1188.66 ;
      RECT 16618.345 1048.035 16618.625 1188.42 ;
      RECT 16617.785 1048.035 16618.065 1188.18 ;
      RECT 16617.225 1048.035 16617.505 1187.94 ;
      RECT 16616.665 1048.035 16616.945 1187.7 ;
      RECT 16616.105 1048.035 16616.385 1187.46 ;
      RECT 16615.545 1048.035 16615.825 1187.22 ;
      RECT 16614.985 1048.035 16615.265 1186.98 ;
      RECT 16614.425 1046.935 16614.705 1186.74 ;
      RECT 16613.865 1048.035 16614.145 1186.5 ;
      RECT 16613.305 1046.935 16613.585 1186.26 ;
      RECT 16574.105 1048.035 16574.385 1191.87 ;
      RECT 16573.545 1048.035 16573.825 1192.11 ;
      RECT 16572.985 1048.035 16573.265 1192.35 ;
      RECT 16572.425 1048.035 16572.705 1192.59 ;
      RECT 16571.865 1048.035 16572.145 1192.83 ;
      RECT 16571.305 1048.035 16571.585 1193.07 ;
      RECT 16570.745 1048.035 16571.025 1193.31 ;
      RECT 16570.185 1048.035 16570.465 1193.55 ;
      RECT 16569.625 1048.035 16569.905 1193.79 ;
      RECT 16569.065 1048.035 16569.345 1194.03 ;
      RECT 16568.505 1048.035 16568.785 1194.27 ;
      RECT 16567.945 1048.035 16568.225 1194.51 ;
      RECT 16567.385 1048.035 16567.665 1194.75 ;
      RECT 16566.825 1048.035 16567.105 1194.75 ;
      RECT 16566.265 1046.935 16566.545 1194.51 ;
      RECT 16565.705 1048.035 16565.985 1194.27 ;
      RECT 16565.145 1046.935 16565.425 1194.03 ;
      RECT 16564.585 1048.035 16564.865 1193.79 ;
      RECT 16564.025 1048.035 16564.305 1193.55 ;
      RECT 16563.465 1048.035 16563.745 1193.31 ;
      RECT 16562.905 1046.935 16563.185 1193.045 ;
      RECT 16562.345 1048.035 16562.625 1192.805 ;
      RECT 16561.785 1046.935 16562.065 1192.565 ;
      RECT 16561.225 1048.035 16561.505 1192.325 ;
      RECT 16552.265 1046.935 16552.545 1186.16 ;
      RECT 16551.705 1048.035 16551.985 1186.4 ;
      RECT 16551.145 1048.035 16551.425 1186.64 ;
      RECT 16550.585 1048.035 16550.865 1186.64 ;
      RECT 16550.025 1048.035 16550.305 1186.4 ;
      RECT 16549.465 1048.035 16549.745 1186.16 ;
      RECT 16548.905 1048.035 16549.185 1185.92 ;
      RECT 16548.345 1048.035 16548.625 1185.68 ;
      RECT 16547.785 1048.035 16548.065 1185.44 ;
      RECT 16547.225 1048.035 16547.505 1185.2 ;
      RECT 16546.665 1048.035 16546.945 1184.96 ;
      RECT 16546.105 1048.035 16546.385 1184.72 ;
      RECT 16545.545 1048.035 16545.825 1184.48 ;
      RECT 16544.985 1046.935 16545.265 1184.24 ;
      RECT 16542.465 1048.035 16542.745 1185.96 ;
      RECT 16541.905 1046.935 16542.185 1185.72 ;
      RECT 16541.345 1048.035 16541.625 1185.48 ;
      RECT 16540.785 1046.935 16541.065 1185.24 ;
      RECT 16540.225 1048.035 16540.505 1185 ;
      RECT 16539.665 1048.035 16539.945 1184.76 ;
      RECT 16539.105 1048.035 16539.385 1184.52 ;
      RECT 16513.065 1048.035 16513.345 1187.305 ;
      RECT 16512.505 1048.035 16512.785 1187.545 ;
      RECT 16511.945 1048.035 16512.225 1187.785 ;
      RECT 16511.385 1048.035 16511.665 1188.025 ;
      RECT 16510.825 1048.035 16511.105 1188.265 ;
      RECT 16510.265 1046.935 16510.545 1188.505 ;
      RECT 16509.705 1048.035 16509.985 1188.745 ;
      RECT 16509.145 1046.935 16509.425 1188.985 ;
      RECT 16508.585 1048.035 16508.865 1189.225 ;
      RECT 16508.025 1048.035 16508.305 1189.465 ;
      RECT 16507.465 1048.035 16507.745 1189.705 ;
      RECT 16506.905 1048.035 16507.185 1189.945 ;
      RECT 16506.345 1048.035 16506.625 1190.185 ;
      RECT 16505.785 1048.035 16506.065 1190.425 ;
      RECT 16505.225 1048.035 16505.505 1190.665 ;
      RECT 16504.665 1048.035 16504.945 1190.665 ;
      RECT 16504.105 1048.035 16504.385 1190.425 ;
      RECT 16503.545 1048.035 16503.825 1190.185 ;
      RECT 16502.985 1048.035 16503.265 1189.945 ;
      RECT 16502.425 1048.035 16502.705 1189.7 ;
      RECT 16501.865 1048.035 16502.145 1189.46 ;
      RECT 16501.305 1048.035 16501.585 1189.22 ;
      RECT 16500.745 1046.935 16501.025 1188.98 ;
      RECT 16500.185 1048.035 16500.465 1188.74 ;
      RECT 16486.745 1046.935 16487.025 1186.22 ;
      RECT 16486.185 1048.035 16486.465 1185.98 ;
      RECT 16485.625 1048.035 16485.905 1185.74 ;
      RECT 16485.065 1048.035 16485.345 1185.5 ;
      RECT 16484.505 1046.935 16484.785 1185.26 ;
      RECT 16483.945 1048.035 16484.225 1185.02 ;
      RECT 16483.385 1046.935 16483.665 1184.78 ;
      RECT 16482.825 1048.035 16483.105 1184.54 ;
      RECT 16482.265 1046.935 16482.545 1184.3 ;
      RECT 16481.705 1048.035 16481.985 1184.06 ;
      RECT 16481.145 1048.035 16481.425 1183.82 ;
      RECT 16480.585 1048.035 16480.865 1183.58 ;
      RECT 16480.025 1048.035 16480.305 1183.34 ;
      RECT 16479.465 1048.035 16479.745 1183.1 ;
      RECT 16478.905 1048.035 16479.185 1182.86 ;
      RECT 16478.345 1048.035 16478.625 1182.62 ;
      RECT 16477.785 1048.035 16478.065 1182.38 ;
      RECT 16477.225 1048.035 16477.505 1182.14 ;
      RECT 16476.665 1048.035 16476.945 1181.9 ;
      RECT 16476.105 1048.035 16476.385 1181.66 ;
      RECT 16475.545 1048.035 16475.825 1181.42 ;
      RECT 16474.985 1046.935 16475.265 1181.18 ;
      RECT 16474.425 1048.035 16474.705 1180.94 ;
      RECT 16473.865 1046.935 16474.145 1180.7 ;
      RECT 16434.105 1048.035 16434.385 1191.17 ;
      RECT 16433.545 1046.935 16433.825 1191.41 ;
      RECT 16432.985 1048.035 16433.265 1191.65 ;
      RECT 16432.425 1048.035 16432.705 1191.89 ;
      RECT 16431.865 1048.035 16432.145 1192.13 ;
      RECT 16431.305 1048.035 16431.585 1192.37 ;
      RECT 16430.745 1048.035 16431.025 1192.61 ;
      RECT 16430.185 1048.035 16430.465 1192.855 ;
      RECT 16429.625 1048.035 16429.905 1193.095 ;
      RECT 16429.065 1048.035 16429.345 1193.335 ;
      RECT 16428.505 1046.935 16428.785 1193.575 ;
      RECT 16427.945 1048.035 16428.225 1193.815 ;
      RECT 16427.385 1046.935 16427.665 1194.055 ;
      RECT 16426.825 1048.035 16427.105 1194.295 ;
      RECT 16426.265 1048.035 16426.545 1194.535 ;
      RECT 16425.705 1048.035 16425.985 1194.775 ;
      RECT 16425.145 1048.035 16425.425 1195.015 ;
      RECT 16424.585 1048.035 16424.865 1195.255 ;
      RECT 16424.025 1048.035 16424.305 1195.495 ;
      RECT 16423.465 1048.035 16423.745 1195.735 ;
      RECT 16422.905 1048.035 16423.185 1195.975 ;
      RECT 16422.345 1048.035 16422.625 1196.215 ;
      RECT 16421.785 1048.035 16422.065 1196.455 ;
      RECT 16421.225 1048.035 16421.505 1196.695 ;
      RECT 16412.265 1048.035 16412.545 1192.28 ;
      RECT 16411.705 1048.035 16411.985 1192.04 ;
      RECT 16411.145 1048.035 16411.425 1191.8 ;
      RECT 16410.585 1046.935 16410.865 1191.56 ;
      RECT 16410.025 1048.035 16410.305 1191.32 ;
      RECT 16409.465 1046.935 16409.745 1191.08 ;
      RECT 16408.905 1048.035 16409.185 1190.84 ;
      RECT 16408.345 1048.035 16408.625 1190.6 ;
      RECT 16407.785 1048.035 16408.065 1190.36 ;
      RECT 16407.225 1046.935 16407.505 1190.12 ;
      RECT 16406.665 1048.035 16406.945 1189.88 ;
      RECT 16406.105 1046.935 16406.385 1189.64 ;
      RECT 16405.545 1048.035 16405.825 1189.4 ;
      RECT 16404.985 1046.935 16405.265 1189.16 ;
      RECT 16402.465 1048.035 16402.745 1181.56 ;
      RECT 16401.905 1048.035 16402.185 1181.32 ;
      RECT 16401.345 1048.035 16401.625 1181.08 ;
      RECT 16400.785 1048.035 16401.065 1180.84 ;
      RECT 16400.225 1048.035 16400.505 1180.6 ;
      RECT 16399.665 1048.035 16399.945 1180.36 ;
      RECT 16399.105 1048.035 16399.385 1180.12 ;
      RECT 16373.065 1048.035 16373.345 1193.995 ;
      RECT 16372.505 1048.035 16372.785 1194.235 ;
      RECT 16371.945 1048.035 16372.225 1194.475 ;
      RECT 16371.385 1048.035 16371.665 1194.715 ;
      RECT 16370.825 1048.035 16371.105 1194.955 ;
      RECT 16370.265 1046.935 16370.545 1194.955 ;
      RECT 16369.705 1048.035 16369.985 1194.715 ;
      RECT 16369.145 1046.935 16369.425 1194.47 ;
      RECT 16368.585 1048.035 16368.865 1194.23 ;
      RECT 16368.025 1046.935 16368.305 1193.99 ;
      RECT 16367.465 1048.035 16367.745 1193.75 ;
      RECT 16366.905 1048.035 16367.185 1193.51 ;
      RECT 16366.345 1048.035 16366.625 1193.27 ;
      RECT 16365.785 1048.035 16366.065 1193.03 ;
      RECT 16365.225 1048.035 16365.505 1192.79 ;
      RECT 16364.665 1048.035 16364.945 1192.55 ;
      RECT 16364.105 1048.035 16364.385 1192.31 ;
      RECT 16363.545 1048.035 16363.825 1192.07 ;
      RECT 16362.985 1046.935 16363.265 1191.83 ;
      RECT 16362.425 1048.035 16362.705 1191.59 ;
      RECT 16361.865 1046.935 16362.145 1191.35 ;
      RECT 16361.305 1048.035 16361.585 1191.11 ;
      RECT 16360.745 1048.035 16361.025 1190.87 ;
      RECT 16360.185 1048.035 16360.465 1190.63 ;
      RECT 16346.745 1048.035 16347.025 1194.03 ;
      RECT 16346.185 1048.035 16346.465 1194.27 ;
      RECT 16345.625 1048.035 16345.905 1194.515 ;
      RECT 16345.065 1048.035 16345.345 1194.755 ;
      RECT 16344.505 1048.035 16344.785 1194.995 ;
      RECT 16343.945 1048.035 16344.225 1194.995 ;
      RECT 16343.385 1048.035 16343.665 1194.755 ;
      RECT 16342.825 1048.035 16343.105 1194.515 ;
      RECT 16342.265 1048.035 16342.545 1187.5 ;
      RECT 16341.705 1048.035 16341.985 1187.26 ;
      RECT 16341.145 1048.035 16341.425 1187.02 ;
      RECT 16340.585 1046.935 16340.865 1186.78 ;
      RECT 16340.025 1048.035 16340.305 1186.54 ;
      RECT 16339.465 1046.935 16339.745 1186.3 ;
      RECT 16338.905 1048.035 16339.185 1186.06 ;
      RECT 16338.345 1048.035 16338.625 1185.82 ;
      RECT 16337.785 1048.035 16338.065 1185.58 ;
      RECT 16337.225 1046.935 16337.505 1185.34 ;
      RECT 16336.665 1048.035 16336.945 1185.1 ;
      RECT 16336.105 1046.935 16336.385 1184.86 ;
      RECT 16335.545 1048.035 16335.825 1184.62 ;
      RECT 16334.985 1046.935 16335.265 1184.38 ;
      RECT 16334.425 1048.035 16334.705 1184.14 ;
      RECT 16333.865 1048.035 16334.145 1183.9 ;
      RECT 16293.545 1048.035 16293.825 1192.795 ;
      RECT 16292.985 1048.035 16293.265 1193.035 ;
      RECT 16292.425 1048.035 16292.705 1193.28 ;
      RECT 16291.865 1048.035 16292.145 1193.52 ;
      RECT 16291.305 1048.035 16291.585 1193.76 ;
      RECT 16290.745 1048.035 16291.025 1194 ;
      RECT 16290.185 1048.035 16290.465 1194.24 ;
      RECT 16289.625 1048.035 16289.905 1194.48 ;
      RECT 16289.065 1048.035 16289.345 1194.72 ;
      RECT 16288.505 1048.035 16288.785 1194.96 ;
      RECT 16287.945 1046.935 16288.225 1195.2 ;
      RECT 16287.385 1048.035 16287.665 1195.44 ;
      RECT 16286.825 1046.935 16287.105 1195.68 ;
      RECT 16286.265 1048.035 16286.545 1195.92 ;
      RECT 16285.705 1046.935 16285.985 1196.16 ;
      RECT 16285.145 1048.035 16285.425 1196.16 ;
      RECT 16284.585 1048.035 16284.865 1195.92 ;
      RECT 16284.025 1048.035 16284.305 1195.68 ;
      RECT 16283.465 1048.035 16283.745 1195.44 ;
      RECT 16282.905 1048.035 16283.185 1195.2 ;
      RECT 16282.345 1048.035 16282.625 1194.96 ;
      RECT 16281.785 1048.035 16282.065 1194.72 ;
      RECT 16281.225 1048.035 16281.505 1194.48 ;
      RECT 16272.265 1046.935 16272.545 1194.51 ;
      RECT 16271.705 1048.035 16271.985 1194.75 ;
      RECT 16271.145 1046.935 16271.425 1194.99 ;
      RECT 16270.585 1048.035 16270.865 1195.205 ;
      RECT 16270.025 1048.035 16270.305 1194.78 ;
      RECT 16269.465 1048.035 16269.745 1194.54 ;
      RECT 16268.905 1048.035 16269.185 1194.3 ;
      RECT 16268.345 1048.035 16268.625 1194.06 ;
      RECT 16267.785 1048.035 16268.065 1193.82 ;
      RECT 16267.225 1048.035 16267.505 1193.58 ;
      RECT 16266.665 1048.035 16266.945 1193.34 ;
      RECT 16266.105 1048.035 16266.385 1193.1 ;
      RECT 16265.545 1048.035 16265.825 1192.86 ;
      RECT 16264.985 1048.035 16265.265 1192.62 ;
      RECT 16262.465 1048.035 16262.745 1191.795 ;
      RECT 16261.905 1048.035 16262.185 1191.555 ;
      RECT 16261.345 1048.035 16261.625 1191.315 ;
      RECT 16260.785 1046.935 16261.065 1191.075 ;
      RECT 16260.225 1048.035 16260.505 1190.835 ;
      RECT 16259.665 1046.935 16259.945 1190.595 ;
      RECT 16259.105 1048.035 16259.385 1190.355 ;
      RECT 16258.545 1048.035 16258.825 1190.115 ;
      RECT 16231.945 1048.035 16232.225 1201.16 ;
      RECT 16231.385 1046.935 16231.665 1201.4 ;
      RECT 16230.825 1048.035 16231.105 1201.64 ;
      RECT 16230.265 1046.935 16230.545 1201.885 ;
      RECT 16229.705 1048.035 16229.985 1202.125 ;
      RECT 16229.145 1046.935 16229.425 1202.365 ;
      RECT 16228.585 1048.035 16228.865 1202.605 ;
      RECT 16228.025 1048.035 16228.305 1202.845 ;
      RECT 16227.465 1048.035 16227.745 1188.465 ;
      RECT 16226.905 1048.035 16227.185 1188.225 ;
      RECT 16226.345 1048.035 16226.625 1187.985 ;
      RECT 16225.785 1048.035 16226.065 1187.745 ;
      RECT 16225.225 1048.035 16225.505 1187.505 ;
      RECT 16224.665 1048.035 16224.945 1187.265 ;
      RECT 16224.105 1048.035 16224.385 1187.025 ;
      RECT 16223.545 1048.035 16223.825 1186.785 ;
      RECT 16222.985 1048.035 16223.265 1186.545 ;
      RECT 16222.425 1048.035 16222.705 1186.305 ;
      RECT 16221.865 1046.935 16222.145 1186.065 ;
      RECT 16221.305 1048.035 16221.585 1185.825 ;
      RECT 16220.745 1046.935 16221.025 1185.585 ;
      RECT 16220.185 1048.035 16220.465 1185.345 ;
      RECT 16206.185 1046.935 16206.465 1191.465 ;
      RECT 16205.625 1048.035 16205.905 1191.225 ;
      RECT 16205.065 1048.035 16205.345 1190.985 ;
      RECT 16204.505 1048.035 16204.785 1190.745 ;
      RECT 16203.945 1048.035 16204.225 1190.505 ;
      RECT 16203.385 1048.035 16203.665 1190.265 ;
      RECT 16202.825 1048.035 16203.105 1190.025 ;
      RECT 16202.265 1048.035 16202.545 1189.785 ;
      RECT 16201.705 1048.035 16201.985 1189.545 ;
      RECT 16201.145 1046.935 16201.425 1189.305 ;
      RECT 16200.585 1048.035 16200.865 1189.065 ;
      RECT 16200.025 1046.935 16200.305 1188.825 ;
      RECT 16199.465 1048.035 16199.745 1188.585 ;
      RECT 16198.905 1048.035 16199.185 1188.345 ;
      RECT 16198.345 1048.035 16198.625 1188.105 ;
      RECT 16197.785 1048.035 16198.065 1187.865 ;
      RECT 16197.225 1048.035 16197.505 1187.625 ;
      RECT 16196.665 1048.035 16196.945 1187.385 ;
      RECT 16196.105 1048.035 16196.385 1187.145 ;
      RECT 16195.545 1048.035 16195.825 1186.905 ;
      RECT 16194.985 1048.035 16195.265 1186.665 ;
      RECT 16194.425 1048.035 16194.705 1186.425 ;
      RECT 16193.865 1048.035 16194.145 1186.185 ;
      RECT 16154.665 1048.035 16154.945 1193.09 ;
      RECT 16154.105 1048.035 16154.385 1193.33 ;
      RECT 16153.545 1048.035 16153.825 1193.57 ;
      RECT 16152.985 1046.935 16153.265 1193.81 ;
      RECT 16152.425 1048.035 16152.705 1194.05 ;
      RECT 16151.865 1046.935 16152.145 1194.29 ;
      RECT 16151.305 1048.035 16151.585 1194.53 ;
      RECT 16150.745 1048.035 16151.025 1194.77 ;
      RECT 16150.185 1048.035 16150.465 1195.01 ;
      RECT 16149.625 1046.935 16149.905 1195.25 ;
      RECT 16149.065 1048.035 16149.345 1195.49 ;
      RECT 16148.505 1046.935 16148.785 1195.73 ;
      RECT 16147.945 1048.035 16148.225 1195.97 ;
      RECT 16147.385 1046.935 16147.665 1196.21 ;
      RECT 16146.825 1048.035 16147.105 1196.45 ;
      RECT 16146.265 1048.035 16146.545 1196.69 ;
      RECT 16145.705 1048.035 16145.985 1196.69 ;
      RECT 16145.145 1048.035 16145.425 1196.45 ;
      RECT 16144.585 1048.035 16144.865 1196.21 ;
      RECT 16144.025 1048.035 16144.305 1195.97 ;
      RECT 16143.465 1048.035 16143.745 1195.73 ;
      RECT 16142.905 1048.035 16143.185 1195.49 ;
      RECT 16142.345 1048.035 16142.625 1195.25 ;
      RECT 16141.785 1048.035 16142.065 1195.01 ;
      RECT 16141.225 1048.035 16141.505 1194.77 ;
      RECT 16132.265 1048.035 16132.545 1194.285 ;
      RECT 16131.705 1046.935 16131.985 1194.045 ;
      RECT 16131.145 1048.035 16131.425 1193.805 ;
      RECT 16130.585 1046.935 16130.865 1193.565 ;
      RECT 16130.025 1048.035 16130.305 1193.325 ;
      RECT 16129.465 1046.935 16129.745 1193.085 ;
      RECT 16128.905 1048.035 16129.185 1192.845 ;
      RECT 16128.345 1048.035 16128.625 1192.605 ;
      RECT 16127.785 1048.035 16128.065 1192.365 ;
      RECT 16127.225 1048.035 16127.505 1192.125 ;
      RECT 16126.665 1048.035 16126.945 1191.885 ;
      RECT 16126.105 1048.035 16126.385 1191.645 ;
      RECT 16125.545 1048.035 16125.825 1191.405 ;
      RECT 16124.985 1048.035 16125.265 1191.165 ;
      RECT 16122.465 1046.935 16122.745 1192.885 ;
      RECT 16121.905 1048.035 16122.185 1192.645 ;
      RECT 16121.345 1046.935 16121.625 1192.405 ;
      RECT 16120.785 1048.035 16121.065 1192.165 ;
      RECT 16120.225 1048.035 16120.505 1191.925 ;
      RECT 16119.665 1048.035 16119.945 1191.685 ;
      RECT 16119.105 1048.035 16119.385 1191.445 ;
      RECT 16118.545 1048.035 16118.825 1191.205 ;
      RECT 16092.505 1048.035 16092.785 1188.855 ;
      RECT 16091.945 1048.035 16092.225 1189.095 ;
      RECT 16091.385 1048.035 16091.665 1189.335 ;
      RECT 16090.825 1048.035 16091.105 1189.58 ;
      RECT 16090.265 1048.035 16090.545 1189.82 ;
      RECT 16089.705 1048.035 16089.985 1190.06 ;
      RECT 16089.145 1048.035 16089.425 1190.06 ;
      RECT 16088.585 1048.035 16088.865 1189.82 ;
      RECT 16088.025 1048.035 16088.305 1189.58 ;
      RECT 16087.465 1046.935 16087.745 1189.34 ;
      RECT 16086.905 1048.035 16087.185 1189.1 ;
      RECT 16086.345 1046.935 16086.625 1188.86 ;
      RECT 16085.785 1048.035 16086.065 1188.62 ;
      RECT 16085.225 1048.035 16085.505 1188.38 ;
      RECT 16084.665 1048.035 16084.945 1188.14 ;
      RECT 16084.105 1046.935 16084.385 1187.9 ;
      RECT 16083.545 1048.035 16083.825 1187.66 ;
      RECT 16082.985 1046.935 16083.265 1187.42 ;
      RECT 16082.425 1048.035 16082.705 1187.18 ;
      RECT 16081.865 1046.935 16082.145 1186.94 ;
      RECT 16081.305 1048.035 16081.585 1186.7 ;
      RECT 16080.745 1048.035 16081.025 1186.46 ;
      RECT 16080.185 1048.035 16080.465 1186.22 ;
      RECT 16079.625 1048.035 16079.905 1185.98 ;
      RECT 16066.185 1048.035 16066.465 1191.78 ;
      RECT 16065.625 1048.035 16065.905 1191.54 ;
      RECT 16065.065 1048.035 16065.345 1191.3 ;
      RECT 16064.505 1048.035 16064.785 1191.06 ;
      RECT 16063.945 1048.035 16064.225 1190.82 ;
      RECT 16063.385 1048.035 16063.665 1190.58 ;
      RECT 16062.825 1048.035 16063.105 1190.34 ;
      RECT 16062.265 1048.035 16062.545 1190.1 ;
      RECT 16061.705 1046.935 16061.985 1189.86 ;
      RECT 16061.145 1048.035 16061.425 1189.62 ;
      RECT 16060.585 1046.935 16060.865 1189.3 ;
      RECT 16060.025 1048.035 16060.305 1189.14 ;
      RECT 16059.465 1046.935 16059.745 1188.9 ;
      RECT 16058.905 1048.035 16059.185 1188.66 ;
      RECT 16058.345 1048.035 16058.625 1188.42 ;
      RECT 16057.785 1048.035 16058.065 1188.18 ;
      RECT 16057.225 1048.035 16057.505 1187.94 ;
      RECT 16056.665 1048.035 16056.945 1187.7 ;
      RECT 16056.105 1048.035 16056.385 1187.46 ;
      RECT 16055.545 1048.035 16055.825 1187.22 ;
      RECT 16054.985 1048.035 16055.265 1186.98 ;
      RECT 16054.425 1046.935 16054.705 1186.74 ;
      RECT 16053.865 1048.035 16054.145 1186.5 ;
      RECT 16053.305 1046.935 16053.585 1186.26 ;
      RECT 16014.105 1048.035 16014.385 1191.87 ;
      RECT 16013.545 1048.035 16013.825 1192.11 ;
      RECT 16012.985 1048.035 16013.265 1192.35 ;
      RECT 16012.425 1048.035 16012.705 1192.59 ;
      RECT 16011.865 1048.035 16012.145 1192.83 ;
      RECT 16011.305 1048.035 16011.585 1193.07 ;
      RECT 16010.745 1048.035 16011.025 1193.31 ;
      RECT 16010.185 1048.035 16010.465 1193.55 ;
      RECT 16009.625 1048.035 16009.905 1193.79 ;
      RECT 16009.065 1048.035 16009.345 1194.03 ;
      RECT 16008.505 1048.035 16008.785 1194.27 ;
      RECT 16007.945 1048.035 16008.225 1194.51 ;
      RECT 16007.385 1048.035 16007.665 1194.75 ;
      RECT 16006.825 1048.035 16007.105 1194.75 ;
      RECT 16006.265 1046.935 16006.545 1194.51 ;
      RECT 16005.705 1048.035 16005.985 1194.27 ;
      RECT 16005.145 1046.935 16005.425 1194.03 ;
      RECT 16004.585 1048.035 16004.865 1193.79 ;
      RECT 16004.025 1048.035 16004.305 1193.55 ;
      RECT 16003.465 1048.035 16003.745 1193.31 ;
      RECT 16002.905 1046.935 16003.185 1193.045 ;
      RECT 16002.345 1048.035 16002.625 1192.805 ;
      RECT 16001.785 1046.935 16002.065 1192.565 ;
      RECT 16001.225 1048.035 16001.505 1192.325 ;
      RECT 15992.265 1046.935 15992.545 1186.16 ;
      RECT 15991.705 1048.035 15991.985 1186.4 ;
      RECT 15991.145 1048.035 15991.425 1186.64 ;
      RECT 15990.585 1048.035 15990.865 1186.64 ;
      RECT 15990.025 1048.035 15990.305 1186.4 ;
      RECT 15989.465 1048.035 15989.745 1186.16 ;
      RECT 15988.905 1048.035 15989.185 1185.92 ;
      RECT 15988.345 1048.035 15988.625 1185.68 ;
      RECT 15987.785 1048.035 15988.065 1185.44 ;
      RECT 15987.225 1048.035 15987.505 1185.2 ;
      RECT 15986.665 1048.035 15986.945 1184.96 ;
      RECT 15986.105 1048.035 15986.385 1184.72 ;
      RECT 15985.545 1048.035 15985.825 1184.48 ;
      RECT 15984.985 1046.935 15985.265 1184.24 ;
      RECT 15982.465 1048.035 15982.745 1185.96 ;
      RECT 15981.905 1046.935 15982.185 1185.72 ;
      RECT 15981.345 1048.035 15981.625 1185.48 ;
      RECT 15980.785 1046.935 15981.065 1185.24 ;
      RECT 15980.225 1048.035 15980.505 1185 ;
      RECT 15979.665 1048.035 15979.945 1184.76 ;
      RECT 15979.105 1048.035 15979.385 1184.52 ;
      RECT 15953.065 1048.035 15953.345 1187.305 ;
      RECT 15952.505 1048.035 15952.785 1187.545 ;
      RECT 15951.945 1048.035 15952.225 1187.785 ;
      RECT 15951.385 1048.035 15951.665 1188.025 ;
      RECT 15950.825 1048.035 15951.105 1188.265 ;
      RECT 15950.265 1046.935 15950.545 1188.505 ;
      RECT 15949.705 1048.035 15949.985 1188.745 ;
      RECT 15949.145 1046.935 15949.425 1188.985 ;
      RECT 15948.585 1048.035 15948.865 1189.225 ;
      RECT 15948.025 1048.035 15948.305 1189.465 ;
      RECT 15947.465 1048.035 15947.745 1189.705 ;
      RECT 15946.905 1048.035 15947.185 1189.945 ;
      RECT 15946.345 1048.035 15946.625 1190.185 ;
      RECT 15945.785 1048.035 15946.065 1190.425 ;
      RECT 15945.225 1048.035 15945.505 1190.665 ;
      RECT 15944.665 1048.035 15944.945 1190.665 ;
      RECT 15944.105 1048.035 15944.385 1190.425 ;
      RECT 15943.545 1048.035 15943.825 1190.185 ;
      RECT 15942.985 1048.035 15943.265 1189.945 ;
      RECT 15942.425 1048.035 15942.705 1189.7 ;
      RECT 15941.865 1048.035 15942.145 1189.46 ;
      RECT 15941.305 1048.035 15941.585 1189.22 ;
      RECT 15940.745 1046.935 15941.025 1188.98 ;
      RECT 15940.185 1048.035 15940.465 1188.74 ;
      RECT 15926.745 1046.935 15927.025 1186.22 ;
      RECT 15926.185 1048.035 15926.465 1185.98 ;
      RECT 15925.625 1048.035 15925.905 1185.74 ;
      RECT 15925.065 1048.035 15925.345 1185.5 ;
      RECT 15924.505 1046.935 15924.785 1185.26 ;
      RECT 15923.945 1048.035 15924.225 1185.02 ;
      RECT 15923.385 1046.935 15923.665 1184.78 ;
      RECT 15922.825 1048.035 15923.105 1184.54 ;
      RECT 15922.265 1046.935 15922.545 1184.3 ;
      RECT 15921.705 1048.035 15921.985 1184.06 ;
      RECT 15921.145 1048.035 15921.425 1183.82 ;
      RECT 15920.585 1048.035 15920.865 1183.58 ;
      RECT 15920.025 1048.035 15920.305 1183.34 ;
      RECT 15919.465 1048.035 15919.745 1183.1 ;
      RECT 15918.905 1048.035 15919.185 1182.86 ;
      RECT 15918.345 1048.035 15918.625 1182.62 ;
      RECT 15917.785 1048.035 15918.065 1182.38 ;
      RECT 15917.225 1048.035 15917.505 1182.14 ;
      RECT 15916.665 1048.035 15916.945 1181.9 ;
      RECT 15916.105 1048.035 15916.385 1181.66 ;
      RECT 15915.545 1048.035 15915.825 1181.42 ;
      RECT 15914.985 1046.935 15915.265 1181.18 ;
      RECT 15914.425 1048.035 15914.705 1180.94 ;
      RECT 15913.865 1046.935 15914.145 1180.7 ;
      RECT 15874.105 1048.035 15874.385 1191.17 ;
      RECT 15873.545 1046.935 15873.825 1191.41 ;
      RECT 15872.985 1048.035 15873.265 1191.65 ;
      RECT 15872.425 1048.035 15872.705 1191.89 ;
      RECT 15871.865 1048.035 15872.145 1192.13 ;
      RECT 15871.305 1048.035 15871.585 1192.37 ;
      RECT 15870.745 1048.035 15871.025 1192.61 ;
      RECT 15870.185 1048.035 15870.465 1192.855 ;
      RECT 15869.625 1048.035 15869.905 1193.095 ;
      RECT 15869.065 1048.035 15869.345 1193.335 ;
      RECT 15868.505 1046.935 15868.785 1193.575 ;
      RECT 15867.945 1048.035 15868.225 1193.815 ;
      RECT 15867.385 1046.935 15867.665 1194.055 ;
      RECT 15866.825 1048.035 15867.105 1194.295 ;
      RECT 15866.265 1048.035 15866.545 1194.535 ;
      RECT 15865.705 1048.035 15865.985 1194.775 ;
      RECT 15865.145 1048.035 15865.425 1195.015 ;
      RECT 15864.585 1048.035 15864.865 1195.255 ;
      RECT 15864.025 1048.035 15864.305 1195.495 ;
      RECT 15863.465 1048.035 15863.745 1195.735 ;
      RECT 15862.905 1048.035 15863.185 1195.975 ;
      RECT 15862.345 1048.035 15862.625 1196.215 ;
      RECT 15861.785 1048.035 15862.065 1196.455 ;
      RECT 15861.225 1048.035 15861.505 1196.695 ;
      RECT 15852.265 1048.035 15852.545 1192.28 ;
      RECT 15851.705 1048.035 15851.985 1192.04 ;
      RECT 15851.145 1048.035 15851.425 1191.8 ;
      RECT 15850.585 1046.935 15850.865 1191.56 ;
      RECT 15850.025 1048.035 15850.305 1191.32 ;
      RECT 15849.465 1046.935 15849.745 1191.08 ;
      RECT 15848.905 1048.035 15849.185 1190.84 ;
      RECT 15848.345 1048.035 15848.625 1190.6 ;
      RECT 15847.785 1048.035 15848.065 1190.36 ;
      RECT 15847.225 1046.935 15847.505 1190.12 ;
      RECT 15846.665 1048.035 15846.945 1189.88 ;
      RECT 15846.105 1046.935 15846.385 1189.64 ;
      RECT 15845.545 1048.035 15845.825 1189.4 ;
      RECT 15844.985 1046.935 15845.265 1189.16 ;
      RECT 15842.465 1048.035 15842.745 1181.56 ;
      RECT 15841.905 1048.035 15842.185 1181.32 ;
      RECT 15841.345 1048.035 15841.625 1181.08 ;
      RECT 15840.785 1048.035 15841.065 1180.84 ;
      RECT 15840.225 1048.035 15840.505 1180.6 ;
      RECT 15839.665 1048.035 15839.945 1180.36 ;
      RECT 15839.105 1048.035 15839.385 1180.12 ;
      RECT 15813.065 1048.035 15813.345 1193.995 ;
      RECT 15812.505 1048.035 15812.785 1194.235 ;
      RECT 15811.945 1048.035 15812.225 1194.475 ;
      RECT 15811.385 1048.035 15811.665 1194.715 ;
      RECT 15810.825 1048.035 15811.105 1194.955 ;
      RECT 15810.265 1046.935 15810.545 1194.955 ;
      RECT 15809.705 1048.035 15809.985 1194.715 ;
      RECT 15809.145 1046.935 15809.425 1194.47 ;
      RECT 15808.585 1048.035 15808.865 1194.23 ;
      RECT 15808.025 1046.935 15808.305 1193.99 ;
      RECT 15807.465 1048.035 15807.745 1193.75 ;
      RECT 15806.905 1048.035 15807.185 1193.51 ;
      RECT 15806.345 1048.035 15806.625 1193.27 ;
      RECT 15805.785 1048.035 15806.065 1193.03 ;
      RECT 15805.225 1048.035 15805.505 1192.79 ;
      RECT 15804.665 1048.035 15804.945 1192.55 ;
      RECT 15804.105 1048.035 15804.385 1192.31 ;
      RECT 15803.545 1048.035 15803.825 1192.07 ;
      RECT 15802.985 1046.935 15803.265 1191.83 ;
      RECT 15802.425 1048.035 15802.705 1191.59 ;
      RECT 15801.865 1046.935 15802.145 1191.35 ;
      RECT 15801.305 1048.035 15801.585 1191.11 ;
      RECT 15800.745 1048.035 15801.025 1190.87 ;
      RECT 15800.185 1048.035 15800.465 1190.63 ;
      RECT 15786.745 1048.035 15787.025 1194.03 ;
      RECT 15786.185 1048.035 15786.465 1194.27 ;
      RECT 15785.625 1048.035 15785.905 1194.515 ;
      RECT 15785.065 1048.035 15785.345 1194.755 ;
      RECT 15784.505 1048.035 15784.785 1194.995 ;
      RECT 15783.945 1048.035 15784.225 1194.995 ;
      RECT 15783.385 1048.035 15783.665 1194.755 ;
      RECT 15782.825 1048.035 15783.105 1194.515 ;
      RECT 15782.265 1048.035 15782.545 1187.5 ;
      RECT 15781.705 1048.035 15781.985 1187.26 ;
      RECT 15781.145 1048.035 15781.425 1187.02 ;
      RECT 15780.585 1046.935 15780.865 1186.78 ;
      RECT 15780.025 1048.035 15780.305 1186.54 ;
      RECT 15779.465 1046.935 15779.745 1186.3 ;
      RECT 15778.905 1048.035 15779.185 1186.06 ;
      RECT 15778.345 1048.035 15778.625 1185.82 ;
      RECT 15777.785 1048.035 15778.065 1185.58 ;
      RECT 15777.225 1046.935 15777.505 1185.34 ;
      RECT 15776.665 1048.035 15776.945 1185.1 ;
      RECT 15776.105 1046.935 15776.385 1184.86 ;
      RECT 15775.545 1048.035 15775.825 1184.62 ;
      RECT 15774.985 1046.935 15775.265 1184.38 ;
      RECT 15774.425 1048.035 15774.705 1184.14 ;
      RECT 15773.865 1048.035 15774.145 1183.9 ;
      RECT 15733.545 1048.035 15733.825 1192.795 ;
      RECT 15732.985 1048.035 15733.265 1193.035 ;
      RECT 15732.425 1048.035 15732.705 1193.28 ;
      RECT 15731.865 1048.035 15732.145 1193.52 ;
      RECT 15731.305 1048.035 15731.585 1193.76 ;
      RECT 15730.745 1048.035 15731.025 1194 ;
      RECT 15730.185 1048.035 15730.465 1194.24 ;
      RECT 15729.625 1048.035 15729.905 1194.48 ;
      RECT 15729.065 1048.035 15729.345 1194.72 ;
      RECT 15728.505 1048.035 15728.785 1194.96 ;
      RECT 15727.945 1046.935 15728.225 1195.2 ;
      RECT 15727.385 1048.035 15727.665 1195.44 ;
      RECT 15726.825 1046.935 15727.105 1195.68 ;
      RECT 15726.265 1048.035 15726.545 1195.92 ;
      RECT 15725.705 1046.935 15725.985 1196.16 ;
      RECT 15725.145 1048.035 15725.425 1196.16 ;
      RECT 15724.585 1048.035 15724.865 1195.92 ;
      RECT 15724.025 1048.035 15724.305 1195.68 ;
      RECT 15723.465 1048.035 15723.745 1195.44 ;
      RECT 15722.905 1048.035 15723.185 1195.2 ;
      RECT 15722.345 1048.035 15722.625 1194.96 ;
      RECT 15721.785 1048.035 15722.065 1194.72 ;
      RECT 15721.225 1048.035 15721.505 1194.48 ;
      RECT 15712.265 1046.935 15712.545 1194.51 ;
      RECT 15711.705 1048.035 15711.985 1194.75 ;
      RECT 15711.145 1046.935 15711.425 1194.99 ;
      RECT 15710.585 1048.035 15710.865 1195.205 ;
      RECT 15710.025 1048.035 15710.305 1194.78 ;
      RECT 15709.465 1048.035 15709.745 1194.54 ;
      RECT 15708.905 1048.035 15709.185 1194.3 ;
      RECT 15708.345 1048.035 15708.625 1194.06 ;
      RECT 15707.785 1048.035 15708.065 1193.82 ;
      RECT 15707.225 1048.035 15707.505 1193.58 ;
      RECT 15706.665 1048.035 15706.945 1193.34 ;
      RECT 15706.105 1048.035 15706.385 1193.1 ;
      RECT 15705.545 1048.035 15705.825 1192.86 ;
      RECT 15704.985 1048.035 15705.265 1192.62 ;
      RECT 15702.465 1048.035 15702.745 1191.795 ;
      RECT 15701.905 1048.035 15702.185 1191.555 ;
      RECT 15701.345 1048.035 15701.625 1191.315 ;
      RECT 15700.785 1046.935 15701.065 1191.075 ;
      RECT 15700.225 1048.035 15700.505 1190.835 ;
      RECT 15699.665 1046.935 15699.945 1190.595 ;
      RECT 15699.105 1048.035 15699.385 1190.355 ;
      RECT 15698.545 1048.035 15698.825 1190.115 ;
      RECT 15671.945 1048.035 15672.225 1201.16 ;
      RECT 15671.385 1046.935 15671.665 1201.4 ;
      RECT 15670.825 1048.035 15671.105 1201.64 ;
      RECT 15670.265 1046.935 15670.545 1201.885 ;
      RECT 15669.705 1048.035 15669.985 1202.125 ;
      RECT 15669.145 1046.935 15669.425 1202.365 ;
      RECT 15668.585 1048.035 15668.865 1202.605 ;
      RECT 15668.025 1048.035 15668.305 1202.845 ;
      RECT 15667.465 1048.035 15667.745 1188.465 ;
      RECT 15666.905 1048.035 15667.185 1188.225 ;
      RECT 15666.345 1048.035 15666.625 1187.985 ;
      RECT 15665.785 1048.035 15666.065 1187.745 ;
      RECT 15665.225 1048.035 15665.505 1187.505 ;
      RECT 15664.665 1048.035 15664.945 1187.265 ;
      RECT 15664.105 1048.035 15664.385 1187.025 ;
      RECT 15663.545 1048.035 15663.825 1186.785 ;
      RECT 15662.985 1048.035 15663.265 1186.545 ;
      RECT 15662.425 1048.035 15662.705 1186.305 ;
      RECT 15661.865 1046.935 15662.145 1186.065 ;
      RECT 15661.305 1048.035 15661.585 1185.825 ;
      RECT 15660.745 1046.935 15661.025 1185.585 ;
      RECT 15660.185 1048.035 15660.465 1185.345 ;
      RECT 15646.185 1046.935 15646.465 1191.465 ;
      RECT 15645.625 1048.035 15645.905 1191.225 ;
      RECT 15645.065 1048.035 15645.345 1190.985 ;
      RECT 15644.505 1048.035 15644.785 1190.745 ;
      RECT 15643.945 1048.035 15644.225 1190.505 ;
      RECT 15643.385 1048.035 15643.665 1190.265 ;
      RECT 15642.825 1048.035 15643.105 1190.025 ;
      RECT 15642.265 1048.035 15642.545 1189.785 ;
      RECT 15641.705 1048.035 15641.985 1189.545 ;
      RECT 15641.145 1046.935 15641.425 1189.305 ;
      RECT 15640.585 1048.035 15640.865 1189.065 ;
      RECT 15640.025 1046.935 15640.305 1188.825 ;
      RECT 15639.465 1048.035 15639.745 1188.585 ;
      RECT 15638.905 1048.035 15639.185 1188.345 ;
      RECT 15638.345 1048.035 15638.625 1188.105 ;
      RECT 15637.785 1048.035 15638.065 1187.865 ;
      RECT 15637.225 1048.035 15637.505 1187.625 ;
      RECT 15636.665 1048.035 15636.945 1187.385 ;
      RECT 15636.105 1048.035 15636.385 1187.145 ;
      RECT 15635.545 1048.035 15635.825 1186.905 ;
      RECT 15634.985 1048.035 15635.265 1186.665 ;
      RECT 15634.425 1048.035 15634.705 1186.425 ;
      RECT 15633.865 1048.035 15634.145 1186.185 ;
      RECT 15594.665 1048.035 15594.945 1193.09 ;
      RECT 15594.105 1048.035 15594.385 1193.33 ;
      RECT 15593.545 1048.035 15593.825 1193.57 ;
      RECT 15592.985 1046.935 15593.265 1193.81 ;
      RECT 15592.425 1048.035 15592.705 1194.05 ;
      RECT 15591.865 1046.935 15592.145 1194.29 ;
      RECT 15591.305 1048.035 15591.585 1194.53 ;
      RECT 15590.745 1048.035 15591.025 1194.77 ;
      RECT 15590.185 1048.035 15590.465 1195.01 ;
      RECT 15589.625 1046.935 15589.905 1195.25 ;
      RECT 15589.065 1048.035 15589.345 1195.49 ;
      RECT 15588.505 1046.935 15588.785 1195.73 ;
      RECT 15587.945 1048.035 15588.225 1195.97 ;
      RECT 15587.385 1046.935 15587.665 1196.21 ;
      RECT 15586.825 1048.035 15587.105 1196.45 ;
      RECT 15586.265 1048.035 15586.545 1196.69 ;
      RECT 15585.705 1048.035 15585.985 1196.69 ;
      RECT 15585.145 1048.035 15585.425 1196.45 ;
      RECT 15584.585 1048.035 15584.865 1196.21 ;
      RECT 15584.025 1048.035 15584.305 1195.97 ;
      RECT 15583.465 1048.035 15583.745 1195.73 ;
      RECT 15582.905 1048.035 15583.185 1195.49 ;
      RECT 15582.345 1048.035 15582.625 1195.25 ;
      RECT 15581.785 1048.035 15582.065 1195.01 ;
      RECT 15581.225 1048.035 15581.505 1194.77 ;
      RECT 15572.265 1048.035 15572.545 1194.285 ;
      RECT 15571.705 1046.935 15571.985 1194.045 ;
      RECT 15571.145 1048.035 15571.425 1193.805 ;
      RECT 15570.585 1046.935 15570.865 1193.565 ;
      RECT 15570.025 1048.035 15570.305 1193.325 ;
      RECT 15569.465 1046.935 15569.745 1193.085 ;
      RECT 15568.905 1048.035 15569.185 1192.845 ;
      RECT 15568.345 1048.035 15568.625 1192.605 ;
      RECT 15567.785 1048.035 15568.065 1192.365 ;
      RECT 15567.225 1048.035 15567.505 1192.125 ;
      RECT 15566.665 1048.035 15566.945 1191.885 ;
      RECT 15566.105 1048.035 15566.385 1191.645 ;
      RECT 15565.545 1048.035 15565.825 1191.405 ;
      RECT 15564.985 1048.035 15565.265 1191.165 ;
      RECT 15562.465 1046.935 15562.745 1192.885 ;
      RECT 15561.905 1048.035 15562.185 1192.645 ;
      RECT 15561.345 1046.935 15561.625 1192.405 ;
      RECT 15560.785 1048.035 15561.065 1192.165 ;
      RECT 15560.225 1048.035 15560.505 1191.925 ;
      RECT 15559.665 1048.035 15559.945 1191.685 ;
      RECT 15559.105 1048.035 15559.385 1191.445 ;
      RECT 15558.545 1048.035 15558.825 1191.205 ;
      RECT 15532.505 1048.035 15532.785 1188.855 ;
      RECT 15531.945 1048.035 15532.225 1189.095 ;
      RECT 15531.385 1048.035 15531.665 1189.335 ;
      RECT 15530.825 1048.035 15531.105 1189.58 ;
      RECT 15530.265 1048.035 15530.545 1189.82 ;
      RECT 15529.705 1048.035 15529.985 1190.06 ;
      RECT 15529.145 1048.035 15529.425 1190.06 ;
      RECT 15528.585 1048.035 15528.865 1189.82 ;
      RECT 15528.025 1048.035 15528.305 1189.58 ;
      RECT 15527.465 1046.935 15527.745 1189.34 ;
      RECT 15526.905 1048.035 15527.185 1189.1 ;
      RECT 15526.345 1046.935 15526.625 1188.86 ;
      RECT 15525.785 1048.035 15526.065 1188.62 ;
      RECT 15525.225 1048.035 15525.505 1188.38 ;
      RECT 15524.665 1048.035 15524.945 1188.14 ;
      RECT 15524.105 1046.935 15524.385 1187.9 ;
      RECT 15523.545 1048.035 15523.825 1187.66 ;
      RECT 15522.985 1046.935 15523.265 1187.42 ;
      RECT 15522.425 1048.035 15522.705 1187.18 ;
      RECT 15521.865 1046.935 15522.145 1186.94 ;
      RECT 15521.305 1048.035 15521.585 1186.7 ;
      RECT 15520.745 1048.035 15521.025 1186.46 ;
      RECT 15520.185 1048.035 15520.465 1186.22 ;
      RECT 15519.625 1048.035 15519.905 1185.98 ;
      RECT 15506.185 1048.035 15506.465 1191.78 ;
      RECT 15505.625 1048.035 15505.905 1191.54 ;
      RECT 15505.065 1048.035 15505.345 1191.3 ;
      RECT 15504.505 1048.035 15504.785 1191.06 ;
      RECT 15503.945 1048.035 15504.225 1190.82 ;
      RECT 15503.385 1048.035 15503.665 1190.58 ;
      RECT 15502.825 1048.035 15503.105 1190.34 ;
      RECT 15502.265 1048.035 15502.545 1190.1 ;
      RECT 15501.705 1046.935 15501.985 1189.86 ;
      RECT 15501.145 1048.035 15501.425 1189.62 ;
      RECT 15500.585 1046.935 15500.865 1189.3 ;
      RECT 15500.025 1048.035 15500.305 1189.14 ;
      RECT 15499.465 1046.935 15499.745 1188.9 ;
      RECT 15498.905 1048.035 15499.185 1188.66 ;
      RECT 15498.345 1048.035 15498.625 1188.42 ;
      RECT 15497.785 1048.035 15498.065 1188.18 ;
      RECT 15497.225 1048.035 15497.505 1187.94 ;
      RECT 15496.665 1048.035 15496.945 1187.7 ;
      RECT 15496.105 1048.035 15496.385 1187.46 ;
      RECT 15495.545 1048.035 15495.825 1187.22 ;
      RECT 15494.985 1048.035 15495.265 1186.98 ;
      RECT 15494.425 1046.935 15494.705 1186.74 ;
      RECT 15493.865 1048.035 15494.145 1186.5 ;
      RECT 15493.305 1046.935 15493.585 1186.26 ;
      RECT 15454.105 1048.035 15454.385 1191.87 ;
      RECT 15453.545 1048.035 15453.825 1192.11 ;
      RECT 15452.985 1048.035 15453.265 1192.35 ;
      RECT 15452.425 1048.035 15452.705 1192.59 ;
      RECT 15451.865 1048.035 15452.145 1192.83 ;
      RECT 15451.305 1048.035 15451.585 1193.07 ;
      RECT 15450.745 1048.035 15451.025 1193.31 ;
      RECT 15450.185 1048.035 15450.465 1193.55 ;
      RECT 15449.625 1048.035 15449.905 1193.79 ;
      RECT 15449.065 1048.035 15449.345 1194.03 ;
      RECT 15448.505 1048.035 15448.785 1194.27 ;
      RECT 15447.945 1048.035 15448.225 1194.51 ;
      RECT 15447.385 1048.035 15447.665 1194.75 ;
      RECT 15446.825 1048.035 15447.105 1194.75 ;
      RECT 15446.265 1046.935 15446.545 1194.51 ;
      RECT 15445.705 1048.035 15445.985 1194.27 ;
      RECT 15445.145 1046.935 15445.425 1194.03 ;
      RECT 15444.585 1048.035 15444.865 1193.79 ;
      RECT 15444.025 1048.035 15444.305 1193.55 ;
      RECT 15443.465 1048.035 15443.745 1193.31 ;
      RECT 15442.905 1046.935 15443.185 1193.045 ;
      RECT 15442.345 1048.035 15442.625 1192.805 ;
      RECT 15441.785 1046.935 15442.065 1192.565 ;
      RECT 15441.225 1048.035 15441.505 1192.325 ;
      RECT 15432.265 1046.935 15432.545 1186.16 ;
      RECT 15431.705 1048.035 15431.985 1186.4 ;
      RECT 15431.145 1048.035 15431.425 1186.64 ;
      RECT 15430.585 1048.035 15430.865 1186.64 ;
      RECT 15430.025 1048.035 15430.305 1186.4 ;
      RECT 15429.465 1048.035 15429.745 1186.16 ;
      RECT 15428.905 1048.035 15429.185 1185.92 ;
      RECT 15428.345 1048.035 15428.625 1185.68 ;
      RECT 15427.785 1048.035 15428.065 1185.44 ;
      RECT 15427.225 1048.035 15427.505 1185.2 ;
      RECT 15426.665 1048.035 15426.945 1184.96 ;
      RECT 15426.105 1048.035 15426.385 1184.72 ;
      RECT 15425.545 1048.035 15425.825 1184.48 ;
      RECT 15424.985 1046.935 15425.265 1184.24 ;
      RECT 15422.465 1048.035 15422.745 1185.96 ;
      RECT 15421.905 1046.935 15422.185 1185.72 ;
      RECT 15421.345 1048.035 15421.625 1185.48 ;
      RECT 15420.785 1046.935 15421.065 1185.24 ;
      RECT 15420.225 1048.035 15420.505 1185 ;
      RECT 15419.665 1048.035 15419.945 1184.76 ;
      RECT 15419.105 1048.035 15419.385 1184.52 ;
      RECT 15393.065 1048.035 15393.345 1187.305 ;
      RECT 15392.505 1048.035 15392.785 1187.545 ;
      RECT 15391.945 1048.035 15392.225 1187.785 ;
      RECT 15391.385 1048.035 15391.665 1188.025 ;
      RECT 15390.825 1048.035 15391.105 1188.265 ;
      RECT 15390.265 1046.935 15390.545 1188.505 ;
      RECT 15389.705 1048.035 15389.985 1188.745 ;
      RECT 15389.145 1046.935 15389.425 1188.985 ;
      RECT 15388.585 1048.035 15388.865 1189.225 ;
      RECT 15388.025 1048.035 15388.305 1189.465 ;
      RECT 15387.465 1048.035 15387.745 1189.705 ;
      RECT 15386.905 1048.035 15387.185 1189.945 ;
      RECT 15386.345 1048.035 15386.625 1190.185 ;
      RECT 15385.785 1048.035 15386.065 1190.425 ;
      RECT 15385.225 1048.035 15385.505 1190.665 ;
      RECT 15384.665 1048.035 15384.945 1190.665 ;
      RECT 15384.105 1048.035 15384.385 1190.425 ;
      RECT 15383.545 1048.035 15383.825 1190.185 ;
      RECT 15382.985 1048.035 15383.265 1189.945 ;
      RECT 15382.425 1048.035 15382.705 1189.7 ;
      RECT 15381.865 1048.035 15382.145 1189.46 ;
      RECT 15381.305 1048.035 15381.585 1189.22 ;
      RECT 15380.745 1046.935 15381.025 1188.98 ;
      RECT 15380.185 1048.035 15380.465 1188.74 ;
      RECT 15366.745 1046.935 15367.025 1186.22 ;
      RECT 15366.185 1048.035 15366.465 1185.98 ;
      RECT 15365.625 1048.035 15365.905 1185.74 ;
      RECT 15365.065 1048.035 15365.345 1185.5 ;
      RECT 15364.505 1046.935 15364.785 1185.26 ;
      RECT 15363.945 1048.035 15364.225 1185.02 ;
      RECT 15363.385 1046.935 15363.665 1184.78 ;
      RECT 15362.825 1048.035 15363.105 1184.54 ;
      RECT 15362.265 1046.935 15362.545 1184.3 ;
      RECT 15361.705 1048.035 15361.985 1184.06 ;
      RECT 15361.145 1048.035 15361.425 1183.82 ;
      RECT 15360.585 1048.035 15360.865 1183.58 ;
      RECT 15360.025 1048.035 15360.305 1183.34 ;
      RECT 15359.465 1048.035 15359.745 1183.1 ;
      RECT 15358.905 1048.035 15359.185 1182.86 ;
      RECT 15358.345 1048.035 15358.625 1182.62 ;
      RECT 15357.785 1048.035 15358.065 1182.38 ;
      RECT 15357.225 1048.035 15357.505 1182.14 ;
      RECT 15356.665 1048.035 15356.945 1181.9 ;
      RECT 15356.105 1048.035 15356.385 1181.66 ;
      RECT 15355.545 1048.035 15355.825 1181.42 ;
      RECT 15354.985 1046.935 15355.265 1181.18 ;
      RECT 15354.425 1048.035 15354.705 1180.94 ;
      RECT 15353.865 1046.935 15354.145 1180.7 ;
      RECT 15314.105 1048.035 15314.385 1191.17 ;
      RECT 15313.545 1046.935 15313.825 1191.41 ;
      RECT 15312.985 1048.035 15313.265 1191.65 ;
      RECT 15312.425 1048.035 15312.705 1191.89 ;
      RECT 15311.865 1048.035 15312.145 1192.13 ;
      RECT 15311.305 1048.035 15311.585 1192.37 ;
      RECT 15310.745 1048.035 15311.025 1192.61 ;
      RECT 15310.185 1048.035 15310.465 1192.855 ;
      RECT 15309.625 1048.035 15309.905 1193.095 ;
      RECT 15309.065 1048.035 15309.345 1193.335 ;
      RECT 15308.505 1046.935 15308.785 1193.575 ;
      RECT 15307.945 1048.035 15308.225 1193.815 ;
      RECT 15307.385 1046.935 15307.665 1194.055 ;
      RECT 15306.825 1048.035 15307.105 1194.295 ;
      RECT 15306.265 1048.035 15306.545 1194.535 ;
      RECT 15305.705 1048.035 15305.985 1194.775 ;
      RECT 15305.145 1048.035 15305.425 1195.015 ;
      RECT 15304.585 1048.035 15304.865 1195.255 ;
      RECT 15304.025 1048.035 15304.305 1195.495 ;
      RECT 15303.465 1048.035 15303.745 1195.735 ;
      RECT 15302.905 1048.035 15303.185 1195.975 ;
      RECT 15302.345 1048.035 15302.625 1196.215 ;
      RECT 15301.785 1048.035 15302.065 1196.455 ;
      RECT 15301.225 1048.035 15301.505 1196.695 ;
      RECT 15292.265 1048.035 15292.545 1192.28 ;
      RECT 15291.705 1048.035 15291.985 1192.04 ;
      RECT 15291.145 1048.035 15291.425 1191.8 ;
      RECT 15290.585 1046.935 15290.865 1191.56 ;
      RECT 15290.025 1048.035 15290.305 1191.32 ;
      RECT 15289.465 1046.935 15289.745 1191.08 ;
      RECT 15288.905 1048.035 15289.185 1190.84 ;
      RECT 15288.345 1048.035 15288.625 1190.6 ;
      RECT 15287.785 1048.035 15288.065 1190.36 ;
      RECT 15287.225 1046.935 15287.505 1190.12 ;
      RECT 15286.665 1048.035 15286.945 1189.88 ;
      RECT 15286.105 1046.935 15286.385 1189.64 ;
      RECT 15285.545 1048.035 15285.825 1189.4 ;
      RECT 15284.985 1046.935 15285.265 1189.16 ;
      RECT 15282.465 1048.035 15282.745 1181.56 ;
      RECT 15281.905 1048.035 15282.185 1181.32 ;
      RECT 15281.345 1048.035 15281.625 1181.08 ;
      RECT 15280.785 1048.035 15281.065 1180.84 ;
      RECT 15280.225 1048.035 15280.505 1180.6 ;
      RECT 15279.665 1048.035 15279.945 1180.36 ;
      RECT 15279.105 1048.035 15279.385 1180.12 ;
      RECT 15253.065 1048.035 15253.345 1193.995 ;
      RECT 15252.505 1048.035 15252.785 1194.235 ;
      RECT 15251.945 1048.035 15252.225 1194.475 ;
      RECT 15251.385 1048.035 15251.665 1194.715 ;
      RECT 15250.825 1048.035 15251.105 1194.955 ;
      RECT 15250.265 1046.935 15250.545 1194.955 ;
      RECT 15249.705 1048.035 15249.985 1194.715 ;
      RECT 15249.145 1046.935 15249.425 1194.47 ;
      RECT 15248.585 1048.035 15248.865 1194.23 ;
      RECT 15248.025 1046.935 15248.305 1193.99 ;
      RECT 15247.465 1048.035 15247.745 1193.75 ;
      RECT 15246.905 1048.035 15247.185 1193.51 ;
      RECT 15246.345 1048.035 15246.625 1193.27 ;
      RECT 15245.785 1048.035 15246.065 1193.03 ;
      RECT 15245.225 1048.035 15245.505 1192.79 ;
      RECT 15244.665 1048.035 15244.945 1192.55 ;
      RECT 15244.105 1048.035 15244.385 1192.31 ;
      RECT 15243.545 1048.035 15243.825 1192.07 ;
      RECT 15242.985 1046.935 15243.265 1191.83 ;
      RECT 15242.425 1048.035 15242.705 1191.59 ;
      RECT 15241.865 1046.935 15242.145 1191.35 ;
      RECT 15241.305 1048.035 15241.585 1191.11 ;
      RECT 15240.745 1048.035 15241.025 1190.87 ;
      RECT 15240.185 1048.035 15240.465 1190.63 ;
      RECT 15226.745 1048.035 15227.025 1194.03 ;
      RECT 15226.185 1048.035 15226.465 1194.27 ;
      RECT 15225.625 1048.035 15225.905 1194.515 ;
      RECT 15225.065 1048.035 15225.345 1194.755 ;
      RECT 15224.505 1048.035 15224.785 1194.995 ;
      RECT 15223.945 1048.035 15224.225 1194.995 ;
      RECT 15223.385 1048.035 15223.665 1194.755 ;
      RECT 15222.825 1048.035 15223.105 1194.515 ;
      RECT 15222.265 1048.035 15222.545 1187.5 ;
      RECT 15221.705 1048.035 15221.985 1187.26 ;
      RECT 15221.145 1048.035 15221.425 1187.02 ;
      RECT 15220.585 1046.935 15220.865 1186.78 ;
      RECT 15220.025 1048.035 15220.305 1186.54 ;
      RECT 15219.465 1046.935 15219.745 1186.3 ;
      RECT 15218.905 1048.035 15219.185 1186.06 ;
      RECT 15218.345 1048.035 15218.625 1185.82 ;
      RECT 15217.785 1048.035 15218.065 1185.58 ;
      RECT 15217.225 1046.935 15217.505 1185.34 ;
      RECT 15216.665 1048.035 15216.945 1185.1 ;
      RECT 15216.105 1046.935 15216.385 1184.86 ;
      RECT 15215.545 1048.035 15215.825 1184.62 ;
      RECT 15214.985 1046.935 15215.265 1184.38 ;
      RECT 15214.425 1048.035 15214.705 1184.14 ;
      RECT 15213.865 1048.035 15214.145 1183.9 ;
      RECT 15173.545 1048.035 15173.825 1192.795 ;
      RECT 15172.985 1048.035 15173.265 1193.035 ;
      RECT 15172.425 1048.035 15172.705 1193.28 ;
      RECT 15171.865 1048.035 15172.145 1193.52 ;
      RECT 15171.305 1048.035 15171.585 1193.76 ;
      RECT 15170.745 1048.035 15171.025 1194 ;
      RECT 15170.185 1048.035 15170.465 1194.24 ;
      RECT 15169.625 1048.035 15169.905 1194.48 ;
      RECT 15169.065 1048.035 15169.345 1194.72 ;
      RECT 15168.505 1048.035 15168.785 1194.96 ;
      RECT 15167.945 1046.935 15168.225 1195.2 ;
      RECT 15167.385 1048.035 15167.665 1195.44 ;
      RECT 15166.825 1046.935 15167.105 1195.68 ;
      RECT 15166.265 1048.035 15166.545 1195.92 ;
      RECT 15165.705 1046.935 15165.985 1196.16 ;
      RECT 15165.145 1048.035 15165.425 1196.16 ;
      RECT 15164.585 1048.035 15164.865 1195.92 ;
      RECT 15164.025 1048.035 15164.305 1195.68 ;
      RECT 15163.465 1048.035 15163.745 1195.44 ;
      RECT 15162.905 1048.035 15163.185 1195.2 ;
      RECT 15162.345 1048.035 15162.625 1194.96 ;
      RECT 15161.785 1048.035 15162.065 1194.72 ;
      RECT 15161.225 1048.035 15161.505 1194.48 ;
      RECT 15152.265 1046.935 15152.545 1194.51 ;
      RECT 15151.705 1048.035 15151.985 1194.75 ;
      RECT 15151.145 1046.935 15151.425 1194.99 ;
      RECT 15150.585 1048.035 15150.865 1195.205 ;
      RECT 15150.025 1048.035 15150.305 1194.78 ;
      RECT 15149.465 1048.035 15149.745 1194.54 ;
      RECT 15148.905 1048.035 15149.185 1194.3 ;
      RECT 15148.345 1048.035 15148.625 1194.06 ;
      RECT 15147.785 1048.035 15148.065 1193.82 ;
      RECT 15147.225 1048.035 15147.505 1193.58 ;
      RECT 15146.665 1048.035 15146.945 1193.34 ;
      RECT 15146.105 1048.035 15146.385 1193.1 ;
      RECT 15145.545 1048.035 15145.825 1192.86 ;
      RECT 15144.985 1048.035 15145.265 1192.62 ;
      RECT 15142.465 1048.035 15142.745 1191.795 ;
      RECT 15141.905 1048.035 15142.185 1191.555 ;
      RECT 15141.345 1048.035 15141.625 1191.315 ;
      RECT 15140.785 1046.935 15141.065 1191.075 ;
      RECT 15140.225 1048.035 15140.505 1190.835 ;
      RECT 15139.665 1046.935 15139.945 1190.595 ;
      RECT 15139.105 1048.035 15139.385 1190.355 ;
      RECT 15138.545 1048.035 15138.825 1190.115 ;
      RECT 15111.945 1048.035 15112.225 1201.16 ;
      RECT 15111.385 1046.935 15111.665 1201.4 ;
      RECT 15110.825 1048.035 15111.105 1201.64 ;
      RECT 15110.265 1046.935 15110.545 1201.885 ;
      RECT 15109.705 1048.035 15109.985 1202.125 ;
      RECT 15109.145 1046.935 15109.425 1202.365 ;
      RECT 15108.585 1048.035 15108.865 1202.605 ;
      RECT 15108.025 1048.035 15108.305 1202.845 ;
      RECT 15107.465 1048.035 15107.745 1188.465 ;
      RECT 15106.905 1048.035 15107.185 1188.225 ;
      RECT 15106.345 1048.035 15106.625 1187.985 ;
      RECT 15105.785 1048.035 15106.065 1187.745 ;
      RECT 15105.225 1048.035 15105.505 1187.505 ;
      RECT 15104.665 1048.035 15104.945 1187.265 ;
      RECT 15104.105 1048.035 15104.385 1187.025 ;
      RECT 15103.545 1048.035 15103.825 1186.785 ;
      RECT 15102.985 1048.035 15103.265 1186.545 ;
      RECT 15102.425 1048.035 15102.705 1186.305 ;
      RECT 15101.865 1046.935 15102.145 1186.065 ;
      RECT 15101.305 1048.035 15101.585 1185.825 ;
      RECT 15100.745 1046.935 15101.025 1185.585 ;
      RECT 15100.185 1048.035 15100.465 1185.345 ;
      RECT 15086.185 1046.935 15086.465 1191.465 ;
      RECT 15085.625 1048.035 15085.905 1191.225 ;
      RECT 15085.065 1048.035 15085.345 1190.985 ;
      RECT 15084.505 1048.035 15084.785 1190.745 ;
      RECT 15083.945 1048.035 15084.225 1190.505 ;
      RECT 15083.385 1048.035 15083.665 1190.265 ;
      RECT 15082.825 1048.035 15083.105 1190.025 ;
      RECT 15082.265 1048.035 15082.545 1189.785 ;
      RECT 15081.705 1048.035 15081.985 1189.545 ;
      RECT 15081.145 1046.935 15081.425 1189.305 ;
      RECT 15080.585 1048.035 15080.865 1189.065 ;
      RECT 15080.025 1046.935 15080.305 1188.825 ;
      RECT 15079.465 1048.035 15079.745 1188.585 ;
      RECT 15078.905 1048.035 15079.185 1188.345 ;
      RECT 15078.345 1048.035 15078.625 1188.105 ;
      RECT 15077.785 1048.035 15078.065 1187.865 ;
      RECT 15077.225 1048.035 15077.505 1187.625 ;
      RECT 15076.665 1048.035 15076.945 1187.385 ;
      RECT 15076.105 1048.035 15076.385 1187.145 ;
      RECT 15075.545 1048.035 15075.825 1186.905 ;
      RECT 15074.985 1048.035 15075.265 1186.665 ;
      RECT 15074.425 1048.035 15074.705 1186.425 ;
      RECT 15073.865 1048.035 15074.145 1186.185 ;
      RECT 15034.665 1048.035 15034.945 1193.09 ;
      RECT 15034.105 1048.035 15034.385 1193.33 ;
      RECT 15033.545 1048.035 15033.825 1193.57 ;
      RECT 15032.985 1046.935 15033.265 1193.81 ;
      RECT 15032.425 1048.035 15032.705 1194.05 ;
      RECT 15031.865 1046.935 15032.145 1194.29 ;
      RECT 15031.305 1048.035 15031.585 1194.53 ;
      RECT 15030.745 1048.035 15031.025 1194.77 ;
      RECT 15030.185 1048.035 15030.465 1195.01 ;
      RECT 15029.625 1046.935 15029.905 1195.25 ;
      RECT 15029.065 1048.035 15029.345 1195.49 ;
      RECT 15028.505 1046.935 15028.785 1195.73 ;
      RECT 15027.945 1048.035 15028.225 1195.97 ;
      RECT 15027.385 1046.935 15027.665 1196.21 ;
      RECT 15026.825 1048.035 15027.105 1196.45 ;
      RECT 15026.265 1048.035 15026.545 1196.69 ;
      RECT 15025.705 1048.035 15025.985 1196.69 ;
      RECT 15025.145 1048.035 15025.425 1196.45 ;
      RECT 15024.585 1048.035 15024.865 1196.21 ;
      RECT 15024.025 1048.035 15024.305 1195.97 ;
      RECT 15023.465 1048.035 15023.745 1195.73 ;
      RECT 15022.905 1048.035 15023.185 1195.49 ;
      RECT 15022.345 1048.035 15022.625 1195.25 ;
      RECT 15021.785 1048.035 15022.065 1195.01 ;
      RECT 15021.225 1048.035 15021.505 1194.77 ;
      RECT 15012.265 1048.035 15012.545 1194.285 ;
      RECT 15011.705 1046.935 15011.985 1194.045 ;
      RECT 15011.145 1048.035 15011.425 1193.805 ;
      RECT 15010.585 1046.935 15010.865 1193.565 ;
      RECT 15010.025 1048.035 15010.305 1193.325 ;
      RECT 15009.465 1046.935 15009.745 1193.085 ;
      RECT 15008.905 1048.035 15009.185 1192.845 ;
      RECT 15008.345 1048.035 15008.625 1192.605 ;
      RECT 15007.785 1048.035 15008.065 1192.365 ;
      RECT 15007.225 1048.035 15007.505 1192.125 ;
      RECT 15006.665 1048.035 15006.945 1191.885 ;
      RECT 15006.105 1048.035 15006.385 1191.645 ;
      RECT 15005.545 1048.035 15005.825 1191.405 ;
      RECT 15004.985 1048.035 15005.265 1191.165 ;
      RECT 15002.465 1046.935 15002.745 1192.885 ;
      RECT 15001.905 1048.035 15002.185 1192.645 ;
      RECT 15001.345 1046.935 15001.625 1192.405 ;
      RECT 15000.785 1048.035 15001.065 1192.165 ;
      RECT 15000.225 1048.035 15000.505 1191.925 ;
      RECT 14999.665 1048.035 14999.945 1191.685 ;
      RECT 14999.105 1048.035 14999.385 1191.445 ;
      RECT 14998.545 1048.035 14998.825 1191.205 ;
      RECT 14972.505 1048.035 14972.785 1188.855 ;
      RECT 14971.945 1048.035 14972.225 1189.095 ;
      RECT 14971.385 1048.035 14971.665 1189.335 ;
      RECT 14970.825 1048.035 14971.105 1189.58 ;
      RECT 14970.265 1048.035 14970.545 1189.82 ;
      RECT 14969.705 1048.035 14969.985 1190.06 ;
      RECT 14969.145 1048.035 14969.425 1190.06 ;
      RECT 14968.585 1048.035 14968.865 1189.82 ;
      RECT 14968.025 1048.035 14968.305 1189.58 ;
      RECT 14967.465 1046.935 14967.745 1189.34 ;
      RECT 14966.905 1048.035 14967.185 1189.1 ;
      RECT 14966.345 1046.935 14966.625 1188.86 ;
      RECT 14965.785 1048.035 14966.065 1188.62 ;
      RECT 14965.225 1048.035 14965.505 1188.38 ;
      RECT 14964.665 1048.035 14964.945 1188.14 ;
      RECT 14964.105 1046.935 14964.385 1187.9 ;
      RECT 14963.545 1048.035 14963.825 1187.66 ;
      RECT 14962.985 1046.935 14963.265 1187.42 ;
      RECT 14962.425 1048.035 14962.705 1187.18 ;
      RECT 14961.865 1046.935 14962.145 1186.94 ;
      RECT 14961.305 1048.035 14961.585 1186.7 ;
      RECT 14960.745 1048.035 14961.025 1186.46 ;
      RECT 14960.185 1048.035 14960.465 1186.22 ;
      RECT 14959.625 1048.035 14959.905 1185.98 ;
      RECT 14946.185 1048.035 14946.465 1191.78 ;
      RECT 14945.625 1048.035 14945.905 1191.54 ;
      RECT 14945.065 1048.035 14945.345 1191.3 ;
      RECT 14944.505 1048.035 14944.785 1191.06 ;
      RECT 14943.945 1048.035 14944.225 1190.82 ;
      RECT 14943.385 1048.035 14943.665 1190.58 ;
      RECT 14942.825 1048.035 14943.105 1190.34 ;
      RECT 14942.265 1048.035 14942.545 1190.1 ;
      RECT 14941.705 1046.935 14941.985 1189.86 ;
      RECT 14941.145 1048.035 14941.425 1189.62 ;
      RECT 14940.585 1046.935 14940.865 1189.3 ;
      RECT 14940.025 1048.035 14940.305 1189.14 ;
      RECT 14939.465 1046.935 14939.745 1188.9 ;
      RECT 14938.905 1048.035 14939.185 1188.66 ;
      RECT 14938.345 1048.035 14938.625 1188.42 ;
      RECT 14937.785 1048.035 14938.065 1188.18 ;
      RECT 14937.225 1048.035 14937.505 1187.94 ;
      RECT 14936.665 1048.035 14936.945 1187.7 ;
      RECT 14936.105 1048.035 14936.385 1187.46 ;
      RECT 14935.545 1048.035 14935.825 1187.22 ;
      RECT 14934.985 1048.035 14935.265 1186.98 ;
      RECT 14934.425 1046.935 14934.705 1186.74 ;
      RECT 14933.865 1048.035 14934.145 1186.5 ;
      RECT 14933.305 1046.935 14933.585 1186.26 ;
      RECT 14894.105 1048.035 14894.385 1191.87 ;
      RECT 14893.545 1048.035 14893.825 1192.11 ;
      RECT 14892.985 1048.035 14893.265 1192.35 ;
      RECT 14892.425 1048.035 14892.705 1192.59 ;
      RECT 14891.865 1048.035 14892.145 1192.83 ;
      RECT 14891.305 1048.035 14891.585 1193.07 ;
      RECT 14890.745 1048.035 14891.025 1193.31 ;
      RECT 14890.185 1048.035 14890.465 1193.55 ;
      RECT 14889.625 1048.035 14889.905 1193.79 ;
      RECT 14889.065 1048.035 14889.345 1194.03 ;
      RECT 14888.505 1048.035 14888.785 1194.27 ;
      RECT 14887.945 1048.035 14888.225 1194.51 ;
      RECT 14887.385 1048.035 14887.665 1194.75 ;
      RECT 14886.825 1048.035 14887.105 1194.75 ;
      RECT 14886.265 1046.935 14886.545 1194.51 ;
      RECT 14885.705 1048.035 14885.985 1194.27 ;
      RECT 14885.145 1046.935 14885.425 1194.03 ;
      RECT 14884.585 1048.035 14884.865 1193.79 ;
      RECT 14884.025 1048.035 14884.305 1193.55 ;
      RECT 14883.465 1048.035 14883.745 1193.31 ;
      RECT 14882.905 1046.935 14883.185 1193.045 ;
      RECT 14882.345 1048.035 14882.625 1192.805 ;
      RECT 14881.785 1046.935 14882.065 1192.565 ;
      RECT 14881.225 1048.035 14881.505 1192.325 ;
      RECT 14872.265 1046.935 14872.545 1186.16 ;
      RECT 14871.705 1048.035 14871.985 1186.4 ;
      RECT 14871.145 1048.035 14871.425 1186.64 ;
      RECT 14870.585 1048.035 14870.865 1186.64 ;
      RECT 14870.025 1048.035 14870.305 1186.4 ;
      RECT 14869.465 1048.035 14869.745 1186.16 ;
      RECT 14868.905 1048.035 14869.185 1185.92 ;
      RECT 14868.345 1048.035 14868.625 1185.68 ;
      RECT 14867.785 1048.035 14868.065 1185.44 ;
      RECT 14867.225 1048.035 14867.505 1185.2 ;
      RECT 14866.665 1048.035 14866.945 1184.96 ;
      RECT 14866.105 1048.035 14866.385 1184.72 ;
      RECT 14865.545 1048.035 14865.825 1184.48 ;
      RECT 14864.985 1046.935 14865.265 1184.24 ;
      RECT 14862.465 1048.035 14862.745 1185.96 ;
      RECT 14861.905 1046.935 14862.185 1185.72 ;
      RECT 14861.345 1048.035 14861.625 1185.48 ;
      RECT 14860.785 1046.935 14861.065 1185.24 ;
      RECT 14860.225 1048.035 14860.505 1185 ;
      RECT 14859.665 1048.035 14859.945 1184.76 ;
      RECT 14859.105 1048.035 14859.385 1184.52 ;
      RECT 14833.065 1048.035 14833.345 1187.305 ;
      RECT 14832.505 1048.035 14832.785 1187.545 ;
      RECT 14831.945 1048.035 14832.225 1187.785 ;
      RECT 14831.385 1048.035 14831.665 1188.025 ;
      RECT 14830.825 1048.035 14831.105 1188.265 ;
      RECT 14830.265 1046.935 14830.545 1188.505 ;
      RECT 14829.705 1048.035 14829.985 1188.745 ;
      RECT 14829.145 1046.935 14829.425 1188.985 ;
      RECT 14828.585 1048.035 14828.865 1189.225 ;
      RECT 14828.025 1048.035 14828.305 1189.465 ;
      RECT 14827.465 1048.035 14827.745 1189.705 ;
      RECT 14826.905 1048.035 14827.185 1189.945 ;
      RECT 14826.345 1048.035 14826.625 1190.185 ;
      RECT 14825.785 1048.035 14826.065 1190.425 ;
      RECT 14825.225 1048.035 14825.505 1190.665 ;
      RECT 14824.665 1048.035 14824.945 1190.665 ;
      RECT 14824.105 1048.035 14824.385 1190.425 ;
      RECT 14823.545 1048.035 14823.825 1190.185 ;
      RECT 14822.985 1048.035 14823.265 1189.945 ;
      RECT 14822.425 1048.035 14822.705 1189.7 ;
      RECT 14821.865 1048.035 14822.145 1189.46 ;
      RECT 14821.305 1048.035 14821.585 1189.22 ;
      RECT 14820.745 1046.935 14821.025 1188.98 ;
      RECT 14820.185 1048.035 14820.465 1188.74 ;
      RECT 14806.745 1046.935 14807.025 1186.22 ;
      RECT 14806.185 1048.035 14806.465 1185.98 ;
      RECT 14805.625 1048.035 14805.905 1185.74 ;
      RECT 14805.065 1048.035 14805.345 1185.5 ;
      RECT 14804.505 1046.935 14804.785 1185.26 ;
      RECT 14803.945 1048.035 14804.225 1185.02 ;
      RECT 14803.385 1046.935 14803.665 1184.78 ;
      RECT 14802.825 1048.035 14803.105 1184.54 ;
      RECT 14802.265 1046.935 14802.545 1184.3 ;
      RECT 14801.705 1048.035 14801.985 1184.06 ;
      RECT 14801.145 1048.035 14801.425 1183.82 ;
      RECT 14800.585 1048.035 14800.865 1183.58 ;
      RECT 14800.025 1048.035 14800.305 1183.34 ;
      RECT 14799.465 1048.035 14799.745 1183.1 ;
      RECT 14798.905 1048.035 14799.185 1182.86 ;
      RECT 14798.345 1048.035 14798.625 1182.62 ;
      RECT 14797.785 1048.035 14798.065 1182.38 ;
      RECT 14797.225 1048.035 14797.505 1182.14 ;
      RECT 14796.665 1048.035 14796.945 1181.9 ;
      RECT 14796.105 1048.035 14796.385 1181.66 ;
      RECT 14795.545 1048.035 14795.825 1181.42 ;
      RECT 14794.985 1046.935 14795.265 1181.18 ;
      RECT 14794.425 1048.035 14794.705 1180.94 ;
      RECT 14793.865 1046.935 14794.145 1180.7 ;
      RECT 14754.105 1048.035 14754.385 1191.17 ;
      RECT 14753.545 1046.935 14753.825 1191.41 ;
      RECT 14752.985 1048.035 14753.265 1191.65 ;
      RECT 14752.425 1048.035 14752.705 1191.89 ;
      RECT 14751.865 1048.035 14752.145 1192.13 ;
      RECT 14751.305 1048.035 14751.585 1192.37 ;
      RECT 14750.745 1048.035 14751.025 1192.61 ;
      RECT 14750.185 1048.035 14750.465 1192.855 ;
      RECT 14749.625 1048.035 14749.905 1193.095 ;
      RECT 14749.065 1048.035 14749.345 1193.335 ;
      RECT 14748.505 1046.935 14748.785 1193.575 ;
      RECT 14747.945 1048.035 14748.225 1193.815 ;
      RECT 14747.385 1046.935 14747.665 1194.055 ;
      RECT 14746.825 1048.035 14747.105 1194.295 ;
      RECT 14746.265 1048.035 14746.545 1194.535 ;
      RECT 14745.705 1048.035 14745.985 1194.775 ;
      RECT 14745.145 1048.035 14745.425 1195.015 ;
      RECT 14744.585 1048.035 14744.865 1195.255 ;
      RECT 14744.025 1048.035 14744.305 1195.495 ;
      RECT 14743.465 1048.035 14743.745 1195.735 ;
      RECT 14742.905 1048.035 14743.185 1195.975 ;
      RECT 14742.345 1048.035 14742.625 1196.215 ;
      RECT 14741.785 1048.035 14742.065 1196.455 ;
      RECT 14741.225 1048.035 14741.505 1196.695 ;
      RECT 14732.265 1048.035 14732.545 1192.28 ;
      RECT 14731.705 1048.035 14731.985 1192.04 ;
      RECT 14731.145 1048.035 14731.425 1191.8 ;
      RECT 14730.585 1046.935 14730.865 1191.56 ;
      RECT 14730.025 1048.035 14730.305 1191.32 ;
      RECT 14729.465 1046.935 14729.745 1191.08 ;
      RECT 14728.905 1048.035 14729.185 1190.84 ;
      RECT 14728.345 1048.035 14728.625 1190.6 ;
      RECT 14727.785 1048.035 14728.065 1190.36 ;
      RECT 14727.225 1046.935 14727.505 1190.12 ;
      RECT 14726.665 1048.035 14726.945 1189.88 ;
      RECT 14726.105 1046.935 14726.385 1189.64 ;
      RECT 14725.545 1048.035 14725.825 1189.4 ;
      RECT 14724.985 1046.935 14725.265 1189.16 ;
      RECT 14722.465 1048.035 14722.745 1181.56 ;
      RECT 14721.905 1048.035 14722.185 1181.32 ;
      RECT 14721.345 1048.035 14721.625 1181.08 ;
      RECT 14720.785 1048.035 14721.065 1180.84 ;
      RECT 14720.225 1048.035 14720.505 1180.6 ;
      RECT 14719.665 1048.035 14719.945 1180.36 ;
      RECT 14719.105 1048.035 14719.385 1180.12 ;
      RECT 14693.065 1048.035 14693.345 1193.995 ;
      RECT 14692.505 1048.035 14692.785 1194.235 ;
      RECT 14691.945 1048.035 14692.225 1194.475 ;
      RECT 14691.385 1048.035 14691.665 1194.715 ;
      RECT 14690.825 1048.035 14691.105 1194.955 ;
      RECT 14690.265 1046.935 14690.545 1194.955 ;
      RECT 14689.705 1048.035 14689.985 1194.715 ;
      RECT 14689.145 1046.935 14689.425 1194.47 ;
      RECT 14688.585 1048.035 14688.865 1194.23 ;
      RECT 14688.025 1046.935 14688.305 1193.99 ;
      RECT 14687.465 1048.035 14687.745 1193.75 ;
      RECT 14686.905 1048.035 14687.185 1193.51 ;
      RECT 14686.345 1048.035 14686.625 1193.27 ;
      RECT 14685.785 1048.035 14686.065 1193.03 ;
      RECT 14685.225 1048.035 14685.505 1192.79 ;
      RECT 14684.665 1048.035 14684.945 1192.55 ;
      RECT 14684.105 1048.035 14684.385 1192.31 ;
      RECT 14683.545 1048.035 14683.825 1192.07 ;
      RECT 14682.985 1046.935 14683.265 1191.83 ;
      RECT 14682.425 1048.035 14682.705 1191.59 ;
      RECT 14681.865 1046.935 14682.145 1191.35 ;
      RECT 14681.305 1048.035 14681.585 1191.11 ;
      RECT 14680.745 1048.035 14681.025 1190.87 ;
      RECT 14680.185 1048.035 14680.465 1190.63 ;
      RECT 14666.745 1048.035 14667.025 1194.03 ;
      RECT 14666.185 1048.035 14666.465 1194.27 ;
      RECT 14665.625 1048.035 14665.905 1194.515 ;
      RECT 14665.065 1048.035 14665.345 1194.755 ;
      RECT 14664.505 1048.035 14664.785 1194.995 ;
      RECT 14663.945 1048.035 14664.225 1194.995 ;
      RECT 14663.385 1048.035 14663.665 1194.755 ;
      RECT 14662.825 1048.035 14663.105 1194.515 ;
      RECT 14662.265 1048.035 14662.545 1187.5 ;
      RECT 14661.705 1048.035 14661.985 1187.26 ;
      RECT 14661.145 1048.035 14661.425 1187.02 ;
      RECT 14660.585 1046.935 14660.865 1186.78 ;
      RECT 14660.025 1048.035 14660.305 1186.54 ;
      RECT 14659.465 1046.935 14659.745 1186.3 ;
      RECT 14658.905 1048.035 14659.185 1186.06 ;
      RECT 14658.345 1048.035 14658.625 1185.82 ;
      RECT 14657.785 1048.035 14658.065 1185.58 ;
      RECT 14657.225 1046.935 14657.505 1185.34 ;
      RECT 14656.665 1048.035 14656.945 1185.1 ;
      RECT 14656.105 1046.935 14656.385 1184.86 ;
      RECT 14655.545 1048.035 14655.825 1184.62 ;
      RECT 14654.985 1046.935 14655.265 1184.38 ;
      RECT 14654.425 1048.035 14654.705 1184.14 ;
      RECT 14653.865 1048.035 14654.145 1183.9 ;
      RECT 14613.545 1048.035 14613.825 1192.795 ;
      RECT 14612.985 1048.035 14613.265 1193.035 ;
      RECT 14612.425 1048.035 14612.705 1193.28 ;
      RECT 14611.865 1048.035 14612.145 1193.52 ;
      RECT 14611.305 1048.035 14611.585 1193.76 ;
      RECT 14610.745 1048.035 14611.025 1194 ;
      RECT 14610.185 1048.035 14610.465 1194.24 ;
      RECT 14609.625 1048.035 14609.905 1194.48 ;
      RECT 14609.065 1048.035 14609.345 1194.72 ;
      RECT 14608.505 1048.035 14608.785 1194.96 ;
      RECT 14607.945 1046.935 14608.225 1195.2 ;
      RECT 14607.385 1048.035 14607.665 1195.44 ;
      RECT 14606.825 1046.935 14607.105 1195.68 ;
      RECT 14606.265 1048.035 14606.545 1195.92 ;
      RECT 14605.705 1046.935 14605.985 1196.16 ;
      RECT 14605.145 1048.035 14605.425 1196.16 ;
      RECT 14604.585 1048.035 14604.865 1195.92 ;
      RECT 14604.025 1048.035 14604.305 1195.68 ;
      RECT 14603.465 1048.035 14603.745 1195.44 ;
      RECT 14602.905 1048.035 14603.185 1195.2 ;
      RECT 14602.345 1048.035 14602.625 1194.96 ;
      RECT 14601.785 1048.035 14602.065 1194.72 ;
      RECT 14601.225 1048.035 14601.505 1194.48 ;
      RECT 14592.265 1046.935 14592.545 1194.51 ;
      RECT 14591.705 1048.035 14591.985 1194.75 ;
      RECT 14591.145 1046.935 14591.425 1194.99 ;
      RECT 14590.585 1048.035 14590.865 1195.205 ;
      RECT 14590.025 1048.035 14590.305 1194.78 ;
      RECT 14589.465 1048.035 14589.745 1194.54 ;
      RECT 14588.905 1048.035 14589.185 1194.3 ;
      RECT 14588.345 1048.035 14588.625 1194.06 ;
      RECT 14587.785 1048.035 14588.065 1193.82 ;
      RECT 14587.225 1048.035 14587.505 1193.58 ;
      RECT 14586.665 1048.035 14586.945 1193.34 ;
      RECT 14586.105 1048.035 14586.385 1193.1 ;
      RECT 14585.545 1048.035 14585.825 1192.86 ;
      RECT 14584.985 1048.035 14585.265 1192.62 ;
      RECT 14582.465 1048.035 14582.745 1191.795 ;
      RECT 14581.905 1048.035 14582.185 1191.555 ;
      RECT 14581.345 1048.035 14581.625 1191.315 ;
      RECT 14580.785 1046.935 14581.065 1191.075 ;
      RECT 14580.225 1048.035 14580.505 1190.835 ;
      RECT 14579.665 1046.935 14579.945 1190.595 ;
      RECT 14579.105 1048.035 14579.385 1190.355 ;
      RECT 14578.545 1048.035 14578.825 1190.115 ;
      RECT 14551.945 1048.035 14552.225 1201.16 ;
      RECT 14551.385 1046.935 14551.665 1201.4 ;
      RECT 14550.825 1048.035 14551.105 1201.64 ;
      RECT 14550.265 1046.935 14550.545 1201.885 ;
      RECT 14549.705 1048.035 14549.985 1202.125 ;
      RECT 14549.145 1046.935 14549.425 1202.365 ;
      RECT 14548.585 1048.035 14548.865 1202.605 ;
      RECT 14548.025 1048.035 14548.305 1202.845 ;
      RECT 14547.465 1048.035 14547.745 1188.465 ;
      RECT 14546.905 1048.035 14547.185 1188.225 ;
      RECT 14546.345 1048.035 14546.625 1187.985 ;
      RECT 14545.785 1048.035 14546.065 1187.745 ;
      RECT 14545.225 1048.035 14545.505 1187.505 ;
      RECT 14544.665 1048.035 14544.945 1187.265 ;
      RECT 14544.105 1048.035 14544.385 1187.025 ;
      RECT 14543.545 1048.035 14543.825 1186.785 ;
      RECT 14542.985 1048.035 14543.265 1186.545 ;
      RECT 14542.425 1048.035 14542.705 1186.305 ;
      RECT 14541.865 1046.935 14542.145 1186.065 ;
      RECT 14541.305 1048.035 14541.585 1185.825 ;
      RECT 14540.745 1046.935 14541.025 1185.585 ;
      RECT 14540.185 1048.035 14540.465 1185.345 ;
      RECT 14526.185 1046.935 14526.465 1191.465 ;
      RECT 14525.625 1048.035 14525.905 1191.225 ;
      RECT 14525.065 1048.035 14525.345 1190.985 ;
      RECT 14524.505 1048.035 14524.785 1190.745 ;
      RECT 14523.945 1048.035 14524.225 1190.505 ;
      RECT 14523.385 1048.035 14523.665 1190.265 ;
      RECT 14522.825 1048.035 14523.105 1190.025 ;
      RECT 14522.265 1048.035 14522.545 1189.785 ;
      RECT 14521.705 1048.035 14521.985 1189.545 ;
      RECT 14521.145 1046.935 14521.425 1189.305 ;
      RECT 14520.585 1048.035 14520.865 1189.065 ;
      RECT 14520.025 1046.935 14520.305 1188.825 ;
      RECT 14519.465 1048.035 14519.745 1188.585 ;
      RECT 14518.905 1048.035 14519.185 1188.345 ;
      RECT 14518.345 1048.035 14518.625 1188.105 ;
      RECT 14517.785 1048.035 14518.065 1187.865 ;
      RECT 14517.225 1048.035 14517.505 1187.625 ;
      RECT 14516.665 1048.035 14516.945 1187.385 ;
      RECT 14516.105 1048.035 14516.385 1187.145 ;
      RECT 14515.545 1048.035 14515.825 1186.905 ;
      RECT 14514.985 1048.035 14515.265 1186.665 ;
      RECT 14514.425 1048.035 14514.705 1186.425 ;
      RECT 14513.865 1048.035 14514.145 1186.185 ;
      RECT 14474.665 1048.035 14474.945 1193.09 ;
      RECT 14474.105 1048.035 14474.385 1193.33 ;
      RECT 14473.545 1048.035 14473.825 1193.57 ;
      RECT 14472.985 1046.935 14473.265 1193.81 ;
      RECT 14472.425 1048.035 14472.705 1194.05 ;
      RECT 14471.865 1046.935 14472.145 1194.29 ;
      RECT 14471.305 1048.035 14471.585 1194.53 ;
      RECT 14470.745 1048.035 14471.025 1194.77 ;
      RECT 14470.185 1048.035 14470.465 1195.01 ;
      RECT 14469.625 1046.935 14469.905 1195.25 ;
      RECT 14469.065 1048.035 14469.345 1195.49 ;
      RECT 14468.505 1046.935 14468.785 1195.73 ;
      RECT 14467.945 1048.035 14468.225 1195.97 ;
      RECT 14467.385 1046.935 14467.665 1196.21 ;
      RECT 14466.825 1048.035 14467.105 1196.45 ;
      RECT 14466.265 1048.035 14466.545 1196.69 ;
      RECT 14465.705 1048.035 14465.985 1196.69 ;
      RECT 14465.145 1048.035 14465.425 1196.45 ;
      RECT 14464.585 1048.035 14464.865 1196.21 ;
      RECT 14464.025 1048.035 14464.305 1195.97 ;
      RECT 14463.465 1048.035 14463.745 1195.73 ;
      RECT 14462.905 1048.035 14463.185 1195.49 ;
      RECT 14462.345 1048.035 14462.625 1195.25 ;
      RECT 14461.785 1048.035 14462.065 1195.01 ;
      RECT 14461.225 1048.035 14461.505 1194.77 ;
      RECT 14452.265 1048.035 14452.545 1194.285 ;
      RECT 14451.705 1046.935 14451.985 1194.045 ;
      RECT 14451.145 1048.035 14451.425 1193.805 ;
      RECT 14450.585 1046.935 14450.865 1193.565 ;
      RECT 14450.025 1048.035 14450.305 1193.325 ;
      RECT 14449.465 1046.935 14449.745 1193.085 ;
      RECT 14448.905 1048.035 14449.185 1192.845 ;
      RECT 14448.345 1048.035 14448.625 1192.605 ;
      RECT 14447.785 1048.035 14448.065 1192.365 ;
      RECT 14447.225 1048.035 14447.505 1192.125 ;
      RECT 14446.665 1048.035 14446.945 1191.885 ;
      RECT 14446.105 1048.035 14446.385 1191.645 ;
      RECT 14445.545 1048.035 14445.825 1191.405 ;
      RECT 14444.985 1048.035 14445.265 1191.165 ;
      RECT 14442.465 1046.935 14442.745 1192.885 ;
      RECT 14441.905 1048.035 14442.185 1192.645 ;
      RECT 14441.345 1046.935 14441.625 1192.405 ;
      RECT 14440.785 1048.035 14441.065 1192.165 ;
      RECT 14440.225 1048.035 14440.505 1191.925 ;
      RECT 14439.665 1048.035 14439.945 1191.685 ;
      RECT 14439.105 1048.035 14439.385 1191.445 ;
      RECT 14438.545 1048.035 14438.825 1191.205 ;
      RECT 14412.505 1048.035 14412.785 1188.855 ;
      RECT 14411.945 1048.035 14412.225 1189.095 ;
      RECT 14411.385 1048.035 14411.665 1189.335 ;
      RECT 14410.825 1048.035 14411.105 1189.58 ;
      RECT 14410.265 1048.035 14410.545 1189.82 ;
      RECT 14409.705 1048.035 14409.985 1190.06 ;
      RECT 14409.145 1048.035 14409.425 1190.06 ;
      RECT 14408.585 1048.035 14408.865 1189.82 ;
      RECT 14408.025 1048.035 14408.305 1189.58 ;
      RECT 14407.465 1046.935 14407.745 1189.34 ;
      RECT 14406.905 1048.035 14407.185 1189.1 ;
      RECT 14406.345 1046.935 14406.625 1188.86 ;
      RECT 14405.785 1048.035 14406.065 1188.62 ;
      RECT 14405.225 1048.035 14405.505 1188.38 ;
      RECT 14404.665 1048.035 14404.945 1188.14 ;
      RECT 14404.105 1046.935 14404.385 1187.9 ;
      RECT 14403.545 1048.035 14403.825 1187.66 ;
      RECT 14402.985 1046.935 14403.265 1187.42 ;
      RECT 14402.425 1048.035 14402.705 1187.18 ;
      RECT 14401.865 1046.935 14402.145 1186.94 ;
      RECT 14401.305 1048.035 14401.585 1186.7 ;
      RECT 14400.745 1048.035 14401.025 1186.46 ;
      RECT 14400.185 1048.035 14400.465 1186.22 ;
      RECT 14399.625 1048.035 14399.905 1185.98 ;
      RECT 14386.185 1048.035 14386.465 1191.78 ;
      RECT 14385.625 1048.035 14385.905 1191.54 ;
      RECT 14385.065 1048.035 14385.345 1191.3 ;
      RECT 14384.505 1048.035 14384.785 1191.06 ;
      RECT 14383.945 1048.035 14384.225 1190.82 ;
      RECT 14383.385 1048.035 14383.665 1190.58 ;
      RECT 14382.825 1048.035 14383.105 1190.34 ;
      RECT 14382.265 1048.035 14382.545 1190.1 ;
      RECT 14381.705 1046.935 14381.985 1189.86 ;
      RECT 14381.145 1048.035 14381.425 1189.62 ;
      RECT 14380.585 1046.935 14380.865 1189.3 ;
      RECT 14380.025 1048.035 14380.305 1189.14 ;
      RECT 14379.465 1046.935 14379.745 1188.9 ;
      RECT 14378.905 1048.035 14379.185 1188.66 ;
      RECT 14378.345 1048.035 14378.625 1188.42 ;
      RECT 14377.785 1048.035 14378.065 1188.18 ;
      RECT 14377.225 1048.035 14377.505 1187.94 ;
      RECT 14376.665 1048.035 14376.945 1187.7 ;
      RECT 14376.105 1048.035 14376.385 1187.46 ;
      RECT 14375.545 1048.035 14375.825 1187.22 ;
      RECT 14374.985 1048.035 14375.265 1186.98 ;
      RECT 14374.425 1046.935 14374.705 1186.74 ;
      RECT 14373.865 1048.035 14374.145 1186.5 ;
      RECT 14373.305 1046.935 14373.585 1186.26 ;
      RECT 14334.105 1048.035 14334.385 1191.87 ;
      RECT 14333.545 1048.035 14333.825 1192.11 ;
      RECT 14332.985 1048.035 14333.265 1192.35 ;
      RECT 14332.425 1048.035 14332.705 1192.59 ;
      RECT 14331.865 1048.035 14332.145 1192.83 ;
      RECT 14331.305 1048.035 14331.585 1193.07 ;
      RECT 14330.745 1048.035 14331.025 1193.31 ;
      RECT 14330.185 1048.035 14330.465 1193.55 ;
      RECT 14329.625 1048.035 14329.905 1193.79 ;
      RECT 14329.065 1048.035 14329.345 1194.03 ;
      RECT 14328.505 1048.035 14328.785 1194.27 ;
      RECT 14327.945 1048.035 14328.225 1194.51 ;
      RECT 14327.385 1048.035 14327.665 1194.75 ;
      RECT 14326.825 1048.035 14327.105 1194.75 ;
      RECT 14326.265 1046.935 14326.545 1194.51 ;
      RECT 14325.705 1048.035 14325.985 1194.27 ;
      RECT 14325.145 1046.935 14325.425 1194.03 ;
      RECT 14324.585 1048.035 14324.865 1193.79 ;
      RECT 14324.025 1048.035 14324.305 1193.55 ;
      RECT 14323.465 1048.035 14323.745 1193.31 ;
      RECT 14322.905 1046.935 14323.185 1193.045 ;
      RECT 14322.345 1048.035 14322.625 1192.805 ;
      RECT 14321.785 1046.935 14322.065 1192.565 ;
      RECT 14321.225 1048.035 14321.505 1192.325 ;
      RECT 14312.265 1046.935 14312.545 1186.16 ;
      RECT 14311.705 1048.035 14311.985 1186.4 ;
      RECT 14311.145 1048.035 14311.425 1186.64 ;
      RECT 14310.585 1048.035 14310.865 1186.64 ;
      RECT 14310.025 1048.035 14310.305 1186.4 ;
      RECT 14309.465 1048.035 14309.745 1186.16 ;
      RECT 14308.905 1048.035 14309.185 1185.92 ;
      RECT 14308.345 1048.035 14308.625 1185.68 ;
      RECT 14307.785 1048.035 14308.065 1185.44 ;
      RECT 14307.225 1048.035 14307.505 1185.2 ;
      RECT 14306.665 1048.035 14306.945 1184.96 ;
      RECT 14306.105 1048.035 14306.385 1184.72 ;
      RECT 14305.545 1048.035 14305.825 1184.48 ;
      RECT 14304.985 1046.935 14305.265 1184.24 ;
      RECT 14302.465 1048.035 14302.745 1185.96 ;
      RECT 14301.905 1046.935 14302.185 1185.72 ;
      RECT 14301.345 1048.035 14301.625 1185.48 ;
      RECT 14300.785 1046.935 14301.065 1185.24 ;
      RECT 14300.225 1048.035 14300.505 1185 ;
      RECT 14299.665 1048.035 14299.945 1184.76 ;
      RECT 14299.105 1048.035 14299.385 1184.52 ;
      RECT 14273.065 1048.035 14273.345 1187.305 ;
      RECT 14272.505 1048.035 14272.785 1187.545 ;
      RECT 14271.945 1048.035 14272.225 1187.785 ;
      RECT 14271.385 1048.035 14271.665 1188.025 ;
      RECT 14270.825 1048.035 14271.105 1188.265 ;
      RECT 14270.265 1046.935 14270.545 1188.505 ;
      RECT 14269.705 1048.035 14269.985 1188.745 ;
      RECT 14269.145 1046.935 14269.425 1188.985 ;
      RECT 14268.585 1048.035 14268.865 1189.225 ;
      RECT 14268.025 1048.035 14268.305 1189.465 ;
      RECT 14267.465 1048.035 14267.745 1189.705 ;
      RECT 14266.905 1048.035 14267.185 1189.945 ;
      RECT 14266.345 1048.035 14266.625 1190.185 ;
      RECT 14265.785 1048.035 14266.065 1190.425 ;
      RECT 14265.225 1048.035 14265.505 1190.665 ;
      RECT 14264.665 1048.035 14264.945 1190.665 ;
      RECT 14264.105 1048.035 14264.385 1190.425 ;
      RECT 14263.545 1048.035 14263.825 1190.185 ;
      RECT 14262.985 1048.035 14263.265 1189.945 ;
      RECT 14262.425 1048.035 14262.705 1189.7 ;
      RECT 14261.865 1048.035 14262.145 1189.46 ;
      RECT 14261.305 1048.035 14261.585 1189.22 ;
      RECT 14260.745 1046.935 14261.025 1188.98 ;
      RECT 14260.185 1048.035 14260.465 1188.74 ;
      RECT 14246.745 1046.935 14247.025 1186.22 ;
      RECT 14246.185 1048.035 14246.465 1185.98 ;
      RECT 14245.625 1048.035 14245.905 1185.74 ;
      RECT 14245.065 1048.035 14245.345 1185.5 ;
      RECT 14244.505 1046.935 14244.785 1185.26 ;
      RECT 14243.945 1048.035 14244.225 1185.02 ;
      RECT 14243.385 1046.935 14243.665 1184.78 ;
      RECT 14242.825 1048.035 14243.105 1184.54 ;
      RECT 14242.265 1046.935 14242.545 1184.3 ;
      RECT 14241.705 1048.035 14241.985 1184.06 ;
      RECT 14241.145 1048.035 14241.425 1183.82 ;
      RECT 14240.585 1048.035 14240.865 1183.58 ;
      RECT 14240.025 1048.035 14240.305 1183.34 ;
      RECT 14239.465 1048.035 14239.745 1183.1 ;
      RECT 14238.905 1048.035 14239.185 1182.86 ;
      RECT 14238.345 1048.035 14238.625 1182.62 ;
      RECT 14237.785 1048.035 14238.065 1182.38 ;
      RECT 14237.225 1048.035 14237.505 1182.14 ;
      RECT 14236.665 1048.035 14236.945 1181.9 ;
      RECT 14236.105 1048.035 14236.385 1181.66 ;
      RECT 14235.545 1048.035 14235.825 1181.42 ;
      RECT 14234.985 1046.935 14235.265 1181.18 ;
      RECT 14234.425 1048.035 14234.705 1180.94 ;
      RECT 14233.865 1046.935 14234.145 1180.7 ;
      RECT 14194.105 1048.035 14194.385 1191.17 ;
      RECT 14193.545 1046.935 14193.825 1191.41 ;
      RECT 14192.985 1048.035 14193.265 1191.65 ;
      RECT 14192.425 1048.035 14192.705 1191.89 ;
      RECT 14191.865 1048.035 14192.145 1192.13 ;
      RECT 14191.305 1048.035 14191.585 1192.37 ;
      RECT 14190.745 1048.035 14191.025 1192.61 ;
      RECT 14190.185 1048.035 14190.465 1192.855 ;
      RECT 14189.625 1048.035 14189.905 1193.095 ;
      RECT 14189.065 1048.035 14189.345 1193.335 ;
      RECT 14188.505 1046.935 14188.785 1193.575 ;
      RECT 14187.945 1048.035 14188.225 1193.815 ;
      RECT 14187.385 1046.935 14187.665 1194.055 ;
      RECT 14186.825 1048.035 14187.105 1194.295 ;
      RECT 14186.265 1048.035 14186.545 1194.535 ;
      RECT 14185.705 1048.035 14185.985 1194.775 ;
      RECT 14185.145 1048.035 14185.425 1195.015 ;
      RECT 14184.585 1048.035 14184.865 1195.255 ;
      RECT 14184.025 1048.035 14184.305 1195.495 ;
      RECT 14183.465 1048.035 14183.745 1195.735 ;
      RECT 14182.905 1048.035 14183.185 1195.975 ;
      RECT 14182.345 1048.035 14182.625 1196.215 ;
      RECT 14181.785 1048.035 14182.065 1196.455 ;
      RECT 14181.225 1048.035 14181.505 1196.695 ;
      RECT 14172.265 1048.035 14172.545 1192.28 ;
      RECT 14171.705 1048.035 14171.985 1192.04 ;
      RECT 14171.145 1048.035 14171.425 1191.8 ;
      RECT 14170.585 1046.935 14170.865 1191.56 ;
      RECT 14170.025 1048.035 14170.305 1191.32 ;
      RECT 14169.465 1046.935 14169.745 1191.08 ;
      RECT 14168.905 1048.035 14169.185 1190.84 ;
      RECT 14168.345 1048.035 14168.625 1190.6 ;
      RECT 14167.785 1048.035 14168.065 1190.36 ;
      RECT 14167.225 1046.935 14167.505 1190.12 ;
      RECT 14166.665 1048.035 14166.945 1189.88 ;
      RECT 14166.105 1046.935 14166.385 1189.64 ;
      RECT 14165.545 1048.035 14165.825 1189.4 ;
      RECT 14164.985 1046.935 14165.265 1189.16 ;
      RECT 14162.465 1048.035 14162.745 1181.56 ;
      RECT 14161.905 1048.035 14162.185 1181.32 ;
      RECT 14161.345 1048.035 14161.625 1181.08 ;
      RECT 14160.785 1048.035 14161.065 1180.84 ;
      RECT 14160.225 1048.035 14160.505 1180.6 ;
      RECT 14159.665 1048.035 14159.945 1180.36 ;
      RECT 14159.105 1048.035 14159.385 1180.12 ;
      RECT 14133.065 1048.035 14133.345 1193.995 ;
      RECT 14132.505 1048.035 14132.785 1194.235 ;
      RECT 14131.945 1048.035 14132.225 1194.475 ;
      RECT 14131.385 1048.035 14131.665 1194.715 ;
      RECT 14130.825 1048.035 14131.105 1194.955 ;
      RECT 14130.265 1046.935 14130.545 1194.955 ;
      RECT 14129.705 1048.035 14129.985 1194.715 ;
      RECT 14129.145 1046.935 14129.425 1194.47 ;
      RECT 14128.585 1048.035 14128.865 1194.23 ;
      RECT 14128.025 1046.935 14128.305 1193.99 ;
      RECT 14127.465 1048.035 14127.745 1193.75 ;
      RECT 14126.905 1048.035 14127.185 1193.51 ;
      RECT 14126.345 1048.035 14126.625 1193.27 ;
      RECT 14125.785 1048.035 14126.065 1193.03 ;
      RECT 14125.225 1048.035 14125.505 1192.79 ;
      RECT 14124.665 1048.035 14124.945 1192.55 ;
      RECT 14124.105 1048.035 14124.385 1192.31 ;
      RECT 14123.545 1048.035 14123.825 1192.07 ;
      RECT 14122.985 1046.935 14123.265 1191.83 ;
      RECT 14122.425 1048.035 14122.705 1191.59 ;
      RECT 14121.865 1046.935 14122.145 1191.35 ;
      RECT 14121.305 1048.035 14121.585 1191.11 ;
      RECT 14120.745 1048.035 14121.025 1190.87 ;
      RECT 14120.185 1048.035 14120.465 1190.63 ;
      RECT 14106.745 1048.035 14107.025 1194.03 ;
      RECT 14106.185 1048.035 14106.465 1194.27 ;
      RECT 14105.625 1048.035 14105.905 1194.515 ;
      RECT 14105.065 1048.035 14105.345 1194.755 ;
      RECT 14104.505 1048.035 14104.785 1194.995 ;
      RECT 14103.945 1048.035 14104.225 1194.995 ;
      RECT 14103.385 1048.035 14103.665 1194.755 ;
      RECT 14102.825 1048.035 14103.105 1194.515 ;
      RECT 14102.265 1048.035 14102.545 1187.5 ;
      RECT 14101.705 1048.035 14101.985 1187.26 ;
      RECT 14101.145 1048.035 14101.425 1187.02 ;
      RECT 14100.585 1046.935 14100.865 1186.78 ;
      RECT 14100.025 1048.035 14100.305 1186.54 ;
      RECT 14099.465 1046.935 14099.745 1186.3 ;
      RECT 14098.905 1048.035 14099.185 1186.06 ;
      RECT 14098.345 1048.035 14098.625 1185.82 ;
      RECT 14097.785 1048.035 14098.065 1185.58 ;
      RECT 14097.225 1046.935 14097.505 1185.34 ;
      RECT 14096.665 1048.035 14096.945 1185.1 ;
      RECT 14096.105 1046.935 14096.385 1184.86 ;
      RECT 14095.545 1048.035 14095.825 1184.62 ;
      RECT 14094.985 1046.935 14095.265 1184.38 ;
      RECT 14094.425 1048.035 14094.705 1184.14 ;
      RECT 14093.865 1048.035 14094.145 1183.9 ;
      RECT 14053.545 1048.035 14053.825 1192.795 ;
      RECT 14052.985 1048.035 14053.265 1193.035 ;
      RECT 14052.425 1048.035 14052.705 1193.28 ;
      RECT 14051.865 1048.035 14052.145 1193.52 ;
      RECT 14051.305 1048.035 14051.585 1193.76 ;
      RECT 14050.745 1048.035 14051.025 1194 ;
      RECT 14050.185 1048.035 14050.465 1194.24 ;
      RECT 14049.625 1048.035 14049.905 1194.48 ;
      RECT 14049.065 1048.035 14049.345 1194.72 ;
      RECT 14048.505 1048.035 14048.785 1194.96 ;
      RECT 14047.945 1046.935 14048.225 1195.2 ;
      RECT 14047.385 1048.035 14047.665 1195.44 ;
      RECT 14046.825 1046.935 14047.105 1195.68 ;
      RECT 14046.265 1048.035 14046.545 1195.92 ;
      RECT 14045.705 1046.935 14045.985 1196.16 ;
      RECT 14045.145 1048.035 14045.425 1196.16 ;
      RECT 14044.585 1048.035 14044.865 1195.92 ;
      RECT 14044.025 1048.035 14044.305 1195.68 ;
      RECT 14043.465 1048.035 14043.745 1195.44 ;
      RECT 14042.905 1048.035 14043.185 1195.2 ;
      RECT 14042.345 1048.035 14042.625 1194.96 ;
      RECT 14041.785 1048.035 14042.065 1194.72 ;
      RECT 14041.225 1048.035 14041.505 1194.48 ;
      RECT 14032.265 1046.935 14032.545 1194.51 ;
      RECT 14031.705 1048.035 14031.985 1194.75 ;
      RECT 14031.145 1046.935 14031.425 1194.99 ;
      RECT 14030.585 1048.035 14030.865 1195.205 ;
      RECT 14030.025 1048.035 14030.305 1194.78 ;
      RECT 14029.465 1048.035 14029.745 1194.54 ;
      RECT 14028.905 1048.035 14029.185 1194.3 ;
      RECT 14028.345 1048.035 14028.625 1194.06 ;
      RECT 14027.785 1048.035 14028.065 1193.82 ;
      RECT 14027.225 1048.035 14027.505 1193.58 ;
      RECT 14026.665 1048.035 14026.945 1193.34 ;
      RECT 14026.105 1048.035 14026.385 1193.1 ;
      RECT 14025.545 1048.035 14025.825 1192.86 ;
      RECT 14024.985 1048.035 14025.265 1192.62 ;
      RECT 14022.465 1048.035 14022.745 1191.795 ;
      RECT 14021.905 1048.035 14022.185 1191.555 ;
      RECT 14021.345 1048.035 14021.625 1191.315 ;
      RECT 14020.785 1046.935 14021.065 1191.075 ;
      RECT 14020.225 1048.035 14020.505 1190.835 ;
      RECT 14019.665 1046.935 14019.945 1190.595 ;
      RECT 14019.105 1048.035 14019.385 1190.355 ;
      RECT 14018.545 1048.035 14018.825 1190.115 ;
      RECT 13991.945 1048.035 13992.225 1201.16 ;
      RECT 13991.385 1046.935 13991.665 1201.4 ;
      RECT 13990.825 1048.035 13991.105 1201.64 ;
      RECT 13990.265 1046.935 13990.545 1201.885 ;
      RECT 13989.705 1048.035 13989.985 1202.125 ;
      RECT 13989.145 1046.935 13989.425 1202.365 ;
      RECT 13988.585 1048.035 13988.865 1202.605 ;
      RECT 13988.025 1048.035 13988.305 1202.845 ;
      RECT 13987.465 1048.035 13987.745 1188.465 ;
      RECT 13986.905 1048.035 13987.185 1188.225 ;
      RECT 13986.345 1048.035 13986.625 1187.985 ;
      RECT 13985.785 1048.035 13986.065 1187.745 ;
      RECT 13985.225 1048.035 13985.505 1187.505 ;
      RECT 13984.665 1048.035 13984.945 1187.265 ;
      RECT 13984.105 1048.035 13984.385 1187.025 ;
      RECT 13983.545 1048.035 13983.825 1186.785 ;
      RECT 13982.985 1048.035 13983.265 1186.545 ;
      RECT 13982.425 1048.035 13982.705 1186.305 ;
      RECT 13981.865 1046.935 13982.145 1186.065 ;
      RECT 13981.305 1048.035 13981.585 1185.825 ;
      RECT 13980.745 1046.935 13981.025 1185.585 ;
      RECT 13980.185 1048.035 13980.465 1185.345 ;
      RECT 13966.185 1046.935 13966.465 1191.465 ;
      RECT 13965.625 1048.035 13965.905 1191.225 ;
      RECT 13965.065 1048.035 13965.345 1190.985 ;
      RECT 13964.505 1048.035 13964.785 1190.745 ;
      RECT 13963.945 1048.035 13964.225 1190.505 ;
      RECT 13963.385 1048.035 13963.665 1190.265 ;
      RECT 13962.825 1048.035 13963.105 1190.025 ;
      RECT 13962.265 1048.035 13962.545 1189.785 ;
      RECT 13961.705 1048.035 13961.985 1189.545 ;
      RECT 13961.145 1046.935 13961.425 1189.305 ;
      RECT 13960.585 1048.035 13960.865 1189.065 ;
      RECT 13960.025 1046.935 13960.305 1188.825 ;
      RECT 13959.465 1048.035 13959.745 1188.585 ;
      RECT 13958.905 1048.035 13959.185 1188.345 ;
      RECT 13958.345 1048.035 13958.625 1188.105 ;
      RECT 13957.785 1048.035 13958.065 1187.865 ;
      RECT 13957.225 1048.035 13957.505 1187.625 ;
      RECT 13956.665 1048.035 13956.945 1187.385 ;
      RECT 13956.105 1048.035 13956.385 1187.145 ;
      RECT 13955.545 1048.035 13955.825 1186.905 ;
      RECT 13954.985 1048.035 13955.265 1186.665 ;
      RECT 13954.425 1048.035 13954.705 1186.425 ;
      RECT 13953.865 1048.035 13954.145 1186.185 ;
      RECT 13914.665 1048.035 13914.945 1193.09 ;
      RECT 13914.105 1048.035 13914.385 1193.33 ;
      RECT 13913.545 1048.035 13913.825 1193.57 ;
      RECT 13912.985 1046.935 13913.265 1193.81 ;
      RECT 13912.425 1048.035 13912.705 1194.05 ;
      RECT 13911.865 1046.935 13912.145 1194.29 ;
      RECT 13911.305 1048.035 13911.585 1194.53 ;
      RECT 13910.745 1048.035 13911.025 1194.77 ;
      RECT 13910.185 1048.035 13910.465 1195.01 ;
      RECT 13909.625 1046.935 13909.905 1195.25 ;
      RECT 13909.065 1048.035 13909.345 1195.49 ;
      RECT 13908.505 1046.935 13908.785 1195.73 ;
      RECT 13907.945 1048.035 13908.225 1195.97 ;
      RECT 13907.385 1046.935 13907.665 1196.21 ;
      RECT 13906.825 1048.035 13907.105 1196.45 ;
      RECT 13906.265 1048.035 13906.545 1196.69 ;
      RECT 13905.705 1048.035 13905.985 1196.69 ;
      RECT 13905.145 1048.035 13905.425 1196.45 ;
      RECT 13904.585 1048.035 13904.865 1196.21 ;
      RECT 13904.025 1048.035 13904.305 1195.97 ;
      RECT 13903.465 1048.035 13903.745 1195.73 ;
      RECT 13902.905 1048.035 13903.185 1195.49 ;
      RECT 13902.345 1048.035 13902.625 1195.25 ;
      RECT 13901.785 1048.035 13902.065 1195.01 ;
      RECT 13901.225 1048.035 13901.505 1194.77 ;
      RECT 13892.265 1048.035 13892.545 1194.285 ;
      RECT 13891.705 1046.935 13891.985 1194.045 ;
      RECT 13891.145 1048.035 13891.425 1193.805 ;
      RECT 13890.585 1046.935 13890.865 1193.565 ;
      RECT 13890.025 1048.035 13890.305 1193.325 ;
      RECT 13889.465 1046.935 13889.745 1193.085 ;
      RECT 13888.905 1048.035 13889.185 1192.845 ;
      RECT 13888.345 1048.035 13888.625 1192.605 ;
      RECT 13887.785 1048.035 13888.065 1192.365 ;
      RECT 13887.225 1048.035 13887.505 1192.125 ;
      RECT 13886.665 1048.035 13886.945 1191.885 ;
      RECT 13886.105 1048.035 13886.385 1191.645 ;
      RECT 13885.545 1048.035 13885.825 1191.405 ;
      RECT 13884.985 1048.035 13885.265 1191.165 ;
      RECT 13882.465 1046.935 13882.745 1192.885 ;
      RECT 13881.905 1048.035 13882.185 1192.645 ;
      RECT 13881.345 1046.935 13881.625 1192.405 ;
      RECT 13880.785 1048.035 13881.065 1192.165 ;
      RECT 13880.225 1048.035 13880.505 1191.925 ;
      RECT 13879.665 1048.035 13879.945 1191.685 ;
      RECT 13879.105 1048.035 13879.385 1191.445 ;
      RECT 13878.545 1048.035 13878.825 1191.205 ;
      RECT 13852.505 1048.035 13852.785 1188.855 ;
      RECT 13851.945 1048.035 13852.225 1189.095 ;
      RECT 13851.385 1048.035 13851.665 1189.335 ;
      RECT 13850.825 1048.035 13851.105 1189.58 ;
      RECT 13850.265 1048.035 13850.545 1189.82 ;
      RECT 13849.705 1048.035 13849.985 1190.06 ;
      RECT 13849.145 1048.035 13849.425 1190.06 ;
      RECT 13848.585 1048.035 13848.865 1189.82 ;
      RECT 13848.025 1048.035 13848.305 1189.58 ;
      RECT 13847.465 1046.935 13847.745 1189.34 ;
      RECT 13846.905 1048.035 13847.185 1189.1 ;
      RECT 13846.345 1046.935 13846.625 1188.86 ;
      RECT 13845.785 1048.035 13846.065 1188.62 ;
      RECT 13845.225 1048.035 13845.505 1188.38 ;
      RECT 13844.665 1048.035 13844.945 1188.14 ;
      RECT 13844.105 1046.935 13844.385 1187.9 ;
      RECT 13843.545 1048.035 13843.825 1187.66 ;
      RECT 13842.985 1046.935 13843.265 1187.42 ;
      RECT 13842.425 1048.035 13842.705 1187.18 ;
      RECT 13841.865 1046.935 13842.145 1186.94 ;
      RECT 13841.305 1048.035 13841.585 1186.7 ;
      RECT 13840.745 1048.035 13841.025 1186.46 ;
      RECT 13840.185 1048.035 13840.465 1186.22 ;
      RECT 13839.625 1048.035 13839.905 1185.98 ;
      RECT 13826.185 1048.035 13826.465 1191.78 ;
      RECT 13825.625 1048.035 13825.905 1191.54 ;
      RECT 13825.065 1048.035 13825.345 1191.3 ;
      RECT 13824.505 1048.035 13824.785 1191.06 ;
      RECT 13823.945 1048.035 13824.225 1190.82 ;
      RECT 13823.385 1048.035 13823.665 1190.58 ;
      RECT 13822.825 1048.035 13823.105 1190.34 ;
      RECT 13822.265 1048.035 13822.545 1190.1 ;
      RECT 13821.705 1046.935 13821.985 1189.86 ;
      RECT 13821.145 1048.035 13821.425 1189.62 ;
      RECT 13820.585 1046.935 13820.865 1189.3 ;
      RECT 13820.025 1048.035 13820.305 1189.14 ;
      RECT 13819.465 1046.935 13819.745 1188.9 ;
      RECT 13818.905 1048.035 13819.185 1188.66 ;
      RECT 13818.345 1048.035 13818.625 1188.42 ;
      RECT 13817.785 1048.035 13818.065 1188.18 ;
      RECT 13817.225 1048.035 13817.505 1187.94 ;
      RECT 13816.665 1048.035 13816.945 1187.7 ;
      RECT 13816.105 1048.035 13816.385 1187.46 ;
      RECT 13815.545 1048.035 13815.825 1187.22 ;
      RECT 13814.985 1048.035 13815.265 1186.98 ;
      RECT 13814.425 1046.935 13814.705 1186.74 ;
      RECT 13813.865 1048.035 13814.145 1186.5 ;
      RECT 13813.305 1046.935 13813.585 1186.26 ;
      RECT 13774.105 1048.035 13774.385 1191.87 ;
      RECT 13773.545 1048.035 13773.825 1192.11 ;
      RECT 13772.985 1048.035 13773.265 1192.35 ;
      RECT 13772.425 1048.035 13772.705 1192.59 ;
      RECT 13771.865 1048.035 13772.145 1192.83 ;
      RECT 13771.305 1048.035 13771.585 1193.07 ;
      RECT 13770.745 1048.035 13771.025 1193.31 ;
      RECT 13770.185 1048.035 13770.465 1193.55 ;
      RECT 13769.625 1048.035 13769.905 1193.79 ;
      RECT 13769.065 1048.035 13769.345 1194.03 ;
      RECT 13768.505 1048.035 13768.785 1194.27 ;
      RECT 13767.945 1048.035 13768.225 1194.51 ;
      RECT 13767.385 1048.035 13767.665 1194.75 ;
      RECT 13766.825 1048.035 13767.105 1194.75 ;
      RECT 13766.265 1046.935 13766.545 1194.51 ;
      RECT 13765.705 1048.035 13765.985 1194.27 ;
      RECT 13765.145 1046.935 13765.425 1194.03 ;
      RECT 13764.585 1048.035 13764.865 1193.79 ;
      RECT 13764.025 1048.035 13764.305 1193.55 ;
      RECT 13763.465 1048.035 13763.745 1193.31 ;
      RECT 13762.905 1046.935 13763.185 1193.045 ;
      RECT 13762.345 1048.035 13762.625 1192.805 ;
      RECT 13761.785 1046.935 13762.065 1192.565 ;
      RECT 13761.225 1048.035 13761.505 1192.325 ;
      RECT 13752.265 1046.935 13752.545 1186.16 ;
      RECT 13751.705 1048.035 13751.985 1186.4 ;
      RECT 13751.145 1048.035 13751.425 1186.64 ;
      RECT 13750.585 1048.035 13750.865 1186.64 ;
      RECT 13750.025 1048.035 13750.305 1186.4 ;
      RECT 13749.465 1048.035 13749.745 1186.16 ;
      RECT 13748.905 1048.035 13749.185 1185.92 ;
      RECT 13748.345 1048.035 13748.625 1185.68 ;
      RECT 13747.785 1048.035 13748.065 1185.44 ;
      RECT 13747.225 1048.035 13747.505 1185.2 ;
      RECT 13746.665 1048.035 13746.945 1184.96 ;
      RECT 13746.105 1048.035 13746.385 1184.72 ;
      RECT 13745.545 1048.035 13745.825 1184.48 ;
      RECT 13744.985 1046.935 13745.265 1184.24 ;
      RECT 13742.465 1048.035 13742.745 1185.96 ;
      RECT 13741.905 1046.935 13742.185 1185.72 ;
      RECT 13741.345 1048.035 13741.625 1185.48 ;
      RECT 13740.785 1046.935 13741.065 1185.24 ;
      RECT 13740.225 1048.035 13740.505 1185 ;
      RECT 13739.665 1048.035 13739.945 1184.76 ;
      RECT 13739.105 1048.035 13739.385 1184.52 ;
      RECT 13713.065 1048.035 13713.345 1187.305 ;
      RECT 13712.505 1048.035 13712.785 1187.545 ;
      RECT 13711.945 1048.035 13712.225 1187.785 ;
      RECT 13711.385 1048.035 13711.665 1188.025 ;
      RECT 13710.825 1048.035 13711.105 1188.265 ;
      RECT 13710.265 1046.935 13710.545 1188.505 ;
      RECT 13709.705 1048.035 13709.985 1188.745 ;
      RECT 13709.145 1046.935 13709.425 1188.985 ;
      RECT 13708.585 1048.035 13708.865 1189.225 ;
      RECT 13708.025 1048.035 13708.305 1189.465 ;
      RECT 13707.465 1048.035 13707.745 1189.705 ;
      RECT 13706.905 1048.035 13707.185 1189.945 ;
      RECT 13706.345 1048.035 13706.625 1190.185 ;
      RECT 13705.785 1048.035 13706.065 1190.425 ;
      RECT 13705.225 1048.035 13705.505 1190.665 ;
      RECT 13704.665 1048.035 13704.945 1190.665 ;
      RECT 13704.105 1048.035 13704.385 1190.425 ;
      RECT 13703.545 1048.035 13703.825 1190.185 ;
      RECT 13702.985 1048.035 13703.265 1189.945 ;
      RECT 13702.425 1048.035 13702.705 1189.7 ;
      RECT 13701.865 1048.035 13702.145 1189.46 ;
      RECT 13701.305 1048.035 13701.585 1189.22 ;
      RECT 13700.745 1046.935 13701.025 1188.98 ;
      RECT 13700.185 1048.035 13700.465 1188.74 ;
      RECT 13686.745 1046.935 13687.025 1186.22 ;
      RECT 13686.185 1048.035 13686.465 1185.98 ;
      RECT 13685.625 1048.035 13685.905 1185.74 ;
      RECT 13685.065 1048.035 13685.345 1185.5 ;
      RECT 13684.505 1046.935 13684.785 1185.26 ;
      RECT 13683.945 1048.035 13684.225 1185.02 ;
      RECT 13683.385 1046.935 13683.665 1184.78 ;
      RECT 13682.825 1048.035 13683.105 1184.54 ;
      RECT 13682.265 1046.935 13682.545 1184.3 ;
      RECT 13681.705 1048.035 13681.985 1184.06 ;
      RECT 13681.145 1048.035 13681.425 1183.82 ;
      RECT 13680.585 1048.035 13680.865 1183.58 ;
      RECT 13680.025 1048.035 13680.305 1183.34 ;
      RECT 13679.465 1048.035 13679.745 1183.1 ;
      RECT 13678.905 1048.035 13679.185 1182.86 ;
      RECT 13678.345 1048.035 13678.625 1182.62 ;
      RECT 13677.785 1048.035 13678.065 1182.38 ;
      RECT 13677.225 1048.035 13677.505 1182.14 ;
      RECT 13676.665 1048.035 13676.945 1181.9 ;
      RECT 13676.105 1048.035 13676.385 1181.66 ;
      RECT 13675.545 1048.035 13675.825 1181.42 ;
      RECT 13674.985 1046.935 13675.265 1181.18 ;
      RECT 13674.425 1048.035 13674.705 1180.94 ;
      RECT 13673.865 1046.935 13674.145 1180.7 ;
      RECT 13634.105 1048.035 13634.385 1191.17 ;
      RECT 13633.545 1046.935 13633.825 1191.41 ;
      RECT 13632.985 1048.035 13633.265 1191.65 ;
      RECT 13632.425 1048.035 13632.705 1191.89 ;
      RECT 13631.865 1048.035 13632.145 1192.13 ;
      RECT 13631.305 1048.035 13631.585 1192.37 ;
      RECT 13630.745 1048.035 13631.025 1192.61 ;
      RECT 13630.185 1048.035 13630.465 1192.855 ;
      RECT 13629.625 1048.035 13629.905 1193.095 ;
      RECT 13629.065 1048.035 13629.345 1193.335 ;
      RECT 13628.505 1046.935 13628.785 1193.575 ;
      RECT 13627.945 1048.035 13628.225 1193.815 ;
      RECT 13627.385 1046.935 13627.665 1194.055 ;
      RECT 13626.825 1048.035 13627.105 1194.295 ;
      RECT 13626.265 1048.035 13626.545 1194.535 ;
      RECT 13625.705 1048.035 13625.985 1194.775 ;
      RECT 13625.145 1048.035 13625.425 1195.015 ;
      RECT 13624.585 1048.035 13624.865 1195.255 ;
      RECT 13624.025 1048.035 13624.305 1195.495 ;
      RECT 13623.465 1048.035 13623.745 1195.735 ;
      RECT 13622.905 1048.035 13623.185 1195.975 ;
      RECT 13622.345 1048.035 13622.625 1196.215 ;
      RECT 13621.785 1048.035 13622.065 1196.455 ;
      RECT 13621.225 1048.035 13621.505 1196.695 ;
      RECT 13612.265 1048.035 13612.545 1192.28 ;
      RECT 13611.705 1048.035 13611.985 1192.04 ;
      RECT 13611.145 1048.035 13611.425 1191.8 ;
      RECT 13610.585 1046.935 13610.865 1191.56 ;
      RECT 13610.025 1048.035 13610.305 1191.32 ;
      RECT 13609.465 1046.935 13609.745 1191.08 ;
      RECT 13608.905 1048.035 13609.185 1190.84 ;
      RECT 13608.345 1048.035 13608.625 1190.6 ;
      RECT 13607.785 1048.035 13608.065 1190.36 ;
      RECT 13607.225 1046.935 13607.505 1190.12 ;
      RECT 13606.665 1048.035 13606.945 1189.88 ;
      RECT 13606.105 1046.935 13606.385 1189.64 ;
      RECT 13605.545 1048.035 13605.825 1189.4 ;
      RECT 13604.985 1046.935 13605.265 1189.16 ;
      RECT 13602.465 1048.035 13602.745 1181.56 ;
      RECT 13601.905 1048.035 13602.185 1181.32 ;
      RECT 13601.345 1048.035 13601.625 1181.08 ;
      RECT 13600.785 1048.035 13601.065 1180.84 ;
      RECT 13600.225 1048.035 13600.505 1180.6 ;
      RECT 13599.665 1048.035 13599.945 1180.36 ;
      RECT 13599.105 1048.035 13599.385 1180.12 ;
      RECT 13573.065 1048.035 13573.345 1193.995 ;
      RECT 13572.505 1048.035 13572.785 1194.235 ;
      RECT 13571.945 1048.035 13572.225 1194.475 ;
      RECT 13571.385 1048.035 13571.665 1194.715 ;
      RECT 13570.825 1048.035 13571.105 1194.955 ;
      RECT 13570.265 1046.935 13570.545 1194.955 ;
      RECT 13569.705 1048.035 13569.985 1194.715 ;
      RECT 13569.145 1046.935 13569.425 1194.47 ;
      RECT 13568.585 1048.035 13568.865 1194.23 ;
      RECT 13568.025 1046.935 13568.305 1193.99 ;
      RECT 13567.465 1048.035 13567.745 1193.75 ;
      RECT 13566.905 1048.035 13567.185 1193.51 ;
      RECT 13566.345 1048.035 13566.625 1193.27 ;
      RECT 13565.785 1048.035 13566.065 1193.03 ;
      RECT 13565.225 1048.035 13565.505 1192.79 ;
      RECT 13564.665 1048.035 13564.945 1192.55 ;
      RECT 13564.105 1048.035 13564.385 1192.31 ;
      RECT 13563.545 1048.035 13563.825 1192.07 ;
      RECT 13562.985 1046.935 13563.265 1191.83 ;
      RECT 13562.425 1048.035 13562.705 1191.59 ;
      RECT 13561.865 1046.935 13562.145 1191.35 ;
      RECT 13561.305 1048.035 13561.585 1191.11 ;
      RECT 13560.745 1048.035 13561.025 1190.87 ;
      RECT 13560.185 1048.035 13560.465 1190.63 ;
      RECT 13546.745 1048.035 13547.025 1194.03 ;
      RECT 13546.185 1048.035 13546.465 1194.27 ;
      RECT 13545.625 1048.035 13545.905 1194.515 ;
      RECT 13545.065 1048.035 13545.345 1194.755 ;
      RECT 13544.505 1048.035 13544.785 1194.995 ;
      RECT 13543.945 1048.035 13544.225 1194.995 ;
      RECT 13543.385 1048.035 13543.665 1194.755 ;
      RECT 13542.825 1048.035 13543.105 1194.515 ;
      RECT 13542.265 1048.035 13542.545 1187.5 ;
      RECT 13541.705 1048.035 13541.985 1187.26 ;
      RECT 13541.145 1048.035 13541.425 1187.02 ;
      RECT 13540.585 1046.935 13540.865 1186.78 ;
      RECT 13540.025 1048.035 13540.305 1186.54 ;
      RECT 13539.465 1046.935 13539.745 1186.3 ;
      RECT 13538.905 1048.035 13539.185 1186.06 ;
      RECT 13538.345 1048.035 13538.625 1185.82 ;
      RECT 13537.785 1048.035 13538.065 1185.58 ;
      RECT 13537.225 1046.935 13537.505 1185.34 ;
      RECT 13536.665 1048.035 13536.945 1185.1 ;
      RECT 13536.105 1046.935 13536.385 1184.86 ;
      RECT 13535.545 1048.035 13535.825 1184.62 ;
      RECT 13534.985 1046.935 13535.265 1184.38 ;
      RECT 13534.425 1048.035 13534.705 1184.14 ;
      RECT 13533.865 1048.035 13534.145 1183.9 ;
      RECT 13493.545 1048.035 13493.825 1192.795 ;
      RECT 13492.985 1048.035 13493.265 1193.035 ;
      RECT 13492.425 1048.035 13492.705 1193.28 ;
      RECT 13491.865 1048.035 13492.145 1193.52 ;
      RECT 13491.305 1048.035 13491.585 1193.76 ;
      RECT 13490.745 1048.035 13491.025 1194 ;
      RECT 13490.185 1048.035 13490.465 1194.24 ;
      RECT 13489.625 1048.035 13489.905 1194.48 ;
      RECT 13489.065 1048.035 13489.345 1194.72 ;
      RECT 13488.505 1048.035 13488.785 1194.96 ;
      RECT 13487.945 1046.935 13488.225 1195.2 ;
      RECT 13487.385 1048.035 13487.665 1195.44 ;
      RECT 13486.825 1046.935 13487.105 1195.68 ;
      RECT 13486.265 1048.035 13486.545 1195.92 ;
      RECT 13485.705 1046.935 13485.985 1196.16 ;
      RECT 13485.145 1048.035 13485.425 1196.16 ;
      RECT 13484.585 1048.035 13484.865 1195.92 ;
      RECT 13484.025 1048.035 13484.305 1195.68 ;
      RECT 13483.465 1048.035 13483.745 1195.44 ;
      RECT 13482.905 1048.035 13483.185 1195.2 ;
      RECT 13482.345 1048.035 13482.625 1194.96 ;
      RECT 13481.785 1048.035 13482.065 1194.72 ;
      RECT 13481.225 1048.035 13481.505 1194.48 ;
      RECT 13472.265 1046.935 13472.545 1194.51 ;
      RECT 13471.705 1048.035 13471.985 1194.75 ;
      RECT 13471.145 1046.935 13471.425 1194.99 ;
      RECT 13470.585 1048.035 13470.865 1195.205 ;
      RECT 13470.025 1048.035 13470.305 1194.78 ;
      RECT 13469.465 1048.035 13469.745 1194.54 ;
      RECT 13468.905 1048.035 13469.185 1194.3 ;
      RECT 13468.345 1048.035 13468.625 1194.06 ;
      RECT 13467.785 1048.035 13468.065 1193.82 ;
      RECT 13467.225 1048.035 13467.505 1193.58 ;
      RECT 13466.665 1048.035 13466.945 1193.34 ;
      RECT 13466.105 1048.035 13466.385 1193.1 ;
      RECT 13465.545 1048.035 13465.825 1192.86 ;
      RECT 13464.985 1048.035 13465.265 1192.62 ;
      RECT 13462.465 1048.035 13462.745 1191.795 ;
      RECT 13461.905 1048.035 13462.185 1191.555 ;
      RECT 13461.345 1048.035 13461.625 1191.315 ;
      RECT 13460.785 1046.935 13461.065 1191.075 ;
      RECT 13460.225 1048.035 13460.505 1190.835 ;
      RECT 13459.665 1046.935 13459.945 1190.595 ;
      RECT 13459.105 1048.035 13459.385 1190.355 ;
      RECT 13458.545 1048.035 13458.825 1190.115 ;
      RECT 13431.945 1048.035 13432.225 1201.16 ;
      RECT 13431.385 1046.935 13431.665 1201.4 ;
      RECT 13430.825 1048.035 13431.105 1201.64 ;
      RECT 13430.265 1046.935 13430.545 1201.885 ;
      RECT 13429.705 1048.035 13429.985 1202.125 ;
      RECT 13429.145 1046.935 13429.425 1202.365 ;
      RECT 13428.585 1048.035 13428.865 1202.605 ;
      RECT 13428.025 1048.035 13428.305 1202.845 ;
      RECT 13427.465 1048.035 13427.745 1188.465 ;
      RECT 13426.905 1048.035 13427.185 1188.225 ;
      RECT 13426.345 1048.035 13426.625 1187.985 ;
      RECT 13425.785 1048.035 13426.065 1187.745 ;
      RECT 13425.225 1048.035 13425.505 1187.505 ;
      RECT 13424.665 1048.035 13424.945 1187.265 ;
      RECT 13424.105 1048.035 13424.385 1187.025 ;
      RECT 13423.545 1048.035 13423.825 1186.785 ;
      RECT 13422.985 1048.035 13423.265 1186.545 ;
      RECT 13422.425 1048.035 13422.705 1186.305 ;
      RECT 13421.865 1046.935 13422.145 1186.065 ;
      RECT 13421.305 1048.035 13421.585 1185.825 ;
      RECT 13420.745 1046.935 13421.025 1185.585 ;
      RECT 13420.185 1048.035 13420.465 1185.345 ;
      RECT 13406.185 1046.935 13406.465 1191.465 ;
      RECT 13405.625 1048.035 13405.905 1191.225 ;
      RECT 13405.065 1048.035 13405.345 1190.985 ;
      RECT 13404.505 1048.035 13404.785 1190.745 ;
      RECT 13403.945 1048.035 13404.225 1190.505 ;
      RECT 13403.385 1048.035 13403.665 1190.265 ;
      RECT 13402.825 1048.035 13403.105 1190.025 ;
      RECT 13402.265 1048.035 13402.545 1189.785 ;
      RECT 13401.705 1048.035 13401.985 1189.545 ;
      RECT 13401.145 1046.935 13401.425 1189.305 ;
      RECT 13400.585 1048.035 13400.865 1189.065 ;
      RECT 13400.025 1046.935 13400.305 1188.825 ;
      RECT 13399.465 1048.035 13399.745 1188.585 ;
      RECT 13398.905 1048.035 13399.185 1188.345 ;
      RECT 13398.345 1048.035 13398.625 1188.105 ;
      RECT 13397.785 1048.035 13398.065 1187.865 ;
      RECT 13397.225 1048.035 13397.505 1187.625 ;
      RECT 13396.665 1048.035 13396.945 1187.385 ;
      RECT 13396.105 1048.035 13396.385 1187.145 ;
      RECT 13395.545 1048.035 13395.825 1186.905 ;
      RECT 13394.985 1048.035 13395.265 1186.665 ;
      RECT 13394.425 1048.035 13394.705 1186.425 ;
      RECT 13393.865 1048.035 13394.145 1186.185 ;
      RECT 13354.665 1048.035 13354.945 1193.09 ;
      RECT 13354.105 1048.035 13354.385 1193.33 ;
      RECT 13353.545 1048.035 13353.825 1193.57 ;
      RECT 13352.985 1046.935 13353.265 1193.81 ;
      RECT 13352.425 1048.035 13352.705 1194.05 ;
      RECT 13351.865 1046.935 13352.145 1194.29 ;
      RECT 13351.305 1048.035 13351.585 1194.53 ;
      RECT 13350.745 1048.035 13351.025 1194.77 ;
      RECT 13350.185 1048.035 13350.465 1195.01 ;
      RECT 13349.625 1046.935 13349.905 1195.25 ;
      RECT 13349.065 1048.035 13349.345 1195.49 ;
      RECT 13348.505 1046.935 13348.785 1195.73 ;
      RECT 13347.945 1048.035 13348.225 1195.97 ;
      RECT 13347.385 1046.935 13347.665 1196.21 ;
      RECT 13346.825 1048.035 13347.105 1196.45 ;
      RECT 13346.265 1048.035 13346.545 1196.69 ;
      RECT 13345.705 1048.035 13345.985 1196.69 ;
      RECT 13345.145 1048.035 13345.425 1196.45 ;
      RECT 13344.585 1048.035 13344.865 1196.21 ;
      RECT 13344.025 1048.035 13344.305 1195.97 ;
      RECT 13343.465 1048.035 13343.745 1195.73 ;
      RECT 13342.905 1048.035 13343.185 1195.49 ;
      RECT 13342.345 1048.035 13342.625 1195.25 ;
      RECT 13341.785 1048.035 13342.065 1195.01 ;
      RECT 13341.225 1048.035 13341.505 1194.77 ;
      RECT 13332.265 1048.035 13332.545 1194.285 ;
      RECT 13331.705 1046.935 13331.985 1194.045 ;
      RECT 13331.145 1048.035 13331.425 1193.805 ;
      RECT 13330.585 1046.935 13330.865 1193.565 ;
      RECT 13330.025 1048.035 13330.305 1193.325 ;
      RECT 13329.465 1046.935 13329.745 1193.085 ;
      RECT 13328.905 1048.035 13329.185 1192.845 ;
      RECT 13328.345 1048.035 13328.625 1192.605 ;
      RECT 13327.785 1048.035 13328.065 1192.365 ;
      RECT 13327.225 1048.035 13327.505 1192.125 ;
      RECT 13326.665 1048.035 13326.945 1191.885 ;
      RECT 13326.105 1048.035 13326.385 1191.645 ;
      RECT 13325.545 1048.035 13325.825 1191.405 ;
      RECT 13324.985 1048.035 13325.265 1191.165 ;
      RECT 13322.465 1046.935 13322.745 1192.885 ;
      RECT 13321.905 1048.035 13322.185 1192.645 ;
      RECT 13321.345 1046.935 13321.625 1192.405 ;
      RECT 13320.785 1048.035 13321.065 1192.165 ;
      RECT 13320.225 1048.035 13320.505 1191.925 ;
      RECT 13319.665 1048.035 13319.945 1191.685 ;
      RECT 13319.105 1048.035 13319.385 1191.445 ;
      RECT 13318.545 1048.035 13318.825 1191.205 ;
      RECT 13292.505 1048.035 13292.785 1188.855 ;
      RECT 13291.945 1048.035 13292.225 1189.095 ;
      RECT 13291.385 1048.035 13291.665 1189.335 ;
      RECT 13290.825 1048.035 13291.105 1189.58 ;
      RECT 13290.265 1048.035 13290.545 1189.82 ;
      RECT 13289.705 1048.035 13289.985 1190.06 ;
      RECT 13289.145 1048.035 13289.425 1190.06 ;
      RECT 13288.585 1048.035 13288.865 1189.82 ;
      RECT 13288.025 1048.035 13288.305 1189.58 ;
      RECT 13287.465 1046.935 13287.745 1189.34 ;
      RECT 13286.905 1048.035 13287.185 1189.1 ;
      RECT 13286.345 1046.935 13286.625 1188.86 ;
      RECT 13285.785 1048.035 13286.065 1188.62 ;
      RECT 13285.225 1048.035 13285.505 1188.38 ;
      RECT 13284.665 1048.035 13284.945 1188.14 ;
      RECT 13284.105 1046.935 13284.385 1187.9 ;
      RECT 13283.545 1048.035 13283.825 1187.66 ;
      RECT 13282.985 1046.935 13283.265 1187.42 ;
      RECT 13282.425 1048.035 13282.705 1187.18 ;
      RECT 13281.865 1046.935 13282.145 1186.94 ;
      RECT 13281.305 1048.035 13281.585 1186.7 ;
      RECT 13280.745 1048.035 13281.025 1186.46 ;
      RECT 13280.185 1048.035 13280.465 1186.22 ;
      RECT 13279.625 1048.035 13279.905 1185.98 ;
      RECT 13266.185 1048.035 13266.465 1191.78 ;
      RECT 13265.625 1048.035 13265.905 1191.54 ;
      RECT 13265.065 1048.035 13265.345 1191.3 ;
      RECT 13264.505 1048.035 13264.785 1191.06 ;
      RECT 13263.945 1048.035 13264.225 1190.82 ;
      RECT 13263.385 1048.035 13263.665 1190.58 ;
      RECT 13262.825 1048.035 13263.105 1190.34 ;
      RECT 13262.265 1048.035 13262.545 1190.1 ;
      RECT 13261.705 1046.935 13261.985 1189.86 ;
      RECT 13261.145 1048.035 13261.425 1189.62 ;
      RECT 13260.585 1046.935 13260.865 1189.3 ;
      RECT 13260.025 1048.035 13260.305 1189.14 ;
      RECT 13259.465 1046.935 13259.745 1188.9 ;
      RECT 13258.905 1048.035 13259.185 1188.66 ;
      RECT 13258.345 1048.035 13258.625 1188.42 ;
      RECT 13257.785 1048.035 13258.065 1188.18 ;
      RECT 13257.225 1048.035 13257.505 1187.94 ;
      RECT 13256.665 1048.035 13256.945 1187.7 ;
      RECT 13256.105 1048.035 13256.385 1187.46 ;
      RECT 13255.545 1048.035 13255.825 1187.22 ;
      RECT 13254.985 1048.035 13255.265 1186.98 ;
      RECT 13254.425 1046.935 13254.705 1186.74 ;
      RECT 13253.865 1048.035 13254.145 1186.5 ;
      RECT 13253.305 1046.935 13253.585 1186.26 ;
      RECT 13214.105 1048.035 13214.385 1191.87 ;
      RECT 13213.545 1048.035 13213.825 1192.11 ;
      RECT 13212.985 1048.035 13213.265 1192.35 ;
      RECT 13212.425 1048.035 13212.705 1192.59 ;
      RECT 13211.865 1048.035 13212.145 1192.83 ;
      RECT 13211.305 1048.035 13211.585 1193.07 ;
      RECT 13210.745 1048.035 13211.025 1193.31 ;
      RECT 13210.185 1048.035 13210.465 1193.55 ;
      RECT 13209.625 1048.035 13209.905 1193.79 ;
      RECT 13209.065 1048.035 13209.345 1194.03 ;
      RECT 13208.505 1048.035 13208.785 1194.27 ;
      RECT 13207.945 1048.035 13208.225 1194.51 ;
      RECT 13207.385 1048.035 13207.665 1194.75 ;
      RECT 13206.825 1048.035 13207.105 1194.75 ;
      RECT 13206.265 1046.935 13206.545 1194.51 ;
      RECT 13205.705 1048.035 13205.985 1194.27 ;
      RECT 13205.145 1046.935 13205.425 1194.03 ;
      RECT 13204.585 1048.035 13204.865 1193.79 ;
      RECT 13204.025 1048.035 13204.305 1193.55 ;
      RECT 13203.465 1048.035 13203.745 1193.31 ;
      RECT 13202.905 1046.935 13203.185 1193.045 ;
      RECT 13202.345 1048.035 13202.625 1192.805 ;
      RECT 13201.785 1046.935 13202.065 1192.565 ;
      RECT 13201.225 1048.035 13201.505 1192.325 ;
      RECT 13192.265 1046.935 13192.545 1186.16 ;
      RECT 13191.705 1048.035 13191.985 1186.4 ;
      RECT 13191.145 1048.035 13191.425 1186.64 ;
      RECT 13190.585 1048.035 13190.865 1186.64 ;
      RECT 13190.025 1048.035 13190.305 1186.4 ;
      RECT 13189.465 1048.035 13189.745 1186.16 ;
      RECT 13188.905 1048.035 13189.185 1185.92 ;
      RECT 13188.345 1048.035 13188.625 1185.68 ;
      RECT 13187.785 1048.035 13188.065 1185.44 ;
      RECT 13187.225 1048.035 13187.505 1185.2 ;
      RECT 13186.665 1048.035 13186.945 1184.96 ;
      RECT 13186.105 1048.035 13186.385 1184.72 ;
      RECT 13185.545 1048.035 13185.825 1184.48 ;
      RECT 13184.985 1046.935 13185.265 1184.24 ;
      RECT 13182.465 1048.035 13182.745 1185.96 ;
      RECT 13181.905 1046.935 13182.185 1185.72 ;
      RECT 13181.345 1048.035 13181.625 1185.48 ;
      RECT 13180.785 1046.935 13181.065 1185.24 ;
      RECT 13180.225 1048.035 13180.505 1185 ;
      RECT 13179.665 1048.035 13179.945 1184.76 ;
      RECT 13179.105 1048.035 13179.385 1184.52 ;
      RECT 13153.065 1048.035 13153.345 1187.305 ;
      RECT 13152.505 1048.035 13152.785 1187.545 ;
      RECT 13151.945 1048.035 13152.225 1187.785 ;
      RECT 13151.385 1048.035 13151.665 1188.025 ;
      RECT 13150.825 1048.035 13151.105 1188.265 ;
      RECT 13150.265 1046.935 13150.545 1188.505 ;
      RECT 13149.705 1048.035 13149.985 1188.745 ;
      RECT 13149.145 1046.935 13149.425 1188.985 ;
      RECT 13148.585 1048.035 13148.865 1189.225 ;
      RECT 13148.025 1048.035 13148.305 1189.465 ;
      RECT 13147.465 1048.035 13147.745 1189.705 ;
      RECT 13146.905 1048.035 13147.185 1189.945 ;
      RECT 13146.345 1048.035 13146.625 1190.185 ;
      RECT 13145.785 1048.035 13146.065 1190.425 ;
      RECT 13145.225 1048.035 13145.505 1190.665 ;
      RECT 13144.665 1048.035 13144.945 1190.665 ;
      RECT 13144.105 1048.035 13144.385 1190.425 ;
      RECT 13143.545 1048.035 13143.825 1190.185 ;
      RECT 13142.985 1048.035 13143.265 1189.945 ;
      RECT 13142.425 1048.035 13142.705 1189.7 ;
      RECT 13141.865 1048.035 13142.145 1189.46 ;
      RECT 13141.305 1048.035 13141.585 1189.22 ;
      RECT 13140.745 1046.935 13141.025 1188.98 ;
      RECT 13140.185 1048.035 13140.465 1188.74 ;
      RECT 13126.745 1046.935 13127.025 1186.22 ;
      RECT 13126.185 1048.035 13126.465 1185.98 ;
      RECT 13125.625 1048.035 13125.905 1185.74 ;
      RECT 13125.065 1048.035 13125.345 1185.5 ;
      RECT 13124.505 1046.935 13124.785 1185.26 ;
      RECT 13123.945 1048.035 13124.225 1185.02 ;
      RECT 13123.385 1046.935 13123.665 1184.78 ;
      RECT 13122.825 1048.035 13123.105 1184.54 ;
      RECT 13122.265 1046.935 13122.545 1184.3 ;
      RECT 13121.705 1048.035 13121.985 1184.06 ;
      RECT 13121.145 1048.035 13121.425 1183.82 ;
      RECT 13120.585 1048.035 13120.865 1183.58 ;
      RECT 13120.025 1048.035 13120.305 1183.34 ;
      RECT 13119.465 1048.035 13119.745 1183.1 ;
      RECT 13118.905 1048.035 13119.185 1182.86 ;
      RECT 13118.345 1048.035 13118.625 1182.62 ;
      RECT 13117.785 1048.035 13118.065 1182.38 ;
      RECT 13117.225 1048.035 13117.505 1182.14 ;
      RECT 13116.665 1048.035 13116.945 1181.9 ;
      RECT 13116.105 1048.035 13116.385 1181.66 ;
      RECT 13115.545 1048.035 13115.825 1181.42 ;
      RECT 13114.985 1046.935 13115.265 1181.18 ;
      RECT 13114.425 1048.035 13114.705 1180.94 ;
      RECT 13113.865 1046.935 13114.145 1180.7 ;
      RECT 13074.105 1048.035 13074.385 1191.17 ;
      RECT 13073.545 1046.935 13073.825 1191.41 ;
      RECT 13072.985 1048.035 13073.265 1191.65 ;
      RECT 13072.425 1048.035 13072.705 1191.89 ;
      RECT 13071.865 1048.035 13072.145 1192.13 ;
      RECT 13071.305 1048.035 13071.585 1192.37 ;
      RECT 13070.745 1048.035 13071.025 1192.61 ;
      RECT 13070.185 1048.035 13070.465 1192.855 ;
      RECT 13069.625 1048.035 13069.905 1193.095 ;
      RECT 13069.065 1048.035 13069.345 1193.335 ;
      RECT 13068.505 1046.935 13068.785 1193.575 ;
      RECT 13067.945 1048.035 13068.225 1193.815 ;
      RECT 13067.385 1046.935 13067.665 1194.055 ;
      RECT 13066.825 1048.035 13067.105 1194.295 ;
      RECT 13066.265 1048.035 13066.545 1194.535 ;
      RECT 13065.705 1048.035 13065.985 1194.775 ;
      RECT 13065.145 1048.035 13065.425 1195.015 ;
      RECT 13064.585 1048.035 13064.865 1195.255 ;
      RECT 13064.025 1048.035 13064.305 1195.495 ;
      RECT 13063.465 1048.035 13063.745 1195.735 ;
      RECT 13062.905 1048.035 13063.185 1195.975 ;
      RECT 13062.345 1048.035 13062.625 1196.215 ;
      RECT 13061.785 1048.035 13062.065 1196.455 ;
      RECT 13061.225 1048.035 13061.505 1196.695 ;
      RECT 13052.265 1048.035 13052.545 1192.28 ;
      RECT 13051.705 1048.035 13051.985 1192.04 ;
      RECT 13051.145 1048.035 13051.425 1191.8 ;
      RECT 13050.585 1046.935 13050.865 1191.56 ;
      RECT 13050.025 1048.035 13050.305 1191.32 ;
      RECT 13049.465 1046.935 13049.745 1191.08 ;
      RECT 13048.905 1048.035 13049.185 1190.84 ;
      RECT 13048.345 1048.035 13048.625 1190.6 ;
      RECT 13047.785 1048.035 13048.065 1190.36 ;
      RECT 13047.225 1046.935 13047.505 1190.12 ;
      RECT 13046.665 1048.035 13046.945 1189.88 ;
      RECT 13046.105 1046.935 13046.385 1189.64 ;
      RECT 13045.545 1048.035 13045.825 1189.4 ;
      RECT 13044.985 1046.935 13045.265 1189.16 ;
      RECT 13042.465 1048.035 13042.745 1181.56 ;
      RECT 13041.905 1048.035 13042.185 1181.32 ;
      RECT 13041.345 1048.035 13041.625 1181.08 ;
      RECT 13040.785 1048.035 13041.065 1180.84 ;
      RECT 13040.225 1048.035 13040.505 1180.6 ;
      RECT 13039.665 1048.035 13039.945 1180.36 ;
      RECT 13039.105 1048.035 13039.385 1180.12 ;
      RECT 13013.065 1048.035 13013.345 1193.995 ;
      RECT 13012.505 1048.035 13012.785 1194.235 ;
      RECT 13011.945 1048.035 13012.225 1194.475 ;
      RECT 13011.385 1048.035 13011.665 1194.715 ;
      RECT 13010.825 1048.035 13011.105 1194.955 ;
      RECT 13010.265 1046.935 13010.545 1194.955 ;
      RECT 13009.705 1048.035 13009.985 1194.715 ;
      RECT 13009.145 1046.935 13009.425 1194.47 ;
      RECT 13008.585 1048.035 13008.865 1194.23 ;
      RECT 13008.025 1046.935 13008.305 1193.99 ;
      RECT 13007.465 1048.035 13007.745 1193.75 ;
      RECT 13006.905 1048.035 13007.185 1193.51 ;
      RECT 13006.345 1048.035 13006.625 1193.27 ;
      RECT 13005.785 1048.035 13006.065 1193.03 ;
      RECT 13005.225 1048.035 13005.505 1192.79 ;
      RECT 13004.665 1048.035 13004.945 1192.55 ;
      RECT 13004.105 1048.035 13004.385 1192.31 ;
      RECT 13003.545 1048.035 13003.825 1192.07 ;
      RECT 13002.985 1046.935 13003.265 1191.83 ;
      RECT 13002.425 1048.035 13002.705 1191.59 ;
      RECT 13001.865 1046.935 13002.145 1191.35 ;
      RECT 13001.305 1048.035 13001.585 1191.11 ;
      RECT 13000.745 1048.035 13001.025 1190.87 ;
      RECT 13000.185 1048.035 13000.465 1190.63 ;
      RECT 12986.745 1048.035 12987.025 1194.03 ;
      RECT 12986.185 1048.035 12986.465 1194.27 ;
      RECT 12985.625 1048.035 12985.905 1194.515 ;
      RECT 12985.065 1048.035 12985.345 1194.755 ;
      RECT 12984.505 1048.035 12984.785 1194.995 ;
      RECT 12983.945 1048.035 12984.225 1194.995 ;
      RECT 12983.385 1048.035 12983.665 1194.755 ;
      RECT 12982.825 1048.035 12983.105 1194.515 ;
      RECT 12982.265 1048.035 12982.545 1187.5 ;
      RECT 12981.705 1048.035 12981.985 1187.26 ;
      RECT 12981.145 1048.035 12981.425 1187.02 ;
      RECT 12980.585 1046.935 12980.865 1186.78 ;
      RECT 12980.025 1048.035 12980.305 1186.54 ;
      RECT 12979.465 1046.935 12979.745 1186.3 ;
      RECT 12978.905 1048.035 12979.185 1186.06 ;
      RECT 12978.345 1048.035 12978.625 1185.82 ;
      RECT 12977.785 1048.035 12978.065 1185.58 ;
      RECT 12977.225 1046.935 12977.505 1185.34 ;
      RECT 12976.665 1048.035 12976.945 1185.1 ;
      RECT 12976.105 1046.935 12976.385 1184.86 ;
      RECT 12975.545 1048.035 12975.825 1184.62 ;
      RECT 12974.985 1046.935 12975.265 1184.38 ;
      RECT 12974.425 1048.035 12974.705 1184.14 ;
      RECT 12973.865 1048.035 12974.145 1183.9 ;
      RECT 12933.545 1048.035 12933.825 1192.795 ;
      RECT 12932.985 1048.035 12933.265 1193.035 ;
      RECT 12932.425 1048.035 12932.705 1193.28 ;
      RECT 12931.865 1048.035 12932.145 1193.52 ;
      RECT 12931.305 1048.035 12931.585 1193.76 ;
      RECT 12930.745 1048.035 12931.025 1194 ;
      RECT 12930.185 1048.035 12930.465 1194.24 ;
      RECT 12929.625 1048.035 12929.905 1194.48 ;
      RECT 12929.065 1048.035 12929.345 1194.72 ;
      RECT 12928.505 1048.035 12928.785 1194.96 ;
      RECT 12927.945 1046.935 12928.225 1195.2 ;
      RECT 12927.385 1048.035 12927.665 1195.44 ;
      RECT 12926.825 1046.935 12927.105 1195.68 ;
      RECT 12926.265 1048.035 12926.545 1195.92 ;
      RECT 12925.705 1046.935 12925.985 1196.16 ;
      RECT 12925.145 1048.035 12925.425 1196.16 ;
      RECT 12924.585 1048.035 12924.865 1195.92 ;
      RECT 12924.025 1048.035 12924.305 1195.68 ;
      RECT 12923.465 1048.035 12923.745 1195.44 ;
      RECT 12922.905 1048.035 12923.185 1195.2 ;
      RECT 12922.345 1048.035 12922.625 1194.96 ;
      RECT 12921.785 1048.035 12922.065 1194.72 ;
      RECT 12921.225 1048.035 12921.505 1194.48 ;
      RECT 12912.265 1046.935 12912.545 1194.51 ;
      RECT 12911.705 1048.035 12911.985 1194.75 ;
      RECT 12911.145 1046.935 12911.425 1194.99 ;
      RECT 12910.585 1048.035 12910.865 1195.205 ;
      RECT 12910.025 1048.035 12910.305 1194.78 ;
      RECT 12909.465 1048.035 12909.745 1194.54 ;
      RECT 12908.905 1048.035 12909.185 1194.3 ;
      RECT 12908.345 1048.035 12908.625 1194.06 ;
      RECT 12907.785 1048.035 12908.065 1193.82 ;
      RECT 12907.225 1048.035 12907.505 1193.58 ;
      RECT 12906.665 1048.035 12906.945 1193.34 ;
      RECT 12906.105 1048.035 12906.385 1193.1 ;
      RECT 12905.545 1048.035 12905.825 1192.86 ;
      RECT 12904.985 1048.035 12905.265 1192.62 ;
      RECT 12902.465 1048.035 12902.745 1191.795 ;
      RECT 12901.905 1048.035 12902.185 1191.555 ;
      RECT 12901.345 1048.035 12901.625 1191.315 ;
      RECT 12900.785 1046.935 12901.065 1191.075 ;
      RECT 12900.225 1048.035 12900.505 1190.835 ;
      RECT 12899.665 1046.935 12899.945 1190.595 ;
      RECT 12899.105 1048.035 12899.385 1190.355 ;
      RECT 12898.545 1048.035 12898.825 1190.115 ;
      RECT 12871.945 1048.035 12872.225 1201.16 ;
      RECT 12871.385 1046.935 12871.665 1201.4 ;
      RECT 12870.825 1048.035 12871.105 1201.64 ;
      RECT 12870.265 1046.935 12870.545 1201.885 ;
      RECT 12869.705 1048.035 12869.985 1202.125 ;
      RECT 12869.145 1046.935 12869.425 1202.365 ;
      RECT 12868.585 1048.035 12868.865 1202.605 ;
      RECT 12868.025 1048.035 12868.305 1202.845 ;
      RECT 12867.465 1048.035 12867.745 1188.465 ;
      RECT 12866.905 1048.035 12867.185 1188.225 ;
      RECT 12866.345 1048.035 12866.625 1187.985 ;
      RECT 12865.785 1048.035 12866.065 1187.745 ;
      RECT 12865.225 1048.035 12865.505 1187.505 ;
      RECT 12864.665 1048.035 12864.945 1187.265 ;
      RECT 12864.105 1048.035 12864.385 1187.025 ;
      RECT 12863.545 1048.035 12863.825 1186.785 ;
      RECT 12862.985 1048.035 12863.265 1186.545 ;
      RECT 12862.425 1048.035 12862.705 1186.305 ;
      RECT 12861.865 1046.935 12862.145 1186.065 ;
      RECT 12861.305 1048.035 12861.585 1185.825 ;
      RECT 12860.745 1046.935 12861.025 1185.585 ;
      RECT 12860.185 1048.035 12860.465 1185.345 ;
      RECT 12846.185 1046.935 12846.465 1191.465 ;
      RECT 12845.625 1048.035 12845.905 1191.225 ;
      RECT 12845.065 1048.035 12845.345 1190.985 ;
      RECT 12844.505 1048.035 12844.785 1190.745 ;
      RECT 12843.945 1048.035 12844.225 1190.505 ;
      RECT 12843.385 1048.035 12843.665 1190.265 ;
      RECT 12842.825 1048.035 12843.105 1190.025 ;
      RECT 12842.265 1048.035 12842.545 1189.785 ;
      RECT 12841.705 1048.035 12841.985 1189.545 ;
      RECT 12841.145 1046.935 12841.425 1189.305 ;
      RECT 12840.585 1048.035 12840.865 1189.065 ;
      RECT 12840.025 1046.935 12840.305 1188.825 ;
      RECT 12839.465 1048.035 12839.745 1188.585 ;
      RECT 12838.905 1048.035 12839.185 1188.345 ;
      RECT 12838.345 1048.035 12838.625 1188.105 ;
      RECT 12837.785 1048.035 12838.065 1187.865 ;
      RECT 12837.225 1048.035 12837.505 1187.625 ;
      RECT 12836.665 1048.035 12836.945 1187.385 ;
      RECT 12836.105 1048.035 12836.385 1187.145 ;
      RECT 12835.545 1048.035 12835.825 1186.905 ;
      RECT 12834.985 1048.035 12835.265 1186.665 ;
      RECT 12834.425 1048.035 12834.705 1186.425 ;
      RECT 12833.865 1048.035 12834.145 1186.185 ;
      RECT 12794.665 1048.035 12794.945 1193.09 ;
      RECT 12794.105 1048.035 12794.385 1193.33 ;
      RECT 12793.545 1048.035 12793.825 1193.57 ;
      RECT 12792.985 1046.935 12793.265 1193.81 ;
      RECT 12792.425 1048.035 12792.705 1194.05 ;
      RECT 12791.865 1046.935 12792.145 1194.29 ;
      RECT 12791.305 1048.035 12791.585 1194.53 ;
      RECT 12790.745 1048.035 12791.025 1194.77 ;
      RECT 12790.185 1048.035 12790.465 1195.01 ;
      RECT 12789.625 1046.935 12789.905 1195.25 ;
      RECT 12789.065 1048.035 12789.345 1195.49 ;
      RECT 12788.505 1046.935 12788.785 1195.73 ;
      RECT 12787.945 1048.035 12788.225 1195.97 ;
      RECT 12787.385 1046.935 12787.665 1196.21 ;
      RECT 12786.825 1048.035 12787.105 1196.45 ;
      RECT 12786.265 1048.035 12786.545 1196.69 ;
      RECT 12785.705 1048.035 12785.985 1196.69 ;
      RECT 12785.145 1048.035 12785.425 1196.45 ;
      RECT 12784.585 1048.035 12784.865 1196.21 ;
      RECT 12784.025 1048.035 12784.305 1195.97 ;
      RECT 12783.465 1048.035 12783.745 1195.73 ;
      RECT 12782.905 1048.035 12783.185 1195.49 ;
      RECT 12782.345 1048.035 12782.625 1195.25 ;
      RECT 12781.785 1048.035 12782.065 1195.01 ;
      RECT 12781.225 1048.035 12781.505 1194.77 ;
      RECT 12772.265 1048.035 12772.545 1194.285 ;
      RECT 12771.705 1046.935 12771.985 1194.045 ;
      RECT 12771.145 1048.035 12771.425 1193.805 ;
      RECT 12770.585 1046.935 12770.865 1193.565 ;
      RECT 12770.025 1048.035 12770.305 1193.325 ;
      RECT 12769.465 1046.935 12769.745 1193.085 ;
      RECT 12768.905 1048.035 12769.185 1192.845 ;
      RECT 12768.345 1048.035 12768.625 1192.605 ;
      RECT 12767.785 1048.035 12768.065 1192.365 ;
      RECT 12767.225 1048.035 12767.505 1192.125 ;
      RECT 12766.665 1048.035 12766.945 1191.885 ;
      RECT 12766.105 1048.035 12766.385 1191.645 ;
      RECT 12765.545 1048.035 12765.825 1191.405 ;
      RECT 12764.985 1048.035 12765.265 1191.165 ;
      RECT 12762.465 1046.935 12762.745 1192.885 ;
      RECT 12761.905 1048.035 12762.185 1192.645 ;
      RECT 12761.345 1046.935 12761.625 1192.405 ;
      RECT 12760.785 1048.035 12761.065 1192.165 ;
      RECT 12760.225 1048.035 12760.505 1191.925 ;
      RECT 12759.665 1048.035 12759.945 1191.685 ;
      RECT 12759.105 1048.035 12759.385 1191.445 ;
      RECT 12758.545 1048.035 12758.825 1191.205 ;
      RECT 12732.505 1048.035 12732.785 1188.855 ;
      RECT 12731.945 1048.035 12732.225 1189.095 ;
      RECT 12731.385 1048.035 12731.665 1189.335 ;
      RECT 12730.825 1048.035 12731.105 1189.58 ;
      RECT 12730.265 1048.035 12730.545 1189.82 ;
      RECT 12729.705 1048.035 12729.985 1190.06 ;
      RECT 12729.145 1048.035 12729.425 1190.06 ;
      RECT 12728.585 1048.035 12728.865 1189.82 ;
      RECT 12728.025 1048.035 12728.305 1189.58 ;
      RECT 12727.465 1046.935 12727.745 1189.34 ;
      RECT 12726.905 1048.035 12727.185 1189.1 ;
      RECT 12726.345 1046.935 12726.625 1188.86 ;
      RECT 12725.785 1048.035 12726.065 1188.62 ;
      RECT 12725.225 1048.035 12725.505 1188.38 ;
      RECT 12724.665 1048.035 12724.945 1188.14 ;
      RECT 12724.105 1046.935 12724.385 1187.9 ;
      RECT 12723.545 1048.035 12723.825 1187.66 ;
      RECT 12722.985 1046.935 12723.265 1187.42 ;
      RECT 12722.425 1048.035 12722.705 1187.18 ;
      RECT 12721.865 1046.935 12722.145 1186.94 ;
      RECT 12721.305 1048.035 12721.585 1186.7 ;
      RECT 12720.745 1048.035 12721.025 1186.46 ;
      RECT 12720.185 1048.035 12720.465 1186.22 ;
      RECT 12719.625 1048.035 12719.905 1185.98 ;
      RECT 12706.185 1048.035 12706.465 1191.78 ;
      RECT 12705.625 1048.035 12705.905 1191.54 ;
      RECT 12705.065 1048.035 12705.345 1191.3 ;
      RECT 12704.505 1048.035 12704.785 1191.06 ;
      RECT 12703.945 1048.035 12704.225 1190.82 ;
      RECT 12703.385 1048.035 12703.665 1190.58 ;
      RECT 12702.825 1048.035 12703.105 1190.34 ;
      RECT 12702.265 1048.035 12702.545 1190.1 ;
      RECT 12701.705 1046.935 12701.985 1189.86 ;
      RECT 12701.145 1048.035 12701.425 1189.62 ;
      RECT 12700.585 1046.935 12700.865 1189.3 ;
      RECT 12700.025 1048.035 12700.305 1189.14 ;
      RECT 12699.465 1046.935 12699.745 1188.9 ;
      RECT 12698.905 1048.035 12699.185 1188.66 ;
      RECT 12698.345 1048.035 12698.625 1188.42 ;
      RECT 12697.785 1048.035 12698.065 1188.18 ;
      RECT 12697.225 1048.035 12697.505 1187.94 ;
      RECT 12696.665 1048.035 12696.945 1187.7 ;
      RECT 12696.105 1048.035 12696.385 1187.46 ;
      RECT 12695.545 1048.035 12695.825 1187.22 ;
      RECT 12694.985 1048.035 12695.265 1186.98 ;
      RECT 12694.425 1046.935 12694.705 1186.74 ;
      RECT 12693.865 1048.035 12694.145 1186.5 ;
      RECT 12693.305 1046.935 12693.585 1186.26 ;
      RECT 12654.105 1048.035 12654.385 1191.87 ;
      RECT 12653.545 1048.035 12653.825 1192.11 ;
      RECT 12652.985 1048.035 12653.265 1192.35 ;
      RECT 12652.425 1048.035 12652.705 1192.59 ;
      RECT 12651.865 1048.035 12652.145 1192.83 ;
      RECT 12651.305 1048.035 12651.585 1193.07 ;
      RECT 12650.745 1048.035 12651.025 1193.31 ;
      RECT 12650.185 1048.035 12650.465 1193.55 ;
      RECT 12649.625 1048.035 12649.905 1193.79 ;
      RECT 12649.065 1048.035 12649.345 1194.03 ;
      RECT 12648.505 1048.035 12648.785 1194.27 ;
      RECT 12647.945 1048.035 12648.225 1194.51 ;
      RECT 12647.385 1048.035 12647.665 1194.75 ;
      RECT 12646.825 1048.035 12647.105 1194.75 ;
      RECT 12646.265 1046.935 12646.545 1194.51 ;
      RECT 12645.705 1048.035 12645.985 1194.27 ;
      RECT 12645.145 1046.935 12645.425 1194.03 ;
      RECT 12644.585 1048.035 12644.865 1193.79 ;
      RECT 12644.025 1048.035 12644.305 1193.55 ;
      RECT 12643.465 1048.035 12643.745 1193.31 ;
      RECT 12642.905 1046.935 12643.185 1193.045 ;
      RECT 12642.345 1048.035 12642.625 1192.805 ;
      RECT 12641.785 1046.935 12642.065 1192.565 ;
      RECT 12641.225 1048.035 12641.505 1192.325 ;
      RECT 12632.265 1046.935 12632.545 1186.16 ;
      RECT 12631.705 1048.035 12631.985 1186.4 ;
      RECT 12631.145 1048.035 12631.425 1186.64 ;
      RECT 12630.585 1048.035 12630.865 1186.64 ;
      RECT 12630.025 1048.035 12630.305 1186.4 ;
      RECT 12629.465 1048.035 12629.745 1186.16 ;
      RECT 12628.905 1048.035 12629.185 1185.92 ;
      RECT 12628.345 1048.035 12628.625 1185.68 ;
      RECT 12627.785 1048.035 12628.065 1185.44 ;
      RECT 12627.225 1048.035 12627.505 1185.2 ;
      RECT 12626.665 1048.035 12626.945 1184.96 ;
      RECT 12626.105 1048.035 12626.385 1184.72 ;
      RECT 12625.545 1048.035 12625.825 1184.48 ;
      RECT 12624.985 1046.935 12625.265 1184.24 ;
      RECT 12622.465 1048.035 12622.745 1185.96 ;
      RECT 12621.905 1046.935 12622.185 1185.72 ;
      RECT 12621.345 1048.035 12621.625 1185.48 ;
      RECT 12620.785 1046.935 12621.065 1185.24 ;
      RECT 12620.225 1048.035 12620.505 1185 ;
      RECT 12619.665 1048.035 12619.945 1184.76 ;
      RECT 12619.105 1048.035 12619.385 1184.52 ;
      RECT 12593.065 1048.035 12593.345 1187.305 ;
      RECT 12592.505 1048.035 12592.785 1187.545 ;
      RECT 12591.945 1048.035 12592.225 1187.785 ;
      RECT 12591.385 1048.035 12591.665 1188.025 ;
      RECT 12590.825 1048.035 12591.105 1188.265 ;
      RECT 12590.265 1046.935 12590.545 1188.505 ;
      RECT 12589.705 1048.035 12589.985 1188.745 ;
      RECT 12589.145 1046.935 12589.425 1188.985 ;
      RECT 12588.585 1048.035 12588.865 1189.225 ;
      RECT 12588.025 1048.035 12588.305 1189.465 ;
      RECT 12587.465 1048.035 12587.745 1189.705 ;
      RECT 12586.905 1048.035 12587.185 1189.945 ;
      RECT 12586.345 1048.035 12586.625 1190.185 ;
      RECT 12585.785 1048.035 12586.065 1190.425 ;
      RECT 12585.225 1048.035 12585.505 1190.665 ;
      RECT 12584.665 1048.035 12584.945 1190.665 ;
      RECT 12584.105 1048.035 12584.385 1190.425 ;
      RECT 12583.545 1048.035 12583.825 1190.185 ;
      RECT 12582.985 1048.035 12583.265 1189.945 ;
      RECT 12582.425 1048.035 12582.705 1189.7 ;
      RECT 12581.865 1048.035 12582.145 1189.46 ;
      RECT 12581.305 1048.035 12581.585 1189.22 ;
      RECT 12580.745 1046.935 12581.025 1188.98 ;
      RECT 12580.185 1048.035 12580.465 1188.74 ;
      RECT 12566.745 1046.935 12567.025 1186.22 ;
      RECT 12566.185 1048.035 12566.465 1185.98 ;
      RECT 12565.625 1048.035 12565.905 1185.74 ;
      RECT 12565.065 1048.035 12565.345 1185.5 ;
      RECT 12564.505 1046.935 12564.785 1185.26 ;
      RECT 12563.945 1048.035 12564.225 1185.02 ;
      RECT 12563.385 1046.935 12563.665 1184.78 ;
      RECT 12562.825 1048.035 12563.105 1184.54 ;
      RECT 12562.265 1046.935 12562.545 1184.3 ;
      RECT 12561.705 1048.035 12561.985 1184.06 ;
      RECT 12561.145 1048.035 12561.425 1183.82 ;
      RECT 12560.585 1048.035 12560.865 1183.58 ;
      RECT 12560.025 1048.035 12560.305 1183.34 ;
      RECT 12559.465 1048.035 12559.745 1183.1 ;
      RECT 12558.905 1048.035 12559.185 1182.86 ;
      RECT 12558.345 1048.035 12558.625 1182.62 ;
      RECT 12557.785 1048.035 12558.065 1182.38 ;
      RECT 12557.225 1048.035 12557.505 1182.14 ;
      RECT 12556.665 1048.035 12556.945 1181.9 ;
      RECT 12556.105 1048.035 12556.385 1181.66 ;
      RECT 12555.545 1048.035 12555.825 1181.42 ;
      RECT 12554.985 1046.935 12555.265 1181.18 ;
      RECT 12554.425 1048.035 12554.705 1180.94 ;
      RECT 12553.865 1046.935 12554.145 1180.7 ;
      RECT 12514.105 1048.035 12514.385 1191.17 ;
      RECT 12513.545 1046.935 12513.825 1191.41 ;
      RECT 12512.985 1048.035 12513.265 1191.65 ;
      RECT 12512.425 1048.035 12512.705 1191.89 ;
      RECT 12511.865 1048.035 12512.145 1192.13 ;
      RECT 12511.305 1048.035 12511.585 1192.37 ;
      RECT 12510.745 1048.035 12511.025 1192.61 ;
      RECT 12510.185 1048.035 12510.465 1192.855 ;
      RECT 12509.625 1048.035 12509.905 1193.095 ;
      RECT 12509.065 1048.035 12509.345 1193.335 ;
      RECT 12508.505 1046.935 12508.785 1193.575 ;
      RECT 12507.945 1048.035 12508.225 1193.815 ;
      RECT 12507.385 1046.935 12507.665 1194.055 ;
      RECT 12506.825 1048.035 12507.105 1194.295 ;
      RECT 12506.265 1048.035 12506.545 1194.535 ;
      RECT 12505.705 1048.035 12505.985 1194.775 ;
      RECT 12505.145 1048.035 12505.425 1195.015 ;
      RECT 12504.585 1048.035 12504.865 1195.255 ;
      RECT 12504.025 1048.035 12504.305 1195.495 ;
      RECT 12503.465 1048.035 12503.745 1195.735 ;
      RECT 12502.905 1048.035 12503.185 1195.975 ;
      RECT 12502.345 1048.035 12502.625 1196.215 ;
      RECT 12501.785 1048.035 12502.065 1196.455 ;
      RECT 12501.225 1048.035 12501.505 1196.695 ;
      RECT 12492.265 1048.035 12492.545 1192.28 ;
      RECT 12491.705 1048.035 12491.985 1192.04 ;
      RECT 12491.145 1048.035 12491.425 1191.8 ;
      RECT 12490.585 1046.935 12490.865 1191.56 ;
      RECT 12490.025 1048.035 12490.305 1191.32 ;
      RECT 12489.465 1046.935 12489.745 1191.08 ;
      RECT 12488.905 1048.035 12489.185 1190.84 ;
      RECT 12488.345 1048.035 12488.625 1190.6 ;
      RECT 12487.785 1048.035 12488.065 1190.36 ;
      RECT 12487.225 1046.935 12487.505 1190.12 ;
      RECT 12486.665 1048.035 12486.945 1189.88 ;
      RECT 12486.105 1046.935 12486.385 1189.64 ;
      RECT 12485.545 1048.035 12485.825 1189.4 ;
      RECT 12484.985 1046.935 12485.265 1189.16 ;
      RECT 12482.465 1048.035 12482.745 1181.56 ;
      RECT 12481.905 1048.035 12482.185 1181.32 ;
      RECT 12481.345 1048.035 12481.625 1181.08 ;
      RECT 12480.785 1048.035 12481.065 1180.84 ;
      RECT 12480.225 1048.035 12480.505 1180.6 ;
      RECT 12479.665 1048.035 12479.945 1180.36 ;
      RECT 12479.105 1048.035 12479.385 1180.12 ;
      RECT 12453.065 1048.035 12453.345 1193.995 ;
      RECT 12452.505 1048.035 12452.785 1194.235 ;
      RECT 12451.945 1048.035 12452.225 1194.475 ;
      RECT 12451.385 1048.035 12451.665 1194.715 ;
      RECT 12450.825 1048.035 12451.105 1194.955 ;
      RECT 12450.265 1046.935 12450.545 1194.955 ;
      RECT 12449.705 1048.035 12449.985 1194.715 ;
      RECT 12449.145 1046.935 12449.425 1194.47 ;
      RECT 12448.585 1048.035 12448.865 1194.23 ;
      RECT 12448.025 1046.935 12448.305 1193.99 ;
      RECT 12447.465 1048.035 12447.745 1193.75 ;
      RECT 12446.905 1048.035 12447.185 1193.51 ;
      RECT 12446.345 1048.035 12446.625 1193.27 ;
      RECT 12445.785 1048.035 12446.065 1193.03 ;
      RECT 12445.225 1048.035 12445.505 1192.79 ;
      RECT 12444.665 1048.035 12444.945 1192.55 ;
      RECT 12444.105 1048.035 12444.385 1192.31 ;
      RECT 12443.545 1048.035 12443.825 1192.07 ;
      RECT 12442.985 1046.935 12443.265 1191.83 ;
      RECT 12442.425 1048.035 12442.705 1191.59 ;
      RECT 12441.865 1046.935 12442.145 1191.35 ;
      RECT 12441.305 1048.035 12441.585 1191.11 ;
      RECT 12440.745 1048.035 12441.025 1190.87 ;
      RECT 12440.185 1048.035 12440.465 1190.63 ;
      RECT 12426.745 1048.035 12427.025 1194.03 ;
      RECT 12426.185 1048.035 12426.465 1194.27 ;
      RECT 12425.625 1048.035 12425.905 1194.515 ;
      RECT 12425.065 1048.035 12425.345 1194.755 ;
      RECT 12424.505 1048.035 12424.785 1194.995 ;
      RECT 12423.945 1048.035 12424.225 1194.995 ;
      RECT 12423.385 1048.035 12423.665 1194.755 ;
      RECT 12422.825 1048.035 12423.105 1194.515 ;
      RECT 12422.265 1048.035 12422.545 1187.5 ;
      RECT 12421.705 1048.035 12421.985 1187.26 ;
      RECT 12421.145 1048.035 12421.425 1187.02 ;
      RECT 12420.585 1046.935 12420.865 1186.78 ;
      RECT 12420.025 1048.035 12420.305 1186.54 ;
      RECT 12419.465 1046.935 12419.745 1186.3 ;
      RECT 12418.905 1048.035 12419.185 1186.06 ;
      RECT 12418.345 1048.035 12418.625 1185.82 ;
      RECT 12417.785 1048.035 12418.065 1185.58 ;
      RECT 12417.225 1046.935 12417.505 1185.34 ;
      RECT 12416.665 1048.035 12416.945 1185.1 ;
      RECT 12416.105 1046.935 12416.385 1184.86 ;
      RECT 12415.545 1048.035 12415.825 1184.62 ;
      RECT 12414.985 1046.935 12415.265 1184.38 ;
      RECT 12414.425 1048.035 12414.705 1184.14 ;
      RECT 12413.865 1048.035 12414.145 1183.9 ;
      RECT 12373.545 1048.035 12373.825 1192.795 ;
      RECT 12372.985 1048.035 12373.265 1193.035 ;
      RECT 12372.425 1048.035 12372.705 1193.28 ;
      RECT 12371.865 1048.035 12372.145 1193.52 ;
      RECT 12371.305 1048.035 12371.585 1193.76 ;
      RECT 12370.745 1048.035 12371.025 1194 ;
      RECT 12370.185 1048.035 12370.465 1194.24 ;
      RECT 12369.625 1048.035 12369.905 1194.48 ;
      RECT 12369.065 1048.035 12369.345 1194.72 ;
      RECT 12368.505 1048.035 12368.785 1194.96 ;
      RECT 12367.945 1046.935 12368.225 1195.2 ;
      RECT 12367.385 1048.035 12367.665 1195.44 ;
      RECT 12366.825 1046.935 12367.105 1195.68 ;
      RECT 12366.265 1048.035 12366.545 1195.92 ;
      RECT 12365.705 1046.935 12365.985 1196.16 ;
      RECT 12365.145 1048.035 12365.425 1196.16 ;
      RECT 12364.585 1048.035 12364.865 1195.92 ;
      RECT 12364.025 1048.035 12364.305 1195.68 ;
      RECT 12363.465 1048.035 12363.745 1195.44 ;
      RECT 12362.905 1048.035 12363.185 1195.2 ;
      RECT 12362.345 1048.035 12362.625 1194.96 ;
      RECT 12361.785 1048.035 12362.065 1194.72 ;
      RECT 12361.225 1048.035 12361.505 1194.48 ;
      RECT 12352.265 1046.935 12352.545 1194.51 ;
      RECT 12351.705 1048.035 12351.985 1194.75 ;
      RECT 12351.145 1046.935 12351.425 1194.99 ;
      RECT 12350.585 1048.035 12350.865 1195.205 ;
      RECT 12350.025 1048.035 12350.305 1194.78 ;
      RECT 12349.465 1048.035 12349.745 1194.54 ;
      RECT 12348.905 1048.035 12349.185 1194.3 ;
      RECT 12348.345 1048.035 12348.625 1194.06 ;
      RECT 12347.785 1048.035 12348.065 1193.82 ;
      RECT 12347.225 1048.035 12347.505 1193.58 ;
      RECT 12346.665 1048.035 12346.945 1193.34 ;
      RECT 12346.105 1048.035 12346.385 1193.1 ;
      RECT 12345.545 1048.035 12345.825 1192.86 ;
      RECT 12344.985 1048.035 12345.265 1192.62 ;
      RECT 12342.465 1048.035 12342.745 1191.795 ;
      RECT 12341.905 1048.035 12342.185 1191.555 ;
      RECT 12341.345 1048.035 12341.625 1191.315 ;
      RECT 12340.785 1046.935 12341.065 1191.075 ;
      RECT 12340.225 1048.035 12340.505 1190.835 ;
      RECT 12339.665 1046.935 12339.945 1190.595 ;
      RECT 12339.105 1048.035 12339.385 1190.355 ;
      RECT 12338.545 1048.035 12338.825 1190.115 ;
      RECT 12311.945 1048.035 12312.225 1201.16 ;
      RECT 12311.385 1046.935 12311.665 1201.4 ;
      RECT 12310.825 1048.035 12311.105 1201.64 ;
      RECT 12310.265 1046.935 12310.545 1201.885 ;
      RECT 12309.705 1048.035 12309.985 1202.125 ;
      RECT 12309.145 1046.935 12309.425 1202.365 ;
      RECT 12308.585 1048.035 12308.865 1202.605 ;
      RECT 12308.025 1048.035 12308.305 1202.845 ;
      RECT 12307.465 1048.035 12307.745 1188.465 ;
      RECT 12306.905 1048.035 12307.185 1188.225 ;
      RECT 12306.345 1048.035 12306.625 1187.985 ;
      RECT 12305.785 1048.035 12306.065 1187.745 ;
      RECT 12305.225 1048.035 12305.505 1187.505 ;
      RECT 12304.665 1048.035 12304.945 1187.265 ;
      RECT 12304.105 1048.035 12304.385 1187.025 ;
      RECT 12303.545 1048.035 12303.825 1186.785 ;
      RECT 12302.985 1048.035 12303.265 1186.545 ;
      RECT 12302.425 1048.035 12302.705 1186.305 ;
      RECT 12301.865 1046.935 12302.145 1186.065 ;
      RECT 12301.305 1048.035 12301.585 1185.825 ;
      RECT 12300.745 1046.935 12301.025 1185.585 ;
      RECT 12300.185 1048.035 12300.465 1185.345 ;
      RECT 12286.185 1046.935 12286.465 1191.465 ;
      RECT 12285.625 1048.035 12285.905 1191.225 ;
      RECT 12285.065 1048.035 12285.345 1190.985 ;
      RECT 12284.505 1048.035 12284.785 1190.745 ;
      RECT 12283.945 1048.035 12284.225 1190.505 ;
      RECT 12283.385 1048.035 12283.665 1190.265 ;
      RECT 12282.825 1048.035 12283.105 1190.025 ;
      RECT 12282.265 1048.035 12282.545 1189.785 ;
      RECT 12281.705 1048.035 12281.985 1189.545 ;
      RECT 12281.145 1046.935 12281.425 1189.305 ;
      RECT 12280.585 1048.035 12280.865 1189.065 ;
      RECT 12280.025 1046.935 12280.305 1188.825 ;
      RECT 12279.465 1048.035 12279.745 1188.585 ;
      RECT 12278.905 1048.035 12279.185 1188.345 ;
      RECT 12278.345 1048.035 12278.625 1188.105 ;
      RECT 12277.785 1048.035 12278.065 1187.865 ;
      RECT 12277.225 1048.035 12277.505 1187.625 ;
      RECT 12276.665 1048.035 12276.945 1187.385 ;
      RECT 12276.105 1048.035 12276.385 1187.145 ;
      RECT 12275.545 1048.035 12275.825 1186.905 ;
      RECT 12274.985 1048.035 12275.265 1186.665 ;
      RECT 12274.425 1048.035 12274.705 1186.425 ;
      RECT 12273.865 1048.035 12274.145 1186.185 ;
      RECT 12234.665 1048.035 12234.945 1193.09 ;
      RECT 12234.105 1048.035 12234.385 1193.33 ;
      RECT 12233.545 1048.035 12233.825 1193.57 ;
      RECT 12232.985 1046.935 12233.265 1193.81 ;
      RECT 12232.425 1048.035 12232.705 1194.05 ;
      RECT 12231.865 1046.935 12232.145 1194.29 ;
      RECT 12231.305 1048.035 12231.585 1194.53 ;
      RECT 12230.745 1048.035 12231.025 1194.77 ;
      RECT 12230.185 1048.035 12230.465 1195.01 ;
      RECT 12229.625 1046.935 12229.905 1195.25 ;
      RECT 12229.065 1048.035 12229.345 1195.49 ;
      RECT 12228.505 1046.935 12228.785 1195.73 ;
      RECT 12227.945 1048.035 12228.225 1195.97 ;
      RECT 12227.385 1046.935 12227.665 1196.21 ;
      RECT 12226.825 1048.035 12227.105 1196.45 ;
      RECT 12226.265 1048.035 12226.545 1196.69 ;
      RECT 12225.705 1048.035 12225.985 1196.69 ;
      RECT 12225.145 1048.035 12225.425 1196.45 ;
      RECT 12224.585 1048.035 12224.865 1196.21 ;
      RECT 12224.025 1048.035 12224.305 1195.97 ;
      RECT 12223.465 1048.035 12223.745 1195.73 ;
      RECT 12222.905 1048.035 12223.185 1195.49 ;
      RECT 12222.345 1048.035 12222.625 1195.25 ;
      RECT 12221.785 1048.035 12222.065 1195.01 ;
      RECT 12221.225 1048.035 12221.505 1194.77 ;
      RECT 12212.265 1048.035 12212.545 1194.285 ;
      RECT 12211.705 1046.935 12211.985 1194.045 ;
      RECT 12211.145 1048.035 12211.425 1193.805 ;
      RECT 12210.585 1046.935 12210.865 1193.565 ;
      RECT 12210.025 1048.035 12210.305 1193.325 ;
      RECT 12209.465 1046.935 12209.745 1193.085 ;
      RECT 12208.905 1048.035 12209.185 1192.845 ;
      RECT 12208.345 1048.035 12208.625 1192.605 ;
      RECT 12207.785 1048.035 12208.065 1192.365 ;
      RECT 12207.225 1048.035 12207.505 1192.125 ;
      RECT 12206.665 1048.035 12206.945 1191.885 ;
      RECT 12206.105 1048.035 12206.385 1191.645 ;
      RECT 12205.545 1048.035 12205.825 1191.405 ;
      RECT 12204.985 1048.035 12205.265 1191.165 ;
      RECT 12202.465 1046.935 12202.745 1192.885 ;
      RECT 12201.905 1048.035 12202.185 1192.645 ;
      RECT 12201.345 1046.935 12201.625 1192.405 ;
      RECT 12200.785 1048.035 12201.065 1192.165 ;
      RECT 12200.225 1048.035 12200.505 1191.925 ;
      RECT 12199.665 1048.035 12199.945 1191.685 ;
      RECT 12199.105 1048.035 12199.385 1191.445 ;
      RECT 12198.545 1048.035 12198.825 1191.205 ;
      RECT 12172.505 1048.035 12172.785 1188.855 ;
      RECT 12171.945 1048.035 12172.225 1189.095 ;
      RECT 12171.385 1048.035 12171.665 1189.335 ;
      RECT 12170.825 1048.035 12171.105 1189.58 ;
      RECT 12170.265 1048.035 12170.545 1189.82 ;
      RECT 12169.705 1048.035 12169.985 1190.06 ;
      RECT 12169.145 1048.035 12169.425 1190.06 ;
      RECT 12168.585 1048.035 12168.865 1189.82 ;
      RECT 12168.025 1048.035 12168.305 1189.58 ;
      RECT 12167.465 1046.935 12167.745 1189.34 ;
      RECT 12166.905 1048.035 12167.185 1189.1 ;
      RECT 12166.345 1046.935 12166.625 1188.86 ;
      RECT 12165.785 1048.035 12166.065 1188.62 ;
      RECT 12165.225 1048.035 12165.505 1188.38 ;
      RECT 12164.665 1048.035 12164.945 1188.14 ;
      RECT 12164.105 1046.935 12164.385 1187.9 ;
      RECT 12163.545 1048.035 12163.825 1187.66 ;
      RECT 12162.985 1046.935 12163.265 1187.42 ;
      RECT 12162.425 1048.035 12162.705 1187.18 ;
      RECT 12161.865 1046.935 12162.145 1186.94 ;
      RECT 12161.305 1048.035 12161.585 1186.7 ;
      RECT 12160.745 1048.035 12161.025 1186.46 ;
      RECT 12160.185 1048.035 12160.465 1186.22 ;
      RECT 12159.625 1048.035 12159.905 1185.98 ;
      RECT 12146.185 1048.035 12146.465 1191.78 ;
      RECT 12145.625 1048.035 12145.905 1191.54 ;
      RECT 12145.065 1048.035 12145.345 1191.3 ;
      RECT 12144.505 1048.035 12144.785 1191.06 ;
      RECT 12143.945 1048.035 12144.225 1190.82 ;
      RECT 12143.385 1048.035 12143.665 1190.58 ;
      RECT 12142.825 1048.035 12143.105 1190.34 ;
      RECT 12142.265 1048.035 12142.545 1190.1 ;
      RECT 12141.705 1046.935 12141.985 1189.86 ;
      RECT 12141.145 1048.035 12141.425 1189.62 ;
      RECT 12140.585 1046.935 12140.865 1189.3 ;
      RECT 12140.025 1048.035 12140.305 1189.14 ;
      RECT 12139.465 1046.935 12139.745 1188.9 ;
      RECT 12138.905 1048.035 12139.185 1188.66 ;
      RECT 12138.345 1048.035 12138.625 1188.42 ;
      RECT 12137.785 1048.035 12138.065 1188.18 ;
      RECT 12137.225 1048.035 12137.505 1187.94 ;
      RECT 12136.665 1048.035 12136.945 1187.7 ;
      RECT 12136.105 1048.035 12136.385 1187.46 ;
      RECT 12135.545 1048.035 12135.825 1187.22 ;
      RECT 12134.985 1048.035 12135.265 1186.98 ;
      RECT 12134.425 1046.935 12134.705 1186.74 ;
      RECT 12133.865 1048.035 12134.145 1186.5 ;
      RECT 12133.305 1046.935 12133.585 1186.26 ;
      RECT 12094.105 1048.035 12094.385 1191.87 ;
      RECT 12093.545 1048.035 12093.825 1192.11 ;
      RECT 12092.985 1048.035 12093.265 1192.35 ;
      RECT 12092.425 1048.035 12092.705 1192.59 ;
      RECT 12091.865 1048.035 12092.145 1192.83 ;
      RECT 12091.305 1048.035 12091.585 1193.07 ;
      RECT 12090.745 1048.035 12091.025 1193.31 ;
      RECT 12090.185 1048.035 12090.465 1193.55 ;
      RECT 12089.625 1048.035 12089.905 1193.79 ;
      RECT 12089.065 1048.035 12089.345 1194.03 ;
      RECT 12088.505 1048.035 12088.785 1194.27 ;
      RECT 12087.945 1048.035 12088.225 1194.51 ;
      RECT 12087.385 1048.035 12087.665 1194.75 ;
      RECT 12086.825 1048.035 12087.105 1194.75 ;
      RECT 12086.265 1046.935 12086.545 1194.51 ;
      RECT 12085.705 1048.035 12085.985 1194.27 ;
      RECT 12085.145 1046.935 12085.425 1194.03 ;
      RECT 12084.585 1048.035 12084.865 1193.79 ;
      RECT 12084.025 1048.035 12084.305 1193.55 ;
      RECT 12083.465 1048.035 12083.745 1193.31 ;
      RECT 12082.905 1046.935 12083.185 1193.045 ;
      RECT 12082.345 1048.035 12082.625 1192.805 ;
      RECT 12081.785 1046.935 12082.065 1192.565 ;
      RECT 12081.225 1048.035 12081.505 1192.325 ;
      RECT 12072.265 1046.935 12072.545 1186.16 ;
      RECT 12071.705 1048.035 12071.985 1186.4 ;
      RECT 12071.145 1048.035 12071.425 1186.64 ;
      RECT 12070.585 1048.035 12070.865 1186.64 ;
      RECT 12070.025 1048.035 12070.305 1186.4 ;
      RECT 12069.465 1048.035 12069.745 1186.16 ;
      RECT 12068.905 1048.035 12069.185 1185.92 ;
      RECT 12068.345 1048.035 12068.625 1185.68 ;
      RECT 12067.785 1048.035 12068.065 1185.44 ;
      RECT 12067.225 1048.035 12067.505 1185.2 ;
      RECT 12066.665 1048.035 12066.945 1184.96 ;
      RECT 12066.105 1048.035 12066.385 1184.72 ;
      RECT 12065.545 1048.035 12065.825 1184.48 ;
      RECT 12064.985 1046.935 12065.265 1184.24 ;
      RECT 12062.465 1048.035 12062.745 1185.96 ;
      RECT 12061.905 1046.935 12062.185 1185.72 ;
      RECT 12061.345 1048.035 12061.625 1185.48 ;
      RECT 12060.785 1046.935 12061.065 1185.24 ;
      RECT 12060.225 1048.035 12060.505 1185 ;
      RECT 12059.665 1048.035 12059.945 1184.76 ;
      RECT 12059.105 1048.035 12059.385 1184.52 ;
      RECT 12033.065 1048.035 12033.345 1187.305 ;
      RECT 12032.505 1048.035 12032.785 1187.545 ;
      RECT 12031.945 1048.035 12032.225 1187.785 ;
      RECT 12031.385 1048.035 12031.665 1188.025 ;
      RECT 12030.825 1048.035 12031.105 1188.265 ;
      RECT 12030.265 1046.935 12030.545 1188.505 ;
      RECT 12029.705 1048.035 12029.985 1188.745 ;
      RECT 12029.145 1046.935 12029.425 1188.985 ;
      RECT 12028.585 1048.035 12028.865 1189.225 ;
      RECT 12028.025 1048.035 12028.305 1189.465 ;
      RECT 12027.465 1048.035 12027.745 1189.705 ;
      RECT 12026.905 1048.035 12027.185 1189.945 ;
      RECT 12026.345 1048.035 12026.625 1190.185 ;
      RECT 12025.785 1048.035 12026.065 1190.425 ;
      RECT 12025.225 1048.035 12025.505 1190.665 ;
      RECT 12024.665 1048.035 12024.945 1190.665 ;
      RECT 12024.105 1048.035 12024.385 1190.425 ;
      RECT 12023.545 1048.035 12023.825 1190.185 ;
      RECT 12022.985 1048.035 12023.265 1189.945 ;
      RECT 12022.425 1048.035 12022.705 1189.7 ;
      RECT 12021.865 1048.035 12022.145 1189.46 ;
      RECT 12021.305 1048.035 12021.585 1189.22 ;
      RECT 12020.745 1046.935 12021.025 1188.98 ;
      RECT 12020.185 1048.035 12020.465 1188.74 ;
      RECT 12006.745 1046.935 12007.025 1186.22 ;
      RECT 12006.185 1048.035 12006.465 1185.98 ;
      RECT 12005.625 1048.035 12005.905 1185.74 ;
      RECT 12005.065 1048.035 12005.345 1185.5 ;
      RECT 12004.505 1046.935 12004.785 1185.26 ;
      RECT 12003.945 1048.035 12004.225 1185.02 ;
      RECT 12003.385 1046.935 12003.665 1184.78 ;
      RECT 12002.825 1048.035 12003.105 1184.54 ;
      RECT 12002.265 1046.935 12002.545 1184.3 ;
      RECT 12001.705 1048.035 12001.985 1184.06 ;
      RECT 12001.145 1048.035 12001.425 1183.82 ;
      RECT 12000.585 1048.035 12000.865 1183.58 ;
      RECT 12000.025 1048.035 12000.305 1183.34 ;
      RECT 11999.465 1048.035 11999.745 1183.1 ;
      RECT 11998.905 1048.035 11999.185 1182.86 ;
      RECT 11998.345 1048.035 11998.625 1182.62 ;
      RECT 11997.785 1048.035 11998.065 1182.38 ;
      RECT 11997.225 1048.035 11997.505 1182.14 ;
      RECT 11996.665 1048.035 11996.945 1181.9 ;
      RECT 11996.105 1048.035 11996.385 1181.66 ;
      RECT 11995.545 1048.035 11995.825 1181.42 ;
      RECT 11994.985 1046.935 11995.265 1181.18 ;
      RECT 11994.425 1048.035 11994.705 1180.94 ;
      RECT 11993.865 1046.935 11994.145 1180.7 ;
      RECT 11954.105 1048.035 11954.385 1191.17 ;
      RECT 11953.545 1046.935 11953.825 1191.41 ;
      RECT 11952.985 1048.035 11953.265 1191.65 ;
      RECT 11952.425 1048.035 11952.705 1191.89 ;
      RECT 11951.865 1048.035 11952.145 1192.13 ;
      RECT 11951.305 1048.035 11951.585 1192.37 ;
      RECT 11950.745 1048.035 11951.025 1192.61 ;
      RECT 11950.185 1048.035 11950.465 1192.855 ;
      RECT 11949.625 1048.035 11949.905 1193.095 ;
      RECT 11949.065 1048.035 11949.345 1193.335 ;
      RECT 11948.505 1046.935 11948.785 1193.575 ;
      RECT 11947.945 1048.035 11948.225 1193.815 ;
      RECT 11947.385 1046.935 11947.665 1194.055 ;
      RECT 11946.825 1048.035 11947.105 1194.295 ;
      RECT 11946.265 1048.035 11946.545 1194.535 ;
      RECT 11945.705 1048.035 11945.985 1194.775 ;
      RECT 11945.145 1048.035 11945.425 1195.015 ;
      RECT 11944.585 1048.035 11944.865 1195.255 ;
      RECT 11944.025 1048.035 11944.305 1195.495 ;
      RECT 11943.465 1048.035 11943.745 1195.735 ;
      RECT 11942.905 1048.035 11943.185 1195.975 ;
      RECT 11942.345 1048.035 11942.625 1196.215 ;
      RECT 11941.785 1048.035 11942.065 1196.455 ;
      RECT 11941.225 1048.035 11941.505 1196.695 ;
      RECT 11932.265 1048.035 11932.545 1192.28 ;
      RECT 11931.705 1048.035 11931.985 1192.04 ;
      RECT 11931.145 1048.035 11931.425 1191.8 ;
      RECT 11930.585 1046.935 11930.865 1191.56 ;
      RECT 11930.025 1048.035 11930.305 1191.32 ;
      RECT 11929.465 1046.935 11929.745 1191.08 ;
      RECT 11928.905 1048.035 11929.185 1190.84 ;
      RECT 11928.345 1048.035 11928.625 1190.6 ;
      RECT 11927.785 1048.035 11928.065 1190.36 ;
      RECT 11927.225 1046.935 11927.505 1190.12 ;
      RECT 11926.665 1048.035 11926.945 1189.88 ;
      RECT 11926.105 1046.935 11926.385 1189.64 ;
      RECT 11925.545 1048.035 11925.825 1189.4 ;
      RECT 11924.985 1046.935 11925.265 1189.16 ;
      RECT 11922.465 1048.035 11922.745 1181.56 ;
      RECT 11921.905 1048.035 11922.185 1181.32 ;
      RECT 11921.345 1048.035 11921.625 1181.08 ;
      RECT 11920.785 1048.035 11921.065 1180.84 ;
      RECT 11920.225 1048.035 11920.505 1180.6 ;
      RECT 11919.665 1048.035 11919.945 1180.36 ;
      RECT 11919.105 1048.035 11919.385 1180.12 ;
      RECT 11893.065 1048.035 11893.345 1193.995 ;
      RECT 11892.505 1048.035 11892.785 1194.235 ;
      RECT 11891.945 1048.035 11892.225 1194.475 ;
      RECT 11891.385 1048.035 11891.665 1194.715 ;
      RECT 11890.825 1048.035 11891.105 1194.955 ;
      RECT 11890.265 1046.935 11890.545 1194.955 ;
      RECT 11889.705 1048.035 11889.985 1194.715 ;
      RECT 11889.145 1046.935 11889.425 1194.47 ;
      RECT 11888.585 1048.035 11888.865 1194.23 ;
      RECT 11888.025 1046.935 11888.305 1193.99 ;
      RECT 11887.465 1048.035 11887.745 1193.75 ;
      RECT 11886.905 1048.035 11887.185 1193.51 ;
      RECT 11886.345 1048.035 11886.625 1193.27 ;
      RECT 11885.785 1048.035 11886.065 1193.03 ;
      RECT 11885.225 1048.035 11885.505 1192.79 ;
      RECT 11884.665 1048.035 11884.945 1192.55 ;
      RECT 11884.105 1048.035 11884.385 1192.31 ;
      RECT 11883.545 1048.035 11883.825 1192.07 ;
      RECT 11882.985 1046.935 11883.265 1191.83 ;
      RECT 11882.425 1048.035 11882.705 1191.59 ;
      RECT 11881.865 1046.935 11882.145 1191.35 ;
      RECT 11881.305 1048.035 11881.585 1191.11 ;
      RECT 11880.745 1048.035 11881.025 1190.87 ;
      RECT 11880.185 1048.035 11880.465 1190.63 ;
      RECT 11866.745 1048.035 11867.025 1194.03 ;
      RECT 11866.185 1048.035 11866.465 1194.27 ;
      RECT 11865.625 1048.035 11865.905 1194.515 ;
      RECT 11865.065 1048.035 11865.345 1194.755 ;
      RECT 11864.505 1048.035 11864.785 1194.995 ;
      RECT 11863.945 1048.035 11864.225 1194.995 ;
      RECT 11863.385 1048.035 11863.665 1194.755 ;
      RECT 11862.825 1048.035 11863.105 1194.515 ;
      RECT 11862.265 1048.035 11862.545 1187.5 ;
      RECT 11861.705 1048.035 11861.985 1187.26 ;
      RECT 11861.145 1048.035 11861.425 1187.02 ;
      RECT 11860.585 1046.935 11860.865 1186.78 ;
      RECT 11860.025 1048.035 11860.305 1186.54 ;
      RECT 11859.465 1046.935 11859.745 1186.3 ;
      RECT 11858.905 1048.035 11859.185 1186.06 ;
      RECT 11858.345 1048.035 11858.625 1185.82 ;
      RECT 11857.785 1048.035 11858.065 1185.58 ;
      RECT 11857.225 1046.935 11857.505 1185.34 ;
      RECT 11856.665 1048.035 11856.945 1185.1 ;
      RECT 11856.105 1046.935 11856.385 1184.86 ;
      RECT 11855.545 1048.035 11855.825 1184.62 ;
      RECT 11854.985 1046.935 11855.265 1184.38 ;
      RECT 11854.425 1048.035 11854.705 1184.14 ;
      RECT 11853.865 1048.035 11854.145 1183.9 ;
      RECT 11813.545 1048.035 11813.825 1192.795 ;
      RECT 11812.985 1048.035 11813.265 1193.035 ;
      RECT 11812.425 1048.035 11812.705 1193.28 ;
      RECT 11811.865 1048.035 11812.145 1193.52 ;
      RECT 11811.305 1048.035 11811.585 1193.76 ;
      RECT 11810.745 1048.035 11811.025 1194 ;
      RECT 11810.185 1048.035 11810.465 1194.24 ;
      RECT 11809.625 1048.035 11809.905 1194.48 ;
      RECT 11809.065 1048.035 11809.345 1194.72 ;
      RECT 11808.505 1048.035 11808.785 1194.96 ;
      RECT 11807.945 1046.935 11808.225 1195.2 ;
      RECT 11807.385 1048.035 11807.665 1195.44 ;
      RECT 11806.825 1046.935 11807.105 1195.68 ;
      RECT 11806.265 1048.035 11806.545 1195.92 ;
      RECT 11805.705 1046.935 11805.985 1196.16 ;
      RECT 11805.145 1048.035 11805.425 1196.16 ;
      RECT 11804.585 1048.035 11804.865 1195.92 ;
      RECT 11804.025 1048.035 11804.305 1195.68 ;
      RECT 11803.465 1048.035 11803.745 1195.44 ;
      RECT 11802.905 1048.035 11803.185 1195.2 ;
      RECT 11802.345 1048.035 11802.625 1194.96 ;
      RECT 11801.785 1048.035 11802.065 1194.72 ;
      RECT 11801.225 1048.035 11801.505 1194.48 ;
      RECT 11792.265 1046.935 11792.545 1194.51 ;
      RECT 11791.705 1048.035 11791.985 1194.75 ;
      RECT 11791.145 1046.935 11791.425 1194.99 ;
      RECT 11790.585 1048.035 11790.865 1195.205 ;
      RECT 11790.025 1048.035 11790.305 1194.78 ;
      RECT 11789.465 1048.035 11789.745 1194.54 ;
      RECT 11788.905 1048.035 11789.185 1194.3 ;
      RECT 11788.345 1048.035 11788.625 1194.06 ;
      RECT 11787.785 1048.035 11788.065 1193.82 ;
      RECT 11787.225 1048.035 11787.505 1193.58 ;
      RECT 11786.665 1048.035 11786.945 1193.34 ;
      RECT 11786.105 1048.035 11786.385 1193.1 ;
      RECT 11785.545 1048.035 11785.825 1192.86 ;
      RECT 11784.985 1048.035 11785.265 1192.62 ;
      RECT 11782.465 1048.035 11782.745 1191.795 ;
      RECT 11781.905 1048.035 11782.185 1191.555 ;
      RECT 11781.345 1048.035 11781.625 1191.315 ;
      RECT 11780.785 1046.935 11781.065 1191.075 ;
      RECT 11780.225 1048.035 11780.505 1190.835 ;
      RECT 11779.665 1046.935 11779.945 1190.595 ;
      RECT 11779.105 1048.035 11779.385 1190.355 ;
      RECT 11778.545 1048.035 11778.825 1190.115 ;
      RECT 11751.945 1048.035 11752.225 1201.16 ;
      RECT 11751.385 1046.935 11751.665 1201.4 ;
      RECT 11750.825 1048.035 11751.105 1201.64 ;
      RECT 11750.265 1046.935 11750.545 1201.885 ;
      RECT 11749.705 1048.035 11749.985 1202.125 ;
      RECT 11749.145 1046.935 11749.425 1202.365 ;
      RECT 11748.585 1048.035 11748.865 1202.605 ;
      RECT 11748.025 1048.035 11748.305 1202.845 ;
      RECT 11747.465 1048.035 11747.745 1188.465 ;
      RECT 11746.905 1048.035 11747.185 1188.225 ;
      RECT 11746.345 1048.035 11746.625 1187.985 ;
      RECT 11745.785 1048.035 11746.065 1187.745 ;
      RECT 11745.225 1048.035 11745.505 1187.505 ;
      RECT 11744.665 1048.035 11744.945 1187.265 ;
      RECT 11744.105 1048.035 11744.385 1187.025 ;
      RECT 11743.545 1048.035 11743.825 1186.785 ;
      RECT 11742.985 1048.035 11743.265 1186.545 ;
      RECT 11742.425 1048.035 11742.705 1186.305 ;
      RECT 11741.865 1046.935 11742.145 1186.065 ;
      RECT 11741.305 1048.035 11741.585 1185.825 ;
      RECT 11740.745 1046.935 11741.025 1185.585 ;
      RECT 11740.185 1048.035 11740.465 1185.345 ;
      RECT 11726.185 1046.935 11726.465 1191.465 ;
      RECT 11725.625 1048.035 11725.905 1191.225 ;
      RECT 11725.065 1048.035 11725.345 1190.985 ;
      RECT 11724.505 1048.035 11724.785 1190.745 ;
      RECT 11723.945 1048.035 11724.225 1190.505 ;
      RECT 11723.385 1048.035 11723.665 1190.265 ;
      RECT 11722.825 1048.035 11723.105 1190.025 ;
      RECT 11722.265 1048.035 11722.545 1189.785 ;
      RECT 11721.705 1048.035 11721.985 1189.545 ;
      RECT 11721.145 1046.935 11721.425 1189.305 ;
      RECT 11720.585 1048.035 11720.865 1189.065 ;
      RECT 11720.025 1046.935 11720.305 1188.825 ;
      RECT 11719.465 1048.035 11719.745 1188.585 ;
      RECT 11718.905 1048.035 11719.185 1188.345 ;
      RECT 11718.345 1048.035 11718.625 1188.105 ;
      RECT 11717.785 1048.035 11718.065 1187.865 ;
      RECT 11717.225 1048.035 11717.505 1187.625 ;
      RECT 11716.665 1048.035 11716.945 1187.385 ;
      RECT 11716.105 1048.035 11716.385 1187.145 ;
      RECT 11715.545 1048.035 11715.825 1186.905 ;
      RECT 11714.985 1048.035 11715.265 1186.665 ;
      RECT 11714.425 1048.035 11714.705 1186.425 ;
      RECT 11713.865 1048.035 11714.145 1186.185 ;
      RECT 11674.665 1048.035 11674.945 1193.09 ;
      RECT 11674.105 1048.035 11674.385 1193.33 ;
      RECT 11673.545 1048.035 11673.825 1193.57 ;
      RECT 11672.985 1046.935 11673.265 1193.81 ;
      RECT 11672.425 1048.035 11672.705 1194.05 ;
      RECT 11671.865 1046.935 11672.145 1194.29 ;
      RECT 11671.305 1048.035 11671.585 1194.53 ;
      RECT 11670.745 1048.035 11671.025 1194.77 ;
      RECT 11670.185 1048.035 11670.465 1195.01 ;
      RECT 11669.625 1046.935 11669.905 1195.25 ;
      RECT 11669.065 1048.035 11669.345 1195.49 ;
      RECT 11668.505 1046.935 11668.785 1195.73 ;
      RECT 11667.945 1048.035 11668.225 1195.97 ;
      RECT 11667.385 1046.935 11667.665 1196.21 ;
      RECT 11666.825 1048.035 11667.105 1196.45 ;
      RECT 11666.265 1048.035 11666.545 1196.69 ;
      RECT 11665.705 1048.035 11665.985 1196.69 ;
      RECT 11665.145 1048.035 11665.425 1196.45 ;
      RECT 11664.585 1048.035 11664.865 1196.21 ;
      RECT 11664.025 1048.035 11664.305 1195.97 ;
      RECT 11663.465 1048.035 11663.745 1195.73 ;
      RECT 11662.905 1048.035 11663.185 1195.49 ;
      RECT 11662.345 1048.035 11662.625 1195.25 ;
      RECT 11661.785 1048.035 11662.065 1195.01 ;
      RECT 11661.225 1048.035 11661.505 1194.77 ;
      RECT 11652.265 1048.035 11652.545 1194.285 ;
      RECT 11651.705 1046.935 11651.985 1194.045 ;
      RECT 11651.145 1048.035 11651.425 1193.805 ;
      RECT 11650.585 1046.935 11650.865 1193.565 ;
      RECT 11650.025 1048.035 11650.305 1193.325 ;
      RECT 11649.465 1046.935 11649.745 1193.085 ;
      RECT 11648.905 1048.035 11649.185 1192.845 ;
      RECT 11648.345 1048.035 11648.625 1192.605 ;
      RECT 11647.785 1048.035 11648.065 1192.365 ;
      RECT 11647.225 1048.035 11647.505 1192.125 ;
      RECT 11646.665 1048.035 11646.945 1191.885 ;
      RECT 11646.105 1048.035 11646.385 1191.645 ;
      RECT 11645.545 1048.035 11645.825 1191.405 ;
      RECT 11644.985 1048.035 11645.265 1191.165 ;
      RECT 11642.465 1046.935 11642.745 1192.885 ;
      RECT 11641.905 1048.035 11642.185 1192.645 ;
      RECT 11641.345 1046.935 11641.625 1192.405 ;
      RECT 11640.785 1048.035 11641.065 1192.165 ;
      RECT 11640.225 1048.035 11640.505 1191.925 ;
      RECT 11639.665 1048.035 11639.945 1191.685 ;
      RECT 11639.105 1048.035 11639.385 1191.445 ;
      RECT 11638.545 1048.035 11638.825 1191.205 ;
      RECT 11612.505 1048.035 11612.785 1188.855 ;
      RECT 11611.945 1048.035 11612.225 1189.095 ;
      RECT 11611.385 1048.035 11611.665 1189.335 ;
      RECT 11610.825 1048.035 11611.105 1189.58 ;
      RECT 11610.265 1048.035 11610.545 1189.82 ;
      RECT 11609.705 1048.035 11609.985 1190.06 ;
      RECT 11609.145 1048.035 11609.425 1190.06 ;
      RECT 11608.585 1048.035 11608.865 1189.82 ;
      RECT 11608.025 1048.035 11608.305 1189.58 ;
      RECT 11607.465 1046.935 11607.745 1189.34 ;
      RECT 11606.905 1048.035 11607.185 1189.1 ;
      RECT 11606.345 1046.935 11606.625 1188.86 ;
      RECT 11605.785 1048.035 11606.065 1188.62 ;
      RECT 11605.225 1048.035 11605.505 1188.38 ;
      RECT 11604.665 1048.035 11604.945 1188.14 ;
      RECT 11604.105 1046.935 11604.385 1187.9 ;
      RECT 11603.545 1048.035 11603.825 1187.66 ;
      RECT 11602.985 1046.935 11603.265 1187.42 ;
      RECT 11602.425 1048.035 11602.705 1187.18 ;
      RECT 11601.865 1046.935 11602.145 1186.94 ;
      RECT 11601.305 1048.035 11601.585 1186.7 ;
      RECT 11600.745 1048.035 11601.025 1186.46 ;
      RECT 11600.185 1048.035 11600.465 1186.22 ;
      RECT 11599.625 1048.035 11599.905 1185.98 ;
      RECT 11586.185 1048.035 11586.465 1191.78 ;
      RECT 11585.625 1048.035 11585.905 1191.54 ;
      RECT 11585.065 1048.035 11585.345 1191.3 ;
      RECT 11584.505 1048.035 11584.785 1191.06 ;
      RECT 11583.945 1048.035 11584.225 1190.82 ;
      RECT 11583.385 1048.035 11583.665 1190.58 ;
      RECT 11582.825 1048.035 11583.105 1190.34 ;
      RECT 11582.265 1048.035 11582.545 1190.1 ;
      RECT 11581.705 1046.935 11581.985 1189.86 ;
      RECT 11581.145 1048.035 11581.425 1189.62 ;
      RECT 11580.585 1046.935 11580.865 1189.3 ;
      RECT 11580.025 1048.035 11580.305 1189.14 ;
      RECT 11579.465 1046.935 11579.745 1188.9 ;
      RECT 11578.905 1048.035 11579.185 1188.66 ;
      RECT 11578.345 1048.035 11578.625 1188.42 ;
      RECT 11577.785 1048.035 11578.065 1188.18 ;
      RECT 11577.225 1048.035 11577.505 1187.94 ;
      RECT 11576.665 1048.035 11576.945 1187.7 ;
      RECT 11576.105 1048.035 11576.385 1187.46 ;
      RECT 11575.545 1048.035 11575.825 1187.22 ;
      RECT 11574.985 1048.035 11575.265 1186.98 ;
      RECT 11574.425 1046.935 11574.705 1186.74 ;
      RECT 11573.865 1048.035 11574.145 1186.5 ;
      RECT 11573.305 1046.935 11573.585 1186.26 ;
      RECT 11534.105 1048.035 11534.385 1191.87 ;
      RECT 11533.545 1048.035 11533.825 1192.11 ;
      RECT 11532.985 1048.035 11533.265 1192.35 ;
      RECT 11532.425 1048.035 11532.705 1192.59 ;
      RECT 11531.865 1048.035 11532.145 1192.83 ;
      RECT 11531.305 1048.035 11531.585 1193.07 ;
      RECT 11530.745 1048.035 11531.025 1193.31 ;
      RECT 11530.185 1048.035 11530.465 1193.55 ;
      RECT 11529.625 1048.035 11529.905 1193.79 ;
      RECT 11529.065 1048.035 11529.345 1194.03 ;
      RECT 11528.505 1048.035 11528.785 1194.27 ;
      RECT 11527.945 1048.035 11528.225 1194.51 ;
      RECT 11527.385 1048.035 11527.665 1194.75 ;
      RECT 11526.825 1048.035 11527.105 1194.75 ;
      RECT 11526.265 1046.935 11526.545 1194.51 ;
      RECT 11525.705 1048.035 11525.985 1194.27 ;
      RECT 11525.145 1046.935 11525.425 1194.03 ;
      RECT 11524.585 1048.035 11524.865 1193.79 ;
      RECT 11524.025 1048.035 11524.305 1193.55 ;
      RECT 11523.465 1048.035 11523.745 1193.31 ;
      RECT 11522.905 1046.935 11523.185 1193.045 ;
      RECT 11522.345 1048.035 11522.625 1192.805 ;
      RECT 11521.785 1046.935 11522.065 1192.565 ;
      RECT 11521.225 1048.035 11521.505 1192.325 ;
      RECT 11512.265 1046.935 11512.545 1186.16 ;
      RECT 11511.705 1048.035 11511.985 1186.4 ;
      RECT 11511.145 1048.035 11511.425 1186.64 ;
      RECT 11510.585 1048.035 11510.865 1186.64 ;
      RECT 11510.025 1048.035 11510.305 1186.4 ;
      RECT 11509.465 1048.035 11509.745 1186.16 ;
      RECT 11508.905 1048.035 11509.185 1185.92 ;
      RECT 11508.345 1048.035 11508.625 1185.68 ;
      RECT 11507.785 1048.035 11508.065 1185.44 ;
      RECT 11507.225 1048.035 11507.505 1185.2 ;
      RECT 11506.665 1048.035 11506.945 1184.96 ;
      RECT 11506.105 1048.035 11506.385 1184.72 ;
      RECT 11505.545 1048.035 11505.825 1184.48 ;
      RECT 11504.985 1046.935 11505.265 1184.24 ;
      RECT 11502.465 1048.035 11502.745 1185.96 ;
      RECT 11501.905 1046.935 11502.185 1185.72 ;
      RECT 11501.345 1048.035 11501.625 1185.48 ;
      RECT 11500.785 1046.935 11501.065 1185.24 ;
      RECT 11500.225 1048.035 11500.505 1185 ;
      RECT 11499.665 1048.035 11499.945 1184.76 ;
      RECT 11499.105 1048.035 11499.385 1184.52 ;
      RECT 11473.065 1048.035 11473.345 1187.305 ;
      RECT 11472.505 1048.035 11472.785 1187.545 ;
      RECT 11471.945 1048.035 11472.225 1187.785 ;
      RECT 11471.385 1048.035 11471.665 1188.025 ;
      RECT 11470.825 1048.035 11471.105 1188.265 ;
      RECT 11470.265 1046.935 11470.545 1188.505 ;
      RECT 11469.705 1048.035 11469.985 1188.745 ;
      RECT 11469.145 1046.935 11469.425 1188.985 ;
      RECT 11468.585 1048.035 11468.865 1189.225 ;
      RECT 11468.025 1048.035 11468.305 1189.465 ;
      RECT 11467.465 1048.035 11467.745 1189.705 ;
      RECT 11466.905 1048.035 11467.185 1189.945 ;
      RECT 11466.345 1048.035 11466.625 1190.185 ;
      RECT 11465.785 1048.035 11466.065 1190.425 ;
      RECT 11465.225 1048.035 11465.505 1190.665 ;
      RECT 11464.665 1048.035 11464.945 1190.665 ;
      RECT 11464.105 1048.035 11464.385 1190.425 ;
      RECT 11463.545 1048.035 11463.825 1190.185 ;
      RECT 11462.985 1048.035 11463.265 1189.945 ;
      RECT 11462.425 1048.035 11462.705 1189.7 ;
      RECT 11461.865 1048.035 11462.145 1189.46 ;
      RECT 11461.305 1048.035 11461.585 1189.22 ;
      RECT 11460.745 1046.935 11461.025 1188.98 ;
      RECT 11460.185 1048.035 11460.465 1188.74 ;
      RECT 11446.745 1046.935 11447.025 1186.22 ;
      RECT 11446.185 1048.035 11446.465 1185.98 ;
      RECT 11445.625 1048.035 11445.905 1185.74 ;
      RECT 11445.065 1048.035 11445.345 1185.5 ;
      RECT 11444.505 1046.935 11444.785 1185.26 ;
      RECT 11443.945 1048.035 11444.225 1185.02 ;
      RECT 11443.385 1046.935 11443.665 1184.78 ;
      RECT 11442.825 1048.035 11443.105 1184.54 ;
      RECT 11442.265 1046.935 11442.545 1184.3 ;
      RECT 11441.705 1048.035 11441.985 1184.06 ;
      RECT 11441.145 1048.035 11441.425 1183.82 ;
      RECT 11440.585 1048.035 11440.865 1183.58 ;
      RECT 11440.025 1048.035 11440.305 1183.34 ;
      RECT 11439.465 1048.035 11439.745 1183.1 ;
      RECT 11438.905 1048.035 11439.185 1182.86 ;
      RECT 11438.345 1048.035 11438.625 1182.62 ;
      RECT 11437.785 1048.035 11438.065 1182.38 ;
      RECT 11437.225 1048.035 11437.505 1182.14 ;
      RECT 11436.665 1048.035 11436.945 1181.9 ;
      RECT 11436.105 1048.035 11436.385 1181.66 ;
      RECT 11435.545 1048.035 11435.825 1181.42 ;
      RECT 11434.985 1046.935 11435.265 1181.18 ;
      RECT 11434.425 1048.035 11434.705 1180.94 ;
      RECT 11433.865 1046.935 11434.145 1180.7 ;
      RECT 11394.105 1048.035 11394.385 1191.17 ;
      RECT 11393.545 1046.935 11393.825 1191.41 ;
      RECT 11392.985 1048.035 11393.265 1191.65 ;
      RECT 11392.425 1048.035 11392.705 1191.89 ;
      RECT 11391.865 1048.035 11392.145 1192.13 ;
      RECT 11391.305 1048.035 11391.585 1192.37 ;
      RECT 11390.745 1048.035 11391.025 1192.61 ;
      RECT 11390.185 1048.035 11390.465 1192.855 ;
      RECT 11389.625 1048.035 11389.905 1193.095 ;
      RECT 11389.065 1048.035 11389.345 1193.335 ;
      RECT 11388.505 1046.935 11388.785 1193.575 ;
      RECT 11387.945 1048.035 11388.225 1193.815 ;
      RECT 11387.385 1046.935 11387.665 1194.055 ;
      RECT 11386.825 1048.035 11387.105 1194.295 ;
      RECT 11386.265 1048.035 11386.545 1194.535 ;
      RECT 11385.705 1048.035 11385.985 1194.775 ;
      RECT 11385.145 1048.035 11385.425 1195.015 ;
      RECT 11384.585 1048.035 11384.865 1195.255 ;
      RECT 11384.025 1048.035 11384.305 1195.495 ;
      RECT 11383.465 1048.035 11383.745 1195.735 ;
      RECT 11382.905 1048.035 11383.185 1195.975 ;
      RECT 11382.345 1048.035 11382.625 1196.215 ;
      RECT 11381.785 1048.035 11382.065 1196.455 ;
      RECT 11381.225 1048.035 11381.505 1196.695 ;
      RECT 11372.265 1048.035 11372.545 1192.28 ;
      RECT 11371.705 1048.035 11371.985 1192.04 ;
      RECT 11371.145 1048.035 11371.425 1191.8 ;
      RECT 11370.585 1046.935 11370.865 1191.56 ;
      RECT 11370.025 1048.035 11370.305 1191.32 ;
      RECT 11369.465 1046.935 11369.745 1191.08 ;
      RECT 11368.905 1048.035 11369.185 1190.84 ;
      RECT 11368.345 1048.035 11368.625 1190.6 ;
      RECT 11367.785 1048.035 11368.065 1190.36 ;
      RECT 11367.225 1046.935 11367.505 1190.12 ;
      RECT 11366.665 1048.035 11366.945 1189.88 ;
      RECT 11366.105 1046.935 11366.385 1189.64 ;
      RECT 11365.545 1048.035 11365.825 1189.4 ;
      RECT 11364.985 1046.935 11365.265 1189.16 ;
      RECT 11362.465 1048.035 11362.745 1181.56 ;
      RECT 11361.905 1048.035 11362.185 1181.32 ;
      RECT 11361.345 1048.035 11361.625 1181.08 ;
      RECT 11360.785 1048.035 11361.065 1180.84 ;
      RECT 11360.225 1048.035 11360.505 1180.6 ;
      RECT 11359.665 1048.035 11359.945 1180.36 ;
      RECT 11359.105 1048.035 11359.385 1180.12 ;
      RECT 11333.065 1048.035 11333.345 1193.995 ;
      RECT 11332.505 1048.035 11332.785 1194.235 ;
      RECT 11331.945 1048.035 11332.225 1194.475 ;
      RECT 11331.385 1048.035 11331.665 1194.715 ;
      RECT 11330.825 1048.035 11331.105 1194.955 ;
      RECT 11330.265 1046.935 11330.545 1194.955 ;
      RECT 11329.705 1048.035 11329.985 1194.715 ;
      RECT 11329.145 1046.935 11329.425 1194.47 ;
      RECT 11328.585 1048.035 11328.865 1194.23 ;
      RECT 11328.025 1046.935 11328.305 1193.99 ;
      RECT 11327.465 1048.035 11327.745 1193.75 ;
      RECT 11326.905 1048.035 11327.185 1193.51 ;
      RECT 11326.345 1048.035 11326.625 1193.27 ;
      RECT 11325.785 1048.035 11326.065 1193.03 ;
      RECT 11325.225 1048.035 11325.505 1192.79 ;
      RECT 11324.665 1048.035 11324.945 1192.55 ;
      RECT 11324.105 1048.035 11324.385 1192.31 ;
      RECT 11323.545 1048.035 11323.825 1192.07 ;
      RECT 11322.985 1046.935 11323.265 1191.83 ;
      RECT 11322.425 1048.035 11322.705 1191.59 ;
      RECT 11321.865 1046.935 11322.145 1191.35 ;
      RECT 11321.305 1048.035 11321.585 1191.11 ;
      RECT 11320.745 1048.035 11321.025 1190.87 ;
      RECT 11320.185 1048.035 11320.465 1190.63 ;
      RECT 11306.745 1048.035 11307.025 1194.03 ;
      RECT 11306.185 1048.035 11306.465 1194.27 ;
      RECT 11305.625 1048.035 11305.905 1194.515 ;
      RECT 11305.065 1048.035 11305.345 1194.755 ;
      RECT 11304.505 1048.035 11304.785 1194.995 ;
      RECT 11303.945 1048.035 11304.225 1194.995 ;
      RECT 11303.385 1048.035 11303.665 1194.755 ;
      RECT 11302.825 1048.035 11303.105 1194.515 ;
      RECT 11302.265 1048.035 11302.545 1187.5 ;
      RECT 11301.705 1048.035 11301.985 1187.26 ;
      RECT 11301.145 1048.035 11301.425 1187.02 ;
      RECT 11300.585 1046.935 11300.865 1186.78 ;
      RECT 11300.025 1048.035 11300.305 1186.54 ;
      RECT 11299.465 1046.935 11299.745 1186.3 ;
      RECT 11298.905 1048.035 11299.185 1186.06 ;
      RECT 11298.345 1048.035 11298.625 1185.82 ;
      RECT 11297.785 1048.035 11298.065 1185.58 ;
      RECT 11297.225 1046.935 11297.505 1185.34 ;
      RECT 11296.665 1048.035 11296.945 1185.1 ;
      RECT 11296.105 1046.935 11296.385 1184.86 ;
      RECT 11295.545 1048.035 11295.825 1184.62 ;
      RECT 11294.985 1046.935 11295.265 1184.38 ;
      RECT 11294.425 1048.035 11294.705 1184.14 ;
      RECT 11293.865 1048.035 11294.145 1183.9 ;
      RECT 11253.545 1048.035 11253.825 1192.795 ;
      RECT 11252.985 1048.035 11253.265 1193.035 ;
      RECT 11252.425 1048.035 11252.705 1193.28 ;
      RECT 11251.865 1048.035 11252.145 1193.52 ;
      RECT 11251.305 1048.035 11251.585 1193.76 ;
      RECT 11250.745 1048.035 11251.025 1194 ;
      RECT 11250.185 1048.035 11250.465 1194.24 ;
      RECT 11249.625 1048.035 11249.905 1194.48 ;
      RECT 11249.065 1048.035 11249.345 1194.72 ;
      RECT 11248.505 1048.035 11248.785 1194.96 ;
      RECT 11247.945 1046.935 11248.225 1195.2 ;
      RECT 11247.385 1048.035 11247.665 1195.44 ;
      RECT 11246.825 1046.935 11247.105 1195.68 ;
      RECT 11246.265 1048.035 11246.545 1195.92 ;
      RECT 11245.705 1046.935 11245.985 1196.16 ;
      RECT 11245.145 1048.035 11245.425 1196.16 ;
      RECT 11244.585 1048.035 11244.865 1195.92 ;
      RECT 11244.025 1048.035 11244.305 1195.68 ;
      RECT 11243.465 1048.035 11243.745 1195.44 ;
      RECT 11242.905 1048.035 11243.185 1195.2 ;
      RECT 11242.345 1048.035 11242.625 1194.96 ;
      RECT 11241.785 1048.035 11242.065 1194.72 ;
      RECT 11241.225 1048.035 11241.505 1194.48 ;
      RECT 11232.265 1046.935 11232.545 1194.51 ;
      RECT 11231.705 1048.035 11231.985 1194.75 ;
      RECT 11231.145 1046.935 11231.425 1194.99 ;
      RECT 11230.585 1048.035 11230.865 1195.205 ;
      RECT 11230.025 1048.035 11230.305 1194.78 ;
      RECT 11229.465 1048.035 11229.745 1194.54 ;
      RECT 11228.905 1048.035 11229.185 1194.3 ;
      RECT 11228.345 1048.035 11228.625 1194.06 ;
      RECT 11227.785 1048.035 11228.065 1193.82 ;
      RECT 11227.225 1048.035 11227.505 1193.58 ;
      RECT 11226.665 1048.035 11226.945 1193.34 ;
      RECT 11226.105 1048.035 11226.385 1193.1 ;
      RECT 11225.545 1048.035 11225.825 1192.86 ;
      RECT 11224.985 1048.035 11225.265 1192.62 ;
      RECT 11222.465 1048.035 11222.745 1191.795 ;
      RECT 11221.905 1048.035 11222.185 1191.555 ;
      RECT 11221.345 1048.035 11221.625 1191.315 ;
      RECT 11220.785 1046.935 11221.065 1191.075 ;
      RECT 11220.225 1048.035 11220.505 1190.835 ;
      RECT 11219.665 1046.935 11219.945 1190.595 ;
      RECT 11219.105 1048.035 11219.385 1190.355 ;
      RECT 11218.545 1048.035 11218.825 1190.115 ;
      RECT 11191.945 1048.035 11192.225 1201.16 ;
      RECT 11191.385 1046.935 11191.665 1201.4 ;
      RECT 11190.825 1048.035 11191.105 1201.64 ;
      RECT 11190.265 1046.935 11190.545 1201.885 ;
      RECT 11189.705 1048.035 11189.985 1202.125 ;
      RECT 11189.145 1046.935 11189.425 1202.365 ;
      RECT 11188.585 1048.035 11188.865 1202.605 ;
      RECT 11188.025 1048.035 11188.305 1202.845 ;
      RECT 11187.465 1048.035 11187.745 1188.465 ;
      RECT 11186.905 1048.035 11187.185 1188.225 ;
      RECT 11186.345 1048.035 11186.625 1187.985 ;
      RECT 11185.785 1048.035 11186.065 1187.745 ;
      RECT 11185.225 1048.035 11185.505 1187.505 ;
      RECT 11184.665 1048.035 11184.945 1187.265 ;
      RECT 11184.105 1048.035 11184.385 1187.025 ;
      RECT 11183.545 1048.035 11183.825 1186.785 ;
      RECT 11182.985 1048.035 11183.265 1186.545 ;
      RECT 11182.425 1048.035 11182.705 1186.305 ;
      RECT 11181.865 1046.935 11182.145 1186.065 ;
      RECT 11181.305 1048.035 11181.585 1185.825 ;
      RECT 11180.745 1046.935 11181.025 1185.585 ;
      RECT 11180.185 1048.035 11180.465 1185.345 ;
      RECT 11166.185 1046.935 11166.465 1191.465 ;
      RECT 11165.625 1048.035 11165.905 1191.225 ;
      RECT 11165.065 1048.035 11165.345 1190.985 ;
      RECT 11164.505 1048.035 11164.785 1190.745 ;
      RECT 11163.945 1048.035 11164.225 1190.505 ;
      RECT 11163.385 1048.035 11163.665 1190.265 ;
      RECT 11162.825 1048.035 11163.105 1190.025 ;
      RECT 11162.265 1048.035 11162.545 1189.785 ;
      RECT 11161.705 1048.035 11161.985 1189.545 ;
      RECT 11161.145 1046.935 11161.425 1189.305 ;
      RECT 11160.585 1048.035 11160.865 1189.065 ;
      RECT 11160.025 1046.935 11160.305 1188.825 ;
      RECT 11159.465 1048.035 11159.745 1188.585 ;
      RECT 11158.905 1048.035 11159.185 1188.345 ;
      RECT 11158.345 1048.035 11158.625 1188.105 ;
      RECT 11157.785 1048.035 11158.065 1187.865 ;
      RECT 11157.225 1048.035 11157.505 1187.625 ;
      RECT 11156.665 1048.035 11156.945 1187.385 ;
      RECT 11156.105 1048.035 11156.385 1187.145 ;
      RECT 11155.545 1048.035 11155.825 1186.905 ;
      RECT 11154.985 1048.035 11155.265 1186.665 ;
      RECT 11154.425 1048.035 11154.705 1186.425 ;
      RECT 11153.865 1048.035 11154.145 1186.185 ;
      RECT 11114.665 1048.035 11114.945 1193.09 ;
      RECT 11114.105 1048.035 11114.385 1193.33 ;
      RECT 11113.545 1048.035 11113.825 1193.57 ;
      RECT 11112.985 1046.935 11113.265 1193.81 ;
      RECT 11112.425 1048.035 11112.705 1194.05 ;
      RECT 11111.865 1046.935 11112.145 1194.29 ;
      RECT 11111.305 1048.035 11111.585 1194.53 ;
      RECT 11110.745 1048.035 11111.025 1194.77 ;
      RECT 11110.185 1048.035 11110.465 1195.01 ;
      RECT 11109.625 1046.935 11109.905 1195.25 ;
      RECT 11109.065 1048.035 11109.345 1195.49 ;
      RECT 11108.505 1046.935 11108.785 1195.73 ;
      RECT 11107.945 1048.035 11108.225 1195.97 ;
      RECT 11107.385 1046.935 11107.665 1196.21 ;
      RECT 11106.825 1048.035 11107.105 1196.45 ;
      RECT 11106.265 1048.035 11106.545 1196.69 ;
      RECT 11105.705 1048.035 11105.985 1196.69 ;
      RECT 11105.145 1048.035 11105.425 1196.45 ;
      RECT 11104.585 1048.035 11104.865 1196.21 ;
      RECT 11104.025 1048.035 11104.305 1195.97 ;
      RECT 11103.465 1048.035 11103.745 1195.73 ;
      RECT 11102.905 1048.035 11103.185 1195.49 ;
      RECT 11102.345 1048.035 11102.625 1195.25 ;
      RECT 11101.785 1048.035 11102.065 1195.01 ;
      RECT 11101.225 1048.035 11101.505 1194.77 ;
      RECT 11092.265 1048.035 11092.545 1194.285 ;
      RECT 11091.705 1046.935 11091.985 1194.045 ;
      RECT 11091.145 1048.035 11091.425 1193.805 ;
      RECT 11090.585 1046.935 11090.865 1193.565 ;
      RECT 11090.025 1048.035 11090.305 1193.325 ;
      RECT 11089.465 1046.935 11089.745 1193.085 ;
      RECT 11088.905 1048.035 11089.185 1192.845 ;
      RECT 11088.345 1048.035 11088.625 1192.605 ;
      RECT 11087.785 1048.035 11088.065 1192.365 ;
      RECT 11087.225 1048.035 11087.505 1192.125 ;
      RECT 11086.665 1048.035 11086.945 1191.885 ;
      RECT 11086.105 1048.035 11086.385 1191.645 ;
      RECT 11085.545 1048.035 11085.825 1191.405 ;
      RECT 11084.985 1048.035 11085.265 1191.165 ;
      RECT 11082.465 1046.935 11082.745 1192.885 ;
      RECT 11081.905 1048.035 11082.185 1192.645 ;
      RECT 11081.345 1046.935 11081.625 1192.405 ;
      RECT 11080.785 1048.035 11081.065 1192.165 ;
      RECT 11080.225 1048.035 11080.505 1191.925 ;
      RECT 11079.665 1048.035 11079.945 1191.685 ;
      RECT 11079.105 1048.035 11079.385 1191.445 ;
      RECT 11078.545 1048.035 11078.825 1191.205 ;
      RECT 11052.505 1048.035 11052.785 1188.855 ;
      RECT 11051.945 1048.035 11052.225 1189.095 ;
      RECT 11051.385 1048.035 11051.665 1189.335 ;
      RECT 11050.825 1048.035 11051.105 1189.58 ;
      RECT 11050.265 1048.035 11050.545 1189.82 ;
      RECT 11049.705 1048.035 11049.985 1190.06 ;
      RECT 11049.145 1048.035 11049.425 1190.06 ;
      RECT 11048.585 1048.035 11048.865 1189.82 ;
      RECT 11048.025 1048.035 11048.305 1189.58 ;
      RECT 11047.465 1046.935 11047.745 1189.34 ;
      RECT 11046.905 1048.035 11047.185 1189.1 ;
      RECT 11046.345 1046.935 11046.625 1188.86 ;
      RECT 11045.785 1048.035 11046.065 1188.62 ;
      RECT 11045.225 1048.035 11045.505 1188.38 ;
      RECT 11044.665 1048.035 11044.945 1188.14 ;
      RECT 11044.105 1046.935 11044.385 1187.9 ;
      RECT 11043.545 1048.035 11043.825 1187.66 ;
      RECT 11042.985 1046.935 11043.265 1187.42 ;
      RECT 11042.425 1048.035 11042.705 1187.18 ;
      RECT 11041.865 1046.935 11042.145 1186.94 ;
      RECT 11041.305 1048.035 11041.585 1186.7 ;
      RECT 11040.745 1048.035 11041.025 1186.46 ;
      RECT 11040.185 1048.035 11040.465 1186.22 ;
      RECT 11039.625 1048.035 11039.905 1185.98 ;
      RECT 11026.185 1048.035 11026.465 1191.78 ;
      RECT 11025.625 1048.035 11025.905 1191.54 ;
      RECT 11025.065 1048.035 11025.345 1191.3 ;
      RECT 11024.505 1048.035 11024.785 1191.06 ;
      RECT 11023.945 1048.035 11024.225 1190.82 ;
      RECT 11023.385 1048.035 11023.665 1190.58 ;
      RECT 11022.825 1048.035 11023.105 1190.34 ;
      RECT 11022.265 1048.035 11022.545 1190.1 ;
      RECT 11021.705 1046.935 11021.985 1189.86 ;
      RECT 11021.145 1048.035 11021.425 1189.62 ;
      RECT 11020.585 1046.935 11020.865 1189.3 ;
      RECT 11020.025 1048.035 11020.305 1189.14 ;
      RECT 11019.465 1046.935 11019.745 1188.9 ;
      RECT 11018.905 1048.035 11019.185 1188.66 ;
      RECT 11018.345 1048.035 11018.625 1188.42 ;
      RECT 11017.785 1048.035 11018.065 1188.18 ;
      RECT 11017.225 1048.035 11017.505 1187.94 ;
      RECT 11016.665 1048.035 11016.945 1187.7 ;
      RECT 11016.105 1048.035 11016.385 1187.46 ;
      RECT 11015.545 1048.035 11015.825 1187.22 ;
      RECT 11014.985 1048.035 11015.265 1186.98 ;
      RECT 11014.425 1046.935 11014.705 1186.74 ;
      RECT 11013.865 1048.035 11014.145 1186.5 ;
      RECT 11013.305 1046.935 11013.585 1186.26 ;
      RECT 10974.105 1048.035 10974.385 1191.87 ;
      RECT 10973.545 1048.035 10973.825 1192.11 ;
      RECT 10972.985 1048.035 10973.265 1192.35 ;
      RECT 10972.425 1048.035 10972.705 1192.59 ;
      RECT 10971.865 1048.035 10972.145 1192.83 ;
      RECT 10971.305 1048.035 10971.585 1193.07 ;
      RECT 10970.745 1048.035 10971.025 1193.31 ;
      RECT 10970.185 1048.035 10970.465 1193.55 ;
      RECT 10969.625 1048.035 10969.905 1193.79 ;
      RECT 10969.065 1048.035 10969.345 1194.03 ;
      RECT 10968.505 1048.035 10968.785 1194.27 ;
      RECT 10967.945 1048.035 10968.225 1194.51 ;
      RECT 10967.385 1048.035 10967.665 1194.75 ;
      RECT 10966.825 1048.035 10967.105 1194.75 ;
      RECT 10966.265 1046.935 10966.545 1194.51 ;
      RECT 10965.705 1048.035 10965.985 1194.27 ;
      RECT 10965.145 1046.935 10965.425 1194.03 ;
      RECT 10964.585 1048.035 10964.865 1193.79 ;
      RECT 10964.025 1048.035 10964.305 1193.55 ;
      RECT 10963.465 1048.035 10963.745 1193.31 ;
      RECT 10962.905 1046.935 10963.185 1193.045 ;
      RECT 10962.345 1048.035 10962.625 1192.805 ;
      RECT 10961.785 1046.935 10962.065 1192.565 ;
      RECT 10961.225 1048.035 10961.505 1192.325 ;
      RECT 10952.265 1046.935 10952.545 1186.16 ;
      RECT 10951.705 1048.035 10951.985 1186.4 ;
      RECT 10951.145 1048.035 10951.425 1186.64 ;
      RECT 10950.585 1048.035 10950.865 1186.64 ;
      RECT 10950.025 1048.035 10950.305 1186.4 ;
      RECT 10949.465 1048.035 10949.745 1186.16 ;
      RECT 10948.905 1048.035 10949.185 1185.92 ;
      RECT 10948.345 1048.035 10948.625 1185.68 ;
      RECT 10947.785 1048.035 10948.065 1185.44 ;
      RECT 10947.225 1048.035 10947.505 1185.2 ;
      RECT 10946.665 1048.035 10946.945 1184.96 ;
      RECT 10946.105 1048.035 10946.385 1184.72 ;
      RECT 10945.545 1048.035 10945.825 1184.48 ;
      RECT 10944.985 1046.935 10945.265 1184.24 ;
      RECT 10942.465 1048.035 10942.745 1185.96 ;
      RECT 10941.905 1046.935 10942.185 1185.72 ;
      RECT 10941.345 1048.035 10941.625 1185.48 ;
      RECT 10940.785 1046.935 10941.065 1185.24 ;
      RECT 10940.225 1048.035 10940.505 1185 ;
      RECT 10939.665 1048.035 10939.945 1184.76 ;
      RECT 10939.105 1048.035 10939.385 1184.52 ;
      RECT 10913.065 1048.035 10913.345 1187.305 ;
      RECT 10912.505 1048.035 10912.785 1187.545 ;
      RECT 10911.945 1048.035 10912.225 1187.785 ;
      RECT 10911.385 1048.035 10911.665 1188.025 ;
      RECT 10910.825 1048.035 10911.105 1188.265 ;
      RECT 10910.265 1046.935 10910.545 1188.505 ;
      RECT 10909.705 1048.035 10909.985 1188.745 ;
      RECT 10909.145 1046.935 10909.425 1188.985 ;
      RECT 10908.585 1048.035 10908.865 1189.225 ;
      RECT 10908.025 1048.035 10908.305 1189.465 ;
      RECT 10907.465 1048.035 10907.745 1189.705 ;
      RECT 10906.905 1048.035 10907.185 1189.945 ;
      RECT 10906.345 1048.035 10906.625 1190.185 ;
      RECT 10905.785 1048.035 10906.065 1190.425 ;
      RECT 10905.225 1048.035 10905.505 1190.665 ;
      RECT 10904.665 1048.035 10904.945 1190.665 ;
      RECT 10904.105 1048.035 10904.385 1190.425 ;
      RECT 10903.545 1048.035 10903.825 1190.185 ;
      RECT 10902.985 1048.035 10903.265 1189.945 ;
      RECT 10902.425 1048.035 10902.705 1189.7 ;
      RECT 10901.865 1048.035 10902.145 1189.46 ;
      RECT 10901.305 1048.035 10901.585 1189.22 ;
      RECT 10900.745 1046.935 10901.025 1188.98 ;
      RECT 10900.185 1048.035 10900.465 1188.74 ;
      RECT 10886.745 1046.935 10887.025 1186.22 ;
      RECT 10886.185 1048.035 10886.465 1185.98 ;
      RECT 10885.625 1048.035 10885.905 1185.74 ;
      RECT 10885.065 1048.035 10885.345 1185.5 ;
      RECT 10884.505 1046.935 10884.785 1185.26 ;
      RECT 10883.945 1048.035 10884.225 1185.02 ;
      RECT 10883.385 1046.935 10883.665 1184.78 ;
      RECT 10882.825 1048.035 10883.105 1184.54 ;
      RECT 10882.265 1046.935 10882.545 1184.3 ;
      RECT 10881.705 1048.035 10881.985 1184.06 ;
      RECT 10881.145 1048.035 10881.425 1183.82 ;
      RECT 10880.585 1048.035 10880.865 1183.58 ;
      RECT 10880.025 1048.035 10880.305 1183.34 ;
      RECT 10879.465 1048.035 10879.745 1183.1 ;
      RECT 10878.905 1048.035 10879.185 1182.86 ;
      RECT 10878.345 1048.035 10878.625 1182.62 ;
      RECT 10877.785 1048.035 10878.065 1182.38 ;
      RECT 10877.225 1048.035 10877.505 1182.14 ;
      RECT 10876.665 1048.035 10876.945 1181.9 ;
      RECT 10876.105 1048.035 10876.385 1181.66 ;
      RECT 10875.545 1048.035 10875.825 1181.42 ;
      RECT 10874.985 1046.935 10875.265 1181.18 ;
      RECT 10874.425 1048.035 10874.705 1180.94 ;
      RECT 10873.865 1046.935 10874.145 1180.7 ;
      RECT 10834.105 1048.035 10834.385 1191.17 ;
      RECT 10833.545 1046.935 10833.825 1191.41 ;
      RECT 10832.985 1048.035 10833.265 1191.65 ;
      RECT 10832.425 1048.035 10832.705 1191.89 ;
      RECT 10831.865 1048.035 10832.145 1192.13 ;
      RECT 10831.305 1048.035 10831.585 1192.37 ;
      RECT 10830.745 1048.035 10831.025 1192.61 ;
      RECT 10830.185 1048.035 10830.465 1192.855 ;
      RECT 10829.625 1048.035 10829.905 1193.095 ;
      RECT 10829.065 1048.035 10829.345 1193.335 ;
      RECT 10828.505 1046.935 10828.785 1193.575 ;
      RECT 10827.945 1048.035 10828.225 1193.815 ;
      RECT 10827.385 1046.935 10827.665 1194.055 ;
      RECT 10826.825 1048.035 10827.105 1194.295 ;
      RECT 10826.265 1048.035 10826.545 1194.535 ;
      RECT 10825.705 1048.035 10825.985 1194.775 ;
      RECT 10825.145 1048.035 10825.425 1195.015 ;
      RECT 10824.585 1048.035 10824.865 1195.255 ;
      RECT 10824.025 1048.035 10824.305 1195.495 ;
      RECT 10823.465 1048.035 10823.745 1195.735 ;
      RECT 10822.905 1048.035 10823.185 1195.975 ;
      RECT 10822.345 1048.035 10822.625 1196.215 ;
      RECT 10821.785 1048.035 10822.065 1196.455 ;
      RECT 10821.225 1048.035 10821.505 1196.695 ;
      RECT 10812.265 1048.035 10812.545 1192.28 ;
      RECT 10811.705 1048.035 10811.985 1192.04 ;
      RECT 10811.145 1048.035 10811.425 1191.8 ;
      RECT 10810.585 1046.935 10810.865 1191.56 ;
      RECT 10810.025 1048.035 10810.305 1191.32 ;
      RECT 10809.465 1046.935 10809.745 1191.08 ;
      RECT 10808.905 1048.035 10809.185 1190.84 ;
      RECT 10808.345 1048.035 10808.625 1190.6 ;
      RECT 10807.785 1048.035 10808.065 1190.36 ;
      RECT 10807.225 1046.935 10807.505 1190.12 ;
      RECT 10806.665 1048.035 10806.945 1189.88 ;
      RECT 10806.105 1046.935 10806.385 1189.64 ;
      RECT 10805.545 1048.035 10805.825 1189.4 ;
      RECT 10804.985 1046.935 10805.265 1189.16 ;
      RECT 10802.465 1048.035 10802.745 1181.56 ;
      RECT 10801.905 1048.035 10802.185 1181.32 ;
      RECT 10801.345 1048.035 10801.625 1181.08 ;
      RECT 10800.785 1048.035 10801.065 1180.84 ;
      RECT 10800.225 1048.035 10800.505 1180.6 ;
      RECT 10799.665 1048.035 10799.945 1180.36 ;
      RECT 10799.105 1048.035 10799.385 1180.12 ;
      RECT 10773.065 1048.035 10773.345 1193.995 ;
      RECT 10772.505 1048.035 10772.785 1194.235 ;
      RECT 10771.945 1048.035 10772.225 1194.475 ;
      RECT 10771.385 1048.035 10771.665 1194.715 ;
      RECT 10770.825 1048.035 10771.105 1194.955 ;
      RECT 10770.265 1046.935 10770.545 1194.955 ;
      RECT 10769.705 1048.035 10769.985 1194.715 ;
      RECT 10769.145 1046.935 10769.425 1194.47 ;
      RECT 10768.585 1048.035 10768.865 1194.23 ;
      RECT 10768.025 1046.935 10768.305 1193.99 ;
      RECT 10767.465 1048.035 10767.745 1193.75 ;
      RECT 10766.905 1048.035 10767.185 1193.51 ;
      RECT 10766.345 1048.035 10766.625 1193.27 ;
      RECT 10765.785 1048.035 10766.065 1193.03 ;
      RECT 10765.225 1048.035 10765.505 1192.79 ;
      RECT 10764.665 1048.035 10764.945 1192.55 ;
      RECT 10764.105 1048.035 10764.385 1192.31 ;
      RECT 10763.545 1048.035 10763.825 1192.07 ;
      RECT 10762.985 1046.935 10763.265 1191.83 ;
      RECT 10762.425 1048.035 10762.705 1191.59 ;
      RECT 10761.865 1046.935 10762.145 1191.35 ;
      RECT 10761.305 1048.035 10761.585 1191.11 ;
      RECT 10760.745 1048.035 10761.025 1190.87 ;
      RECT 10760.185 1048.035 10760.465 1190.63 ;
      RECT 10746.745 1048.035 10747.025 1194.03 ;
      RECT 10746.185 1048.035 10746.465 1194.27 ;
      RECT 10745.625 1048.035 10745.905 1194.515 ;
      RECT 10745.065 1048.035 10745.345 1194.755 ;
      RECT 10744.505 1048.035 10744.785 1194.995 ;
      RECT 10743.945 1048.035 10744.225 1194.995 ;
      RECT 10743.385 1048.035 10743.665 1194.755 ;
      RECT 10742.825 1048.035 10743.105 1194.515 ;
      RECT 10742.265 1048.035 10742.545 1187.5 ;
      RECT 10741.705 1048.035 10741.985 1187.26 ;
      RECT 10741.145 1048.035 10741.425 1187.02 ;
      RECT 10740.585 1046.935 10740.865 1186.78 ;
      RECT 10740.025 1048.035 10740.305 1186.54 ;
      RECT 10739.465 1046.935 10739.745 1186.3 ;
      RECT 10738.905 1048.035 10739.185 1186.06 ;
      RECT 10738.345 1048.035 10738.625 1185.82 ;
      RECT 10737.785 1048.035 10738.065 1185.58 ;
      RECT 10737.225 1046.935 10737.505 1185.34 ;
      RECT 10736.665 1048.035 10736.945 1185.1 ;
      RECT 10736.105 1046.935 10736.385 1184.86 ;
      RECT 10735.545 1048.035 10735.825 1184.62 ;
      RECT 10734.985 1046.935 10735.265 1184.38 ;
      RECT 10734.425 1048.035 10734.705 1184.14 ;
      RECT 10733.865 1048.035 10734.145 1183.9 ;
      RECT 10693.545 1048.035 10693.825 1192.795 ;
      RECT 10692.985 1048.035 10693.265 1193.035 ;
      RECT 10692.425 1048.035 10692.705 1193.28 ;
      RECT 10691.865 1048.035 10692.145 1193.52 ;
      RECT 10691.305 1048.035 10691.585 1193.76 ;
      RECT 10690.745 1048.035 10691.025 1194 ;
      RECT 10690.185 1048.035 10690.465 1194.24 ;
      RECT 10689.625 1048.035 10689.905 1194.48 ;
      RECT 10689.065 1048.035 10689.345 1194.72 ;
      RECT 10688.505 1048.035 10688.785 1194.96 ;
      RECT 10687.945 1046.935 10688.225 1195.2 ;
      RECT 10687.385 1048.035 10687.665 1195.44 ;
      RECT 10686.825 1046.935 10687.105 1195.68 ;
      RECT 10686.265 1048.035 10686.545 1195.92 ;
      RECT 10685.705 1046.935 10685.985 1196.16 ;
      RECT 10685.145 1048.035 10685.425 1196.16 ;
      RECT 10684.585 1048.035 10684.865 1195.92 ;
      RECT 10684.025 1048.035 10684.305 1195.68 ;
      RECT 10683.465 1048.035 10683.745 1195.44 ;
      RECT 10682.905 1048.035 10683.185 1195.2 ;
      RECT 10682.345 1048.035 10682.625 1194.96 ;
      RECT 10681.785 1048.035 10682.065 1194.72 ;
      RECT 10681.225 1048.035 10681.505 1194.48 ;
      RECT 10672.265 1046.935 10672.545 1194.51 ;
      RECT 10671.705 1048.035 10671.985 1194.75 ;
      RECT 10671.145 1046.935 10671.425 1194.99 ;
      RECT 10670.585 1048.035 10670.865 1195.205 ;
      RECT 10670.025 1048.035 10670.305 1194.78 ;
      RECT 10669.465 1048.035 10669.745 1194.54 ;
      RECT 10668.905 1048.035 10669.185 1194.3 ;
      RECT 10668.345 1048.035 10668.625 1194.06 ;
      RECT 10667.785 1048.035 10668.065 1193.82 ;
      RECT 10667.225 1048.035 10667.505 1193.58 ;
      RECT 10666.665 1048.035 10666.945 1193.34 ;
      RECT 10666.105 1048.035 10666.385 1193.1 ;
      RECT 10665.545 1048.035 10665.825 1192.86 ;
      RECT 10664.985 1048.035 10665.265 1192.62 ;
      RECT 10662.465 1048.035 10662.745 1191.795 ;
      RECT 10661.905 1048.035 10662.185 1191.555 ;
      RECT 10661.345 1048.035 10661.625 1191.315 ;
      RECT 10660.785 1046.935 10661.065 1191.075 ;
      RECT 10660.225 1048.035 10660.505 1190.835 ;
      RECT 10659.665 1046.935 10659.945 1190.595 ;
      RECT 10659.105 1048.035 10659.385 1190.355 ;
      RECT 10658.545 1048.035 10658.825 1190.115 ;
      RECT 10631.945 1048.035 10632.225 1201.16 ;
      RECT 10631.385 1046.935 10631.665 1201.4 ;
      RECT 10630.825 1048.035 10631.105 1201.64 ;
      RECT 10630.265 1046.935 10630.545 1201.885 ;
      RECT 10629.705 1048.035 10629.985 1202.125 ;
      RECT 10629.145 1046.935 10629.425 1202.365 ;
      RECT 10628.585 1048.035 10628.865 1202.605 ;
      RECT 10628.025 1048.035 10628.305 1202.845 ;
      RECT 10627.465 1048.035 10627.745 1188.465 ;
      RECT 10626.905 1048.035 10627.185 1188.225 ;
      RECT 10626.345 1048.035 10626.625 1187.985 ;
      RECT 10625.785 1048.035 10626.065 1187.745 ;
      RECT 10625.225 1048.035 10625.505 1187.505 ;
      RECT 10624.665 1048.035 10624.945 1187.265 ;
      RECT 10624.105 1048.035 10624.385 1187.025 ;
      RECT 10623.545 1048.035 10623.825 1186.785 ;
      RECT 10622.985 1048.035 10623.265 1186.545 ;
      RECT 10622.425 1048.035 10622.705 1186.305 ;
      RECT 10621.865 1046.935 10622.145 1186.065 ;
      RECT 10621.305 1048.035 10621.585 1185.825 ;
      RECT 10620.745 1046.935 10621.025 1185.585 ;
      RECT 10620.185 1048.035 10620.465 1185.345 ;
      RECT 10606.185 1046.935 10606.465 1191.465 ;
      RECT 10605.625 1048.035 10605.905 1191.225 ;
      RECT 10605.065 1048.035 10605.345 1190.985 ;
      RECT 10604.505 1048.035 10604.785 1190.745 ;
      RECT 10603.945 1048.035 10604.225 1190.505 ;
      RECT 10603.385 1048.035 10603.665 1190.265 ;
      RECT 10602.825 1048.035 10603.105 1190.025 ;
      RECT 10602.265 1048.035 10602.545 1189.785 ;
      RECT 10601.705 1048.035 10601.985 1189.545 ;
      RECT 10601.145 1046.935 10601.425 1189.305 ;
      RECT 10600.585 1048.035 10600.865 1189.065 ;
      RECT 10600.025 1046.935 10600.305 1188.825 ;
      RECT 10599.465 1048.035 10599.745 1188.585 ;
      RECT 10598.905 1048.035 10599.185 1188.345 ;
      RECT 10598.345 1048.035 10598.625 1188.105 ;
      RECT 10597.785 1048.035 10598.065 1187.865 ;
      RECT 10597.225 1048.035 10597.505 1187.625 ;
      RECT 10596.665 1048.035 10596.945 1187.385 ;
      RECT 10596.105 1048.035 10596.385 1187.145 ;
      RECT 10595.545 1048.035 10595.825 1186.905 ;
      RECT 10594.985 1048.035 10595.265 1186.665 ;
      RECT 10594.425 1048.035 10594.705 1186.425 ;
      RECT 10593.865 1048.035 10594.145 1186.185 ;
      RECT 10554.665 1048.035 10554.945 1193.09 ;
      RECT 10554.105 1048.035 10554.385 1193.33 ;
      RECT 10553.545 1048.035 10553.825 1193.57 ;
      RECT 10552.985 1046.935 10553.265 1193.81 ;
      RECT 10552.425 1048.035 10552.705 1194.05 ;
      RECT 10551.865 1046.935 10552.145 1194.29 ;
      RECT 10551.305 1048.035 10551.585 1194.53 ;
      RECT 10550.745 1048.035 10551.025 1194.77 ;
      RECT 10550.185 1048.035 10550.465 1195.01 ;
      RECT 10549.625 1046.935 10549.905 1195.25 ;
      RECT 10549.065 1048.035 10549.345 1195.49 ;
      RECT 10548.505 1046.935 10548.785 1195.73 ;
      RECT 10547.945 1048.035 10548.225 1195.97 ;
      RECT 10547.385 1046.935 10547.665 1196.21 ;
      RECT 10546.825 1048.035 10547.105 1196.45 ;
      RECT 10546.265 1048.035 10546.545 1196.69 ;
      RECT 10545.705 1048.035 10545.985 1196.69 ;
      RECT 10545.145 1048.035 10545.425 1196.45 ;
      RECT 10544.585 1048.035 10544.865 1196.21 ;
      RECT 10544.025 1048.035 10544.305 1195.97 ;
      RECT 10543.465 1048.035 10543.745 1195.73 ;
      RECT 10542.905 1048.035 10543.185 1195.49 ;
      RECT 10542.345 1048.035 10542.625 1195.25 ;
      RECT 10541.785 1048.035 10542.065 1195.01 ;
      RECT 10541.225 1048.035 10541.505 1194.77 ;
      RECT 10532.265 1048.035 10532.545 1194.285 ;
      RECT 10531.705 1046.935 10531.985 1194.045 ;
      RECT 10531.145 1048.035 10531.425 1193.805 ;
      RECT 10530.585 1046.935 10530.865 1193.565 ;
      RECT 10530.025 1048.035 10530.305 1193.325 ;
      RECT 10529.465 1046.935 10529.745 1193.085 ;
      RECT 10528.905 1048.035 10529.185 1192.845 ;
      RECT 10528.345 1048.035 10528.625 1192.605 ;
      RECT 10527.785 1048.035 10528.065 1192.365 ;
      RECT 10527.225 1048.035 10527.505 1192.125 ;
      RECT 10526.665 1048.035 10526.945 1191.885 ;
      RECT 10526.105 1048.035 10526.385 1191.645 ;
      RECT 10525.545 1048.035 10525.825 1191.405 ;
      RECT 10524.985 1048.035 10525.265 1191.165 ;
      RECT 10522.465 1046.935 10522.745 1192.885 ;
      RECT 10521.905 1048.035 10522.185 1192.645 ;
      RECT 10521.345 1046.935 10521.625 1192.405 ;
      RECT 10520.785 1048.035 10521.065 1192.165 ;
      RECT 10520.225 1048.035 10520.505 1191.925 ;
      RECT 10519.665 1048.035 10519.945 1191.685 ;
      RECT 10519.105 1048.035 10519.385 1191.445 ;
      RECT 10518.545 1048.035 10518.825 1191.205 ;
      RECT 10492.505 1048.035 10492.785 1188.855 ;
      RECT 10491.945 1048.035 10492.225 1189.095 ;
      RECT 10491.385 1048.035 10491.665 1189.335 ;
      RECT 10490.825 1048.035 10491.105 1189.58 ;
      RECT 10490.265 1048.035 10490.545 1189.82 ;
      RECT 10489.705 1048.035 10489.985 1190.06 ;
      RECT 10489.145 1048.035 10489.425 1190.06 ;
      RECT 10488.585 1048.035 10488.865 1189.82 ;
      RECT 10488.025 1048.035 10488.305 1189.58 ;
      RECT 10487.465 1046.935 10487.745 1189.34 ;
      RECT 10486.905 1048.035 10487.185 1189.1 ;
      RECT 10486.345 1046.935 10486.625 1188.86 ;
      RECT 10485.785 1048.035 10486.065 1188.62 ;
      RECT 10485.225 1048.035 10485.505 1188.38 ;
      RECT 10484.665 1048.035 10484.945 1188.14 ;
      RECT 10484.105 1046.935 10484.385 1187.9 ;
      RECT 10483.545 1048.035 10483.825 1187.66 ;
      RECT 10482.985 1046.935 10483.265 1187.42 ;
      RECT 10482.425 1048.035 10482.705 1187.18 ;
      RECT 10481.865 1046.935 10482.145 1186.94 ;
      RECT 10481.305 1048.035 10481.585 1186.7 ;
      RECT 10480.745 1048.035 10481.025 1186.46 ;
      RECT 10480.185 1048.035 10480.465 1186.22 ;
      RECT 10479.625 1048.035 10479.905 1185.98 ;
      RECT 10466.185 1048.035 10466.465 1191.78 ;
      RECT 10465.625 1048.035 10465.905 1191.54 ;
      RECT 10465.065 1048.035 10465.345 1191.3 ;
      RECT 10464.505 1048.035 10464.785 1191.06 ;
      RECT 10463.945 1048.035 10464.225 1190.82 ;
      RECT 10463.385 1048.035 10463.665 1190.58 ;
      RECT 10462.825 1048.035 10463.105 1190.34 ;
      RECT 10462.265 1048.035 10462.545 1190.1 ;
      RECT 10461.705 1046.935 10461.985 1189.86 ;
      RECT 10461.145 1048.035 10461.425 1189.62 ;
      RECT 10460.585 1046.935 10460.865 1189.3 ;
      RECT 10460.025 1048.035 10460.305 1189.14 ;
      RECT 10459.465 1046.935 10459.745 1188.9 ;
      RECT 10458.905 1048.035 10459.185 1188.66 ;
      RECT 10458.345 1048.035 10458.625 1188.42 ;
      RECT 10457.785 1048.035 10458.065 1188.18 ;
      RECT 10457.225 1048.035 10457.505 1187.94 ;
      RECT 10456.665 1048.035 10456.945 1187.7 ;
      RECT 10456.105 1048.035 10456.385 1187.46 ;
      RECT 10455.545 1048.035 10455.825 1187.22 ;
      RECT 10454.985 1048.035 10455.265 1186.98 ;
      RECT 10454.425 1046.935 10454.705 1186.74 ;
      RECT 10453.865 1048.035 10454.145 1186.5 ;
      RECT 10453.305 1046.935 10453.585 1186.26 ;
      RECT 10414.105 1048.035 10414.385 1191.87 ;
      RECT 10413.545 1048.035 10413.825 1192.11 ;
      RECT 10412.985 1048.035 10413.265 1192.35 ;
      RECT 10412.425 1048.035 10412.705 1192.59 ;
      RECT 10411.865 1048.035 10412.145 1192.83 ;
      RECT 10411.305 1048.035 10411.585 1193.07 ;
      RECT 10410.745 1048.035 10411.025 1193.31 ;
      RECT 10410.185 1048.035 10410.465 1193.55 ;
      RECT 10409.625 1048.035 10409.905 1193.79 ;
      RECT 10409.065 1048.035 10409.345 1194.03 ;
      RECT 10408.505 1048.035 10408.785 1194.27 ;
      RECT 10407.945 1048.035 10408.225 1194.51 ;
      RECT 10407.385 1048.035 10407.665 1194.75 ;
      RECT 10406.825 1048.035 10407.105 1194.75 ;
      RECT 10406.265 1046.935 10406.545 1194.51 ;
      RECT 10405.705 1048.035 10405.985 1194.27 ;
      RECT 10405.145 1046.935 10405.425 1194.03 ;
      RECT 10404.585 1048.035 10404.865 1193.79 ;
      RECT 10404.025 1048.035 10404.305 1193.55 ;
      RECT 10403.465 1048.035 10403.745 1193.31 ;
      RECT 10402.905 1046.935 10403.185 1193.045 ;
      RECT 10402.345 1048.035 10402.625 1192.805 ;
      RECT 10401.785 1046.935 10402.065 1192.565 ;
      RECT 10401.225 1048.035 10401.505 1192.325 ;
      RECT 10392.265 1046.935 10392.545 1186.16 ;
      RECT 10391.705 1048.035 10391.985 1186.4 ;
      RECT 10391.145 1048.035 10391.425 1186.64 ;
      RECT 10390.585 1048.035 10390.865 1186.64 ;
      RECT 10390.025 1048.035 10390.305 1186.4 ;
      RECT 10389.465 1048.035 10389.745 1186.16 ;
      RECT 10388.905 1048.035 10389.185 1185.92 ;
      RECT 10388.345 1048.035 10388.625 1185.68 ;
      RECT 10387.785 1048.035 10388.065 1185.44 ;
      RECT 10387.225 1048.035 10387.505 1185.2 ;
      RECT 10386.665 1048.035 10386.945 1184.96 ;
      RECT 10386.105 1048.035 10386.385 1184.72 ;
      RECT 10385.545 1048.035 10385.825 1184.48 ;
      RECT 10384.985 1046.935 10385.265 1184.24 ;
      RECT 10382.465 1048.035 10382.745 1185.96 ;
      RECT 10381.905 1046.935 10382.185 1185.72 ;
      RECT 10381.345 1048.035 10381.625 1185.48 ;
      RECT 10380.785 1046.935 10381.065 1185.24 ;
      RECT 10380.225 1048.035 10380.505 1185 ;
      RECT 10379.665 1048.035 10379.945 1184.76 ;
      RECT 10379.105 1048.035 10379.385 1184.52 ;
      RECT 10353.065 1048.035 10353.345 1187.305 ;
      RECT 10352.505 1048.035 10352.785 1187.545 ;
      RECT 10351.945 1048.035 10352.225 1187.785 ;
      RECT 10351.385 1048.035 10351.665 1188.025 ;
      RECT 10350.825 1048.035 10351.105 1188.265 ;
      RECT 10350.265 1046.935 10350.545 1188.505 ;
      RECT 10349.705 1048.035 10349.985 1188.745 ;
      RECT 10349.145 1046.935 10349.425 1188.985 ;
      RECT 10348.585 1048.035 10348.865 1189.225 ;
      RECT 10348.025 1048.035 10348.305 1189.465 ;
      RECT 10347.465 1048.035 10347.745 1189.705 ;
      RECT 10346.905 1048.035 10347.185 1189.945 ;
      RECT 10346.345 1048.035 10346.625 1190.185 ;
      RECT 10345.785 1048.035 10346.065 1190.425 ;
      RECT 10345.225 1048.035 10345.505 1190.665 ;
      RECT 10344.665 1048.035 10344.945 1190.665 ;
      RECT 10344.105 1048.035 10344.385 1190.425 ;
      RECT 10343.545 1048.035 10343.825 1190.185 ;
      RECT 10342.985 1048.035 10343.265 1189.945 ;
      RECT 10342.425 1048.035 10342.705 1189.7 ;
      RECT 10341.865 1048.035 10342.145 1189.46 ;
      RECT 10341.305 1048.035 10341.585 1189.22 ;
      RECT 10340.745 1046.935 10341.025 1188.98 ;
      RECT 10340.185 1048.035 10340.465 1188.74 ;
      RECT 10326.745 1046.935 10327.025 1186.22 ;
      RECT 10326.185 1048.035 10326.465 1185.98 ;
      RECT 10325.625 1048.035 10325.905 1185.74 ;
      RECT 10325.065 1048.035 10325.345 1185.5 ;
      RECT 10324.505 1046.935 10324.785 1185.26 ;
      RECT 10323.945 1048.035 10324.225 1185.02 ;
      RECT 10323.385 1046.935 10323.665 1184.78 ;
      RECT 10322.825 1048.035 10323.105 1184.54 ;
      RECT 10322.265 1046.935 10322.545 1184.3 ;
      RECT 10321.705 1048.035 10321.985 1184.06 ;
      RECT 10321.145 1048.035 10321.425 1183.82 ;
      RECT 10320.585 1048.035 10320.865 1183.58 ;
      RECT 10320.025 1048.035 10320.305 1183.34 ;
      RECT 10319.465 1048.035 10319.745 1183.1 ;
      RECT 10318.905 1048.035 10319.185 1182.86 ;
      RECT 10318.345 1048.035 10318.625 1182.62 ;
      RECT 10317.785 1048.035 10318.065 1182.38 ;
      RECT 10317.225 1048.035 10317.505 1182.14 ;
      RECT 10316.665 1048.035 10316.945 1181.9 ;
      RECT 10316.105 1048.035 10316.385 1181.66 ;
      RECT 10315.545 1048.035 10315.825 1181.42 ;
      RECT 10314.985 1046.935 10315.265 1181.18 ;
      RECT 10314.425 1048.035 10314.705 1180.94 ;
      RECT 10313.865 1046.935 10314.145 1180.7 ;
      RECT 10274.105 1048.035 10274.385 1191.17 ;
      RECT 10273.545 1046.935 10273.825 1191.41 ;
      RECT 10272.985 1048.035 10273.265 1191.65 ;
      RECT 10272.425 1048.035 10272.705 1191.89 ;
      RECT 10271.865 1048.035 10272.145 1192.13 ;
      RECT 10271.305 1048.035 10271.585 1192.37 ;
      RECT 10270.745 1048.035 10271.025 1192.61 ;
      RECT 10270.185 1048.035 10270.465 1192.855 ;
      RECT 10269.625 1048.035 10269.905 1193.095 ;
      RECT 10269.065 1048.035 10269.345 1193.335 ;
      RECT 10268.505 1046.935 10268.785 1193.575 ;
      RECT 10267.945 1048.035 10268.225 1193.815 ;
      RECT 10267.385 1046.935 10267.665 1194.055 ;
      RECT 10266.825 1048.035 10267.105 1194.295 ;
      RECT 10266.265 1048.035 10266.545 1194.535 ;
      RECT 10265.705 1048.035 10265.985 1194.775 ;
      RECT 10265.145 1048.035 10265.425 1195.015 ;
      RECT 10264.585 1048.035 10264.865 1195.255 ;
      RECT 10264.025 1048.035 10264.305 1195.495 ;
      RECT 10263.465 1048.035 10263.745 1195.735 ;
      RECT 10262.905 1048.035 10263.185 1195.975 ;
      RECT 10262.345 1048.035 10262.625 1196.215 ;
      RECT 10261.785 1048.035 10262.065 1196.455 ;
      RECT 10261.225 1048.035 10261.505 1196.695 ;
      RECT 10252.265 1048.035 10252.545 1192.28 ;
      RECT 10251.705 1048.035 10251.985 1192.04 ;
      RECT 10251.145 1048.035 10251.425 1191.8 ;
      RECT 10250.585 1046.935 10250.865 1191.56 ;
      RECT 10250.025 1048.035 10250.305 1191.32 ;
      RECT 10249.465 1046.935 10249.745 1191.08 ;
      RECT 10248.905 1048.035 10249.185 1190.84 ;
      RECT 10248.345 1048.035 10248.625 1190.6 ;
      RECT 10247.785 1048.035 10248.065 1190.36 ;
      RECT 10247.225 1046.935 10247.505 1190.12 ;
      RECT 10246.665 1048.035 10246.945 1189.88 ;
      RECT 10246.105 1046.935 10246.385 1189.64 ;
      RECT 10245.545 1048.035 10245.825 1189.4 ;
      RECT 10244.985 1046.935 10245.265 1189.16 ;
      RECT 10242.465 1048.035 10242.745 1181.56 ;
      RECT 10241.905 1048.035 10242.185 1181.32 ;
      RECT 10241.345 1048.035 10241.625 1181.08 ;
      RECT 10240.785 1048.035 10241.065 1180.84 ;
      RECT 10240.225 1048.035 10240.505 1180.6 ;
      RECT 10239.665 1048.035 10239.945 1180.36 ;
      RECT 10239.105 1048.035 10239.385 1180.12 ;
      RECT 10213.065 1048.035 10213.345 1193.995 ;
      RECT 10212.505 1048.035 10212.785 1194.235 ;
      RECT 10211.945 1048.035 10212.225 1194.475 ;
      RECT 10211.385 1048.035 10211.665 1194.715 ;
      RECT 10210.825 1048.035 10211.105 1194.955 ;
      RECT 10210.265 1046.935 10210.545 1194.955 ;
      RECT 10209.705 1048.035 10209.985 1194.715 ;
      RECT 10209.145 1046.935 10209.425 1194.47 ;
      RECT 10208.585 1048.035 10208.865 1194.23 ;
      RECT 10208.025 1046.935 10208.305 1193.99 ;
      RECT 10207.465 1048.035 10207.745 1193.75 ;
      RECT 10206.905 1048.035 10207.185 1193.51 ;
      RECT 10206.345 1048.035 10206.625 1193.27 ;
      RECT 10205.785 1048.035 10206.065 1193.03 ;
      RECT 10205.225 1048.035 10205.505 1192.79 ;
      RECT 10204.665 1048.035 10204.945 1192.55 ;
      RECT 10204.105 1048.035 10204.385 1192.31 ;
      RECT 10203.545 1048.035 10203.825 1192.07 ;
      RECT 10202.985 1046.935 10203.265 1191.83 ;
      RECT 10202.425 1048.035 10202.705 1191.59 ;
      RECT 10201.865 1046.935 10202.145 1191.35 ;
      RECT 10201.305 1048.035 10201.585 1191.11 ;
      RECT 10200.745 1048.035 10201.025 1190.87 ;
      RECT 10200.185 1048.035 10200.465 1190.63 ;
      RECT 10186.745 1048.035 10187.025 1194.03 ;
      RECT 10186.185 1048.035 10186.465 1194.27 ;
      RECT 10185.625 1048.035 10185.905 1194.515 ;
      RECT 10185.065 1048.035 10185.345 1194.755 ;
      RECT 10184.505 1048.035 10184.785 1194.995 ;
      RECT 10183.945 1048.035 10184.225 1194.995 ;
      RECT 10183.385 1048.035 10183.665 1194.755 ;
      RECT 10182.825 1048.035 10183.105 1194.515 ;
      RECT 10182.265 1048.035 10182.545 1187.5 ;
      RECT 10181.705 1048.035 10181.985 1187.26 ;
      RECT 10181.145 1048.035 10181.425 1187.02 ;
      RECT 10180.585 1046.935 10180.865 1186.78 ;
      RECT 10180.025 1048.035 10180.305 1186.54 ;
      RECT 10179.465 1046.935 10179.745 1186.3 ;
      RECT 10178.905 1048.035 10179.185 1186.06 ;
      RECT 10178.345 1048.035 10178.625 1185.82 ;
      RECT 10177.785 1048.035 10178.065 1185.58 ;
      RECT 10177.225 1046.935 10177.505 1185.34 ;
      RECT 10176.665 1048.035 10176.945 1185.1 ;
      RECT 10176.105 1046.935 10176.385 1184.86 ;
      RECT 10175.545 1048.035 10175.825 1184.62 ;
      RECT 10174.985 1046.935 10175.265 1184.38 ;
      RECT 10174.425 1048.035 10174.705 1184.14 ;
      RECT 10173.865 1048.035 10174.145 1183.9 ;
      RECT 10133.545 1048.035 10133.825 1192.795 ;
      RECT 10132.985 1048.035 10133.265 1193.035 ;
      RECT 10132.425 1048.035 10132.705 1193.28 ;
      RECT 10131.865 1048.035 10132.145 1193.52 ;
      RECT 10131.305 1048.035 10131.585 1193.76 ;
      RECT 10130.745 1048.035 10131.025 1194 ;
      RECT 10130.185 1048.035 10130.465 1194.24 ;
      RECT 10129.625 1048.035 10129.905 1194.48 ;
      RECT 10129.065 1048.035 10129.345 1194.72 ;
      RECT 10128.505 1048.035 10128.785 1194.96 ;
      RECT 10127.945 1046.935 10128.225 1195.2 ;
      RECT 10127.385 1048.035 10127.665 1195.44 ;
      RECT 10126.825 1046.935 10127.105 1195.68 ;
      RECT 10126.265 1048.035 10126.545 1195.92 ;
      RECT 10125.705 1046.935 10125.985 1196.16 ;
      RECT 10125.145 1048.035 10125.425 1196.16 ;
      RECT 10124.585 1048.035 10124.865 1195.92 ;
      RECT 10124.025 1048.035 10124.305 1195.68 ;
      RECT 10123.465 1048.035 10123.745 1195.44 ;
      RECT 10122.905 1048.035 10123.185 1195.2 ;
      RECT 10122.345 1048.035 10122.625 1194.96 ;
      RECT 10121.785 1048.035 10122.065 1194.72 ;
      RECT 10121.225 1048.035 10121.505 1194.48 ;
      RECT 10112.265 1046.935 10112.545 1194.51 ;
      RECT 10111.705 1048.035 10111.985 1194.75 ;
      RECT 10111.145 1046.935 10111.425 1194.99 ;
      RECT 10110.585 1048.035 10110.865 1195.205 ;
      RECT 10110.025 1048.035 10110.305 1194.78 ;
      RECT 10109.465 1048.035 10109.745 1194.54 ;
      RECT 10108.905 1048.035 10109.185 1194.3 ;
      RECT 10108.345 1048.035 10108.625 1194.06 ;
      RECT 10107.785 1048.035 10108.065 1193.82 ;
      RECT 10107.225 1048.035 10107.505 1193.58 ;
      RECT 10106.665 1048.035 10106.945 1193.34 ;
      RECT 10106.105 1048.035 10106.385 1193.1 ;
      RECT 10105.545 1048.035 10105.825 1192.86 ;
      RECT 10104.985 1048.035 10105.265 1192.62 ;
      RECT 10102.465 1048.035 10102.745 1191.795 ;
      RECT 10101.905 1048.035 10102.185 1191.555 ;
      RECT 10101.345 1048.035 10101.625 1191.315 ;
      RECT 10100.785 1046.935 10101.065 1191.075 ;
      RECT 10100.225 1048.035 10100.505 1190.835 ;
      RECT 10099.665 1046.935 10099.945 1190.595 ;
      RECT 10099.105 1048.035 10099.385 1190.355 ;
      RECT 10098.545 1048.035 10098.825 1190.115 ;
      RECT 10071.945 1048.035 10072.225 1201.16 ;
      RECT 10071.385 1046.935 10071.665 1201.4 ;
      RECT 10070.825 1048.035 10071.105 1201.64 ;
      RECT 10070.265 1046.935 10070.545 1201.885 ;
      RECT 10069.705 1048.035 10069.985 1202.125 ;
      RECT 10069.145 1046.935 10069.425 1202.365 ;
      RECT 10068.585 1048.035 10068.865 1202.605 ;
      RECT 10068.025 1048.035 10068.305 1202.845 ;
      RECT 10067.465 1048.035 10067.745 1188.465 ;
      RECT 10066.905 1048.035 10067.185 1188.225 ;
      RECT 10066.345 1048.035 10066.625 1187.985 ;
      RECT 10065.785 1048.035 10066.065 1187.745 ;
      RECT 10065.225 1048.035 10065.505 1187.505 ;
      RECT 10064.665 1048.035 10064.945 1187.265 ;
      RECT 10064.105 1048.035 10064.385 1187.025 ;
      RECT 10063.545 1048.035 10063.825 1186.785 ;
      RECT 10062.985 1048.035 10063.265 1186.545 ;
      RECT 10062.425 1048.035 10062.705 1186.305 ;
      RECT 10061.865 1046.935 10062.145 1186.065 ;
      RECT 10061.305 1048.035 10061.585 1185.825 ;
      RECT 10060.745 1046.935 10061.025 1185.585 ;
      RECT 10060.185 1048.035 10060.465 1185.345 ;
      RECT 10046.185 1046.935 10046.465 1191.465 ;
      RECT 10045.625 1048.035 10045.905 1191.225 ;
      RECT 10045.065 1048.035 10045.345 1190.985 ;
      RECT 10044.505 1048.035 10044.785 1190.745 ;
      RECT 10043.945 1048.035 10044.225 1190.505 ;
      RECT 10043.385 1048.035 10043.665 1190.265 ;
      RECT 10042.825 1048.035 10043.105 1190.025 ;
      RECT 10042.265 1048.035 10042.545 1189.785 ;
      RECT 10041.705 1048.035 10041.985 1189.545 ;
      RECT 10041.145 1046.935 10041.425 1189.305 ;
      RECT 10040.585 1048.035 10040.865 1189.065 ;
      RECT 10040.025 1046.935 10040.305 1188.825 ;
      RECT 10039.465 1048.035 10039.745 1188.585 ;
      RECT 10038.905 1048.035 10039.185 1188.345 ;
      RECT 10038.345 1048.035 10038.625 1188.105 ;
      RECT 10037.785 1048.035 10038.065 1187.865 ;
      RECT 10037.225 1048.035 10037.505 1187.625 ;
      RECT 10036.665 1048.035 10036.945 1187.385 ;
      RECT 10036.105 1048.035 10036.385 1187.145 ;
      RECT 10035.545 1048.035 10035.825 1186.905 ;
      RECT 10034.985 1048.035 10035.265 1186.665 ;
      RECT 10034.425 1048.035 10034.705 1186.425 ;
      RECT 10033.865 1048.035 10034.145 1186.185 ;
      RECT 9994.665 1048.035 9994.945 1193.09 ;
      RECT 9994.105 1048.035 9994.385 1193.33 ;
      RECT 9993.545 1048.035 9993.825 1193.57 ;
      RECT 9992.985 1046.935 9993.265 1193.81 ;
      RECT 9992.425 1048.035 9992.705 1194.05 ;
      RECT 9991.865 1046.935 9992.145 1194.29 ;
      RECT 9991.305 1048.035 9991.585 1194.53 ;
      RECT 9990.745 1048.035 9991.025 1194.77 ;
      RECT 9990.185 1048.035 9990.465 1195.01 ;
      RECT 9989.625 1046.935 9989.905 1195.25 ;
      RECT 9989.065 1048.035 9989.345 1195.49 ;
      RECT 9988.505 1046.935 9988.785 1195.73 ;
      RECT 9987.945 1048.035 9988.225 1195.97 ;
      RECT 9987.385 1046.935 9987.665 1196.21 ;
      RECT 9986.825 1048.035 9987.105 1196.45 ;
      RECT 9986.265 1048.035 9986.545 1196.69 ;
      RECT 9985.705 1048.035 9985.985 1196.69 ;
      RECT 9985.145 1048.035 9985.425 1196.45 ;
      RECT 9984.585 1048.035 9984.865 1196.21 ;
      RECT 9984.025 1048.035 9984.305 1195.97 ;
      RECT 9983.465 1048.035 9983.745 1195.73 ;
      RECT 9982.905 1048.035 9983.185 1195.49 ;
      RECT 9982.345 1048.035 9982.625 1195.25 ;
      RECT 9981.785 1048.035 9982.065 1195.01 ;
      RECT 9981.225 1048.035 9981.505 1194.77 ;
      RECT 9972.265 1048.035 9972.545 1194.285 ;
      RECT 9971.705 1046.935 9971.985 1194.045 ;
      RECT 9971.145 1048.035 9971.425 1193.805 ;
      RECT 9970.585 1046.935 9970.865 1193.565 ;
      RECT 9970.025 1048.035 9970.305 1193.325 ;
      RECT 9969.465 1046.935 9969.745 1193.085 ;
      RECT 9968.905 1048.035 9969.185 1192.845 ;
      RECT 9968.345 1048.035 9968.625 1192.605 ;
      RECT 9967.785 1048.035 9968.065 1192.365 ;
      RECT 9967.225 1048.035 9967.505 1192.125 ;
      RECT 9966.665 1048.035 9966.945 1191.885 ;
      RECT 9966.105 1048.035 9966.385 1191.645 ;
      RECT 9965.545 1048.035 9965.825 1191.405 ;
      RECT 9964.985 1048.035 9965.265 1191.165 ;
      RECT 9962.465 1046.935 9962.745 1192.885 ;
      RECT 9961.905 1048.035 9962.185 1192.645 ;
      RECT 9961.345 1046.935 9961.625 1192.405 ;
      RECT 9960.785 1048.035 9961.065 1192.165 ;
      RECT 9960.225 1048.035 9960.505 1191.925 ;
      RECT 9959.665 1048.035 9959.945 1191.685 ;
      RECT 9959.105 1048.035 9959.385 1191.445 ;
      RECT 9958.545 1048.035 9958.825 1191.205 ;
      RECT 9932.505 1048.035 9932.785 1188.855 ;
      RECT 9931.945 1048.035 9932.225 1189.095 ;
      RECT 9931.385 1048.035 9931.665 1189.335 ;
      RECT 9930.825 1048.035 9931.105 1189.58 ;
      RECT 9930.265 1048.035 9930.545 1189.82 ;
      RECT 9929.705 1048.035 9929.985 1190.06 ;
      RECT 9929.145 1048.035 9929.425 1190.06 ;
      RECT 9928.585 1048.035 9928.865 1189.82 ;
      RECT 9928.025 1048.035 9928.305 1189.58 ;
      RECT 9927.465 1046.935 9927.745 1189.34 ;
      RECT 9926.905 1048.035 9927.185 1189.1 ;
      RECT 9926.345 1046.935 9926.625 1188.86 ;
      RECT 9925.785 1048.035 9926.065 1188.62 ;
      RECT 9925.225 1048.035 9925.505 1188.38 ;
      RECT 9924.665 1048.035 9924.945 1188.14 ;
      RECT 9924.105 1046.935 9924.385 1187.9 ;
      RECT 9923.545 1048.035 9923.825 1187.66 ;
      RECT 9922.985 1046.935 9923.265 1187.42 ;
      RECT 9922.425 1048.035 9922.705 1187.18 ;
      RECT 9921.865 1046.935 9922.145 1186.94 ;
      RECT 9921.305 1048.035 9921.585 1186.7 ;
      RECT 9920.745 1048.035 9921.025 1186.46 ;
      RECT 9920.185 1048.035 9920.465 1186.22 ;
      RECT 9919.625 1048.035 9919.905 1185.98 ;
      RECT 9906.185 1048.035 9906.465 1191.78 ;
      RECT 9905.625 1048.035 9905.905 1191.54 ;
      RECT 9905.065 1048.035 9905.345 1191.3 ;
      RECT 9904.505 1048.035 9904.785 1191.06 ;
      RECT 9903.945 1048.035 9904.225 1190.82 ;
      RECT 9903.385 1048.035 9903.665 1190.58 ;
      RECT 9902.825 1048.035 9903.105 1190.34 ;
      RECT 9902.265 1048.035 9902.545 1190.1 ;
      RECT 9901.705 1046.935 9901.985 1189.86 ;
      RECT 9901.145 1048.035 9901.425 1189.62 ;
      RECT 9900.585 1046.935 9900.865 1189.3 ;
      RECT 9900.025 1048.035 9900.305 1189.14 ;
      RECT 9899.465 1046.935 9899.745 1188.9 ;
      RECT 9898.905 1048.035 9899.185 1188.66 ;
      RECT 9898.345 1048.035 9898.625 1188.42 ;
      RECT 9897.785 1048.035 9898.065 1188.18 ;
      RECT 9897.225 1048.035 9897.505 1187.94 ;
      RECT 9896.665 1048.035 9896.945 1187.7 ;
      RECT 9896.105 1048.035 9896.385 1187.46 ;
      RECT 9895.545 1048.035 9895.825 1187.22 ;
      RECT 9894.985 1048.035 9895.265 1186.98 ;
      RECT 9894.425 1046.935 9894.705 1186.74 ;
      RECT 9893.865 1048.035 9894.145 1186.5 ;
      RECT 9893.305 1046.935 9893.585 1186.26 ;
      RECT 9854.105 1048.035 9854.385 1191.87 ;
      RECT 9853.545 1048.035 9853.825 1192.11 ;
      RECT 9852.985 1048.035 9853.265 1192.35 ;
      RECT 9852.425 1048.035 9852.705 1192.59 ;
      RECT 9851.865 1048.035 9852.145 1192.83 ;
      RECT 9851.305 1048.035 9851.585 1193.07 ;
      RECT 9850.745 1048.035 9851.025 1193.31 ;
      RECT 9850.185 1048.035 9850.465 1193.55 ;
      RECT 9849.625 1048.035 9849.905 1193.79 ;
      RECT 9849.065 1048.035 9849.345 1194.03 ;
      RECT 9848.505 1048.035 9848.785 1194.27 ;
      RECT 9847.945 1048.035 9848.225 1194.51 ;
      RECT 9847.385 1048.035 9847.665 1194.75 ;
      RECT 9846.825 1048.035 9847.105 1194.75 ;
      RECT 9846.265 1046.935 9846.545 1194.51 ;
      RECT 9845.705 1048.035 9845.985 1194.27 ;
      RECT 9845.145 1046.935 9845.425 1194.03 ;
      RECT 9844.585 1048.035 9844.865 1193.79 ;
      RECT 9844.025 1048.035 9844.305 1193.55 ;
      RECT 9843.465 1048.035 9843.745 1193.31 ;
      RECT 9842.905 1046.935 9843.185 1193.045 ;
      RECT 9842.345 1048.035 9842.625 1192.805 ;
      RECT 9841.785 1046.935 9842.065 1192.565 ;
      RECT 9841.225 1048.035 9841.505 1192.325 ;
      RECT 9832.265 1046.935 9832.545 1186.16 ;
      RECT 9831.705 1048.035 9831.985 1186.4 ;
      RECT 9831.145 1048.035 9831.425 1186.64 ;
      RECT 9830.585 1048.035 9830.865 1186.64 ;
      RECT 9830.025 1048.035 9830.305 1186.4 ;
      RECT 9829.465 1048.035 9829.745 1186.16 ;
      RECT 9828.905 1048.035 9829.185 1185.92 ;
      RECT 9828.345 1048.035 9828.625 1185.68 ;
      RECT 9827.785 1048.035 9828.065 1185.44 ;
      RECT 9827.225 1048.035 9827.505 1185.2 ;
      RECT 9826.665 1048.035 9826.945 1184.96 ;
      RECT 9826.105 1048.035 9826.385 1184.72 ;
      RECT 9825.545 1048.035 9825.825 1184.48 ;
      RECT 9824.985 1046.935 9825.265 1184.24 ;
      RECT 9822.465 1048.035 9822.745 1185.96 ;
      RECT 9821.905 1046.935 9822.185 1185.72 ;
      RECT 9821.345 1048.035 9821.625 1185.48 ;
      RECT 9820.785 1046.935 9821.065 1185.24 ;
      RECT 9820.225 1048.035 9820.505 1185 ;
      RECT 9819.665 1048.035 9819.945 1184.76 ;
      RECT 9819.105 1048.035 9819.385 1184.52 ;
      RECT 9793.065 1048.035 9793.345 1187.305 ;
      RECT 9792.505 1048.035 9792.785 1187.545 ;
      RECT 9791.945 1048.035 9792.225 1187.785 ;
      RECT 9791.385 1048.035 9791.665 1188.025 ;
      RECT 9790.825 1048.035 9791.105 1188.265 ;
      RECT 9790.265 1046.935 9790.545 1188.505 ;
      RECT 9789.705 1048.035 9789.985 1188.745 ;
      RECT 9789.145 1046.935 9789.425 1188.985 ;
      RECT 9788.585 1048.035 9788.865 1189.225 ;
      RECT 9788.025 1048.035 9788.305 1189.465 ;
      RECT 9787.465 1048.035 9787.745 1189.705 ;
      RECT 9786.905 1048.035 9787.185 1189.945 ;
      RECT 9786.345 1048.035 9786.625 1190.185 ;
      RECT 9785.785 1048.035 9786.065 1190.425 ;
      RECT 9785.225 1048.035 9785.505 1190.665 ;
      RECT 9784.665 1048.035 9784.945 1190.665 ;
      RECT 9784.105 1048.035 9784.385 1190.425 ;
      RECT 9783.545 1048.035 9783.825 1190.185 ;
      RECT 9782.985 1048.035 9783.265 1189.945 ;
      RECT 9782.425 1048.035 9782.705 1189.7 ;
      RECT 9781.865 1048.035 9782.145 1189.46 ;
      RECT 9781.305 1048.035 9781.585 1189.22 ;
      RECT 9780.745 1046.935 9781.025 1188.98 ;
      RECT 9780.185 1048.035 9780.465 1188.74 ;
      RECT 9766.745 1046.935 9767.025 1186.22 ;
      RECT 9766.185 1048.035 9766.465 1185.98 ;
      RECT 9765.625 1048.035 9765.905 1185.74 ;
      RECT 9765.065 1048.035 9765.345 1185.5 ;
      RECT 9764.505 1046.935 9764.785 1185.26 ;
      RECT 9763.945 1048.035 9764.225 1185.02 ;
      RECT 9763.385 1046.935 9763.665 1184.78 ;
      RECT 9762.825 1048.035 9763.105 1184.54 ;
      RECT 9762.265 1046.935 9762.545 1184.3 ;
      RECT 9761.705 1048.035 9761.985 1184.06 ;
      RECT 9761.145 1048.035 9761.425 1183.82 ;
      RECT 9760.585 1048.035 9760.865 1183.58 ;
      RECT 9760.025 1048.035 9760.305 1183.34 ;
      RECT 9759.465 1048.035 9759.745 1183.1 ;
      RECT 9758.905 1048.035 9759.185 1182.86 ;
      RECT 9758.345 1048.035 9758.625 1182.62 ;
      RECT 9757.785 1048.035 9758.065 1182.38 ;
      RECT 9757.225 1048.035 9757.505 1182.14 ;
      RECT 9756.665 1048.035 9756.945 1181.9 ;
      RECT 9756.105 1048.035 9756.385 1181.66 ;
      RECT 9755.545 1048.035 9755.825 1181.42 ;
      RECT 9754.985 1046.935 9755.265 1181.18 ;
      RECT 9754.425 1048.035 9754.705 1180.94 ;
      RECT 9753.865 1046.935 9754.145 1180.7 ;
      RECT 9714.105 1048.035 9714.385 1191.17 ;
      RECT 9713.545 1046.935 9713.825 1191.41 ;
      RECT 9712.985 1048.035 9713.265 1191.65 ;
      RECT 9712.425 1048.035 9712.705 1191.89 ;
      RECT 9711.865 1048.035 9712.145 1192.13 ;
      RECT 9711.305 1048.035 9711.585 1192.37 ;
      RECT 9710.745 1048.035 9711.025 1192.61 ;
      RECT 9710.185 1048.035 9710.465 1192.855 ;
      RECT 9709.625 1048.035 9709.905 1193.095 ;
      RECT 9709.065 1048.035 9709.345 1193.335 ;
      RECT 9708.505 1046.935 9708.785 1193.575 ;
      RECT 9707.945 1048.035 9708.225 1193.815 ;
      RECT 9707.385 1046.935 9707.665 1194.055 ;
      RECT 9706.825 1048.035 9707.105 1194.295 ;
      RECT 9706.265 1048.035 9706.545 1194.535 ;
      RECT 9705.705 1048.035 9705.985 1194.775 ;
      RECT 9705.145 1048.035 9705.425 1195.015 ;
      RECT 9704.585 1048.035 9704.865 1195.255 ;
      RECT 9704.025 1048.035 9704.305 1195.495 ;
      RECT 9703.465 1048.035 9703.745 1195.735 ;
      RECT 9702.905 1048.035 9703.185 1195.975 ;
      RECT 9702.345 1048.035 9702.625 1196.215 ;
      RECT 9701.785 1048.035 9702.065 1196.455 ;
      RECT 9701.225 1048.035 9701.505 1196.695 ;
      RECT 9692.265 1048.035 9692.545 1192.28 ;
      RECT 9691.705 1048.035 9691.985 1192.04 ;
      RECT 9691.145 1048.035 9691.425 1191.8 ;
      RECT 9690.585 1046.935 9690.865 1191.56 ;
      RECT 9690.025 1048.035 9690.305 1191.32 ;
      RECT 9689.465 1046.935 9689.745 1191.08 ;
      RECT 9688.905 1048.035 9689.185 1190.84 ;
      RECT 9688.345 1048.035 9688.625 1190.6 ;
      RECT 9687.785 1048.035 9688.065 1190.36 ;
      RECT 9687.225 1046.935 9687.505 1190.12 ;
      RECT 9686.665 1048.035 9686.945 1189.88 ;
      RECT 9686.105 1046.935 9686.385 1189.64 ;
      RECT 9685.545 1048.035 9685.825 1189.4 ;
      RECT 9684.985 1046.935 9685.265 1189.16 ;
      RECT 9682.465 1048.035 9682.745 1181.56 ;
      RECT 9681.905 1048.035 9682.185 1181.32 ;
      RECT 9681.345 1048.035 9681.625 1181.08 ;
      RECT 9680.785 1048.035 9681.065 1180.84 ;
      RECT 9680.225 1048.035 9680.505 1180.6 ;
      RECT 9679.665 1048.035 9679.945 1180.36 ;
      RECT 9679.105 1048.035 9679.385 1180.12 ;
      RECT 9653.065 1048.035 9653.345 1193.995 ;
      RECT 9652.505 1048.035 9652.785 1194.235 ;
      RECT 9651.945 1048.035 9652.225 1194.475 ;
      RECT 9651.385 1048.035 9651.665 1194.715 ;
      RECT 9650.825 1048.035 9651.105 1194.955 ;
      RECT 9650.265 1046.935 9650.545 1194.955 ;
      RECT 9649.705 1048.035 9649.985 1194.715 ;
      RECT 9649.145 1046.935 9649.425 1194.47 ;
      RECT 9648.585 1048.035 9648.865 1194.23 ;
      RECT 9648.025 1046.935 9648.305 1193.99 ;
      RECT 9647.465 1048.035 9647.745 1193.75 ;
      RECT 9646.905 1048.035 9647.185 1193.51 ;
      RECT 9646.345 1048.035 9646.625 1193.27 ;
      RECT 9645.785 1048.035 9646.065 1193.03 ;
      RECT 9645.225 1048.035 9645.505 1192.79 ;
      RECT 9644.665 1048.035 9644.945 1192.55 ;
      RECT 9644.105 1048.035 9644.385 1192.31 ;
      RECT 9643.545 1048.035 9643.825 1192.07 ;
      RECT 9642.985 1046.935 9643.265 1191.83 ;
      RECT 9642.425 1048.035 9642.705 1191.59 ;
      RECT 9641.865 1046.935 9642.145 1191.35 ;
      RECT 9641.305 1048.035 9641.585 1191.11 ;
      RECT 9640.745 1048.035 9641.025 1190.87 ;
      RECT 9640.185 1048.035 9640.465 1190.63 ;
      RECT 9626.745 1048.035 9627.025 1194.03 ;
      RECT 9626.185 1048.035 9626.465 1194.27 ;
      RECT 9625.625 1048.035 9625.905 1194.515 ;
      RECT 9625.065 1048.035 9625.345 1194.755 ;
      RECT 9624.505 1048.035 9624.785 1194.995 ;
      RECT 9623.945 1048.035 9624.225 1194.995 ;
      RECT 9623.385 1048.035 9623.665 1194.755 ;
      RECT 9622.825 1048.035 9623.105 1194.515 ;
      RECT 9622.265 1048.035 9622.545 1187.5 ;
      RECT 9621.705 1048.035 9621.985 1187.26 ;
      RECT 9621.145 1048.035 9621.425 1187.02 ;
      RECT 9620.585 1046.935 9620.865 1186.78 ;
      RECT 9620.025 1048.035 9620.305 1186.54 ;
      RECT 9619.465 1046.935 9619.745 1186.3 ;
      RECT 9618.905 1048.035 9619.185 1186.06 ;
      RECT 9618.345 1048.035 9618.625 1185.82 ;
      RECT 9617.785 1048.035 9618.065 1185.58 ;
      RECT 9617.225 1046.935 9617.505 1185.34 ;
      RECT 9616.665 1048.035 9616.945 1185.1 ;
      RECT 9616.105 1046.935 9616.385 1184.86 ;
      RECT 9615.545 1048.035 9615.825 1184.62 ;
      RECT 9614.985 1046.935 9615.265 1184.38 ;
      RECT 9614.425 1048.035 9614.705 1184.14 ;
      RECT 9613.865 1048.035 9614.145 1183.9 ;
      RECT 9573.545 1048.035 9573.825 1192.795 ;
      RECT 9572.985 1048.035 9573.265 1193.035 ;
      RECT 9572.425 1048.035 9572.705 1193.28 ;
      RECT 9571.865 1048.035 9572.145 1193.52 ;
      RECT 9571.305 1048.035 9571.585 1193.76 ;
      RECT 9570.745 1048.035 9571.025 1194 ;
      RECT 9570.185 1048.035 9570.465 1194.24 ;
      RECT 9569.625 1048.035 9569.905 1194.48 ;
      RECT 9569.065 1048.035 9569.345 1194.72 ;
      RECT 9568.505 1048.035 9568.785 1194.96 ;
      RECT 9567.945 1046.935 9568.225 1195.2 ;
      RECT 9567.385 1048.035 9567.665 1195.44 ;
      RECT 9566.825 1046.935 9567.105 1195.68 ;
      RECT 9566.265 1048.035 9566.545 1195.92 ;
      RECT 9565.705 1046.935 9565.985 1196.16 ;
      RECT 9565.145 1048.035 9565.425 1196.16 ;
      RECT 9564.585 1048.035 9564.865 1195.92 ;
      RECT 9564.025 1048.035 9564.305 1195.68 ;
      RECT 9563.465 1048.035 9563.745 1195.44 ;
      RECT 9562.905 1048.035 9563.185 1195.2 ;
      RECT 9562.345 1048.035 9562.625 1194.96 ;
      RECT 9561.785 1048.035 9562.065 1194.72 ;
      RECT 9561.225 1048.035 9561.505 1194.48 ;
      RECT 9552.265 1046.935 9552.545 1194.51 ;
      RECT 9551.705 1048.035 9551.985 1194.75 ;
      RECT 9551.145 1046.935 9551.425 1194.99 ;
      RECT 9550.585 1048.035 9550.865 1195.205 ;
      RECT 9550.025 1048.035 9550.305 1194.78 ;
      RECT 9549.465 1048.035 9549.745 1194.54 ;
      RECT 9548.905 1048.035 9549.185 1194.3 ;
      RECT 9548.345 1048.035 9548.625 1194.06 ;
      RECT 9547.785 1048.035 9548.065 1193.82 ;
      RECT 9547.225 1048.035 9547.505 1193.58 ;
      RECT 9546.665 1048.035 9546.945 1193.34 ;
      RECT 9546.105 1048.035 9546.385 1193.1 ;
      RECT 9545.545 1048.035 9545.825 1192.86 ;
      RECT 9544.985 1048.035 9545.265 1192.62 ;
      RECT 9542.465 1048.035 9542.745 1191.795 ;
      RECT 9541.905 1048.035 9542.185 1191.555 ;
      RECT 9541.345 1048.035 9541.625 1191.315 ;
      RECT 9540.785 1046.935 9541.065 1191.075 ;
      RECT 9540.225 1048.035 9540.505 1190.835 ;
      RECT 9539.665 1046.935 9539.945 1190.595 ;
      RECT 9539.105 1048.035 9539.385 1190.355 ;
      RECT 9538.545 1048.035 9538.825 1190.115 ;
      RECT 9511.945 1048.035 9512.225 1201.16 ;
      RECT 9511.385 1046.935 9511.665 1201.4 ;
      RECT 9510.825 1048.035 9511.105 1201.64 ;
      RECT 9510.265 1046.935 9510.545 1201.885 ;
      RECT 9509.705 1048.035 9509.985 1202.125 ;
      RECT 9509.145 1046.935 9509.425 1202.365 ;
      RECT 9508.585 1048.035 9508.865 1202.605 ;
      RECT 9508.025 1048.035 9508.305 1202.845 ;
      RECT 9507.465 1048.035 9507.745 1188.465 ;
      RECT 9506.905 1048.035 9507.185 1188.225 ;
      RECT 9506.345 1048.035 9506.625 1187.985 ;
      RECT 9505.785 1048.035 9506.065 1187.745 ;
      RECT 9505.225 1048.035 9505.505 1187.505 ;
      RECT 9504.665 1048.035 9504.945 1187.265 ;
      RECT 9504.105 1048.035 9504.385 1187.025 ;
      RECT 9503.545 1048.035 9503.825 1186.785 ;
      RECT 9502.985 1048.035 9503.265 1186.545 ;
      RECT 9502.425 1048.035 9502.705 1186.305 ;
      RECT 9501.865 1046.935 9502.145 1186.065 ;
      RECT 9501.305 1048.035 9501.585 1185.825 ;
      RECT 9500.745 1046.935 9501.025 1185.585 ;
      RECT 9500.185 1048.035 9500.465 1185.345 ;
      RECT 9486.185 1046.935 9486.465 1191.465 ;
      RECT 9485.625 1048.035 9485.905 1191.225 ;
      RECT 9485.065 1048.035 9485.345 1190.985 ;
      RECT 9484.505 1048.035 9484.785 1190.745 ;
      RECT 9483.945 1048.035 9484.225 1190.505 ;
      RECT 9483.385 1048.035 9483.665 1190.265 ;
      RECT 9482.825 1048.035 9483.105 1190.025 ;
      RECT 9482.265 1048.035 9482.545 1189.785 ;
      RECT 9481.705 1048.035 9481.985 1189.545 ;
      RECT 9481.145 1046.935 9481.425 1189.305 ;
      RECT 9480.585 1048.035 9480.865 1189.065 ;
      RECT 9480.025 1046.935 9480.305 1188.825 ;
      RECT 9479.465 1048.035 9479.745 1188.585 ;
      RECT 9478.905 1048.035 9479.185 1188.345 ;
      RECT 9478.345 1048.035 9478.625 1188.105 ;
      RECT 9477.785 1048.035 9478.065 1187.865 ;
      RECT 9477.225 1048.035 9477.505 1187.625 ;
      RECT 9476.665 1048.035 9476.945 1187.385 ;
      RECT 9476.105 1048.035 9476.385 1187.145 ;
      RECT 9475.545 1048.035 9475.825 1186.905 ;
      RECT 9474.985 1048.035 9475.265 1186.665 ;
      RECT 9474.425 1048.035 9474.705 1186.425 ;
      RECT 9473.865 1048.035 9474.145 1186.185 ;
      RECT 9434.665 1048.035 9434.945 1193.09 ;
      RECT 9434.105 1048.035 9434.385 1193.33 ;
      RECT 9433.545 1048.035 9433.825 1193.57 ;
      RECT 9432.985 1046.935 9433.265 1193.81 ;
      RECT 9432.425 1048.035 9432.705 1194.05 ;
      RECT 9431.865 1046.935 9432.145 1194.29 ;
      RECT 9431.305 1048.035 9431.585 1194.53 ;
      RECT 9430.745 1048.035 9431.025 1194.77 ;
      RECT 9430.185 1048.035 9430.465 1195.01 ;
      RECT 9429.625 1046.935 9429.905 1195.25 ;
      RECT 9429.065 1048.035 9429.345 1195.49 ;
      RECT 9428.505 1046.935 9428.785 1195.73 ;
      RECT 9427.945 1048.035 9428.225 1195.97 ;
      RECT 9427.385 1046.935 9427.665 1196.21 ;
      RECT 9426.825 1048.035 9427.105 1196.45 ;
      RECT 9426.265 1048.035 9426.545 1196.69 ;
      RECT 9425.705 1048.035 9425.985 1196.69 ;
      RECT 9425.145 1048.035 9425.425 1196.45 ;
      RECT 9424.585 1048.035 9424.865 1196.21 ;
      RECT 9424.025 1048.035 9424.305 1195.97 ;
      RECT 9423.465 1048.035 9423.745 1195.73 ;
      RECT 9422.905 1048.035 9423.185 1195.49 ;
      RECT 9422.345 1048.035 9422.625 1195.25 ;
      RECT 9421.785 1048.035 9422.065 1195.01 ;
      RECT 9421.225 1048.035 9421.505 1194.77 ;
      RECT 9412.265 1048.035 9412.545 1194.285 ;
      RECT 9411.705 1046.935 9411.985 1194.045 ;
      RECT 9411.145 1048.035 9411.425 1193.805 ;
      RECT 9410.585 1046.935 9410.865 1193.565 ;
      RECT 9410.025 1048.035 9410.305 1193.325 ;
      RECT 9409.465 1046.935 9409.745 1193.085 ;
      RECT 9408.905 1048.035 9409.185 1192.845 ;
      RECT 9408.345 1048.035 9408.625 1192.605 ;
      RECT 9407.785 1048.035 9408.065 1192.365 ;
      RECT 9407.225 1048.035 9407.505 1192.125 ;
      RECT 9406.665 1048.035 9406.945 1191.885 ;
      RECT 9406.105 1048.035 9406.385 1191.645 ;
      RECT 9405.545 1048.035 9405.825 1191.405 ;
      RECT 9404.985 1048.035 9405.265 1191.165 ;
      RECT 9402.465 1046.935 9402.745 1192.885 ;
      RECT 9401.905 1048.035 9402.185 1192.645 ;
      RECT 9401.345 1046.935 9401.625 1192.405 ;
      RECT 9400.785 1048.035 9401.065 1192.165 ;
      RECT 9400.225 1048.035 9400.505 1191.925 ;
      RECT 9399.665 1048.035 9399.945 1191.685 ;
      RECT 9399.105 1048.035 9399.385 1191.445 ;
      RECT 9398.545 1048.035 9398.825 1191.205 ;
      RECT 9372.505 1048.035 9372.785 1188.855 ;
      RECT 9371.945 1048.035 9372.225 1189.095 ;
      RECT 9371.385 1048.035 9371.665 1189.335 ;
      RECT 9370.825 1048.035 9371.105 1189.58 ;
      RECT 9370.265 1048.035 9370.545 1189.82 ;
      RECT 9369.705 1048.035 9369.985 1190.06 ;
      RECT 9369.145 1048.035 9369.425 1190.06 ;
      RECT 9368.585 1048.035 9368.865 1189.82 ;
      RECT 9368.025 1048.035 9368.305 1189.58 ;
      RECT 9367.465 1046.935 9367.745 1189.34 ;
      RECT 9366.905 1048.035 9367.185 1189.1 ;
      RECT 9366.345 1046.935 9366.625 1188.86 ;
      RECT 9365.785 1048.035 9366.065 1188.62 ;
      RECT 9365.225 1048.035 9365.505 1188.38 ;
      RECT 9364.665 1048.035 9364.945 1188.14 ;
      RECT 9364.105 1046.935 9364.385 1187.9 ;
      RECT 9363.545 1048.035 9363.825 1187.66 ;
      RECT 9362.985 1046.935 9363.265 1187.42 ;
      RECT 9362.425 1048.035 9362.705 1187.18 ;
      RECT 9361.865 1046.935 9362.145 1186.94 ;
      RECT 9361.305 1048.035 9361.585 1186.7 ;
      RECT 9360.745 1048.035 9361.025 1186.46 ;
      RECT 9360.185 1048.035 9360.465 1186.22 ;
      RECT 9359.625 1048.035 9359.905 1185.98 ;
      RECT 9346.185 1048.035 9346.465 1191.78 ;
      RECT 9345.625 1048.035 9345.905 1191.54 ;
      RECT 9345.065 1048.035 9345.345 1191.3 ;
      RECT 9344.505 1048.035 9344.785 1191.06 ;
      RECT 9343.945 1048.035 9344.225 1190.82 ;
      RECT 9343.385 1048.035 9343.665 1190.58 ;
      RECT 9342.825 1048.035 9343.105 1190.34 ;
      RECT 9342.265 1048.035 9342.545 1190.1 ;
      RECT 9341.705 1046.935 9341.985 1189.86 ;
      RECT 9341.145 1048.035 9341.425 1189.62 ;
      RECT 9340.585 1046.935 9340.865 1189.3 ;
      RECT 9340.025 1048.035 9340.305 1189.14 ;
      RECT 9339.465 1046.935 9339.745 1188.9 ;
      RECT 9338.905 1048.035 9339.185 1188.66 ;
      RECT 9338.345 1048.035 9338.625 1188.42 ;
      RECT 9337.785 1048.035 9338.065 1188.18 ;
      RECT 9337.225 1048.035 9337.505 1187.94 ;
      RECT 9336.665 1048.035 9336.945 1187.7 ;
      RECT 9336.105 1048.035 9336.385 1187.46 ;
      RECT 9335.545 1048.035 9335.825 1187.22 ;
      RECT 9334.985 1048.035 9335.265 1186.98 ;
      RECT 9334.425 1046.935 9334.705 1186.74 ;
      RECT 9333.865 1048.035 9334.145 1186.5 ;
      RECT 9333.305 1046.935 9333.585 1186.26 ;
      RECT 9294.105 1048.035 9294.385 1191.87 ;
      RECT 9293.545 1048.035 9293.825 1192.11 ;
      RECT 9292.985 1048.035 9293.265 1192.35 ;
      RECT 9292.425 1048.035 9292.705 1192.59 ;
      RECT 9291.865 1048.035 9292.145 1192.83 ;
      RECT 9291.305 1048.035 9291.585 1193.07 ;
      RECT 9290.745 1048.035 9291.025 1193.31 ;
      RECT 9290.185 1048.035 9290.465 1193.55 ;
      RECT 9289.625 1048.035 9289.905 1193.79 ;
      RECT 9289.065 1048.035 9289.345 1194.03 ;
      RECT 9288.505 1048.035 9288.785 1194.27 ;
      RECT 9287.945 1048.035 9288.225 1194.51 ;
      RECT 9287.385 1048.035 9287.665 1194.75 ;
      RECT 9286.825 1048.035 9287.105 1194.75 ;
      RECT 9286.265 1046.935 9286.545 1194.51 ;
      RECT 9285.705 1048.035 9285.985 1194.27 ;
      RECT 9285.145 1046.935 9285.425 1194.03 ;
      RECT 9284.585 1048.035 9284.865 1193.79 ;
      RECT 9284.025 1048.035 9284.305 1193.55 ;
      RECT 9283.465 1048.035 9283.745 1193.31 ;
      RECT 9282.905 1046.935 9283.185 1193.045 ;
      RECT 9282.345 1048.035 9282.625 1192.805 ;
      RECT 9281.785 1046.935 9282.065 1192.565 ;
      RECT 9281.225 1048.035 9281.505 1192.325 ;
      RECT 9272.265 1046.935 9272.545 1186.16 ;
      RECT 9271.705 1048.035 9271.985 1186.4 ;
      RECT 9271.145 1048.035 9271.425 1186.64 ;
      RECT 9270.585 1048.035 9270.865 1186.64 ;
      RECT 9270.025 1048.035 9270.305 1186.4 ;
      RECT 9269.465 1048.035 9269.745 1186.16 ;
      RECT 9268.905 1048.035 9269.185 1185.92 ;
      RECT 9268.345 1048.035 9268.625 1185.68 ;
      RECT 9267.785 1048.035 9268.065 1185.44 ;
      RECT 9267.225 1048.035 9267.505 1185.2 ;
      RECT 9266.665 1048.035 9266.945 1184.96 ;
      RECT 9266.105 1048.035 9266.385 1184.72 ;
      RECT 9265.545 1048.035 9265.825 1184.48 ;
      RECT 9264.985 1046.935 9265.265 1184.24 ;
      RECT 9262.465 1048.035 9262.745 1185.96 ;
      RECT 9261.905 1046.935 9262.185 1185.72 ;
      RECT 9261.345 1048.035 9261.625 1185.48 ;
      RECT 9260.785 1046.935 9261.065 1185.24 ;
      RECT 9260.225 1048.035 9260.505 1185 ;
      RECT 9259.665 1048.035 9259.945 1184.76 ;
      RECT 9259.105 1048.035 9259.385 1184.52 ;
      RECT 9233.065 1048.035 9233.345 1187.305 ;
      RECT 9232.505 1048.035 9232.785 1187.545 ;
      RECT 9231.945 1048.035 9232.225 1187.785 ;
      RECT 9231.385 1048.035 9231.665 1188.025 ;
      RECT 9230.825 1048.035 9231.105 1188.265 ;
      RECT 9230.265 1046.935 9230.545 1188.505 ;
      RECT 9229.705 1048.035 9229.985 1188.745 ;
      RECT 9229.145 1046.935 9229.425 1188.985 ;
      RECT 9228.585 1048.035 9228.865 1189.225 ;
      RECT 9228.025 1048.035 9228.305 1189.465 ;
      RECT 9227.465 1048.035 9227.745 1189.705 ;
      RECT 9226.905 1048.035 9227.185 1189.945 ;
      RECT 9226.345 1048.035 9226.625 1190.185 ;
      RECT 9225.785 1048.035 9226.065 1190.425 ;
      RECT 9225.225 1048.035 9225.505 1190.665 ;
      RECT 9224.665 1048.035 9224.945 1190.665 ;
      RECT 9224.105 1048.035 9224.385 1190.425 ;
      RECT 9223.545 1048.035 9223.825 1190.185 ;
      RECT 9222.985 1048.035 9223.265 1189.945 ;
      RECT 9222.425 1048.035 9222.705 1189.7 ;
      RECT 9221.865 1048.035 9222.145 1189.46 ;
      RECT 9221.305 1048.035 9221.585 1189.22 ;
      RECT 9220.745 1046.935 9221.025 1188.98 ;
      RECT 9220.185 1048.035 9220.465 1188.74 ;
      RECT 9206.745 1046.935 9207.025 1186.22 ;
      RECT 9206.185 1048.035 9206.465 1185.98 ;
      RECT 9205.625 1048.035 9205.905 1185.74 ;
      RECT 9205.065 1048.035 9205.345 1185.5 ;
      RECT 9204.505 1046.935 9204.785 1185.26 ;
      RECT 9203.945 1048.035 9204.225 1185.02 ;
      RECT 9203.385 1046.935 9203.665 1184.78 ;
      RECT 9202.825 1048.035 9203.105 1184.54 ;
      RECT 9202.265 1046.935 9202.545 1184.3 ;
      RECT 9201.705 1048.035 9201.985 1184.06 ;
      RECT 9201.145 1048.035 9201.425 1183.82 ;
      RECT 9200.585 1048.035 9200.865 1183.58 ;
      RECT 9200.025 1048.035 9200.305 1183.34 ;
      RECT 9199.465 1048.035 9199.745 1183.1 ;
      RECT 9198.905 1048.035 9199.185 1182.86 ;
      RECT 9198.345 1048.035 9198.625 1182.62 ;
      RECT 9197.785 1048.035 9198.065 1182.38 ;
      RECT 9197.225 1048.035 9197.505 1182.14 ;
      RECT 9196.665 1048.035 9196.945 1181.9 ;
      RECT 9196.105 1048.035 9196.385 1181.66 ;
      RECT 9195.545 1048.035 9195.825 1181.42 ;
      RECT 9194.985 1046.935 9195.265 1181.18 ;
      RECT 9194.425 1048.035 9194.705 1180.94 ;
      RECT 9193.865 1046.935 9194.145 1180.7 ;
      RECT 9154.105 1048.035 9154.385 1191.17 ;
      RECT 9153.545 1046.935 9153.825 1191.41 ;
      RECT 9152.985 1048.035 9153.265 1191.65 ;
      RECT 9152.425 1048.035 9152.705 1191.89 ;
      RECT 9151.865 1048.035 9152.145 1192.13 ;
      RECT 9151.305 1048.035 9151.585 1192.37 ;
      RECT 9150.745 1048.035 9151.025 1192.61 ;
      RECT 9150.185 1048.035 9150.465 1192.855 ;
      RECT 9149.625 1048.035 9149.905 1193.095 ;
      RECT 9149.065 1048.035 9149.345 1193.335 ;
      RECT 9148.505 1046.935 9148.785 1193.575 ;
      RECT 9147.945 1048.035 9148.225 1193.815 ;
      RECT 9147.385 1046.935 9147.665 1194.055 ;
      RECT 9146.825 1048.035 9147.105 1194.295 ;
      RECT 9146.265 1048.035 9146.545 1194.535 ;
      RECT 9145.705 1048.035 9145.985 1194.775 ;
      RECT 9145.145 1048.035 9145.425 1195.015 ;
      RECT 9144.585 1048.035 9144.865 1195.255 ;
      RECT 9144.025 1048.035 9144.305 1195.495 ;
      RECT 9143.465 1048.035 9143.745 1195.735 ;
      RECT 9142.905 1048.035 9143.185 1195.975 ;
      RECT 9142.345 1048.035 9142.625 1196.215 ;
      RECT 9141.785 1048.035 9142.065 1196.455 ;
      RECT 9141.225 1048.035 9141.505 1196.695 ;
      RECT 9132.265 1048.035 9132.545 1192.28 ;
      RECT 9131.705 1048.035 9131.985 1192.04 ;
      RECT 9131.145 1048.035 9131.425 1191.8 ;
      RECT 9130.585 1046.935 9130.865 1191.56 ;
      RECT 9130.025 1048.035 9130.305 1191.32 ;
      RECT 9129.465 1046.935 9129.745 1191.08 ;
      RECT 9128.905 1048.035 9129.185 1190.84 ;
      RECT 9128.345 1048.035 9128.625 1190.6 ;
      RECT 9127.785 1048.035 9128.065 1190.36 ;
      RECT 9127.225 1046.935 9127.505 1190.12 ;
      RECT 9126.665 1048.035 9126.945 1189.88 ;
      RECT 9126.105 1046.935 9126.385 1189.64 ;
      RECT 9125.545 1048.035 9125.825 1189.4 ;
      RECT 9124.985 1046.935 9125.265 1189.16 ;
      RECT 9122.465 1048.035 9122.745 1181.56 ;
      RECT 9121.905 1048.035 9122.185 1181.32 ;
      RECT 9121.345 1048.035 9121.625 1181.08 ;
      RECT 9120.785 1048.035 9121.065 1180.84 ;
      RECT 9120.225 1048.035 9120.505 1180.6 ;
      RECT 9119.665 1048.035 9119.945 1180.36 ;
      RECT 9119.105 1048.035 9119.385 1180.12 ;
      RECT 9093.065 1048.035 9093.345 1193.995 ;
      RECT 9092.505 1048.035 9092.785 1194.235 ;
      RECT 9091.945 1048.035 9092.225 1194.475 ;
      RECT 9091.385 1048.035 9091.665 1194.715 ;
      RECT 9090.825 1048.035 9091.105 1194.955 ;
      RECT 9090.265 1046.935 9090.545 1194.955 ;
      RECT 9089.705 1048.035 9089.985 1194.715 ;
      RECT 9089.145 1046.935 9089.425 1194.47 ;
      RECT 9088.585 1048.035 9088.865 1194.23 ;
      RECT 9088.025 1046.935 9088.305 1193.99 ;
      RECT 9087.465 1048.035 9087.745 1193.75 ;
      RECT 9086.905 1048.035 9087.185 1193.51 ;
      RECT 9086.345 1048.035 9086.625 1193.27 ;
      RECT 9085.785 1048.035 9086.065 1193.03 ;
      RECT 9085.225 1048.035 9085.505 1192.79 ;
      RECT 9084.665 1048.035 9084.945 1192.55 ;
      RECT 9084.105 1048.035 9084.385 1192.31 ;
      RECT 9083.545 1048.035 9083.825 1192.07 ;
      RECT 9082.985 1046.935 9083.265 1191.83 ;
      RECT 9082.425 1048.035 9082.705 1191.59 ;
      RECT 9081.865 1046.935 9082.145 1191.35 ;
      RECT 9081.305 1048.035 9081.585 1191.11 ;
      RECT 9080.745 1048.035 9081.025 1190.87 ;
      RECT 9080.185 1048.035 9080.465 1190.63 ;
      RECT 9066.745 1048.035 9067.025 1194.03 ;
      RECT 9066.185 1048.035 9066.465 1194.27 ;
      RECT 9065.625 1048.035 9065.905 1194.515 ;
      RECT 9065.065 1048.035 9065.345 1194.755 ;
      RECT 9064.505 1048.035 9064.785 1194.995 ;
      RECT 9063.945 1048.035 9064.225 1194.995 ;
      RECT 9063.385 1048.035 9063.665 1194.755 ;
      RECT 9062.825 1048.035 9063.105 1194.515 ;
      RECT 9062.265 1048.035 9062.545 1187.5 ;
      RECT 9061.705 1048.035 9061.985 1187.26 ;
      RECT 9061.145 1048.035 9061.425 1187.02 ;
      RECT 9060.585 1046.935 9060.865 1186.78 ;
      RECT 9060.025 1048.035 9060.305 1186.54 ;
      RECT 9059.465 1046.935 9059.745 1186.3 ;
      RECT 9058.905 1048.035 9059.185 1186.06 ;
      RECT 9058.345 1048.035 9058.625 1185.82 ;
      RECT 9057.785 1048.035 9058.065 1185.58 ;
      RECT 9057.225 1046.935 9057.505 1185.34 ;
      RECT 9056.665 1048.035 9056.945 1185.1 ;
      RECT 9056.105 1046.935 9056.385 1184.86 ;
      RECT 9055.545 1048.035 9055.825 1184.62 ;
      RECT 9054.985 1046.935 9055.265 1184.38 ;
      RECT 9054.425 1048.035 9054.705 1184.14 ;
      RECT 9053.865 1048.035 9054.145 1183.9 ;
      RECT 9013.545 1048.035 9013.825 1192.795 ;
      RECT 9012.985 1048.035 9013.265 1193.035 ;
      RECT 9012.425 1048.035 9012.705 1193.28 ;
      RECT 9011.865 1048.035 9012.145 1193.52 ;
      RECT 9011.305 1048.035 9011.585 1193.76 ;
      RECT 9010.745 1048.035 9011.025 1194 ;
      RECT 9010.185 1048.035 9010.465 1194.24 ;
      RECT 9009.625 1048.035 9009.905 1194.48 ;
      RECT 9009.065 1048.035 9009.345 1194.72 ;
      RECT 9008.505 1048.035 9008.785 1194.96 ;
      RECT 9007.945 1046.935 9008.225 1195.2 ;
      RECT 9007.385 1048.035 9007.665 1195.44 ;
      RECT 9006.825 1046.935 9007.105 1195.68 ;
      RECT 9006.265 1048.035 9006.545 1195.92 ;
      RECT 9005.705 1046.935 9005.985 1196.16 ;
      RECT 9005.145 1048.035 9005.425 1196.16 ;
      RECT 9004.585 1048.035 9004.865 1195.92 ;
      RECT 9004.025 1048.035 9004.305 1195.68 ;
      RECT 9003.465 1048.035 9003.745 1195.44 ;
      RECT 9002.905 1048.035 9003.185 1195.2 ;
      RECT 9002.345 1048.035 9002.625 1194.96 ;
      RECT 9001.785 1048.035 9002.065 1194.72 ;
      RECT 9001.225 1048.035 9001.505 1194.48 ;
      RECT 8992.265 1046.935 8992.545 1194.51 ;
      RECT 8991.705 1048.035 8991.985 1194.75 ;
      RECT 8991.145 1046.935 8991.425 1194.99 ;
      RECT 8990.585 1048.035 8990.865 1195.205 ;
      RECT 8990.025 1048.035 8990.305 1194.78 ;
      RECT 8989.465 1048.035 8989.745 1194.54 ;
      RECT 8988.905 1048.035 8989.185 1194.3 ;
      RECT 8988.345 1048.035 8988.625 1194.06 ;
      RECT 8987.785 1048.035 8988.065 1193.82 ;
      RECT 8987.225 1048.035 8987.505 1193.58 ;
      RECT 8986.665 1048.035 8986.945 1193.34 ;
      RECT 8986.105 1048.035 8986.385 1193.1 ;
      RECT 8985.545 1048.035 8985.825 1192.86 ;
      RECT 8984.985 1048.035 8985.265 1192.62 ;
      RECT 8982.465 1048.035 8982.745 1191.795 ;
      RECT 8981.905 1048.035 8982.185 1191.555 ;
      RECT 8981.345 1048.035 8981.625 1191.315 ;
      RECT 8980.785 1046.935 8981.065 1191.075 ;
      RECT 8980.225 1048.035 8980.505 1190.835 ;
      RECT 8979.665 1046.935 8979.945 1190.595 ;
      RECT 8979.105 1048.035 8979.385 1190.355 ;
      RECT 8978.545 1048.035 8978.825 1190.115 ;
      RECT 8951.945 1048.035 8952.225 1201.16 ;
      RECT 8951.385 1046.935 8951.665 1201.4 ;
      RECT 8950.825 1048.035 8951.105 1201.64 ;
      RECT 8950.265 1046.935 8950.545 1201.885 ;
      RECT 8949.705 1048.035 8949.985 1202.125 ;
      RECT 8949.145 1046.935 8949.425 1202.365 ;
      RECT 8948.585 1048.035 8948.865 1202.605 ;
      RECT 8948.025 1048.035 8948.305 1202.845 ;
      RECT 8947.465 1048.035 8947.745 1188.465 ;
      RECT 8946.905 1048.035 8947.185 1188.225 ;
      RECT 8946.345 1048.035 8946.625 1187.985 ;
      RECT 8945.785 1048.035 8946.065 1187.745 ;
      RECT 8945.225 1048.035 8945.505 1187.505 ;
      RECT 8944.665 1048.035 8944.945 1187.265 ;
      RECT 8944.105 1048.035 8944.385 1187.025 ;
      RECT 8943.545 1048.035 8943.825 1186.785 ;
      RECT 8942.985 1048.035 8943.265 1186.545 ;
      RECT 8942.425 1048.035 8942.705 1186.305 ;
      RECT 8941.865 1046.935 8942.145 1186.065 ;
      RECT 8941.305 1048.035 8941.585 1185.825 ;
      RECT 8940.745 1046.935 8941.025 1185.585 ;
      RECT 8940.185 1048.035 8940.465 1185.345 ;
      RECT 8926.185 1046.935 8926.465 1191.465 ;
      RECT 8925.625 1048.035 8925.905 1191.225 ;
      RECT 8925.065 1048.035 8925.345 1190.985 ;
      RECT 8924.505 1048.035 8924.785 1190.745 ;
      RECT 8923.945 1048.035 8924.225 1190.505 ;
      RECT 8923.385 1048.035 8923.665 1190.265 ;
      RECT 8922.825 1048.035 8923.105 1190.025 ;
      RECT 8922.265 1048.035 8922.545 1189.785 ;
      RECT 8921.705 1048.035 8921.985 1189.545 ;
      RECT 8921.145 1046.935 8921.425 1189.305 ;
      RECT 8920.585 1048.035 8920.865 1189.065 ;
      RECT 8920.025 1046.935 8920.305 1188.825 ;
      RECT 8919.465 1048.035 8919.745 1188.585 ;
      RECT 8918.905 1048.035 8919.185 1188.345 ;
      RECT 8918.345 1048.035 8918.625 1188.105 ;
      RECT 8917.785 1048.035 8918.065 1187.865 ;
      RECT 8917.225 1048.035 8917.505 1187.625 ;
      RECT 8916.665 1048.035 8916.945 1187.385 ;
      RECT 8916.105 1048.035 8916.385 1187.145 ;
      RECT 8915.545 1048.035 8915.825 1186.905 ;
      RECT 8914.985 1048.035 8915.265 1186.665 ;
      RECT 8914.425 1048.035 8914.705 1186.425 ;
      RECT 8913.865 1048.035 8914.145 1186.185 ;
      RECT 8874.665 1048.035 8874.945 1193.09 ;
      RECT 8874.105 1048.035 8874.385 1193.33 ;
      RECT 8873.545 1048.035 8873.825 1193.57 ;
      RECT 8872.985 1046.935 8873.265 1193.81 ;
      RECT 8872.425 1048.035 8872.705 1194.05 ;
      RECT 8871.865 1046.935 8872.145 1194.29 ;
      RECT 8871.305 1048.035 8871.585 1194.53 ;
      RECT 8870.745 1048.035 8871.025 1194.77 ;
      RECT 8870.185 1048.035 8870.465 1195.01 ;
      RECT 8869.625 1046.935 8869.905 1195.25 ;
      RECT 8869.065 1048.035 8869.345 1195.49 ;
      RECT 8868.505 1046.935 8868.785 1195.73 ;
      RECT 8867.945 1048.035 8868.225 1195.97 ;
      RECT 8867.385 1046.935 8867.665 1196.21 ;
      RECT 8866.825 1048.035 8867.105 1196.45 ;
      RECT 8866.265 1048.035 8866.545 1196.69 ;
      RECT 8865.705 1048.035 8865.985 1196.69 ;
      RECT 8865.145 1048.035 8865.425 1196.45 ;
      RECT 8864.585 1048.035 8864.865 1196.21 ;
      RECT 8864.025 1048.035 8864.305 1195.97 ;
      RECT 8863.465 1048.035 8863.745 1195.73 ;
      RECT 8862.905 1048.035 8863.185 1195.49 ;
      RECT 8862.345 1048.035 8862.625 1195.25 ;
      RECT 8861.785 1048.035 8862.065 1195.01 ;
      RECT 8861.225 1048.035 8861.505 1194.77 ;
      RECT 8852.265 1048.035 8852.545 1194.285 ;
      RECT 8851.705 1046.935 8851.985 1194.045 ;
      RECT 8851.145 1048.035 8851.425 1193.805 ;
      RECT 8850.585 1046.935 8850.865 1193.565 ;
      RECT 8850.025 1048.035 8850.305 1193.325 ;
      RECT 8849.465 1046.935 8849.745 1193.085 ;
      RECT 8848.905 1048.035 8849.185 1192.845 ;
      RECT 8848.345 1048.035 8848.625 1192.605 ;
      RECT 8847.785 1048.035 8848.065 1192.365 ;
      RECT 8847.225 1048.035 8847.505 1192.125 ;
      RECT 8846.665 1048.035 8846.945 1191.885 ;
      RECT 8846.105 1048.035 8846.385 1191.645 ;
      RECT 8845.545 1048.035 8845.825 1191.405 ;
      RECT 8844.985 1048.035 8845.265 1191.165 ;
      RECT 8842.465 1046.935 8842.745 1192.885 ;
      RECT 8841.905 1048.035 8842.185 1192.645 ;
      RECT 8841.345 1046.935 8841.625 1192.405 ;
      RECT 8840.785 1048.035 8841.065 1192.165 ;
      RECT 8840.225 1048.035 8840.505 1191.925 ;
      RECT 8839.665 1048.035 8839.945 1191.685 ;
      RECT 8839.105 1048.035 8839.385 1191.445 ;
      RECT 8838.545 1048.035 8838.825 1191.205 ;
      RECT 8812.505 1048.035 8812.785 1188.855 ;
      RECT 8811.945 1048.035 8812.225 1189.095 ;
      RECT 8811.385 1048.035 8811.665 1189.335 ;
      RECT 8810.825 1048.035 8811.105 1189.58 ;
      RECT 8810.265 1048.035 8810.545 1189.82 ;
      RECT 8809.705 1048.035 8809.985 1190.06 ;
      RECT 8809.145 1048.035 8809.425 1190.06 ;
      RECT 8808.585 1048.035 8808.865 1189.82 ;
      RECT 8808.025 1048.035 8808.305 1189.58 ;
      RECT 8807.465 1046.935 8807.745 1189.34 ;
      RECT 8806.905 1048.035 8807.185 1189.1 ;
      RECT 8806.345 1046.935 8806.625 1188.86 ;
      RECT 8805.785 1048.035 8806.065 1188.62 ;
      RECT 8805.225 1048.035 8805.505 1188.38 ;
      RECT 8804.665 1048.035 8804.945 1188.14 ;
      RECT 8804.105 1046.935 8804.385 1187.9 ;
      RECT 8803.545 1048.035 8803.825 1187.66 ;
      RECT 8802.985 1046.935 8803.265 1187.42 ;
      RECT 8802.425 1048.035 8802.705 1187.18 ;
      RECT 8801.865 1046.935 8802.145 1186.94 ;
      RECT 8801.305 1048.035 8801.585 1186.7 ;
      RECT 8800.745 1048.035 8801.025 1186.46 ;
      RECT 8800.185 1048.035 8800.465 1186.22 ;
      RECT 8799.625 1048.035 8799.905 1185.98 ;
      RECT 8786.185 1048.035 8786.465 1191.78 ;
      RECT 8785.625 1048.035 8785.905 1191.54 ;
      RECT 8785.065 1048.035 8785.345 1191.3 ;
      RECT 8784.505 1048.035 8784.785 1191.06 ;
      RECT 8783.945 1048.035 8784.225 1190.82 ;
      RECT 8783.385 1048.035 8783.665 1190.58 ;
      RECT 8782.825 1048.035 8783.105 1190.34 ;
      RECT 8782.265 1048.035 8782.545 1190.1 ;
      RECT 8781.705 1046.935 8781.985 1189.86 ;
      RECT 8781.145 1048.035 8781.425 1189.62 ;
      RECT 8780.585 1046.935 8780.865 1189.3 ;
      RECT 8780.025 1048.035 8780.305 1189.14 ;
      RECT 8779.465 1046.935 8779.745 1188.9 ;
      RECT 8778.905 1048.035 8779.185 1188.66 ;
      RECT 8778.345 1048.035 8778.625 1188.42 ;
      RECT 8777.785 1048.035 8778.065 1188.18 ;
      RECT 8777.225 1048.035 8777.505 1187.94 ;
      RECT 8776.665 1048.035 8776.945 1187.7 ;
      RECT 8776.105 1048.035 8776.385 1187.46 ;
      RECT 8775.545 1048.035 8775.825 1187.22 ;
      RECT 8774.985 1048.035 8775.265 1186.98 ;
      RECT 8774.425 1046.935 8774.705 1186.74 ;
      RECT 8773.865 1048.035 8774.145 1186.5 ;
      RECT 8773.305 1046.935 8773.585 1186.26 ;
      RECT 8734.105 1048.035 8734.385 1191.87 ;
      RECT 8733.545 1048.035 8733.825 1192.11 ;
      RECT 8732.985 1048.035 8733.265 1192.35 ;
      RECT 8732.425 1048.035 8732.705 1192.59 ;
      RECT 8731.865 1048.035 8732.145 1192.83 ;
      RECT 8731.305 1048.035 8731.585 1193.07 ;
      RECT 8730.745 1048.035 8731.025 1193.31 ;
      RECT 8730.185 1048.035 8730.465 1193.55 ;
      RECT 8729.625 1048.035 8729.905 1193.79 ;
      RECT 8729.065 1048.035 8729.345 1194.03 ;
      RECT 8728.505 1048.035 8728.785 1194.27 ;
      RECT 8727.945 1048.035 8728.225 1194.51 ;
      RECT 8727.385 1048.035 8727.665 1194.75 ;
      RECT 8726.825 1048.035 8727.105 1194.75 ;
      RECT 8726.265 1046.935 8726.545 1194.51 ;
      RECT 8725.705 1048.035 8725.985 1194.27 ;
      RECT 8725.145 1046.935 8725.425 1194.03 ;
      RECT 8724.585 1048.035 8724.865 1193.79 ;
      RECT 8724.025 1048.035 8724.305 1193.55 ;
      RECT 8723.465 1048.035 8723.745 1193.31 ;
      RECT 8722.905 1046.935 8723.185 1193.045 ;
      RECT 8722.345 1048.035 8722.625 1192.805 ;
      RECT 8721.785 1046.935 8722.065 1192.565 ;
      RECT 8721.225 1048.035 8721.505 1192.325 ;
      RECT 8712.265 1046.935 8712.545 1186.16 ;
      RECT 8711.705 1048.035 8711.985 1186.4 ;
      RECT 8711.145 1048.035 8711.425 1186.64 ;
      RECT 8710.585 1048.035 8710.865 1186.64 ;
      RECT 8710.025 1048.035 8710.305 1186.4 ;
      RECT 8709.465 1048.035 8709.745 1186.16 ;
      RECT 8708.905 1048.035 8709.185 1185.92 ;
      RECT 8708.345 1048.035 8708.625 1185.68 ;
      RECT 8707.785 1048.035 8708.065 1185.44 ;
      RECT 8707.225 1048.035 8707.505 1185.2 ;
      RECT 8706.665 1048.035 8706.945 1184.96 ;
      RECT 8706.105 1048.035 8706.385 1184.72 ;
      RECT 8705.545 1048.035 8705.825 1184.48 ;
      RECT 8704.985 1046.935 8705.265 1184.24 ;
      RECT 8702.465 1048.035 8702.745 1185.96 ;
      RECT 8701.905 1046.935 8702.185 1185.72 ;
      RECT 8701.345 1048.035 8701.625 1185.48 ;
      RECT 8700.785 1046.935 8701.065 1185.24 ;
      RECT 8700.225 1048.035 8700.505 1185 ;
      RECT 8699.665 1048.035 8699.945 1184.76 ;
      RECT 8699.105 1048.035 8699.385 1184.52 ;
      RECT 8673.065 1048.035 8673.345 1187.305 ;
      RECT 8672.505 1048.035 8672.785 1187.545 ;
      RECT 8671.945 1048.035 8672.225 1187.785 ;
      RECT 8671.385 1048.035 8671.665 1188.025 ;
      RECT 8670.825 1048.035 8671.105 1188.265 ;
      RECT 8670.265 1046.935 8670.545 1188.505 ;
      RECT 8669.705 1048.035 8669.985 1188.745 ;
      RECT 8669.145 1046.935 8669.425 1188.985 ;
      RECT 8668.585 1048.035 8668.865 1189.225 ;
      RECT 8668.025 1048.035 8668.305 1189.465 ;
      RECT 8667.465 1048.035 8667.745 1189.705 ;
      RECT 8666.905 1048.035 8667.185 1189.945 ;
      RECT 8666.345 1048.035 8666.625 1190.185 ;
      RECT 8665.785 1048.035 8666.065 1190.425 ;
      RECT 8665.225 1048.035 8665.505 1190.665 ;
      RECT 8664.665 1048.035 8664.945 1190.665 ;
      RECT 8664.105 1048.035 8664.385 1190.425 ;
      RECT 8663.545 1048.035 8663.825 1190.185 ;
      RECT 8662.985 1048.035 8663.265 1189.945 ;
      RECT 8662.425 1048.035 8662.705 1189.7 ;
      RECT 8661.865 1048.035 8662.145 1189.46 ;
      RECT 8661.305 1048.035 8661.585 1189.22 ;
      RECT 8660.745 1046.935 8661.025 1188.98 ;
      RECT 8660.185 1048.035 8660.465 1188.74 ;
      RECT 8646.745 1046.935 8647.025 1186.22 ;
      RECT 8646.185 1048.035 8646.465 1185.98 ;
      RECT 8645.625 1048.035 8645.905 1185.74 ;
      RECT 8645.065 1048.035 8645.345 1185.5 ;
      RECT 8644.505 1046.935 8644.785 1185.26 ;
      RECT 8643.945 1048.035 8644.225 1185.02 ;
      RECT 8643.385 1046.935 8643.665 1184.78 ;
      RECT 8642.825 1048.035 8643.105 1184.54 ;
      RECT 8642.265 1046.935 8642.545 1184.3 ;
      RECT 8641.705 1048.035 8641.985 1184.06 ;
      RECT 8641.145 1048.035 8641.425 1183.82 ;
      RECT 8640.585 1048.035 8640.865 1183.58 ;
      RECT 8640.025 1048.035 8640.305 1183.34 ;
      RECT 8639.465 1048.035 8639.745 1183.1 ;
      RECT 8638.905 1048.035 8639.185 1182.86 ;
      RECT 8638.345 1048.035 8638.625 1182.62 ;
      RECT 8637.785 1048.035 8638.065 1182.38 ;
      RECT 8637.225 1048.035 8637.505 1182.14 ;
      RECT 8636.665 1048.035 8636.945 1181.9 ;
      RECT 8636.105 1048.035 8636.385 1181.66 ;
      RECT 8635.545 1048.035 8635.825 1181.42 ;
      RECT 8634.985 1046.935 8635.265 1181.18 ;
      RECT 8634.425 1048.035 8634.705 1180.94 ;
      RECT 8633.865 1046.935 8634.145 1180.7 ;
      RECT 8594.105 1048.035 8594.385 1191.17 ;
      RECT 8593.545 1046.935 8593.825 1191.41 ;
      RECT 8592.985 1048.035 8593.265 1191.65 ;
      RECT 8592.425 1048.035 8592.705 1191.89 ;
      RECT 8591.865 1048.035 8592.145 1192.13 ;
      RECT 8591.305 1048.035 8591.585 1192.37 ;
      RECT 8590.745 1048.035 8591.025 1192.61 ;
      RECT 8590.185 1048.035 8590.465 1192.855 ;
      RECT 8589.625 1048.035 8589.905 1193.095 ;
      RECT 8589.065 1048.035 8589.345 1193.335 ;
      RECT 8588.505 1046.935 8588.785 1193.575 ;
      RECT 8587.945 1048.035 8588.225 1193.815 ;
      RECT 8587.385 1046.935 8587.665 1194.055 ;
      RECT 8586.825 1048.035 8587.105 1194.295 ;
      RECT 8586.265 1048.035 8586.545 1194.535 ;
      RECT 8585.705 1048.035 8585.985 1194.775 ;
      RECT 8585.145 1048.035 8585.425 1195.015 ;
      RECT 8584.585 1048.035 8584.865 1195.255 ;
      RECT 8584.025 1048.035 8584.305 1195.495 ;
      RECT 8583.465 1048.035 8583.745 1195.735 ;
      RECT 8582.905 1048.035 8583.185 1195.975 ;
      RECT 8582.345 1048.035 8582.625 1196.215 ;
      RECT 8581.785 1048.035 8582.065 1196.455 ;
      RECT 8581.225 1048.035 8581.505 1196.695 ;
      RECT 8572.265 1048.035 8572.545 1192.28 ;
      RECT 8571.705 1048.035 8571.985 1192.04 ;
      RECT 8571.145 1048.035 8571.425 1191.8 ;
      RECT 8570.585 1046.935 8570.865 1191.56 ;
      RECT 8570.025 1048.035 8570.305 1191.32 ;
      RECT 8569.465 1046.935 8569.745 1191.08 ;
      RECT 8568.905 1048.035 8569.185 1190.84 ;
      RECT 8568.345 1048.035 8568.625 1190.6 ;
      RECT 8567.785 1048.035 8568.065 1190.36 ;
      RECT 8567.225 1046.935 8567.505 1190.12 ;
      RECT 8566.665 1048.035 8566.945 1189.88 ;
      RECT 8566.105 1046.935 8566.385 1189.64 ;
      RECT 8565.545 1048.035 8565.825 1189.4 ;
      RECT 8564.985 1046.935 8565.265 1189.16 ;
      RECT 8562.465 1048.035 8562.745 1181.56 ;
      RECT 8561.905 1048.035 8562.185 1181.32 ;
      RECT 8561.345 1048.035 8561.625 1181.08 ;
      RECT 8560.785 1048.035 8561.065 1180.84 ;
      RECT 8560.225 1048.035 8560.505 1180.6 ;
      RECT 8559.665 1048.035 8559.945 1180.36 ;
      RECT 8559.105 1048.035 8559.385 1180.12 ;
      RECT 8533.065 1048.035 8533.345 1193.995 ;
      RECT 8532.505 1048.035 8532.785 1194.235 ;
      RECT 8531.945 1048.035 8532.225 1194.475 ;
      RECT 8531.385 1048.035 8531.665 1194.715 ;
      RECT 8530.825 1048.035 8531.105 1194.955 ;
      RECT 8530.265 1046.935 8530.545 1194.955 ;
      RECT 8529.705 1048.035 8529.985 1194.715 ;
      RECT 8529.145 1046.935 8529.425 1194.47 ;
      RECT 8528.585 1048.035 8528.865 1194.23 ;
      RECT 8528.025 1046.935 8528.305 1193.99 ;
      RECT 8527.465 1048.035 8527.745 1193.75 ;
      RECT 8526.905 1048.035 8527.185 1193.51 ;
      RECT 8526.345 1048.035 8526.625 1193.27 ;
      RECT 8525.785 1048.035 8526.065 1193.03 ;
      RECT 8525.225 1048.035 8525.505 1192.79 ;
      RECT 8524.665 1048.035 8524.945 1192.55 ;
      RECT 8524.105 1048.035 8524.385 1192.31 ;
      RECT 8523.545 1048.035 8523.825 1192.07 ;
      RECT 8522.985 1046.935 8523.265 1191.83 ;
      RECT 8522.425 1048.035 8522.705 1191.59 ;
      RECT 8521.865 1046.935 8522.145 1191.35 ;
      RECT 8521.305 1048.035 8521.585 1191.11 ;
      RECT 8520.745 1048.035 8521.025 1190.87 ;
      RECT 8520.185 1048.035 8520.465 1190.63 ;
      RECT 8506.745 1048.035 8507.025 1194.03 ;
      RECT 8506.185 1048.035 8506.465 1194.27 ;
      RECT 8505.625 1048.035 8505.905 1194.515 ;
      RECT 8505.065 1048.035 8505.345 1194.755 ;
      RECT 8504.505 1048.035 8504.785 1194.995 ;
      RECT 8503.945 1048.035 8504.225 1194.995 ;
      RECT 8503.385 1048.035 8503.665 1194.755 ;
      RECT 8502.825 1048.035 8503.105 1194.515 ;
      RECT 8502.265 1048.035 8502.545 1187.5 ;
      RECT 8501.705 1048.035 8501.985 1187.26 ;
      RECT 8501.145 1048.035 8501.425 1187.02 ;
      RECT 8500.585 1046.935 8500.865 1186.78 ;
      RECT 8500.025 1048.035 8500.305 1186.54 ;
      RECT 8499.465 1046.935 8499.745 1186.3 ;
      RECT 8498.905 1048.035 8499.185 1186.06 ;
      RECT 8498.345 1048.035 8498.625 1185.82 ;
      RECT 8497.785 1048.035 8498.065 1185.58 ;
      RECT 8497.225 1046.935 8497.505 1185.34 ;
      RECT 8496.665 1048.035 8496.945 1185.1 ;
      RECT 8496.105 1046.935 8496.385 1184.86 ;
      RECT 8495.545 1048.035 8495.825 1184.62 ;
      RECT 8494.985 1046.935 8495.265 1184.38 ;
      RECT 8494.425 1048.035 8494.705 1184.14 ;
      RECT 8493.865 1048.035 8494.145 1183.9 ;
      RECT 8453.545 1048.035 8453.825 1192.795 ;
      RECT 8452.985 1048.035 8453.265 1193.035 ;
      RECT 8452.425 1048.035 8452.705 1193.28 ;
      RECT 8451.865 1048.035 8452.145 1193.52 ;
      RECT 8451.305 1048.035 8451.585 1193.76 ;
      RECT 8450.745 1048.035 8451.025 1194 ;
      RECT 8450.185 1048.035 8450.465 1194.24 ;
      RECT 8449.625 1048.035 8449.905 1194.48 ;
      RECT 8449.065 1048.035 8449.345 1194.72 ;
      RECT 8448.505 1048.035 8448.785 1194.96 ;
      RECT 8447.945 1046.935 8448.225 1195.2 ;
      RECT 8447.385 1048.035 8447.665 1195.44 ;
      RECT 8446.825 1046.935 8447.105 1195.68 ;
      RECT 8446.265 1048.035 8446.545 1195.92 ;
      RECT 8445.705 1046.935 8445.985 1196.16 ;
      RECT 8445.145 1048.035 8445.425 1196.16 ;
      RECT 8444.585 1048.035 8444.865 1195.92 ;
      RECT 8444.025 1048.035 8444.305 1195.68 ;
      RECT 8443.465 1048.035 8443.745 1195.44 ;
      RECT 8442.905 1048.035 8443.185 1195.2 ;
      RECT 8442.345 1048.035 8442.625 1194.96 ;
      RECT 8441.785 1048.035 8442.065 1194.72 ;
      RECT 8441.225 1048.035 8441.505 1194.48 ;
      RECT 8432.265 1046.935 8432.545 1194.51 ;
      RECT 8431.705 1048.035 8431.985 1194.75 ;
      RECT 8431.145 1046.935 8431.425 1194.99 ;
      RECT 8430.585 1048.035 8430.865 1195.205 ;
      RECT 8430.025 1048.035 8430.305 1194.78 ;
      RECT 8429.465 1048.035 8429.745 1194.54 ;
      RECT 8428.905 1048.035 8429.185 1194.3 ;
      RECT 8428.345 1048.035 8428.625 1194.06 ;
      RECT 8427.785 1048.035 8428.065 1193.82 ;
      RECT 8427.225 1048.035 8427.505 1193.58 ;
      RECT 8426.665 1048.035 8426.945 1193.34 ;
      RECT 8426.105 1048.035 8426.385 1193.1 ;
      RECT 8425.545 1048.035 8425.825 1192.86 ;
      RECT 8424.985 1048.035 8425.265 1192.62 ;
      RECT 8422.465 1048.035 8422.745 1191.795 ;
      RECT 8421.905 1048.035 8422.185 1191.555 ;
      RECT 8421.345 1048.035 8421.625 1191.315 ;
      RECT 8420.785 1046.935 8421.065 1191.075 ;
      RECT 8420.225 1048.035 8420.505 1190.835 ;
      RECT 8419.665 1046.935 8419.945 1190.595 ;
      RECT 8419.105 1048.035 8419.385 1190.355 ;
      RECT 8418.545 1048.035 8418.825 1190.115 ;
      RECT 8391.945 1048.035 8392.225 1201.16 ;
      RECT 8391.385 1046.935 8391.665 1201.4 ;
      RECT 8390.825 1048.035 8391.105 1201.64 ;
      RECT 8390.265 1046.935 8390.545 1201.885 ;
      RECT 8389.705 1048.035 8389.985 1202.125 ;
      RECT 8389.145 1046.935 8389.425 1202.365 ;
      RECT 8388.585 1048.035 8388.865 1202.605 ;
      RECT 8388.025 1048.035 8388.305 1202.845 ;
      RECT 8387.465 1048.035 8387.745 1188.465 ;
      RECT 8386.905 1048.035 8387.185 1188.225 ;
      RECT 8386.345 1048.035 8386.625 1187.985 ;
      RECT 8385.785 1048.035 8386.065 1187.745 ;
      RECT 8385.225 1048.035 8385.505 1187.505 ;
      RECT 8384.665 1048.035 8384.945 1187.265 ;
      RECT 8384.105 1048.035 8384.385 1187.025 ;
      RECT 8383.545 1048.035 8383.825 1186.785 ;
      RECT 8382.985 1048.035 8383.265 1186.545 ;
      RECT 8382.425 1048.035 8382.705 1186.305 ;
      RECT 8381.865 1046.935 8382.145 1186.065 ;
      RECT 8381.305 1048.035 8381.585 1185.825 ;
      RECT 8380.745 1046.935 8381.025 1185.585 ;
      RECT 8380.185 1048.035 8380.465 1185.345 ;
      RECT 8366.185 1046.935 8366.465 1191.465 ;
      RECT 8365.625 1048.035 8365.905 1191.225 ;
      RECT 8365.065 1048.035 8365.345 1190.985 ;
      RECT 8364.505 1048.035 8364.785 1190.745 ;
      RECT 8363.945 1048.035 8364.225 1190.505 ;
      RECT 8363.385 1048.035 8363.665 1190.265 ;
      RECT 8362.825 1048.035 8363.105 1190.025 ;
      RECT 8362.265 1048.035 8362.545 1189.785 ;
      RECT 8361.705 1048.035 8361.985 1189.545 ;
      RECT 8361.145 1046.935 8361.425 1189.305 ;
      RECT 8360.585 1048.035 8360.865 1189.065 ;
      RECT 8360.025 1046.935 8360.305 1188.825 ;
      RECT 8359.465 1048.035 8359.745 1188.585 ;
      RECT 8358.905 1048.035 8359.185 1188.345 ;
      RECT 8358.345 1048.035 8358.625 1188.105 ;
      RECT 8357.785 1048.035 8358.065 1187.865 ;
      RECT 8357.225 1048.035 8357.505 1187.625 ;
      RECT 8356.665 1048.035 8356.945 1187.385 ;
      RECT 8356.105 1048.035 8356.385 1187.145 ;
      RECT 8355.545 1048.035 8355.825 1186.905 ;
      RECT 8354.985 1048.035 8355.265 1186.665 ;
      RECT 8354.425 1048.035 8354.705 1186.425 ;
      RECT 8353.865 1048.035 8354.145 1186.185 ;
      RECT 8314.665 1048.035 8314.945 1193.09 ;
      RECT 8314.105 1048.035 8314.385 1193.33 ;
      RECT 8313.545 1048.035 8313.825 1193.57 ;
      RECT 8312.985 1046.935 8313.265 1193.81 ;
      RECT 8312.425 1048.035 8312.705 1194.05 ;
      RECT 8311.865 1046.935 8312.145 1194.29 ;
      RECT 8311.305 1048.035 8311.585 1194.53 ;
      RECT 8310.745 1048.035 8311.025 1194.77 ;
      RECT 8310.185 1048.035 8310.465 1195.01 ;
      RECT 8309.625 1046.935 8309.905 1195.25 ;
      RECT 8309.065 1048.035 8309.345 1195.49 ;
      RECT 8308.505 1046.935 8308.785 1195.73 ;
      RECT 8307.945 1048.035 8308.225 1195.97 ;
      RECT 8307.385 1046.935 8307.665 1196.21 ;
      RECT 8306.825 1048.035 8307.105 1196.45 ;
      RECT 8306.265 1048.035 8306.545 1196.69 ;
      RECT 8305.705 1048.035 8305.985 1196.69 ;
      RECT 8305.145 1048.035 8305.425 1196.45 ;
      RECT 8304.585 1048.035 8304.865 1196.21 ;
      RECT 8304.025 1048.035 8304.305 1195.97 ;
      RECT 8303.465 1048.035 8303.745 1195.73 ;
      RECT 8302.905 1048.035 8303.185 1195.49 ;
      RECT 8302.345 1048.035 8302.625 1195.25 ;
      RECT 8301.785 1048.035 8302.065 1195.01 ;
      RECT 8301.225 1048.035 8301.505 1194.77 ;
      RECT 8292.265 1048.035 8292.545 1194.285 ;
      RECT 8291.705 1046.935 8291.985 1194.045 ;
      RECT 8291.145 1048.035 8291.425 1193.805 ;
      RECT 8290.585 1046.935 8290.865 1193.565 ;
      RECT 8290.025 1048.035 8290.305 1193.325 ;
      RECT 8289.465 1046.935 8289.745 1193.085 ;
      RECT 8288.905 1048.035 8289.185 1192.845 ;
      RECT 8288.345 1048.035 8288.625 1192.605 ;
      RECT 8287.785 1048.035 8288.065 1192.365 ;
      RECT 8287.225 1048.035 8287.505 1192.125 ;
      RECT 8286.665 1048.035 8286.945 1191.885 ;
      RECT 8286.105 1048.035 8286.385 1191.645 ;
      RECT 8285.545 1048.035 8285.825 1191.405 ;
      RECT 8284.985 1048.035 8285.265 1191.165 ;
      RECT 8282.465 1046.935 8282.745 1192.885 ;
      RECT 8281.905 1048.035 8282.185 1192.645 ;
      RECT 8281.345 1046.935 8281.625 1192.405 ;
      RECT 8280.785 1048.035 8281.065 1192.165 ;
      RECT 8280.225 1048.035 8280.505 1191.925 ;
      RECT 8279.665 1048.035 8279.945 1191.685 ;
      RECT 8279.105 1048.035 8279.385 1191.445 ;
      RECT 8278.545 1048.035 8278.825 1191.205 ;
      RECT 8252.505 1048.035 8252.785 1188.855 ;
      RECT 8251.945 1048.035 8252.225 1189.095 ;
      RECT 8251.385 1048.035 8251.665 1189.335 ;
      RECT 8250.825 1048.035 8251.105 1189.58 ;
      RECT 8250.265 1048.035 8250.545 1189.82 ;
      RECT 8249.705 1048.035 8249.985 1190.06 ;
      RECT 8249.145 1048.035 8249.425 1190.06 ;
      RECT 8248.585 1048.035 8248.865 1189.82 ;
      RECT 8248.025 1048.035 8248.305 1189.58 ;
      RECT 8247.465 1046.935 8247.745 1189.34 ;
      RECT 8246.905 1048.035 8247.185 1189.1 ;
      RECT 8246.345 1046.935 8246.625 1188.86 ;
      RECT 8245.785 1048.035 8246.065 1188.62 ;
      RECT 8245.225 1048.035 8245.505 1188.38 ;
      RECT 8244.665 1048.035 8244.945 1188.14 ;
      RECT 8244.105 1046.935 8244.385 1187.9 ;
      RECT 8243.545 1048.035 8243.825 1187.66 ;
      RECT 8242.985 1046.935 8243.265 1187.42 ;
      RECT 8242.425 1048.035 8242.705 1187.18 ;
      RECT 8241.865 1046.935 8242.145 1186.94 ;
      RECT 8241.305 1048.035 8241.585 1186.7 ;
      RECT 8240.745 1048.035 8241.025 1186.46 ;
      RECT 8240.185 1048.035 8240.465 1186.22 ;
      RECT 8239.625 1048.035 8239.905 1185.98 ;
      RECT 8226.185 1048.035 8226.465 1191.78 ;
      RECT 8225.625 1048.035 8225.905 1191.54 ;
      RECT 8225.065 1048.035 8225.345 1191.3 ;
      RECT 8224.505 1048.035 8224.785 1191.06 ;
      RECT 8223.945 1048.035 8224.225 1190.82 ;
      RECT 8223.385 1048.035 8223.665 1190.58 ;
      RECT 8222.825 1048.035 8223.105 1190.34 ;
      RECT 8222.265 1048.035 8222.545 1190.1 ;
      RECT 8221.705 1046.935 8221.985 1189.86 ;
      RECT 8221.145 1048.035 8221.425 1189.62 ;
      RECT 8220.585 1046.935 8220.865 1189.3 ;
      RECT 8220.025 1048.035 8220.305 1189.14 ;
      RECT 8219.465 1046.935 8219.745 1188.9 ;
      RECT 8218.905 1048.035 8219.185 1188.66 ;
      RECT 8218.345 1048.035 8218.625 1188.42 ;
      RECT 8217.785 1048.035 8218.065 1188.18 ;
      RECT 8217.225 1048.035 8217.505 1187.94 ;
      RECT 8216.665 1048.035 8216.945 1187.7 ;
      RECT 8216.105 1048.035 8216.385 1187.46 ;
      RECT 8215.545 1048.035 8215.825 1187.22 ;
      RECT 8214.985 1048.035 8215.265 1186.98 ;
      RECT 8214.425 1046.935 8214.705 1186.74 ;
      RECT 8213.865 1048.035 8214.145 1186.5 ;
      RECT 8213.305 1046.935 8213.585 1186.26 ;
      RECT 8174.105 1048.035 8174.385 1191.87 ;
      RECT 8173.545 1048.035 8173.825 1192.11 ;
      RECT 8172.985 1048.035 8173.265 1192.35 ;
      RECT 8172.425 1048.035 8172.705 1192.59 ;
      RECT 8171.865 1048.035 8172.145 1192.83 ;
      RECT 8171.305 1048.035 8171.585 1193.07 ;
      RECT 8170.745 1048.035 8171.025 1193.31 ;
      RECT 8170.185 1048.035 8170.465 1193.55 ;
      RECT 8169.625 1048.035 8169.905 1193.79 ;
      RECT 8169.065 1048.035 8169.345 1194.03 ;
      RECT 8168.505 1048.035 8168.785 1194.27 ;
      RECT 8167.945 1048.035 8168.225 1194.51 ;
      RECT 8167.385 1048.035 8167.665 1194.75 ;
      RECT 8166.825 1048.035 8167.105 1194.75 ;
      RECT 8166.265 1046.935 8166.545 1194.51 ;
      RECT 8165.705 1048.035 8165.985 1194.27 ;
      RECT 8165.145 1046.935 8165.425 1194.03 ;
      RECT 8164.585 1048.035 8164.865 1193.79 ;
      RECT 8164.025 1048.035 8164.305 1193.55 ;
      RECT 8163.465 1048.035 8163.745 1193.31 ;
      RECT 8162.905 1046.935 8163.185 1193.045 ;
      RECT 8162.345 1048.035 8162.625 1192.805 ;
      RECT 8161.785 1046.935 8162.065 1192.565 ;
      RECT 8161.225 1048.035 8161.505 1192.325 ;
      RECT 8152.265 1046.935 8152.545 1186.16 ;
      RECT 8151.705 1048.035 8151.985 1186.4 ;
      RECT 8151.145 1048.035 8151.425 1186.64 ;
      RECT 8150.585 1048.035 8150.865 1186.64 ;
      RECT 8150.025 1048.035 8150.305 1186.4 ;
      RECT 8149.465 1048.035 8149.745 1186.16 ;
      RECT 8148.905 1048.035 8149.185 1185.92 ;
      RECT 8148.345 1048.035 8148.625 1185.68 ;
      RECT 8147.785 1048.035 8148.065 1185.44 ;
      RECT 8147.225 1048.035 8147.505 1185.2 ;
      RECT 8146.665 1048.035 8146.945 1184.96 ;
      RECT 8146.105 1048.035 8146.385 1184.72 ;
      RECT 8145.545 1048.035 8145.825 1184.48 ;
      RECT 8144.985 1046.935 8145.265 1184.24 ;
      RECT 8142.465 1048.035 8142.745 1185.96 ;
      RECT 8141.905 1046.935 8142.185 1185.72 ;
      RECT 8141.345 1048.035 8141.625 1185.48 ;
      RECT 8140.785 1046.935 8141.065 1185.24 ;
      RECT 8140.225 1048.035 8140.505 1185 ;
      RECT 8139.665 1048.035 8139.945 1184.76 ;
      RECT 8139.105 1048.035 8139.385 1184.52 ;
      RECT 8113.065 1048.035 8113.345 1187.305 ;
      RECT 8112.505 1048.035 8112.785 1187.545 ;
      RECT 8111.945 1048.035 8112.225 1187.785 ;
      RECT 8111.385 1048.035 8111.665 1188.025 ;
      RECT 8110.825 1048.035 8111.105 1188.265 ;
      RECT 8110.265 1046.935 8110.545 1188.505 ;
      RECT 8109.705 1048.035 8109.985 1188.745 ;
      RECT 8109.145 1046.935 8109.425 1188.985 ;
      RECT 8108.585 1048.035 8108.865 1189.225 ;
      RECT 8108.025 1048.035 8108.305 1189.465 ;
      RECT 8107.465 1048.035 8107.745 1189.705 ;
      RECT 8106.905 1048.035 8107.185 1189.945 ;
      RECT 8106.345 1048.035 8106.625 1190.185 ;
      RECT 8105.785 1048.035 8106.065 1190.425 ;
      RECT 8105.225 1048.035 8105.505 1190.665 ;
      RECT 8104.665 1048.035 8104.945 1190.665 ;
      RECT 8104.105 1048.035 8104.385 1190.425 ;
      RECT 8103.545 1048.035 8103.825 1190.185 ;
      RECT 8102.985 1048.035 8103.265 1189.945 ;
      RECT 8102.425 1048.035 8102.705 1189.7 ;
      RECT 8101.865 1048.035 8102.145 1189.46 ;
      RECT 8101.305 1048.035 8101.585 1189.22 ;
      RECT 8100.745 1046.935 8101.025 1188.98 ;
      RECT 8100.185 1048.035 8100.465 1188.74 ;
      RECT 8086.745 1046.935 8087.025 1186.22 ;
      RECT 8086.185 1048.035 8086.465 1185.98 ;
      RECT 8085.625 1048.035 8085.905 1185.74 ;
      RECT 8085.065 1048.035 8085.345 1185.5 ;
      RECT 8084.505 1046.935 8084.785 1185.26 ;
      RECT 8083.945 1048.035 8084.225 1185.02 ;
      RECT 8083.385 1046.935 8083.665 1184.78 ;
      RECT 8082.825 1048.035 8083.105 1184.54 ;
      RECT 8082.265 1046.935 8082.545 1184.3 ;
      RECT 8081.705 1048.035 8081.985 1184.06 ;
      RECT 8081.145 1048.035 8081.425 1183.82 ;
      RECT 8080.585 1048.035 8080.865 1183.58 ;
      RECT 8080.025 1048.035 8080.305 1183.34 ;
      RECT 8079.465 1048.035 8079.745 1183.1 ;
      RECT 8078.905 1048.035 8079.185 1182.86 ;
      RECT 8078.345 1048.035 8078.625 1182.62 ;
      RECT 8077.785 1048.035 8078.065 1182.38 ;
      RECT 8077.225 1048.035 8077.505 1182.14 ;
      RECT 8076.665 1048.035 8076.945 1181.9 ;
      RECT 8076.105 1048.035 8076.385 1181.66 ;
      RECT 8075.545 1048.035 8075.825 1181.42 ;
      RECT 8074.985 1046.935 8075.265 1181.18 ;
      RECT 8074.425 1048.035 8074.705 1180.94 ;
      RECT 8073.865 1046.935 8074.145 1180.7 ;
      RECT 8034.105 1048.035 8034.385 1191.17 ;
      RECT 8033.545 1046.935 8033.825 1191.41 ;
      RECT 8032.985 1048.035 8033.265 1191.65 ;
      RECT 8032.425 1048.035 8032.705 1191.89 ;
      RECT 8031.865 1048.035 8032.145 1192.13 ;
      RECT 8031.305 1048.035 8031.585 1192.37 ;
      RECT 8030.745 1048.035 8031.025 1192.61 ;
      RECT 8030.185 1048.035 8030.465 1192.855 ;
      RECT 8029.625 1048.035 8029.905 1193.095 ;
      RECT 8029.065 1048.035 8029.345 1193.335 ;
      RECT 8028.505 1046.935 8028.785 1193.575 ;
      RECT 8027.945 1048.035 8028.225 1193.815 ;
      RECT 8027.385 1046.935 8027.665 1194.055 ;
      RECT 8026.825 1048.035 8027.105 1194.295 ;
      RECT 8026.265 1048.035 8026.545 1194.535 ;
      RECT 8025.705 1048.035 8025.985 1194.775 ;
      RECT 8025.145 1048.035 8025.425 1195.015 ;
      RECT 8024.585 1048.035 8024.865 1195.255 ;
      RECT 8024.025 1048.035 8024.305 1195.495 ;
      RECT 8023.465 1048.035 8023.745 1195.735 ;
      RECT 8022.905 1048.035 8023.185 1195.975 ;
      RECT 8022.345 1048.035 8022.625 1196.215 ;
      RECT 8021.785 1048.035 8022.065 1196.455 ;
      RECT 8021.225 1048.035 8021.505 1196.695 ;
      RECT 8012.265 1048.035 8012.545 1192.28 ;
      RECT 8011.705 1048.035 8011.985 1192.04 ;
      RECT 8011.145 1048.035 8011.425 1191.8 ;
      RECT 8010.585 1046.935 8010.865 1191.56 ;
      RECT 8010.025 1048.035 8010.305 1191.32 ;
      RECT 8009.465 1046.935 8009.745 1191.08 ;
      RECT 8008.905 1048.035 8009.185 1190.84 ;
      RECT 8008.345 1048.035 8008.625 1190.6 ;
      RECT 8007.785 1048.035 8008.065 1190.36 ;
      RECT 8007.225 1046.935 8007.505 1190.12 ;
      RECT 8006.665 1048.035 8006.945 1189.88 ;
      RECT 8006.105 1046.935 8006.385 1189.64 ;
      RECT 8005.545 1048.035 8005.825 1189.4 ;
      RECT 8004.985 1046.935 8005.265 1189.16 ;
      RECT 8002.465 1048.035 8002.745 1181.56 ;
      RECT 8001.905 1048.035 8002.185 1181.32 ;
      RECT 8001.345 1048.035 8001.625 1181.08 ;
      RECT 8000.785 1048.035 8001.065 1180.84 ;
      RECT 8000.225 1048.035 8000.505 1180.6 ;
      RECT 7999.665 1048.035 7999.945 1180.36 ;
      RECT 7999.105 1048.035 7999.385 1180.12 ;
      RECT 7973.065 1048.035 7973.345 1193.995 ;
      RECT 7972.505 1048.035 7972.785 1194.235 ;
      RECT 7971.945 1048.035 7972.225 1194.475 ;
      RECT 7971.385 1048.035 7971.665 1194.715 ;
      RECT 7970.825 1048.035 7971.105 1194.955 ;
      RECT 7970.265 1046.935 7970.545 1194.955 ;
      RECT 7969.705 1048.035 7969.985 1194.715 ;
      RECT 7969.145 1046.935 7969.425 1194.47 ;
      RECT 7968.585 1048.035 7968.865 1194.23 ;
      RECT 7968.025 1046.935 7968.305 1193.99 ;
      RECT 7967.465 1048.035 7967.745 1193.75 ;
      RECT 7966.905 1048.035 7967.185 1193.51 ;
      RECT 7966.345 1048.035 7966.625 1193.27 ;
      RECT 7965.785 1048.035 7966.065 1193.03 ;
      RECT 7965.225 1048.035 7965.505 1192.79 ;
      RECT 7964.665 1048.035 7964.945 1192.55 ;
      RECT 7964.105 1048.035 7964.385 1192.31 ;
      RECT 7963.545 1048.035 7963.825 1192.07 ;
      RECT 7962.985 1046.935 7963.265 1191.83 ;
      RECT 7962.425 1048.035 7962.705 1191.59 ;
      RECT 7961.865 1046.935 7962.145 1191.35 ;
      RECT 7961.305 1048.035 7961.585 1191.11 ;
      RECT 7960.745 1048.035 7961.025 1190.87 ;
      RECT 7960.185 1048.035 7960.465 1190.63 ;
      RECT 7946.745 1048.035 7947.025 1194.03 ;
      RECT 7946.185 1048.035 7946.465 1194.27 ;
      RECT 7945.625 1048.035 7945.905 1194.515 ;
      RECT 7945.065 1048.035 7945.345 1194.755 ;
      RECT 7944.505 1048.035 7944.785 1194.995 ;
      RECT 7943.945 1048.035 7944.225 1194.995 ;
      RECT 7943.385 1048.035 7943.665 1194.755 ;
      RECT 7942.825 1048.035 7943.105 1194.515 ;
      RECT 7942.265 1048.035 7942.545 1187.5 ;
      RECT 7941.705 1048.035 7941.985 1187.26 ;
      RECT 7941.145 1048.035 7941.425 1187.02 ;
      RECT 7940.585 1046.935 7940.865 1186.78 ;
      RECT 7940.025 1048.035 7940.305 1186.54 ;
      RECT 7939.465 1046.935 7939.745 1186.3 ;
      RECT 7938.905 1048.035 7939.185 1186.06 ;
      RECT 7938.345 1048.035 7938.625 1185.82 ;
      RECT 7937.785 1048.035 7938.065 1185.58 ;
      RECT 7937.225 1046.935 7937.505 1185.34 ;
      RECT 7936.665 1048.035 7936.945 1185.1 ;
      RECT 7936.105 1046.935 7936.385 1184.86 ;
      RECT 7935.545 1048.035 7935.825 1184.62 ;
      RECT 7934.985 1046.935 7935.265 1184.38 ;
      RECT 7934.425 1048.035 7934.705 1184.14 ;
      RECT 7933.865 1048.035 7934.145 1183.9 ;
      RECT 7893.545 1048.035 7893.825 1192.795 ;
      RECT 7892.985 1048.035 7893.265 1193.035 ;
      RECT 7892.425 1048.035 7892.705 1193.28 ;
      RECT 7891.865 1048.035 7892.145 1193.52 ;
      RECT 7891.305 1048.035 7891.585 1193.76 ;
      RECT 7890.745 1048.035 7891.025 1194 ;
      RECT 7890.185 1048.035 7890.465 1194.24 ;
      RECT 7889.625 1048.035 7889.905 1194.48 ;
      RECT 7889.065 1048.035 7889.345 1194.72 ;
      RECT 7888.505 1048.035 7888.785 1194.96 ;
      RECT 7887.945 1046.935 7888.225 1195.2 ;
      RECT 7887.385 1048.035 7887.665 1195.44 ;
      RECT 7886.825 1046.935 7887.105 1195.68 ;
      RECT 7886.265 1048.035 7886.545 1195.92 ;
      RECT 7885.705 1046.935 7885.985 1196.16 ;
      RECT 7885.145 1048.035 7885.425 1196.16 ;
      RECT 7884.585 1048.035 7884.865 1195.92 ;
      RECT 7884.025 1048.035 7884.305 1195.68 ;
      RECT 7883.465 1048.035 7883.745 1195.44 ;
      RECT 7882.905 1048.035 7883.185 1195.2 ;
      RECT 7882.345 1048.035 7882.625 1194.96 ;
      RECT 7881.785 1048.035 7882.065 1194.72 ;
      RECT 7881.225 1048.035 7881.505 1194.48 ;
      RECT 7872.265 1046.935 7872.545 1194.51 ;
      RECT 7871.705 1048.035 7871.985 1194.75 ;
      RECT 7871.145 1046.935 7871.425 1194.99 ;
      RECT 7870.585 1048.035 7870.865 1195.205 ;
      RECT 7870.025 1048.035 7870.305 1194.78 ;
      RECT 7869.465 1048.035 7869.745 1194.54 ;
      RECT 7868.905 1048.035 7869.185 1194.3 ;
      RECT 7868.345 1048.035 7868.625 1194.06 ;
      RECT 7867.785 1048.035 7868.065 1193.82 ;
      RECT 7867.225 1048.035 7867.505 1193.58 ;
      RECT 7866.665 1048.035 7866.945 1193.34 ;
      RECT 7866.105 1048.035 7866.385 1193.1 ;
      RECT 7865.545 1048.035 7865.825 1192.86 ;
      RECT 7864.985 1048.035 7865.265 1192.62 ;
      RECT 7862.465 1048.035 7862.745 1191.795 ;
      RECT 7861.905 1048.035 7862.185 1191.555 ;
      RECT 7861.345 1048.035 7861.625 1191.315 ;
      RECT 7860.785 1046.935 7861.065 1191.075 ;
      RECT 7860.225 1048.035 7860.505 1190.835 ;
      RECT 7859.665 1046.935 7859.945 1190.595 ;
      RECT 7859.105 1048.035 7859.385 1190.355 ;
      RECT 7858.545 1048.035 7858.825 1190.115 ;
      RECT 7831.945 1048.035 7832.225 1201.16 ;
      RECT 7831.385 1046.935 7831.665 1201.4 ;
      RECT 7830.825 1048.035 7831.105 1201.64 ;
      RECT 7830.265 1046.935 7830.545 1201.885 ;
      RECT 7829.705 1048.035 7829.985 1202.125 ;
      RECT 7829.145 1046.935 7829.425 1202.365 ;
      RECT 7828.585 1048.035 7828.865 1202.605 ;
      RECT 7828.025 1048.035 7828.305 1202.845 ;
      RECT 7827.465 1048.035 7827.745 1188.465 ;
      RECT 7826.905 1048.035 7827.185 1188.225 ;
      RECT 7826.345 1048.035 7826.625 1187.985 ;
      RECT 7825.785 1048.035 7826.065 1187.745 ;
      RECT 7825.225 1048.035 7825.505 1187.505 ;
      RECT 7824.665 1048.035 7824.945 1187.265 ;
      RECT 7824.105 1048.035 7824.385 1187.025 ;
      RECT 7823.545 1048.035 7823.825 1186.785 ;
      RECT 7822.985 1048.035 7823.265 1186.545 ;
      RECT 7822.425 1048.035 7822.705 1186.305 ;
      RECT 7821.865 1046.935 7822.145 1186.065 ;
      RECT 7821.305 1048.035 7821.585 1185.825 ;
      RECT 7820.745 1046.935 7821.025 1185.585 ;
      RECT 7820.185 1048.035 7820.465 1185.345 ;
      RECT 7806.185 1046.935 7806.465 1191.465 ;
      RECT 7805.625 1048.035 7805.905 1191.225 ;
      RECT 7805.065 1048.035 7805.345 1190.985 ;
      RECT 7804.505 1048.035 7804.785 1190.745 ;
      RECT 7803.945 1048.035 7804.225 1190.505 ;
      RECT 7803.385 1048.035 7803.665 1190.265 ;
      RECT 7802.825 1048.035 7803.105 1190.025 ;
      RECT 7802.265 1048.035 7802.545 1189.785 ;
      RECT 7801.705 1048.035 7801.985 1189.545 ;
      RECT 7801.145 1046.935 7801.425 1189.305 ;
      RECT 7800.585 1048.035 7800.865 1189.065 ;
      RECT 7800.025 1046.935 7800.305 1188.825 ;
      RECT 7799.465 1048.035 7799.745 1188.585 ;
      RECT 7798.905 1048.035 7799.185 1188.345 ;
      RECT 7798.345 1048.035 7798.625 1188.105 ;
      RECT 7797.785 1048.035 7798.065 1187.865 ;
      RECT 7797.225 1048.035 7797.505 1187.625 ;
      RECT 7796.665 1048.035 7796.945 1187.385 ;
      RECT 7796.105 1048.035 7796.385 1187.145 ;
      RECT 7795.545 1048.035 7795.825 1186.905 ;
      RECT 7794.985 1048.035 7795.265 1186.665 ;
      RECT 7794.425 1048.035 7794.705 1186.425 ;
      RECT 7793.865 1048.035 7794.145 1186.185 ;
      RECT 7754.665 1048.035 7754.945 1193.09 ;
      RECT 7754.105 1048.035 7754.385 1193.33 ;
      RECT 7753.545 1048.035 7753.825 1193.57 ;
      RECT 7752.985 1046.935 7753.265 1193.81 ;
      RECT 7752.425 1048.035 7752.705 1194.05 ;
      RECT 7751.865 1046.935 7752.145 1194.29 ;
      RECT 7751.305 1048.035 7751.585 1194.53 ;
      RECT 7750.745 1048.035 7751.025 1194.77 ;
      RECT 7750.185 1048.035 7750.465 1195.01 ;
      RECT 7749.625 1046.935 7749.905 1195.25 ;
      RECT 7749.065 1048.035 7749.345 1195.49 ;
      RECT 7748.505 1046.935 7748.785 1195.73 ;
      RECT 7747.945 1048.035 7748.225 1195.97 ;
      RECT 7747.385 1046.935 7747.665 1196.21 ;
      RECT 7746.825 1048.035 7747.105 1196.45 ;
      RECT 7746.265 1048.035 7746.545 1196.69 ;
      RECT 7745.705 1048.035 7745.985 1196.69 ;
      RECT 7745.145 1048.035 7745.425 1196.45 ;
      RECT 7744.585 1048.035 7744.865 1196.21 ;
      RECT 7744.025 1048.035 7744.305 1195.97 ;
      RECT 7743.465 1048.035 7743.745 1195.73 ;
      RECT 7742.905 1048.035 7743.185 1195.49 ;
      RECT 7742.345 1048.035 7742.625 1195.25 ;
      RECT 7741.785 1048.035 7742.065 1195.01 ;
      RECT 7741.225 1048.035 7741.505 1194.77 ;
      RECT 7732.265 1048.035 7732.545 1194.285 ;
      RECT 7731.705 1046.935 7731.985 1194.045 ;
      RECT 7731.145 1048.035 7731.425 1193.805 ;
      RECT 7730.585 1046.935 7730.865 1193.565 ;
      RECT 7730.025 1048.035 7730.305 1193.325 ;
      RECT 7729.465 1046.935 7729.745 1193.085 ;
      RECT 7728.905 1048.035 7729.185 1192.845 ;
      RECT 7728.345 1048.035 7728.625 1192.605 ;
      RECT 7727.785 1048.035 7728.065 1192.365 ;
      RECT 7727.225 1048.035 7727.505 1192.125 ;
      RECT 7726.665 1048.035 7726.945 1191.885 ;
      RECT 7726.105 1048.035 7726.385 1191.645 ;
      RECT 7725.545 1048.035 7725.825 1191.405 ;
      RECT 7724.985 1048.035 7725.265 1191.165 ;
      RECT 7722.465 1046.935 7722.745 1192.885 ;
      RECT 7721.905 1048.035 7722.185 1192.645 ;
      RECT 7721.345 1046.935 7721.625 1192.405 ;
      RECT 7720.785 1048.035 7721.065 1192.165 ;
      RECT 7720.225 1048.035 7720.505 1191.925 ;
      RECT 7719.665 1048.035 7719.945 1191.685 ;
      RECT 7719.105 1048.035 7719.385 1191.445 ;
      RECT 7718.545 1048.035 7718.825 1191.205 ;
      RECT 7692.505 1048.035 7692.785 1188.855 ;
      RECT 7691.945 1048.035 7692.225 1189.095 ;
      RECT 7691.385 1048.035 7691.665 1189.335 ;
      RECT 7690.825 1048.035 7691.105 1189.58 ;
      RECT 7690.265 1048.035 7690.545 1189.82 ;
      RECT 7689.705 1048.035 7689.985 1190.06 ;
      RECT 7689.145 1048.035 7689.425 1190.06 ;
      RECT 7688.585 1048.035 7688.865 1189.82 ;
      RECT 7688.025 1048.035 7688.305 1189.58 ;
      RECT 7687.465 1046.935 7687.745 1189.34 ;
      RECT 7686.905 1048.035 7687.185 1189.1 ;
      RECT 7686.345 1046.935 7686.625 1188.86 ;
      RECT 7685.785 1048.035 7686.065 1188.62 ;
      RECT 7685.225 1048.035 7685.505 1188.38 ;
      RECT 7684.665 1048.035 7684.945 1188.14 ;
      RECT 7684.105 1046.935 7684.385 1187.9 ;
      RECT 7683.545 1048.035 7683.825 1187.66 ;
      RECT 7682.985 1046.935 7683.265 1187.42 ;
      RECT 7682.425 1048.035 7682.705 1187.18 ;
      RECT 7681.865 1046.935 7682.145 1186.94 ;
      RECT 7681.305 1048.035 7681.585 1186.7 ;
      RECT 7680.745 1048.035 7681.025 1186.46 ;
      RECT 7680.185 1048.035 7680.465 1186.22 ;
      RECT 7679.625 1048.035 7679.905 1185.98 ;
      RECT 7666.185 1048.035 7666.465 1191.78 ;
      RECT 7665.625 1048.035 7665.905 1191.54 ;
      RECT 7665.065 1048.035 7665.345 1191.3 ;
      RECT 7664.505 1048.035 7664.785 1191.06 ;
      RECT 7663.945 1048.035 7664.225 1190.82 ;
      RECT 7663.385 1048.035 7663.665 1190.58 ;
      RECT 7662.825 1048.035 7663.105 1190.34 ;
      RECT 7662.265 1048.035 7662.545 1190.1 ;
      RECT 7661.705 1046.935 7661.985 1189.86 ;
      RECT 7661.145 1048.035 7661.425 1189.62 ;
      RECT 7660.585 1046.935 7660.865 1189.3 ;
      RECT 7660.025 1048.035 7660.305 1189.14 ;
      RECT 7659.465 1046.935 7659.745 1188.9 ;
      RECT 7658.905 1048.035 7659.185 1188.66 ;
      RECT 7658.345 1048.035 7658.625 1188.42 ;
      RECT 7657.785 1048.035 7658.065 1188.18 ;
      RECT 7657.225 1048.035 7657.505 1187.94 ;
      RECT 7656.665 1048.035 7656.945 1187.7 ;
      RECT 7656.105 1048.035 7656.385 1187.46 ;
      RECT 7655.545 1048.035 7655.825 1187.22 ;
      RECT 7654.985 1048.035 7655.265 1186.98 ;
      RECT 7654.425 1046.935 7654.705 1186.74 ;
      RECT 7653.865 1048.035 7654.145 1186.5 ;
      RECT 7653.305 1046.935 7653.585 1186.26 ;
      RECT 7614.105 1048.035 7614.385 1191.87 ;
      RECT 7613.545 1048.035 7613.825 1192.11 ;
      RECT 7612.985 1048.035 7613.265 1192.35 ;
      RECT 7612.425 1048.035 7612.705 1192.59 ;
      RECT 7611.865 1048.035 7612.145 1192.83 ;
      RECT 7611.305 1048.035 7611.585 1193.07 ;
      RECT 7610.745 1048.035 7611.025 1193.31 ;
      RECT 7610.185 1048.035 7610.465 1193.55 ;
      RECT 7609.625 1048.035 7609.905 1193.79 ;
      RECT 7609.065 1048.035 7609.345 1194.03 ;
      RECT 7608.505 1048.035 7608.785 1194.27 ;
      RECT 7607.945 1048.035 7608.225 1194.51 ;
      RECT 7607.385 1048.035 7607.665 1194.75 ;
      RECT 7606.825 1048.035 7607.105 1194.75 ;
      RECT 7606.265 1046.935 7606.545 1194.51 ;
      RECT 7605.705 1048.035 7605.985 1194.27 ;
      RECT 7605.145 1046.935 7605.425 1194.03 ;
      RECT 7604.585 1048.035 7604.865 1193.79 ;
      RECT 7604.025 1048.035 7604.305 1193.55 ;
      RECT 7603.465 1048.035 7603.745 1193.31 ;
      RECT 7602.905 1046.935 7603.185 1193.045 ;
      RECT 7602.345 1048.035 7602.625 1192.805 ;
      RECT 7601.785 1046.935 7602.065 1192.565 ;
      RECT 7601.225 1048.035 7601.505 1192.325 ;
      RECT 7592.265 1046.935 7592.545 1186.16 ;
      RECT 7591.705 1048.035 7591.985 1186.4 ;
      RECT 7591.145 1048.035 7591.425 1186.64 ;
      RECT 7590.585 1048.035 7590.865 1186.64 ;
      RECT 7590.025 1048.035 7590.305 1186.4 ;
      RECT 7589.465 1048.035 7589.745 1186.16 ;
      RECT 7588.905 1048.035 7589.185 1185.92 ;
      RECT 7588.345 1048.035 7588.625 1185.68 ;
      RECT 7587.785 1048.035 7588.065 1185.44 ;
      RECT 7587.225 1048.035 7587.505 1185.2 ;
      RECT 7586.665 1048.035 7586.945 1184.96 ;
      RECT 7586.105 1048.035 7586.385 1184.72 ;
      RECT 7585.545 1048.035 7585.825 1184.48 ;
      RECT 7584.985 1046.935 7585.265 1184.24 ;
      RECT 7582.465 1048.035 7582.745 1185.96 ;
      RECT 7581.905 1046.935 7582.185 1185.72 ;
      RECT 7581.345 1048.035 7581.625 1185.48 ;
      RECT 7580.785 1046.935 7581.065 1185.24 ;
      RECT 7580.225 1048.035 7580.505 1185 ;
      RECT 7579.665 1048.035 7579.945 1184.76 ;
      RECT 7579.105 1048.035 7579.385 1184.52 ;
      RECT 7553.065 1048.035 7553.345 1187.305 ;
      RECT 7552.505 1048.035 7552.785 1187.545 ;
      RECT 7551.945 1048.035 7552.225 1187.785 ;
      RECT 7551.385 1048.035 7551.665 1188.025 ;
      RECT 7550.825 1048.035 7551.105 1188.265 ;
      RECT 7550.265 1046.935 7550.545 1188.505 ;
      RECT 7549.705 1048.035 7549.985 1188.745 ;
      RECT 7549.145 1046.935 7549.425 1188.985 ;
      RECT 7548.585 1048.035 7548.865 1189.225 ;
      RECT 7548.025 1048.035 7548.305 1189.465 ;
      RECT 7547.465 1048.035 7547.745 1189.705 ;
      RECT 7546.905 1048.035 7547.185 1189.945 ;
      RECT 7546.345 1048.035 7546.625 1190.185 ;
      RECT 7545.785 1048.035 7546.065 1190.425 ;
      RECT 7545.225 1048.035 7545.505 1190.665 ;
      RECT 7544.665 1048.035 7544.945 1190.665 ;
      RECT 7544.105 1048.035 7544.385 1190.425 ;
      RECT 7543.545 1048.035 7543.825 1190.185 ;
      RECT 7542.985 1048.035 7543.265 1189.945 ;
      RECT 7542.425 1048.035 7542.705 1189.7 ;
      RECT 7541.865 1048.035 7542.145 1189.46 ;
      RECT 7541.305 1048.035 7541.585 1189.22 ;
      RECT 7540.745 1046.935 7541.025 1188.98 ;
      RECT 7540.185 1048.035 7540.465 1188.74 ;
      RECT 7526.745 1046.935 7527.025 1186.22 ;
      RECT 7526.185 1048.035 7526.465 1185.98 ;
      RECT 7525.625 1048.035 7525.905 1185.74 ;
      RECT 7525.065 1048.035 7525.345 1185.5 ;
      RECT 7524.505 1046.935 7524.785 1185.26 ;
      RECT 7523.945 1048.035 7524.225 1185.02 ;
      RECT 7523.385 1046.935 7523.665 1184.78 ;
      RECT 7522.825 1048.035 7523.105 1184.54 ;
      RECT 7522.265 1046.935 7522.545 1184.3 ;
      RECT 7521.705 1048.035 7521.985 1184.06 ;
      RECT 7521.145 1048.035 7521.425 1183.82 ;
      RECT 7520.585 1048.035 7520.865 1183.58 ;
      RECT 7520.025 1048.035 7520.305 1183.34 ;
      RECT 7519.465 1048.035 7519.745 1183.1 ;
      RECT 7518.905 1048.035 7519.185 1182.86 ;
      RECT 7518.345 1048.035 7518.625 1182.62 ;
      RECT 7517.785 1048.035 7518.065 1182.38 ;
      RECT 7517.225 1048.035 7517.505 1182.14 ;
      RECT 7516.665 1048.035 7516.945 1181.9 ;
      RECT 7516.105 1048.035 7516.385 1181.66 ;
      RECT 7515.545 1048.035 7515.825 1181.42 ;
      RECT 7514.985 1046.935 7515.265 1181.18 ;
      RECT 7514.425 1048.035 7514.705 1180.94 ;
      RECT 7513.865 1046.935 7514.145 1180.7 ;
      RECT 7474.105 1048.035 7474.385 1191.17 ;
      RECT 7473.545 1046.935 7473.825 1191.41 ;
      RECT 7472.985 1048.035 7473.265 1191.65 ;
      RECT 7472.425 1048.035 7472.705 1191.89 ;
      RECT 7471.865 1048.035 7472.145 1192.13 ;
      RECT 7471.305 1048.035 7471.585 1192.37 ;
      RECT 7470.745 1048.035 7471.025 1192.61 ;
      RECT 7470.185 1048.035 7470.465 1192.855 ;
      RECT 7469.625 1048.035 7469.905 1193.095 ;
      RECT 7469.065 1048.035 7469.345 1193.335 ;
      RECT 7468.505 1046.935 7468.785 1193.575 ;
      RECT 7467.945 1048.035 7468.225 1193.815 ;
      RECT 7467.385 1046.935 7467.665 1194.055 ;
      RECT 7466.825 1048.035 7467.105 1194.295 ;
      RECT 7466.265 1048.035 7466.545 1194.535 ;
      RECT 7465.705 1048.035 7465.985 1194.775 ;
      RECT 7465.145 1048.035 7465.425 1195.015 ;
      RECT 7464.585 1048.035 7464.865 1195.255 ;
      RECT 7464.025 1048.035 7464.305 1195.495 ;
      RECT 7463.465 1048.035 7463.745 1195.735 ;
      RECT 7462.905 1048.035 7463.185 1195.975 ;
      RECT 7462.345 1048.035 7462.625 1196.215 ;
      RECT 7461.785 1048.035 7462.065 1196.455 ;
      RECT 7461.225 1048.035 7461.505 1196.695 ;
      RECT 7452.265 1048.035 7452.545 1192.28 ;
      RECT 7451.705 1048.035 7451.985 1192.04 ;
      RECT 7451.145 1048.035 7451.425 1191.8 ;
      RECT 7450.585 1046.935 7450.865 1191.56 ;
      RECT 7450.025 1048.035 7450.305 1191.32 ;
      RECT 7449.465 1046.935 7449.745 1191.08 ;
      RECT 7448.905 1048.035 7449.185 1190.84 ;
      RECT 7448.345 1048.035 7448.625 1190.6 ;
      RECT 7447.785 1048.035 7448.065 1190.36 ;
      RECT 7447.225 1046.935 7447.505 1190.12 ;
      RECT 7446.665 1048.035 7446.945 1189.88 ;
      RECT 7446.105 1046.935 7446.385 1189.64 ;
      RECT 7445.545 1048.035 7445.825 1189.4 ;
      RECT 7444.985 1046.935 7445.265 1189.16 ;
      RECT 7442.465 1048.035 7442.745 1181.56 ;
      RECT 7441.905 1048.035 7442.185 1181.32 ;
      RECT 7441.345 1048.035 7441.625 1181.08 ;
      RECT 7440.785 1048.035 7441.065 1180.84 ;
      RECT 7440.225 1048.035 7440.505 1180.6 ;
      RECT 7439.665 1048.035 7439.945 1180.36 ;
      RECT 7439.105 1048.035 7439.385 1180.12 ;
      RECT 7413.065 1048.035 7413.345 1193.995 ;
      RECT 7412.505 1048.035 7412.785 1194.235 ;
      RECT 7411.945 1048.035 7412.225 1194.475 ;
      RECT 7411.385 1048.035 7411.665 1194.715 ;
      RECT 7410.825 1048.035 7411.105 1194.955 ;
      RECT 7410.265 1046.935 7410.545 1194.955 ;
      RECT 7409.705 1048.035 7409.985 1194.715 ;
      RECT 7409.145 1046.935 7409.425 1194.47 ;
      RECT 7408.585 1048.035 7408.865 1194.23 ;
      RECT 7408.025 1046.935 7408.305 1193.99 ;
      RECT 7407.465 1048.035 7407.745 1193.75 ;
      RECT 7406.905 1048.035 7407.185 1193.51 ;
      RECT 7406.345 1048.035 7406.625 1193.27 ;
      RECT 7405.785 1048.035 7406.065 1193.03 ;
      RECT 7405.225 1048.035 7405.505 1192.79 ;
      RECT 7404.665 1048.035 7404.945 1192.55 ;
      RECT 7404.105 1048.035 7404.385 1192.31 ;
      RECT 7403.545 1048.035 7403.825 1192.07 ;
      RECT 7402.985 1046.935 7403.265 1191.83 ;
      RECT 7402.425 1048.035 7402.705 1191.59 ;
      RECT 7401.865 1046.935 7402.145 1191.35 ;
      RECT 7401.305 1048.035 7401.585 1191.11 ;
      RECT 7400.745 1048.035 7401.025 1190.87 ;
      RECT 7400.185 1048.035 7400.465 1190.63 ;
      RECT 7386.745 1048.035 7387.025 1194.03 ;
      RECT 7386.185 1048.035 7386.465 1194.27 ;
      RECT 7385.625 1048.035 7385.905 1194.515 ;
      RECT 7385.065 1048.035 7385.345 1194.755 ;
      RECT 7384.505 1048.035 7384.785 1194.995 ;
      RECT 7383.945 1048.035 7384.225 1194.995 ;
      RECT 7383.385 1048.035 7383.665 1194.755 ;
      RECT 7382.825 1048.035 7383.105 1194.515 ;
      RECT 7382.265 1048.035 7382.545 1187.5 ;
      RECT 7381.705 1048.035 7381.985 1187.26 ;
      RECT 7381.145 1048.035 7381.425 1187.02 ;
      RECT 7380.585 1046.935 7380.865 1186.78 ;
      RECT 7380.025 1048.035 7380.305 1186.54 ;
      RECT 7379.465 1046.935 7379.745 1186.3 ;
      RECT 7378.905 1048.035 7379.185 1186.06 ;
      RECT 7378.345 1048.035 7378.625 1185.82 ;
      RECT 7377.785 1048.035 7378.065 1185.58 ;
      RECT 7377.225 1046.935 7377.505 1185.34 ;
      RECT 7376.665 1048.035 7376.945 1185.1 ;
      RECT 7376.105 1046.935 7376.385 1184.86 ;
      RECT 7375.545 1048.035 7375.825 1184.62 ;
      RECT 7374.985 1046.935 7375.265 1184.38 ;
      RECT 7374.425 1048.035 7374.705 1184.14 ;
      RECT 7373.865 1048.035 7374.145 1183.9 ;
      RECT 7333.545 1048.035 7333.825 1192.795 ;
      RECT 7332.985 1048.035 7333.265 1193.035 ;
      RECT 7332.425 1048.035 7332.705 1193.28 ;
      RECT 7331.865 1048.035 7332.145 1193.52 ;
      RECT 7331.305 1048.035 7331.585 1193.76 ;
      RECT 7330.745 1048.035 7331.025 1194 ;
      RECT 7330.185 1048.035 7330.465 1194.24 ;
      RECT 7329.625 1048.035 7329.905 1194.48 ;
      RECT 7329.065 1048.035 7329.345 1194.72 ;
      RECT 7328.505 1048.035 7328.785 1194.96 ;
      RECT 7327.945 1046.935 7328.225 1195.2 ;
      RECT 7327.385 1048.035 7327.665 1195.44 ;
      RECT 7326.825 1046.935 7327.105 1195.68 ;
      RECT 7326.265 1048.035 7326.545 1195.92 ;
      RECT 7325.705 1046.935 7325.985 1196.16 ;
      RECT 7325.145 1048.035 7325.425 1196.16 ;
      RECT 7324.585 1048.035 7324.865 1195.92 ;
      RECT 7324.025 1048.035 7324.305 1195.68 ;
      RECT 7323.465 1048.035 7323.745 1195.44 ;
      RECT 7322.905 1048.035 7323.185 1195.2 ;
      RECT 7322.345 1048.035 7322.625 1194.96 ;
      RECT 7321.785 1048.035 7322.065 1194.72 ;
      RECT 7321.225 1048.035 7321.505 1194.48 ;
      RECT 7312.265 1046.935 7312.545 1194.51 ;
      RECT 7311.705 1048.035 7311.985 1194.75 ;
      RECT 7311.145 1046.935 7311.425 1194.99 ;
      RECT 7310.585 1048.035 7310.865 1195.205 ;
      RECT 7310.025 1048.035 7310.305 1194.78 ;
      RECT 7309.465 1048.035 7309.745 1194.54 ;
      RECT 7308.905 1048.035 7309.185 1194.3 ;
      RECT 7308.345 1048.035 7308.625 1194.06 ;
      RECT 7307.785 1048.035 7308.065 1193.82 ;
      RECT 7307.225 1048.035 7307.505 1193.58 ;
      RECT 7306.665 1048.035 7306.945 1193.34 ;
      RECT 7306.105 1048.035 7306.385 1193.1 ;
      RECT 7305.545 1048.035 7305.825 1192.86 ;
      RECT 7304.985 1048.035 7305.265 1192.62 ;
      RECT 7302.465 1048.035 7302.745 1191.795 ;
      RECT 7301.905 1048.035 7302.185 1191.555 ;
      RECT 7301.345 1048.035 7301.625 1191.315 ;
      RECT 7300.785 1046.935 7301.065 1191.075 ;
      RECT 7300.225 1048.035 7300.505 1190.835 ;
      RECT 7299.665 1046.935 7299.945 1190.595 ;
      RECT 7299.105 1048.035 7299.385 1190.355 ;
      RECT 7298.545 1048.035 7298.825 1190.115 ;
      RECT 7271.945 1048.035 7272.225 1201.16 ;
      RECT 7271.385 1046.935 7271.665 1201.4 ;
      RECT 7270.825 1048.035 7271.105 1201.64 ;
      RECT 7270.265 1046.935 7270.545 1201.885 ;
      RECT 7269.705 1048.035 7269.985 1202.125 ;
      RECT 7269.145 1046.935 7269.425 1202.365 ;
      RECT 7268.585 1048.035 7268.865 1202.605 ;
      RECT 7268.025 1048.035 7268.305 1202.845 ;
      RECT 7267.465 1048.035 7267.745 1188.465 ;
      RECT 7266.905 1048.035 7267.185 1188.225 ;
      RECT 7266.345 1048.035 7266.625 1187.985 ;
      RECT 7265.785 1048.035 7266.065 1187.745 ;
      RECT 7265.225 1048.035 7265.505 1187.505 ;
      RECT 7264.665 1048.035 7264.945 1187.265 ;
      RECT 7264.105 1048.035 7264.385 1187.025 ;
      RECT 7263.545 1048.035 7263.825 1186.785 ;
      RECT 7262.985 1048.035 7263.265 1186.545 ;
      RECT 7262.425 1048.035 7262.705 1186.305 ;
      RECT 7261.865 1046.935 7262.145 1186.065 ;
      RECT 7261.305 1048.035 7261.585 1185.825 ;
      RECT 7260.745 1046.935 7261.025 1185.585 ;
      RECT 7260.185 1048.035 7260.465 1185.345 ;
      RECT 7246.185 1046.935 7246.465 1191.465 ;
      RECT 7245.625 1048.035 7245.905 1191.225 ;
      RECT 7245.065 1048.035 7245.345 1190.985 ;
      RECT 7244.505 1048.035 7244.785 1190.745 ;
      RECT 7243.945 1048.035 7244.225 1190.505 ;
      RECT 7243.385 1048.035 7243.665 1190.265 ;
      RECT 7242.825 1048.035 7243.105 1190.025 ;
      RECT 7242.265 1048.035 7242.545 1189.785 ;
      RECT 7241.705 1048.035 7241.985 1189.545 ;
      RECT 7241.145 1046.935 7241.425 1189.305 ;
      RECT 7240.585 1048.035 7240.865 1189.065 ;
      RECT 7240.025 1046.935 7240.305 1188.825 ;
      RECT 7239.465 1048.035 7239.745 1188.585 ;
      RECT 7238.905 1048.035 7239.185 1188.345 ;
      RECT 7238.345 1048.035 7238.625 1188.105 ;
      RECT 7237.785 1048.035 7238.065 1187.865 ;
      RECT 7237.225 1048.035 7237.505 1187.625 ;
      RECT 7236.665 1048.035 7236.945 1187.385 ;
      RECT 7236.105 1048.035 7236.385 1187.145 ;
      RECT 7235.545 1048.035 7235.825 1186.905 ;
      RECT 7234.985 1048.035 7235.265 1186.665 ;
      RECT 7234.425 1048.035 7234.705 1186.425 ;
      RECT 7233.865 1048.035 7234.145 1186.185 ;
      RECT 7194.665 1048.035 7194.945 1193.09 ;
      RECT 7194.105 1048.035 7194.385 1193.33 ;
      RECT 7193.545 1048.035 7193.825 1193.57 ;
      RECT 7192.985 1046.935 7193.265 1193.81 ;
      RECT 7192.425 1048.035 7192.705 1194.05 ;
      RECT 7191.865 1046.935 7192.145 1194.29 ;
      RECT 7191.305 1048.035 7191.585 1194.53 ;
      RECT 7190.745 1048.035 7191.025 1194.77 ;
      RECT 7190.185 1048.035 7190.465 1195.01 ;
      RECT 7189.625 1046.935 7189.905 1195.25 ;
      RECT 7189.065 1048.035 7189.345 1195.49 ;
      RECT 7188.505 1046.935 7188.785 1195.73 ;
      RECT 7187.945 1048.035 7188.225 1195.97 ;
      RECT 7187.385 1046.935 7187.665 1196.21 ;
      RECT 7186.825 1048.035 7187.105 1196.45 ;
      RECT 7186.265 1048.035 7186.545 1196.69 ;
      RECT 7185.705 1048.035 7185.985 1196.69 ;
      RECT 7185.145 1048.035 7185.425 1196.45 ;
      RECT 7184.585 1048.035 7184.865 1196.21 ;
      RECT 7184.025 1048.035 7184.305 1195.97 ;
      RECT 7183.465 1048.035 7183.745 1195.73 ;
      RECT 7182.905 1048.035 7183.185 1195.49 ;
      RECT 7182.345 1048.035 7182.625 1195.25 ;
      RECT 7181.785 1048.035 7182.065 1195.01 ;
      RECT 7181.225 1048.035 7181.505 1194.77 ;
      RECT 7172.265 1048.035 7172.545 1194.285 ;
      RECT 7171.705 1046.935 7171.985 1194.045 ;
      RECT 7171.145 1048.035 7171.425 1193.805 ;
      RECT 7170.585 1046.935 7170.865 1193.565 ;
      RECT 7170.025 1048.035 7170.305 1193.325 ;
      RECT 7169.465 1046.935 7169.745 1193.085 ;
      RECT 7168.905 1048.035 7169.185 1192.845 ;
      RECT 7168.345 1048.035 7168.625 1192.605 ;
      RECT 7167.785 1048.035 7168.065 1192.365 ;
      RECT 7167.225 1048.035 7167.505 1192.125 ;
      RECT 7166.665 1048.035 7166.945 1191.885 ;
      RECT 7166.105 1048.035 7166.385 1191.645 ;
      RECT 7165.545 1048.035 7165.825 1191.405 ;
      RECT 7164.985 1048.035 7165.265 1191.165 ;
      RECT 7162.465 1046.935 7162.745 1192.885 ;
      RECT 7161.905 1048.035 7162.185 1192.645 ;
      RECT 7161.345 1046.935 7161.625 1192.405 ;
      RECT 7160.785 1048.035 7161.065 1192.165 ;
      RECT 7160.225 1048.035 7160.505 1191.925 ;
      RECT 7159.665 1048.035 7159.945 1191.685 ;
      RECT 7159.105 1048.035 7159.385 1191.445 ;
      RECT 7158.545 1048.035 7158.825 1191.205 ;
      RECT 7132.505 1048.035 7132.785 1188.855 ;
      RECT 7131.945 1048.035 7132.225 1189.095 ;
      RECT 7131.385 1048.035 7131.665 1189.335 ;
      RECT 7130.825 1048.035 7131.105 1189.58 ;
      RECT 7130.265 1048.035 7130.545 1189.82 ;
      RECT 7129.705 1048.035 7129.985 1190.06 ;
      RECT 7129.145 1048.035 7129.425 1190.06 ;
      RECT 7128.585 1048.035 7128.865 1189.82 ;
      RECT 7128.025 1048.035 7128.305 1189.58 ;
      RECT 7127.465 1046.935 7127.745 1189.34 ;
      RECT 7126.905 1048.035 7127.185 1189.1 ;
      RECT 7126.345 1046.935 7126.625 1188.86 ;
      RECT 7125.785 1048.035 7126.065 1188.62 ;
      RECT 7125.225 1048.035 7125.505 1188.38 ;
      RECT 7124.665 1048.035 7124.945 1188.14 ;
      RECT 7124.105 1046.935 7124.385 1187.9 ;
      RECT 7123.545 1048.035 7123.825 1187.66 ;
      RECT 7122.985 1046.935 7123.265 1187.42 ;
      RECT 7122.425 1048.035 7122.705 1187.18 ;
      RECT 7121.865 1046.935 7122.145 1186.94 ;
      RECT 7121.305 1048.035 7121.585 1186.7 ;
      RECT 7120.745 1048.035 7121.025 1186.46 ;
      RECT 7120.185 1048.035 7120.465 1186.22 ;
      RECT 7119.625 1048.035 7119.905 1185.98 ;
      RECT 7106.185 1048.035 7106.465 1191.78 ;
      RECT 7105.625 1048.035 7105.905 1191.54 ;
      RECT 7105.065 1048.035 7105.345 1191.3 ;
      RECT 7104.505 1048.035 7104.785 1191.06 ;
      RECT 7103.945 1048.035 7104.225 1190.82 ;
      RECT 7103.385 1048.035 7103.665 1190.58 ;
      RECT 7102.825 1048.035 7103.105 1190.34 ;
      RECT 7102.265 1048.035 7102.545 1190.1 ;
      RECT 7101.705 1046.935 7101.985 1189.86 ;
      RECT 7101.145 1048.035 7101.425 1189.62 ;
      RECT 7100.585 1046.935 7100.865 1189.3 ;
      RECT 7100.025 1048.035 7100.305 1189.14 ;
      RECT 7099.465 1046.935 7099.745 1188.9 ;
      RECT 7098.905 1048.035 7099.185 1188.66 ;
      RECT 7098.345 1048.035 7098.625 1188.42 ;
      RECT 7097.785 1048.035 7098.065 1188.18 ;
      RECT 7097.225 1048.035 7097.505 1187.94 ;
      RECT 7096.665 1048.035 7096.945 1187.7 ;
      RECT 7096.105 1048.035 7096.385 1187.46 ;
      RECT 7095.545 1048.035 7095.825 1187.22 ;
      RECT 7094.985 1048.035 7095.265 1186.98 ;
      RECT 7094.425 1046.935 7094.705 1186.74 ;
      RECT 7093.865 1048.035 7094.145 1186.5 ;
      RECT 7093.305 1046.935 7093.585 1186.26 ;
      RECT 7054.105 1048.035 7054.385 1191.87 ;
      RECT 7053.545 1048.035 7053.825 1192.11 ;
      RECT 7052.985 1048.035 7053.265 1192.35 ;
      RECT 7052.425 1048.035 7052.705 1192.59 ;
      RECT 7051.865 1048.035 7052.145 1192.83 ;
      RECT 7051.305 1048.035 7051.585 1193.07 ;
      RECT 7050.745 1048.035 7051.025 1193.31 ;
      RECT 7050.185 1048.035 7050.465 1193.55 ;
      RECT 7049.625 1048.035 7049.905 1193.79 ;
      RECT 7049.065 1048.035 7049.345 1194.03 ;
      RECT 7048.505 1048.035 7048.785 1194.27 ;
      RECT 7047.945 1048.035 7048.225 1194.51 ;
      RECT 7047.385 1048.035 7047.665 1194.75 ;
      RECT 7046.825 1048.035 7047.105 1194.75 ;
      RECT 7046.265 1046.935 7046.545 1194.51 ;
      RECT 7045.705 1048.035 7045.985 1194.27 ;
      RECT 7045.145 1046.935 7045.425 1194.03 ;
      RECT 7044.585 1048.035 7044.865 1193.79 ;
      RECT 7044.025 1048.035 7044.305 1193.55 ;
      RECT 7043.465 1048.035 7043.745 1193.31 ;
      RECT 7042.905 1046.935 7043.185 1193.045 ;
      RECT 7042.345 1048.035 7042.625 1192.805 ;
      RECT 7041.785 1046.935 7042.065 1192.565 ;
      RECT 7041.225 1048.035 7041.505 1192.325 ;
      RECT 7032.265 1046.935 7032.545 1186.16 ;
      RECT 7031.705 1048.035 7031.985 1186.4 ;
      RECT 7031.145 1048.035 7031.425 1186.64 ;
      RECT 7030.585 1048.035 7030.865 1186.64 ;
      RECT 7030.025 1048.035 7030.305 1186.4 ;
      RECT 7029.465 1048.035 7029.745 1186.16 ;
      RECT 7028.905 1048.035 7029.185 1185.92 ;
      RECT 7028.345 1048.035 7028.625 1185.68 ;
      RECT 7027.785 1048.035 7028.065 1185.44 ;
      RECT 7027.225 1048.035 7027.505 1185.2 ;
      RECT 7026.665 1048.035 7026.945 1184.96 ;
      RECT 7026.105 1048.035 7026.385 1184.72 ;
      RECT 7025.545 1048.035 7025.825 1184.48 ;
      RECT 7024.985 1046.935 7025.265 1184.24 ;
      RECT 7022.465 1048.035 7022.745 1185.96 ;
      RECT 7021.905 1046.935 7022.185 1185.72 ;
      RECT 7021.345 1048.035 7021.625 1185.48 ;
      RECT 7020.785 1046.935 7021.065 1185.24 ;
      RECT 7020.225 1048.035 7020.505 1185 ;
      RECT 7019.665 1048.035 7019.945 1184.76 ;
      RECT 7019.105 1048.035 7019.385 1184.52 ;
      RECT 6993.065 1048.035 6993.345 1187.305 ;
      RECT 6992.505 1048.035 6992.785 1187.545 ;
      RECT 6991.945 1048.035 6992.225 1187.785 ;
      RECT 6991.385 1048.035 6991.665 1188.025 ;
      RECT 6990.825 1048.035 6991.105 1188.265 ;
      RECT 6990.265 1046.935 6990.545 1188.505 ;
      RECT 6989.705 1048.035 6989.985 1188.745 ;
      RECT 6989.145 1046.935 6989.425 1188.985 ;
      RECT 6988.585 1048.035 6988.865 1189.225 ;
      RECT 6988.025 1048.035 6988.305 1189.465 ;
      RECT 6987.465 1048.035 6987.745 1189.705 ;
      RECT 6986.905 1048.035 6987.185 1189.945 ;
      RECT 6986.345 1048.035 6986.625 1190.185 ;
      RECT 6985.785 1048.035 6986.065 1190.425 ;
      RECT 6985.225 1048.035 6985.505 1190.665 ;
      RECT 6984.665 1048.035 6984.945 1190.665 ;
      RECT 6984.105 1048.035 6984.385 1190.425 ;
      RECT 6983.545 1048.035 6983.825 1190.185 ;
      RECT 6982.985 1048.035 6983.265 1189.945 ;
      RECT 6982.425 1048.035 6982.705 1189.7 ;
      RECT 6981.865 1048.035 6982.145 1189.46 ;
      RECT 6981.305 1048.035 6981.585 1189.22 ;
      RECT 6980.745 1046.935 6981.025 1188.98 ;
      RECT 6980.185 1048.035 6980.465 1188.74 ;
      RECT 6966.745 1046.935 6967.025 1186.22 ;
      RECT 6966.185 1048.035 6966.465 1185.98 ;
      RECT 6965.625 1048.035 6965.905 1185.74 ;
      RECT 6965.065 1048.035 6965.345 1185.5 ;
      RECT 6964.505 1046.935 6964.785 1185.26 ;
      RECT 6963.945 1048.035 6964.225 1185.02 ;
      RECT 6963.385 1046.935 6963.665 1184.78 ;
      RECT 6962.825 1048.035 6963.105 1184.54 ;
      RECT 6962.265 1046.935 6962.545 1184.3 ;
      RECT 6961.705 1048.035 6961.985 1184.06 ;
      RECT 6961.145 1048.035 6961.425 1183.82 ;
      RECT 6960.585 1048.035 6960.865 1183.58 ;
      RECT 6960.025 1048.035 6960.305 1183.34 ;
      RECT 6959.465 1048.035 6959.745 1183.1 ;
      RECT 6958.905 1048.035 6959.185 1182.86 ;
      RECT 6958.345 1048.035 6958.625 1182.62 ;
      RECT 6957.785 1048.035 6958.065 1182.38 ;
      RECT 6957.225 1048.035 6957.505 1182.14 ;
      RECT 6956.665 1048.035 6956.945 1181.9 ;
      RECT 6956.105 1048.035 6956.385 1181.66 ;
      RECT 6955.545 1048.035 6955.825 1181.42 ;
      RECT 6954.985 1046.935 6955.265 1181.18 ;
      RECT 6954.425 1048.035 6954.705 1180.94 ;
      RECT 6953.865 1046.935 6954.145 1180.7 ;
      RECT 6914.105 1048.035 6914.385 1191.17 ;
      RECT 6913.545 1046.935 6913.825 1191.41 ;
      RECT 6912.985 1048.035 6913.265 1191.65 ;
      RECT 6912.425 1048.035 6912.705 1191.89 ;
      RECT 6911.865 1048.035 6912.145 1192.13 ;
      RECT 6911.305 1048.035 6911.585 1192.37 ;
      RECT 6910.745 1048.035 6911.025 1192.61 ;
      RECT 6910.185 1048.035 6910.465 1192.855 ;
      RECT 6909.625 1048.035 6909.905 1193.095 ;
      RECT 6909.065 1048.035 6909.345 1193.335 ;
      RECT 6908.505 1046.935 6908.785 1193.575 ;
      RECT 6907.945 1048.035 6908.225 1193.815 ;
      RECT 6907.385 1046.935 6907.665 1194.055 ;
      RECT 6906.825 1048.035 6907.105 1194.295 ;
      RECT 6906.265 1048.035 6906.545 1194.535 ;
      RECT 6905.705 1048.035 6905.985 1194.775 ;
      RECT 6905.145 1048.035 6905.425 1195.015 ;
      RECT 6904.585 1048.035 6904.865 1195.255 ;
      RECT 6904.025 1048.035 6904.305 1195.495 ;
      RECT 6903.465 1048.035 6903.745 1195.735 ;
      RECT 6902.905 1048.035 6903.185 1195.975 ;
      RECT 6902.345 1048.035 6902.625 1196.215 ;
      RECT 6901.785 1048.035 6902.065 1196.455 ;
      RECT 6901.225 1048.035 6901.505 1196.695 ;
      RECT 6892.265 1048.035 6892.545 1192.28 ;
      RECT 6891.705 1048.035 6891.985 1192.04 ;
      RECT 6891.145 1048.035 6891.425 1191.8 ;
      RECT 6890.585 1046.935 6890.865 1191.56 ;
      RECT 6890.025 1048.035 6890.305 1191.32 ;
      RECT 6889.465 1046.935 6889.745 1191.08 ;
      RECT 6888.905 1048.035 6889.185 1190.84 ;
      RECT 6888.345 1048.035 6888.625 1190.6 ;
      RECT 6887.785 1048.035 6888.065 1190.36 ;
      RECT 6887.225 1046.935 6887.505 1190.12 ;
      RECT 6886.665 1048.035 6886.945 1189.88 ;
      RECT 6886.105 1046.935 6886.385 1189.64 ;
      RECT 6885.545 1048.035 6885.825 1189.4 ;
      RECT 6884.985 1046.935 6885.265 1189.16 ;
      RECT 6882.465 1048.035 6882.745 1181.56 ;
      RECT 6881.905 1048.035 6882.185 1181.32 ;
      RECT 6881.345 1048.035 6881.625 1181.08 ;
      RECT 6880.785 1048.035 6881.065 1180.84 ;
      RECT 6880.225 1048.035 6880.505 1180.6 ;
      RECT 6879.665 1048.035 6879.945 1180.36 ;
      RECT 6879.105 1048.035 6879.385 1180.12 ;
      RECT 6853.065 1048.035 6853.345 1193.995 ;
      RECT 6852.505 1048.035 6852.785 1194.235 ;
      RECT 6851.945 1048.035 6852.225 1194.475 ;
      RECT 6851.385 1048.035 6851.665 1194.715 ;
      RECT 6850.825 1048.035 6851.105 1194.955 ;
      RECT 6850.265 1046.935 6850.545 1194.955 ;
      RECT 6849.705 1048.035 6849.985 1194.715 ;
      RECT 6849.145 1046.935 6849.425 1194.47 ;
      RECT 6848.585 1048.035 6848.865 1194.23 ;
      RECT 6848.025 1046.935 6848.305 1193.99 ;
      RECT 6847.465 1048.035 6847.745 1193.75 ;
      RECT 6846.905 1048.035 6847.185 1193.51 ;
      RECT 6846.345 1048.035 6846.625 1193.27 ;
      RECT 6845.785 1048.035 6846.065 1193.03 ;
      RECT 6845.225 1048.035 6845.505 1192.79 ;
      RECT 6844.665 1048.035 6844.945 1192.55 ;
      RECT 6844.105 1048.035 6844.385 1192.31 ;
      RECT 6843.545 1048.035 6843.825 1192.07 ;
      RECT 6842.985 1046.935 6843.265 1191.83 ;
      RECT 6842.425 1048.035 6842.705 1191.59 ;
      RECT 6841.865 1046.935 6842.145 1191.35 ;
      RECT 6841.305 1048.035 6841.585 1191.11 ;
      RECT 6840.745 1048.035 6841.025 1190.87 ;
      RECT 6840.185 1048.035 6840.465 1190.63 ;
      RECT 6826.745 1048.035 6827.025 1194.03 ;
      RECT 6826.185 1048.035 6826.465 1194.27 ;
      RECT 6825.625 1048.035 6825.905 1194.515 ;
      RECT 6825.065 1048.035 6825.345 1194.755 ;
      RECT 6824.505 1048.035 6824.785 1194.995 ;
      RECT 6823.945 1048.035 6824.225 1194.995 ;
      RECT 6823.385 1048.035 6823.665 1194.755 ;
      RECT 6822.825 1048.035 6823.105 1194.515 ;
      RECT 6822.265 1048.035 6822.545 1187.5 ;
      RECT 6821.705 1048.035 6821.985 1187.26 ;
      RECT 6821.145 1048.035 6821.425 1187.02 ;
      RECT 6820.585 1046.935 6820.865 1186.78 ;
      RECT 6820.025 1048.035 6820.305 1186.54 ;
      RECT 6819.465 1046.935 6819.745 1186.3 ;
      RECT 6818.905 1048.035 6819.185 1186.06 ;
      RECT 6818.345 1048.035 6818.625 1185.82 ;
      RECT 6817.785 1048.035 6818.065 1185.58 ;
      RECT 6817.225 1046.935 6817.505 1185.34 ;
      RECT 6816.665 1048.035 6816.945 1185.1 ;
      RECT 6816.105 1046.935 6816.385 1184.86 ;
      RECT 6815.545 1048.035 6815.825 1184.62 ;
      RECT 6814.985 1046.935 6815.265 1184.38 ;
      RECT 6814.425 1048.035 6814.705 1184.14 ;
      RECT 6813.865 1048.035 6814.145 1183.9 ;
      RECT 6773.545 1048.035 6773.825 1192.795 ;
      RECT 6772.985 1048.035 6773.265 1193.035 ;
      RECT 6772.425 1048.035 6772.705 1193.28 ;
      RECT 6771.865 1048.035 6772.145 1193.52 ;
      RECT 6771.305 1048.035 6771.585 1193.76 ;
      RECT 6770.745 1048.035 6771.025 1194 ;
      RECT 6770.185 1048.035 6770.465 1194.24 ;
      RECT 6769.625 1048.035 6769.905 1194.48 ;
      RECT 6769.065 1048.035 6769.345 1194.72 ;
      RECT 6768.505 1048.035 6768.785 1194.96 ;
      RECT 6767.945 1046.935 6768.225 1195.2 ;
      RECT 6767.385 1048.035 6767.665 1195.44 ;
      RECT 6766.825 1046.935 6767.105 1195.68 ;
      RECT 6766.265 1048.035 6766.545 1195.92 ;
      RECT 6765.705 1046.935 6765.985 1196.16 ;
      RECT 6765.145 1048.035 6765.425 1196.16 ;
      RECT 6764.585 1048.035 6764.865 1195.92 ;
      RECT 6764.025 1048.035 6764.305 1195.68 ;
      RECT 6763.465 1048.035 6763.745 1195.44 ;
      RECT 6762.905 1048.035 6763.185 1195.2 ;
      RECT 6762.345 1048.035 6762.625 1194.96 ;
      RECT 6761.785 1048.035 6762.065 1194.72 ;
      RECT 6761.225 1048.035 6761.505 1194.48 ;
      RECT 6752.265 1046.935 6752.545 1194.51 ;
      RECT 6751.705 1048.035 6751.985 1194.75 ;
      RECT 6751.145 1046.935 6751.425 1194.99 ;
      RECT 6750.585 1048.035 6750.865 1195.205 ;
      RECT 6750.025 1048.035 6750.305 1194.78 ;
      RECT 6749.465 1048.035 6749.745 1194.54 ;
      RECT 6748.905 1048.035 6749.185 1194.3 ;
      RECT 6748.345 1048.035 6748.625 1194.06 ;
      RECT 6747.785 1048.035 6748.065 1193.82 ;
      RECT 6747.225 1048.035 6747.505 1193.58 ;
      RECT 6746.665 1048.035 6746.945 1193.34 ;
      RECT 6746.105 1048.035 6746.385 1193.1 ;
      RECT 6745.545 1048.035 6745.825 1192.86 ;
      RECT 6744.985 1048.035 6745.265 1192.62 ;
      RECT 6742.465 1048.035 6742.745 1191.795 ;
      RECT 6741.905 1048.035 6742.185 1191.555 ;
      RECT 6741.345 1048.035 6741.625 1191.315 ;
      RECT 6740.785 1046.935 6741.065 1191.075 ;
      RECT 6740.225 1048.035 6740.505 1190.835 ;
      RECT 6739.665 1046.935 6739.945 1190.595 ;
      RECT 6739.105 1048.035 6739.385 1190.355 ;
      RECT 6738.545 1048.035 6738.825 1190.115 ;
      RECT 6711.945 1048.035 6712.225 1201.16 ;
      RECT 6711.385 1046.935 6711.665 1201.4 ;
      RECT 6710.825 1048.035 6711.105 1201.64 ;
      RECT 6710.265 1046.935 6710.545 1201.885 ;
      RECT 6709.705 1048.035 6709.985 1202.125 ;
      RECT 6709.145 1046.935 6709.425 1202.365 ;
      RECT 6708.585 1048.035 6708.865 1202.605 ;
      RECT 6708.025 1048.035 6708.305 1202.845 ;
      RECT 6707.465 1048.035 6707.745 1188.465 ;
      RECT 6706.905 1048.035 6707.185 1188.225 ;
      RECT 6706.345 1048.035 6706.625 1187.985 ;
      RECT 6705.785 1048.035 6706.065 1187.745 ;
      RECT 6705.225 1048.035 6705.505 1187.505 ;
      RECT 6704.665 1048.035 6704.945 1187.265 ;
      RECT 6704.105 1048.035 6704.385 1187.025 ;
      RECT 6703.545 1048.035 6703.825 1186.785 ;
      RECT 6702.985 1048.035 6703.265 1186.545 ;
      RECT 6702.425 1048.035 6702.705 1186.305 ;
      RECT 6701.865 1046.935 6702.145 1186.065 ;
      RECT 6701.305 1048.035 6701.585 1185.825 ;
      RECT 6700.745 1046.935 6701.025 1185.585 ;
      RECT 6700.185 1048.035 6700.465 1185.345 ;
      RECT 6686.185 1046.935 6686.465 1191.465 ;
      RECT 6685.625 1048.035 6685.905 1191.225 ;
      RECT 6685.065 1048.035 6685.345 1190.985 ;
      RECT 6684.505 1048.035 6684.785 1190.745 ;
      RECT 6683.945 1048.035 6684.225 1190.505 ;
      RECT 6683.385 1048.035 6683.665 1190.265 ;
      RECT 6682.825 1048.035 6683.105 1190.025 ;
      RECT 6682.265 1048.035 6682.545 1189.785 ;
      RECT 6681.705 1048.035 6681.985 1189.545 ;
      RECT 6681.145 1046.935 6681.425 1189.305 ;
      RECT 6680.585 1048.035 6680.865 1189.065 ;
      RECT 6680.025 1046.935 6680.305 1188.825 ;
      RECT 6679.465 1048.035 6679.745 1188.585 ;
      RECT 6678.905 1048.035 6679.185 1188.345 ;
      RECT 6678.345 1048.035 6678.625 1188.105 ;
      RECT 6677.785 1048.035 6678.065 1187.865 ;
      RECT 6677.225 1048.035 6677.505 1187.625 ;
      RECT 6676.665 1048.035 6676.945 1187.385 ;
      RECT 6676.105 1048.035 6676.385 1187.145 ;
      RECT 6675.545 1048.035 6675.825 1186.905 ;
      RECT 6674.985 1048.035 6675.265 1186.665 ;
      RECT 6674.425 1048.035 6674.705 1186.425 ;
      RECT 6673.865 1048.035 6674.145 1186.185 ;
      RECT 6634.665 1048.035 6634.945 1193.09 ;
      RECT 6634.105 1048.035 6634.385 1193.33 ;
      RECT 6633.545 1048.035 6633.825 1193.57 ;
      RECT 6632.985 1046.935 6633.265 1193.81 ;
      RECT 6632.425 1048.035 6632.705 1194.05 ;
      RECT 6631.865 1046.935 6632.145 1194.29 ;
      RECT 6631.305 1048.035 6631.585 1194.53 ;
      RECT 6630.745 1048.035 6631.025 1194.77 ;
      RECT 6630.185 1048.035 6630.465 1195.01 ;
      RECT 6629.625 1046.935 6629.905 1195.25 ;
      RECT 6629.065 1048.035 6629.345 1195.49 ;
      RECT 6628.505 1046.935 6628.785 1195.73 ;
      RECT 6627.945 1048.035 6628.225 1195.97 ;
      RECT 6627.385 1046.935 6627.665 1196.21 ;
      RECT 6626.825 1048.035 6627.105 1196.45 ;
      RECT 6626.265 1048.035 6626.545 1196.69 ;
      RECT 6625.705 1048.035 6625.985 1196.69 ;
      RECT 6625.145 1048.035 6625.425 1196.45 ;
      RECT 6624.585 1048.035 6624.865 1196.21 ;
      RECT 6624.025 1048.035 6624.305 1195.97 ;
      RECT 6623.465 1048.035 6623.745 1195.73 ;
      RECT 6622.905 1048.035 6623.185 1195.49 ;
      RECT 6622.345 1048.035 6622.625 1195.25 ;
      RECT 6621.785 1048.035 6622.065 1195.01 ;
      RECT 6621.225 1048.035 6621.505 1194.77 ;
      RECT 6612.265 1048.035 6612.545 1194.285 ;
      RECT 6611.705 1046.935 6611.985 1194.045 ;
      RECT 6611.145 1048.035 6611.425 1193.805 ;
      RECT 6610.585 1046.935 6610.865 1193.565 ;
      RECT 6610.025 1048.035 6610.305 1193.325 ;
      RECT 6609.465 1046.935 6609.745 1193.085 ;
      RECT 6608.905 1048.035 6609.185 1192.845 ;
      RECT 6608.345 1048.035 6608.625 1192.605 ;
      RECT 6607.785 1048.035 6608.065 1192.365 ;
      RECT 6607.225 1048.035 6607.505 1192.125 ;
      RECT 6606.665 1048.035 6606.945 1191.885 ;
      RECT 6606.105 1048.035 6606.385 1191.645 ;
      RECT 6605.545 1048.035 6605.825 1191.405 ;
      RECT 6604.985 1048.035 6605.265 1191.165 ;
      RECT 6602.465 1046.935 6602.745 1192.885 ;
      RECT 6601.905 1048.035 6602.185 1192.645 ;
      RECT 6601.345 1046.935 6601.625 1192.405 ;
      RECT 6600.785 1048.035 6601.065 1192.165 ;
      RECT 6600.225 1048.035 6600.505 1191.925 ;
      RECT 6599.665 1048.035 6599.945 1191.685 ;
      RECT 6599.105 1048.035 6599.385 1191.445 ;
      RECT 6598.545 1048.035 6598.825 1191.205 ;
      RECT 6572.505 1048.035 6572.785 1188.855 ;
      RECT 6571.945 1048.035 6572.225 1189.095 ;
      RECT 6571.385 1048.035 6571.665 1189.335 ;
      RECT 6570.825 1048.035 6571.105 1189.58 ;
      RECT 6570.265 1048.035 6570.545 1189.82 ;
      RECT 6569.705 1048.035 6569.985 1190.06 ;
      RECT 6569.145 1048.035 6569.425 1190.06 ;
      RECT 6568.585 1048.035 6568.865 1189.82 ;
      RECT 6568.025 1048.035 6568.305 1189.58 ;
      RECT 6567.465 1046.935 6567.745 1189.34 ;
      RECT 6566.905 1048.035 6567.185 1189.1 ;
      RECT 6566.345 1046.935 6566.625 1188.86 ;
      RECT 6565.785 1048.035 6566.065 1188.62 ;
      RECT 6565.225 1048.035 6565.505 1188.38 ;
      RECT 6564.665 1048.035 6564.945 1188.14 ;
      RECT 6564.105 1046.935 6564.385 1187.9 ;
      RECT 6563.545 1048.035 6563.825 1187.66 ;
      RECT 6562.985 1046.935 6563.265 1187.42 ;
      RECT 6562.425 1048.035 6562.705 1187.18 ;
      RECT 6561.865 1046.935 6562.145 1186.94 ;
      RECT 6561.305 1048.035 6561.585 1186.7 ;
      RECT 6560.745 1048.035 6561.025 1186.46 ;
      RECT 6560.185 1048.035 6560.465 1186.22 ;
      RECT 6559.625 1048.035 6559.905 1185.98 ;
      RECT 6546.185 1048.035 6546.465 1191.78 ;
      RECT 6545.625 1048.035 6545.905 1191.54 ;
      RECT 6545.065 1048.035 6545.345 1191.3 ;
      RECT 6544.505 1048.035 6544.785 1191.06 ;
      RECT 6543.945 1048.035 6544.225 1190.82 ;
      RECT 6543.385 1048.035 6543.665 1190.58 ;
      RECT 6542.825 1048.035 6543.105 1190.34 ;
      RECT 6542.265 1048.035 6542.545 1190.1 ;
      RECT 6541.705 1046.935 6541.985 1189.86 ;
      RECT 6541.145 1048.035 6541.425 1189.62 ;
      RECT 6540.585 1046.935 6540.865 1189.3 ;
      RECT 6540.025 1048.035 6540.305 1189.14 ;
      RECT 6539.465 1046.935 6539.745 1188.9 ;
      RECT 6538.905 1048.035 6539.185 1188.66 ;
      RECT 6538.345 1048.035 6538.625 1188.42 ;
      RECT 6537.785 1048.035 6538.065 1188.18 ;
      RECT 6537.225 1048.035 6537.505 1187.94 ;
      RECT 6536.665 1048.035 6536.945 1187.7 ;
      RECT 6536.105 1048.035 6536.385 1187.46 ;
      RECT 6535.545 1048.035 6535.825 1187.22 ;
      RECT 6534.985 1048.035 6535.265 1186.98 ;
      RECT 6534.425 1046.935 6534.705 1186.74 ;
      RECT 6533.865 1048.035 6534.145 1186.5 ;
      RECT 6533.305 1046.935 6533.585 1186.26 ;
      RECT 6494.105 1048.035 6494.385 1191.87 ;
      RECT 6493.545 1048.035 6493.825 1192.11 ;
      RECT 6492.985 1048.035 6493.265 1192.35 ;
      RECT 6492.425 1048.035 6492.705 1192.59 ;
      RECT 6491.865 1048.035 6492.145 1192.83 ;
      RECT 6491.305 1048.035 6491.585 1193.07 ;
      RECT 6490.745 1048.035 6491.025 1193.31 ;
      RECT 6490.185 1048.035 6490.465 1193.55 ;
      RECT 6489.625 1048.035 6489.905 1193.79 ;
      RECT 6489.065 1048.035 6489.345 1194.03 ;
      RECT 6488.505 1048.035 6488.785 1194.27 ;
      RECT 6487.945 1048.035 6488.225 1194.51 ;
      RECT 6487.385 1048.035 6487.665 1194.75 ;
      RECT 6486.825 1048.035 6487.105 1194.75 ;
      RECT 6486.265 1046.935 6486.545 1194.51 ;
      RECT 6485.705 1048.035 6485.985 1194.27 ;
      RECT 6485.145 1046.935 6485.425 1194.03 ;
      RECT 6484.585 1048.035 6484.865 1193.79 ;
      RECT 6484.025 1048.035 6484.305 1193.55 ;
      RECT 6483.465 1048.035 6483.745 1193.31 ;
      RECT 6482.905 1046.935 6483.185 1193.045 ;
      RECT 6482.345 1048.035 6482.625 1192.805 ;
      RECT 6481.785 1046.935 6482.065 1192.565 ;
      RECT 6481.225 1048.035 6481.505 1192.325 ;
      RECT 6472.265 1046.935 6472.545 1186.16 ;
      RECT 6471.705 1048.035 6471.985 1186.4 ;
      RECT 6471.145 1048.035 6471.425 1186.64 ;
      RECT 6470.585 1048.035 6470.865 1186.64 ;
      RECT 6470.025 1048.035 6470.305 1186.4 ;
      RECT 6469.465 1048.035 6469.745 1186.16 ;
      RECT 6468.905 1048.035 6469.185 1185.92 ;
      RECT 6468.345 1048.035 6468.625 1185.68 ;
      RECT 6467.785 1048.035 6468.065 1185.44 ;
      RECT 6467.225 1048.035 6467.505 1185.2 ;
      RECT 6466.665 1048.035 6466.945 1184.96 ;
      RECT 6466.105 1048.035 6466.385 1184.72 ;
      RECT 6465.545 1048.035 6465.825 1184.48 ;
      RECT 6464.985 1046.935 6465.265 1184.24 ;
      RECT 6462.465 1048.035 6462.745 1185.96 ;
      RECT 6461.905 1046.935 6462.185 1185.72 ;
      RECT 6461.345 1048.035 6461.625 1185.48 ;
      RECT 6460.785 1046.935 6461.065 1185.24 ;
      RECT 6460.225 1048.035 6460.505 1185 ;
      RECT 6459.665 1048.035 6459.945 1184.76 ;
      RECT 6459.105 1048.035 6459.385 1184.52 ;
      RECT 6433.065 1048.035 6433.345 1187.305 ;
      RECT 6432.505 1048.035 6432.785 1187.545 ;
      RECT 6431.945 1048.035 6432.225 1187.785 ;
      RECT 6431.385 1048.035 6431.665 1188.025 ;
      RECT 6430.825 1048.035 6431.105 1188.265 ;
      RECT 6430.265 1046.935 6430.545 1188.505 ;
      RECT 6429.705 1048.035 6429.985 1188.745 ;
      RECT 6429.145 1046.935 6429.425 1188.985 ;
      RECT 6428.585 1048.035 6428.865 1189.225 ;
      RECT 6428.025 1048.035 6428.305 1189.465 ;
      RECT 6427.465 1048.035 6427.745 1189.705 ;
      RECT 6426.905 1048.035 6427.185 1189.945 ;
      RECT 6426.345 1048.035 6426.625 1190.185 ;
      RECT 6425.785 1048.035 6426.065 1190.425 ;
      RECT 6425.225 1048.035 6425.505 1190.665 ;
      RECT 6424.665 1048.035 6424.945 1190.665 ;
      RECT 6424.105 1048.035 6424.385 1190.425 ;
      RECT 6423.545 1048.035 6423.825 1190.185 ;
      RECT 6422.985 1048.035 6423.265 1189.945 ;
      RECT 6422.425 1048.035 6422.705 1189.7 ;
      RECT 6421.865 1048.035 6422.145 1189.46 ;
      RECT 6421.305 1048.035 6421.585 1189.22 ;
      RECT 6420.745 1046.935 6421.025 1188.98 ;
      RECT 6420.185 1048.035 6420.465 1188.74 ;
      RECT 6406.745 1046.935 6407.025 1186.22 ;
      RECT 6406.185 1048.035 6406.465 1185.98 ;
      RECT 6405.625 1048.035 6405.905 1185.74 ;
      RECT 6405.065 1048.035 6405.345 1185.5 ;
      RECT 6404.505 1046.935 6404.785 1185.26 ;
      RECT 6403.945 1048.035 6404.225 1185.02 ;
      RECT 6403.385 1046.935 6403.665 1184.78 ;
      RECT 6402.825 1048.035 6403.105 1184.54 ;
      RECT 6402.265 1046.935 6402.545 1184.3 ;
      RECT 6401.705 1048.035 6401.985 1184.06 ;
      RECT 6401.145 1048.035 6401.425 1183.82 ;
      RECT 6400.585 1048.035 6400.865 1183.58 ;
      RECT 6400.025 1048.035 6400.305 1183.34 ;
      RECT 6399.465 1048.035 6399.745 1183.1 ;
      RECT 6398.905 1048.035 6399.185 1182.86 ;
      RECT 6398.345 1048.035 6398.625 1182.62 ;
      RECT 6397.785 1048.035 6398.065 1182.38 ;
      RECT 6397.225 1048.035 6397.505 1182.14 ;
      RECT 6396.665 1048.035 6396.945 1181.9 ;
      RECT 6396.105 1048.035 6396.385 1181.66 ;
      RECT 6395.545 1048.035 6395.825 1181.42 ;
      RECT 6394.985 1046.935 6395.265 1181.18 ;
      RECT 6394.425 1048.035 6394.705 1180.94 ;
      RECT 6393.865 1046.935 6394.145 1180.7 ;
      RECT 6354.105 1048.035 6354.385 1191.17 ;
      RECT 6353.545 1046.935 6353.825 1191.41 ;
      RECT 6352.985 1048.035 6353.265 1191.65 ;
      RECT 6352.425 1048.035 6352.705 1191.89 ;
      RECT 6351.865 1048.035 6352.145 1192.13 ;
      RECT 6351.305 1048.035 6351.585 1192.37 ;
      RECT 6350.745 1048.035 6351.025 1192.61 ;
      RECT 6350.185 1048.035 6350.465 1192.855 ;
      RECT 6349.625 1048.035 6349.905 1193.095 ;
      RECT 6349.065 1048.035 6349.345 1193.335 ;
      RECT 6348.505 1046.935 6348.785 1193.575 ;
      RECT 6347.945 1048.035 6348.225 1193.815 ;
      RECT 6347.385 1046.935 6347.665 1194.055 ;
      RECT 6346.825 1048.035 6347.105 1194.295 ;
      RECT 6346.265 1048.035 6346.545 1194.535 ;
      RECT 6345.705 1048.035 6345.985 1194.775 ;
      RECT 6345.145 1048.035 6345.425 1195.015 ;
      RECT 6344.585 1048.035 6344.865 1195.255 ;
      RECT 6344.025 1048.035 6344.305 1195.495 ;
      RECT 6343.465 1048.035 6343.745 1195.735 ;
      RECT 6342.905 1048.035 6343.185 1195.975 ;
      RECT 6342.345 1048.035 6342.625 1196.215 ;
      RECT 6341.785 1048.035 6342.065 1196.455 ;
      RECT 6341.225 1048.035 6341.505 1196.695 ;
      RECT 6332.265 1048.035 6332.545 1192.28 ;
      RECT 6331.705 1048.035 6331.985 1192.04 ;
      RECT 6331.145 1048.035 6331.425 1191.8 ;
      RECT 6330.585 1046.935 6330.865 1191.56 ;
      RECT 6330.025 1048.035 6330.305 1191.32 ;
      RECT 6329.465 1046.935 6329.745 1191.08 ;
      RECT 6328.905 1048.035 6329.185 1190.84 ;
      RECT 6328.345 1048.035 6328.625 1190.6 ;
      RECT 6327.785 1048.035 6328.065 1190.36 ;
      RECT 6327.225 1046.935 6327.505 1190.12 ;
      RECT 6326.665 1048.035 6326.945 1189.88 ;
      RECT 6326.105 1046.935 6326.385 1189.64 ;
      RECT 6325.545 1048.035 6325.825 1189.4 ;
      RECT 6324.985 1046.935 6325.265 1189.16 ;
      RECT 6322.465 1048.035 6322.745 1181.56 ;
      RECT 6321.905 1048.035 6322.185 1181.32 ;
      RECT 6321.345 1048.035 6321.625 1181.08 ;
      RECT 6320.785 1048.035 6321.065 1180.84 ;
      RECT 6320.225 1048.035 6320.505 1180.6 ;
      RECT 6319.665 1048.035 6319.945 1180.36 ;
      RECT 6319.105 1048.035 6319.385 1180.12 ;
      RECT 6293.065 1048.035 6293.345 1193.995 ;
      RECT 6292.505 1048.035 6292.785 1194.235 ;
      RECT 6291.945 1048.035 6292.225 1194.475 ;
      RECT 6291.385 1048.035 6291.665 1194.715 ;
      RECT 6290.825 1048.035 6291.105 1194.955 ;
      RECT 6290.265 1046.935 6290.545 1194.955 ;
      RECT 6289.705 1048.035 6289.985 1194.715 ;
      RECT 6289.145 1046.935 6289.425 1194.47 ;
      RECT 6288.585 1048.035 6288.865 1194.23 ;
      RECT 6288.025 1046.935 6288.305 1193.99 ;
      RECT 6287.465 1048.035 6287.745 1193.75 ;
      RECT 6286.905 1048.035 6287.185 1193.51 ;
      RECT 6286.345 1048.035 6286.625 1193.27 ;
      RECT 6285.785 1048.035 6286.065 1193.03 ;
      RECT 6285.225 1048.035 6285.505 1192.79 ;
      RECT 6284.665 1048.035 6284.945 1192.55 ;
      RECT 6284.105 1048.035 6284.385 1192.31 ;
      RECT 6283.545 1048.035 6283.825 1192.07 ;
      RECT 6282.985 1046.935 6283.265 1191.83 ;
      RECT 6282.425 1048.035 6282.705 1191.59 ;
      RECT 6281.865 1046.935 6282.145 1191.35 ;
      RECT 6281.305 1048.035 6281.585 1191.11 ;
      RECT 6280.745 1048.035 6281.025 1190.87 ;
      RECT 6280.185 1048.035 6280.465 1190.63 ;
      RECT 6266.745 1048.035 6267.025 1194.03 ;
      RECT 6266.185 1048.035 6266.465 1194.27 ;
      RECT 6265.625 1048.035 6265.905 1194.515 ;
      RECT 6265.065 1048.035 6265.345 1194.755 ;
      RECT 6264.505 1048.035 6264.785 1194.995 ;
      RECT 6263.945 1048.035 6264.225 1194.995 ;
      RECT 6263.385 1048.035 6263.665 1194.755 ;
      RECT 6262.825 1048.035 6263.105 1194.515 ;
      RECT 6262.265 1048.035 6262.545 1187.5 ;
      RECT 6261.705 1048.035 6261.985 1187.26 ;
      RECT 6261.145 1048.035 6261.425 1187.02 ;
      RECT 6260.585 1046.935 6260.865 1186.78 ;
      RECT 6260.025 1048.035 6260.305 1186.54 ;
      RECT 6259.465 1046.935 6259.745 1186.3 ;
      RECT 6258.905 1048.035 6259.185 1186.06 ;
      RECT 6258.345 1048.035 6258.625 1185.82 ;
      RECT 6257.785 1048.035 6258.065 1185.58 ;
      RECT 6257.225 1046.935 6257.505 1185.34 ;
      RECT 6256.665 1048.035 6256.945 1185.1 ;
      RECT 6256.105 1046.935 6256.385 1184.86 ;
      RECT 6255.545 1048.035 6255.825 1184.62 ;
      RECT 6254.985 1046.935 6255.265 1184.38 ;
      RECT 6254.425 1048.035 6254.705 1184.14 ;
      RECT 6253.865 1048.035 6254.145 1183.9 ;
      RECT 6213.545 1048.035 6213.825 1192.795 ;
      RECT 6212.985 1048.035 6213.265 1193.035 ;
      RECT 6212.425 1048.035 6212.705 1193.28 ;
      RECT 6211.865 1048.035 6212.145 1193.52 ;
      RECT 6211.305 1048.035 6211.585 1193.76 ;
      RECT 6210.745 1048.035 6211.025 1194 ;
      RECT 6210.185 1048.035 6210.465 1194.24 ;
      RECT 6209.625 1048.035 6209.905 1194.48 ;
      RECT 6209.065 1048.035 6209.345 1194.72 ;
      RECT 6208.505 1048.035 6208.785 1194.96 ;
      RECT 6207.945 1046.935 6208.225 1195.2 ;
      RECT 6207.385 1048.035 6207.665 1195.44 ;
      RECT 6206.825 1046.935 6207.105 1195.68 ;
      RECT 6206.265 1048.035 6206.545 1195.92 ;
      RECT 6205.705 1046.935 6205.985 1196.16 ;
      RECT 6205.145 1048.035 6205.425 1196.16 ;
      RECT 6204.585 1048.035 6204.865 1195.92 ;
      RECT 6204.025 1048.035 6204.305 1195.68 ;
      RECT 6203.465 1048.035 6203.745 1195.44 ;
      RECT 6202.905 1048.035 6203.185 1195.2 ;
      RECT 6202.345 1048.035 6202.625 1194.96 ;
      RECT 6201.785 1048.035 6202.065 1194.72 ;
      RECT 6201.225 1048.035 6201.505 1194.48 ;
      RECT 6192.265 1046.935 6192.545 1194.51 ;
      RECT 6191.705 1048.035 6191.985 1194.75 ;
      RECT 6191.145 1046.935 6191.425 1194.99 ;
      RECT 6190.585 1048.035 6190.865 1195.205 ;
      RECT 6190.025 1048.035 6190.305 1194.78 ;
      RECT 6189.465 1048.035 6189.745 1194.54 ;
      RECT 6188.905 1048.035 6189.185 1194.3 ;
      RECT 6188.345 1048.035 6188.625 1194.06 ;
      RECT 6187.785 1048.035 6188.065 1193.82 ;
      RECT 6187.225 1048.035 6187.505 1193.58 ;
      RECT 6186.665 1048.035 6186.945 1193.34 ;
      RECT 6186.105 1048.035 6186.385 1193.1 ;
      RECT 6185.545 1048.035 6185.825 1192.86 ;
      RECT 6184.985 1048.035 6185.265 1192.62 ;
      RECT 6182.465 1048.035 6182.745 1191.795 ;
      RECT 6181.905 1048.035 6182.185 1191.555 ;
      RECT 6181.345 1048.035 6181.625 1191.315 ;
      RECT 6180.785 1046.935 6181.065 1191.075 ;
      RECT 6180.225 1048.035 6180.505 1190.835 ;
      RECT 6179.665 1046.935 6179.945 1190.595 ;
      RECT 6179.105 1048.035 6179.385 1190.355 ;
      RECT 6178.545 1048.035 6178.825 1190.115 ;
      RECT 6151.945 1048.035 6152.225 1201.16 ;
      RECT 6151.385 1046.935 6151.665 1201.4 ;
      RECT 6150.825 1048.035 6151.105 1201.64 ;
      RECT 6150.265 1046.935 6150.545 1201.885 ;
      RECT 6149.705 1048.035 6149.985 1202.125 ;
      RECT 6149.145 1046.935 6149.425 1202.365 ;
      RECT 6148.585 1048.035 6148.865 1202.605 ;
      RECT 6148.025 1048.035 6148.305 1202.845 ;
      RECT 6147.465 1048.035 6147.745 1188.465 ;
      RECT 6146.905 1048.035 6147.185 1188.225 ;
      RECT 6146.345 1048.035 6146.625 1187.985 ;
      RECT 6145.785 1048.035 6146.065 1187.745 ;
      RECT 6145.225 1048.035 6145.505 1187.505 ;
      RECT 6144.665 1048.035 6144.945 1187.265 ;
      RECT 6144.105 1048.035 6144.385 1187.025 ;
      RECT 6143.545 1048.035 6143.825 1186.785 ;
      RECT 6142.985 1048.035 6143.265 1186.545 ;
      RECT 6142.425 1048.035 6142.705 1186.305 ;
      RECT 6141.865 1046.935 6142.145 1186.065 ;
      RECT 6141.305 1048.035 6141.585 1185.825 ;
      RECT 6140.745 1046.935 6141.025 1185.585 ;
      RECT 6140.185 1048.035 6140.465 1185.345 ;
      RECT 6126.185 1046.935 6126.465 1191.465 ;
      RECT 6125.625 1048.035 6125.905 1191.225 ;
      RECT 6125.065 1048.035 6125.345 1190.985 ;
      RECT 6124.505 1048.035 6124.785 1190.745 ;
      RECT 6123.945 1048.035 6124.225 1190.505 ;
      RECT 6123.385 1048.035 6123.665 1190.265 ;
      RECT 6122.825 1048.035 6123.105 1190.025 ;
      RECT 6122.265 1048.035 6122.545 1189.785 ;
      RECT 6121.705 1048.035 6121.985 1189.545 ;
      RECT 6121.145 1046.935 6121.425 1189.305 ;
      RECT 6120.585 1048.035 6120.865 1189.065 ;
      RECT 6120.025 1046.935 6120.305 1188.825 ;
      RECT 6119.465 1048.035 6119.745 1188.585 ;
      RECT 6118.905 1048.035 6119.185 1188.345 ;
      RECT 6118.345 1048.035 6118.625 1188.105 ;
      RECT 6117.785 1048.035 6118.065 1187.865 ;
      RECT 6117.225 1048.035 6117.505 1187.625 ;
      RECT 6116.665 1048.035 6116.945 1187.385 ;
      RECT 6116.105 1048.035 6116.385 1187.145 ;
      RECT 6115.545 1048.035 6115.825 1186.905 ;
      RECT 6114.985 1048.035 6115.265 1186.665 ;
      RECT 6114.425 1048.035 6114.705 1186.425 ;
      RECT 6113.865 1048.035 6114.145 1186.185 ;
      RECT 6074.665 1048.035 6074.945 1193.09 ;
      RECT 6074.105 1048.035 6074.385 1193.33 ;
      RECT 6073.545 1048.035 6073.825 1193.57 ;
      RECT 6072.985 1046.935 6073.265 1193.81 ;
      RECT 6072.425 1048.035 6072.705 1194.05 ;
      RECT 6071.865 1046.935 6072.145 1194.29 ;
      RECT 6071.305 1048.035 6071.585 1194.53 ;
      RECT 6070.745 1048.035 6071.025 1194.77 ;
      RECT 6070.185 1048.035 6070.465 1195.01 ;
      RECT 6069.625 1046.935 6069.905 1195.25 ;
      RECT 6069.065 1048.035 6069.345 1195.49 ;
      RECT 6068.505 1046.935 6068.785 1195.73 ;
      RECT 6067.945 1048.035 6068.225 1195.97 ;
      RECT 6067.385 1046.935 6067.665 1196.21 ;
      RECT 6066.825 1048.035 6067.105 1196.45 ;
      RECT 6066.265 1048.035 6066.545 1196.69 ;
      RECT 6065.705 1048.035 6065.985 1196.69 ;
      RECT 6065.145 1048.035 6065.425 1196.45 ;
      RECT 6064.585 1048.035 6064.865 1196.21 ;
      RECT 6064.025 1048.035 6064.305 1195.97 ;
      RECT 6063.465 1048.035 6063.745 1195.73 ;
      RECT 6062.905 1048.035 6063.185 1195.49 ;
      RECT 6062.345 1048.035 6062.625 1195.25 ;
      RECT 6061.785 1048.035 6062.065 1195.01 ;
      RECT 6061.225 1048.035 6061.505 1194.77 ;
      RECT 6052.265 1048.035 6052.545 1194.285 ;
      RECT 6051.705 1046.935 6051.985 1194.045 ;
      RECT 6051.145 1048.035 6051.425 1193.805 ;
      RECT 6050.585 1046.935 6050.865 1193.565 ;
      RECT 6050.025 1048.035 6050.305 1193.325 ;
      RECT 6049.465 1046.935 6049.745 1193.085 ;
      RECT 6048.905 1048.035 6049.185 1192.845 ;
      RECT 6048.345 1048.035 6048.625 1192.605 ;
      RECT 6047.785 1048.035 6048.065 1192.365 ;
      RECT 6047.225 1048.035 6047.505 1192.125 ;
      RECT 6046.665 1048.035 6046.945 1191.885 ;
      RECT 6046.105 1048.035 6046.385 1191.645 ;
      RECT 6045.545 1048.035 6045.825 1191.405 ;
      RECT 6044.985 1048.035 6045.265 1191.165 ;
      RECT 6042.465 1046.935 6042.745 1192.885 ;
      RECT 6041.905 1048.035 6042.185 1192.645 ;
      RECT 6041.345 1046.935 6041.625 1192.405 ;
      RECT 6040.785 1048.035 6041.065 1192.165 ;
      RECT 6040.225 1048.035 6040.505 1191.925 ;
      RECT 6039.665 1048.035 6039.945 1191.685 ;
      RECT 6039.105 1048.035 6039.385 1191.445 ;
      RECT 6038.545 1048.035 6038.825 1191.205 ;
      RECT 6012.505 1048.035 6012.785 1188.855 ;
      RECT 6011.945 1048.035 6012.225 1189.095 ;
      RECT 6011.385 1048.035 6011.665 1189.335 ;
      RECT 6010.825 1048.035 6011.105 1189.58 ;
      RECT 6010.265 1048.035 6010.545 1189.82 ;
      RECT 6009.705 1048.035 6009.985 1190.06 ;
      RECT 6009.145 1048.035 6009.425 1190.06 ;
      RECT 6008.585 1048.035 6008.865 1189.82 ;
      RECT 6008.025 1048.035 6008.305 1189.58 ;
      RECT 6007.465 1046.935 6007.745 1189.34 ;
      RECT 6006.905 1048.035 6007.185 1189.1 ;
      RECT 6006.345 1046.935 6006.625 1188.86 ;
      RECT 6005.785 1048.035 6006.065 1188.62 ;
      RECT 6005.225 1048.035 6005.505 1188.38 ;
      RECT 6004.665 1048.035 6004.945 1188.14 ;
      RECT 6004.105 1046.935 6004.385 1187.9 ;
      RECT 6003.545 1048.035 6003.825 1187.66 ;
      RECT 6002.985 1046.935 6003.265 1187.42 ;
      RECT 6002.425 1048.035 6002.705 1187.18 ;
      RECT 6001.865 1046.935 6002.145 1186.94 ;
      RECT 6001.305 1048.035 6001.585 1186.7 ;
      RECT 6000.745 1048.035 6001.025 1186.46 ;
      RECT 6000.185 1048.035 6000.465 1186.22 ;
      RECT 5999.625 1048.035 5999.905 1185.98 ;
      RECT 5986.185 1048.035 5986.465 1191.78 ;
      RECT 5985.625 1048.035 5985.905 1191.54 ;
      RECT 5985.065 1048.035 5985.345 1191.3 ;
      RECT 5984.505 1048.035 5984.785 1191.06 ;
      RECT 5983.945 1048.035 5984.225 1190.82 ;
      RECT 5983.385 1048.035 5983.665 1190.58 ;
      RECT 5982.825 1048.035 5983.105 1190.34 ;
      RECT 5982.265 1048.035 5982.545 1190.1 ;
      RECT 5981.705 1046.935 5981.985 1189.86 ;
      RECT 5981.145 1048.035 5981.425 1189.62 ;
      RECT 5980.585 1046.935 5980.865 1189.3 ;
      RECT 5980.025 1048.035 5980.305 1189.14 ;
      RECT 5979.465 1046.935 5979.745 1188.9 ;
      RECT 5978.905 1048.035 5979.185 1188.66 ;
      RECT 5978.345 1048.035 5978.625 1188.42 ;
      RECT 5977.785 1048.035 5978.065 1188.18 ;
      RECT 5977.225 1048.035 5977.505 1187.94 ;
      RECT 5976.665 1048.035 5976.945 1187.7 ;
      RECT 5976.105 1048.035 5976.385 1187.46 ;
      RECT 5975.545 1048.035 5975.825 1187.22 ;
      RECT 5974.985 1048.035 5975.265 1186.98 ;
      RECT 5974.425 1046.935 5974.705 1186.74 ;
      RECT 5973.865 1048.035 5974.145 1186.5 ;
      RECT 5973.305 1046.935 5973.585 1186.26 ;
      RECT 5934.105 1048.035 5934.385 1191.87 ;
      RECT 5933.545 1048.035 5933.825 1192.11 ;
      RECT 5932.985 1048.035 5933.265 1192.35 ;
      RECT 5932.425 1048.035 5932.705 1192.59 ;
      RECT 5931.865 1048.035 5932.145 1192.83 ;
      RECT 5931.305 1048.035 5931.585 1193.07 ;
      RECT 5930.745 1048.035 5931.025 1193.31 ;
      RECT 5930.185 1048.035 5930.465 1193.55 ;
      RECT 5929.625 1048.035 5929.905 1193.79 ;
      RECT 5929.065 1048.035 5929.345 1194.03 ;
      RECT 5928.505 1048.035 5928.785 1194.27 ;
      RECT 5927.945 1048.035 5928.225 1194.51 ;
      RECT 5927.385 1048.035 5927.665 1194.75 ;
      RECT 5926.825 1048.035 5927.105 1194.75 ;
      RECT 5926.265 1046.935 5926.545 1194.51 ;
      RECT 5925.705 1048.035 5925.985 1194.27 ;
      RECT 5925.145 1046.935 5925.425 1194.03 ;
      RECT 5924.585 1048.035 5924.865 1193.79 ;
      RECT 5924.025 1048.035 5924.305 1193.55 ;
      RECT 5923.465 1048.035 5923.745 1193.31 ;
      RECT 5922.905 1046.935 5923.185 1193.045 ;
      RECT 5922.345 1048.035 5922.625 1192.805 ;
      RECT 5921.785 1046.935 5922.065 1192.565 ;
      RECT 5921.225 1048.035 5921.505 1192.325 ;
      RECT 5912.265 1046.935 5912.545 1186.16 ;
      RECT 5911.705 1048.035 5911.985 1186.4 ;
      RECT 5911.145 1048.035 5911.425 1186.64 ;
      RECT 5910.585 1048.035 5910.865 1186.64 ;
      RECT 5910.025 1048.035 5910.305 1186.4 ;
      RECT 5909.465 1048.035 5909.745 1186.16 ;
      RECT 5908.905 1048.035 5909.185 1185.92 ;
      RECT 5908.345 1048.035 5908.625 1185.68 ;
      RECT 5907.785 1048.035 5908.065 1185.44 ;
      RECT 5907.225 1048.035 5907.505 1185.2 ;
      RECT 5906.665 1048.035 5906.945 1184.96 ;
      RECT 5906.105 1048.035 5906.385 1184.72 ;
      RECT 5905.545 1048.035 5905.825 1184.48 ;
      RECT 5904.985 1046.935 5905.265 1184.24 ;
      RECT 5902.465 1048.035 5902.745 1185.96 ;
      RECT 5901.905 1046.935 5902.185 1185.72 ;
      RECT 5901.345 1048.035 5901.625 1185.48 ;
      RECT 5900.785 1046.935 5901.065 1185.24 ;
      RECT 5900.225 1048.035 5900.505 1185 ;
      RECT 5899.665 1048.035 5899.945 1184.76 ;
      RECT 5899.105 1048.035 5899.385 1184.52 ;
      RECT 5873.065 1048.035 5873.345 1187.305 ;
      RECT 5872.505 1048.035 5872.785 1187.545 ;
      RECT 5871.945 1048.035 5872.225 1187.785 ;
      RECT 5871.385 1048.035 5871.665 1188.025 ;
      RECT 5870.825 1048.035 5871.105 1188.265 ;
      RECT 5870.265 1046.935 5870.545 1188.505 ;
      RECT 5869.705 1048.035 5869.985 1188.745 ;
      RECT 5869.145 1046.935 5869.425 1188.985 ;
      RECT 5868.585 1048.035 5868.865 1189.225 ;
      RECT 5868.025 1048.035 5868.305 1189.465 ;
      RECT 5867.465 1048.035 5867.745 1189.705 ;
      RECT 5866.905 1048.035 5867.185 1189.945 ;
      RECT 5866.345 1048.035 5866.625 1190.185 ;
      RECT 5865.785 1048.035 5866.065 1190.425 ;
      RECT 5865.225 1048.035 5865.505 1190.665 ;
      RECT 5864.665 1048.035 5864.945 1190.665 ;
      RECT 5864.105 1048.035 5864.385 1190.425 ;
      RECT 5863.545 1048.035 5863.825 1190.185 ;
      RECT 5862.985 1048.035 5863.265 1189.945 ;
      RECT 5862.425 1048.035 5862.705 1189.7 ;
      RECT 5861.865 1048.035 5862.145 1189.46 ;
      RECT 5861.305 1048.035 5861.585 1189.22 ;
      RECT 5860.745 1046.935 5861.025 1188.98 ;
      RECT 5860.185 1048.035 5860.465 1188.74 ;
      RECT 5846.745 1046.935 5847.025 1186.22 ;
      RECT 5846.185 1048.035 5846.465 1185.98 ;
      RECT 5845.625 1048.035 5845.905 1185.74 ;
      RECT 5845.065 1048.035 5845.345 1185.5 ;
      RECT 5844.505 1046.935 5844.785 1185.26 ;
      RECT 5843.945 1048.035 5844.225 1185.02 ;
      RECT 5843.385 1046.935 5843.665 1184.78 ;
      RECT 5842.825 1048.035 5843.105 1184.54 ;
      RECT 5842.265 1046.935 5842.545 1184.3 ;
      RECT 5841.705 1048.035 5841.985 1184.06 ;
      RECT 5841.145 1048.035 5841.425 1183.82 ;
      RECT 5840.585 1048.035 5840.865 1183.58 ;
      RECT 5840.025 1048.035 5840.305 1183.34 ;
      RECT 5839.465 1048.035 5839.745 1183.1 ;
      RECT 5838.905 1048.035 5839.185 1182.86 ;
      RECT 5838.345 1048.035 5838.625 1182.62 ;
      RECT 5837.785 1048.035 5838.065 1182.38 ;
      RECT 5837.225 1048.035 5837.505 1182.14 ;
      RECT 5836.665 1048.035 5836.945 1181.9 ;
      RECT 5836.105 1048.035 5836.385 1181.66 ;
      RECT 5835.545 1048.035 5835.825 1181.42 ;
      RECT 5834.985 1046.935 5835.265 1181.18 ;
      RECT 5834.425 1048.035 5834.705 1180.94 ;
      RECT 5833.865 1046.935 5834.145 1180.7 ;
      RECT 5794.105 1048.035 5794.385 1191.17 ;
      RECT 5793.545 1046.935 5793.825 1191.41 ;
      RECT 5792.985 1048.035 5793.265 1191.65 ;
      RECT 5792.425 1048.035 5792.705 1191.89 ;
      RECT 5791.865 1048.035 5792.145 1192.13 ;
      RECT 5791.305 1048.035 5791.585 1192.37 ;
      RECT 5790.745 1048.035 5791.025 1192.61 ;
      RECT 5790.185 1048.035 5790.465 1192.855 ;
      RECT 5789.625 1048.035 5789.905 1193.095 ;
      RECT 5789.065 1048.035 5789.345 1193.335 ;
      RECT 5788.505 1046.935 5788.785 1193.575 ;
      RECT 5787.945 1048.035 5788.225 1193.815 ;
      RECT 5787.385 1046.935 5787.665 1194.055 ;
      RECT 5786.825 1048.035 5787.105 1194.295 ;
      RECT 5786.265 1048.035 5786.545 1194.535 ;
      RECT 5785.705 1048.035 5785.985 1194.775 ;
      RECT 5785.145 1048.035 5785.425 1195.015 ;
      RECT 5784.585 1048.035 5784.865 1195.255 ;
      RECT 5784.025 1048.035 5784.305 1195.495 ;
      RECT 5783.465 1048.035 5783.745 1195.735 ;
      RECT 5782.905 1048.035 5783.185 1195.975 ;
      RECT 5782.345 1048.035 5782.625 1196.215 ;
      RECT 5781.785 1048.035 5782.065 1196.455 ;
      RECT 5781.225 1048.035 5781.505 1196.695 ;
      RECT 5772.265 1048.035 5772.545 1192.28 ;
      RECT 5771.705 1048.035 5771.985 1192.04 ;
      RECT 5771.145 1048.035 5771.425 1191.8 ;
      RECT 5770.585 1046.935 5770.865 1191.56 ;
      RECT 5770.025 1048.035 5770.305 1191.32 ;
      RECT 5769.465 1046.935 5769.745 1191.08 ;
      RECT 5768.905 1048.035 5769.185 1190.84 ;
      RECT 5768.345 1048.035 5768.625 1190.6 ;
      RECT 5767.785 1048.035 5768.065 1190.36 ;
      RECT 5767.225 1046.935 5767.505 1190.12 ;
      RECT 5766.665 1048.035 5766.945 1189.88 ;
      RECT 5766.105 1046.935 5766.385 1189.64 ;
      RECT 5765.545 1048.035 5765.825 1189.4 ;
      RECT 5764.985 1046.935 5765.265 1189.16 ;
      RECT 5762.465 1048.035 5762.745 1181.56 ;
      RECT 5761.905 1048.035 5762.185 1181.32 ;
      RECT 5761.345 1048.035 5761.625 1181.08 ;
      RECT 5760.785 1048.035 5761.065 1180.84 ;
      RECT 5760.225 1048.035 5760.505 1180.6 ;
      RECT 5759.665 1048.035 5759.945 1180.36 ;
      RECT 5759.105 1048.035 5759.385 1180.12 ;
      RECT 5733.065 1048.035 5733.345 1193.995 ;
      RECT 5732.505 1048.035 5732.785 1194.235 ;
      RECT 5731.945 1048.035 5732.225 1194.475 ;
      RECT 5731.385 1048.035 5731.665 1194.715 ;
      RECT 5730.825 1048.035 5731.105 1194.955 ;
      RECT 5730.265 1046.935 5730.545 1194.955 ;
      RECT 5729.705 1048.035 5729.985 1194.715 ;
      RECT 5729.145 1046.935 5729.425 1194.47 ;
      RECT 5728.585 1048.035 5728.865 1194.23 ;
      RECT 5728.025 1046.935 5728.305 1193.99 ;
      RECT 5727.465 1048.035 5727.745 1193.75 ;
      RECT 5726.905 1048.035 5727.185 1193.51 ;
      RECT 5726.345 1048.035 5726.625 1193.27 ;
      RECT 5725.785 1048.035 5726.065 1193.03 ;
      RECT 5725.225 1048.035 5725.505 1192.79 ;
      RECT 5724.665 1048.035 5724.945 1192.55 ;
      RECT 5724.105 1048.035 5724.385 1192.31 ;
      RECT 5723.545 1048.035 5723.825 1192.07 ;
      RECT 5722.985 1046.935 5723.265 1191.83 ;
      RECT 5722.425 1048.035 5722.705 1191.59 ;
      RECT 5721.865 1046.935 5722.145 1191.35 ;
      RECT 5721.305 1048.035 5721.585 1191.11 ;
      RECT 5720.745 1048.035 5721.025 1190.87 ;
      RECT 5720.185 1048.035 5720.465 1190.63 ;
      RECT 5706.745 1048.035 5707.025 1194.03 ;
      RECT 5706.185 1048.035 5706.465 1194.27 ;
      RECT 5705.625 1048.035 5705.905 1194.515 ;
      RECT 5705.065 1048.035 5705.345 1194.755 ;
      RECT 5704.505 1048.035 5704.785 1194.995 ;
      RECT 5703.945 1048.035 5704.225 1194.995 ;
      RECT 5703.385 1048.035 5703.665 1194.755 ;
      RECT 5702.825 1048.035 5703.105 1194.515 ;
      RECT 5702.265 1048.035 5702.545 1187.5 ;
      RECT 5701.705 1048.035 5701.985 1187.26 ;
      RECT 5701.145 1048.035 5701.425 1187.02 ;
      RECT 5700.585 1046.935 5700.865 1186.78 ;
      RECT 5700.025 1048.035 5700.305 1186.54 ;
      RECT 5699.465 1046.935 5699.745 1186.3 ;
      RECT 5698.905 1048.035 5699.185 1186.06 ;
      RECT 5698.345 1048.035 5698.625 1185.82 ;
      RECT 5697.785 1048.035 5698.065 1185.58 ;
      RECT 5697.225 1046.935 5697.505 1185.34 ;
      RECT 5696.665 1048.035 5696.945 1185.1 ;
      RECT 5696.105 1046.935 5696.385 1184.86 ;
      RECT 5695.545 1048.035 5695.825 1184.62 ;
      RECT 5694.985 1046.935 5695.265 1184.38 ;
      RECT 5694.425 1048.035 5694.705 1184.14 ;
      RECT 5693.865 1048.035 5694.145 1183.9 ;
      RECT 5653.545 1048.035 5653.825 1192.795 ;
      RECT 5652.985 1048.035 5653.265 1193.035 ;
      RECT 5652.425 1048.035 5652.705 1193.28 ;
      RECT 5651.865 1048.035 5652.145 1193.52 ;
      RECT 5651.305 1048.035 5651.585 1193.76 ;
      RECT 5650.745 1048.035 5651.025 1194 ;
      RECT 5650.185 1048.035 5650.465 1194.24 ;
      RECT 5649.625 1048.035 5649.905 1194.48 ;
      RECT 5649.065 1048.035 5649.345 1194.72 ;
      RECT 5648.505 1048.035 5648.785 1194.96 ;
      RECT 5647.945 1046.935 5648.225 1195.2 ;
      RECT 5647.385 1048.035 5647.665 1195.44 ;
      RECT 5646.825 1046.935 5647.105 1195.68 ;
      RECT 5646.265 1048.035 5646.545 1195.92 ;
      RECT 5645.705 1046.935 5645.985 1196.16 ;
      RECT 5645.145 1048.035 5645.425 1196.16 ;
      RECT 5644.585 1048.035 5644.865 1195.92 ;
      RECT 5644.025 1048.035 5644.305 1195.68 ;
      RECT 5643.465 1048.035 5643.745 1195.44 ;
      RECT 5642.905 1048.035 5643.185 1195.2 ;
      RECT 5642.345 1048.035 5642.625 1194.96 ;
      RECT 5641.785 1048.035 5642.065 1194.72 ;
      RECT 5641.225 1048.035 5641.505 1194.48 ;
      RECT 5632.265 1046.935 5632.545 1194.51 ;
      RECT 5631.705 1048.035 5631.985 1194.75 ;
      RECT 5631.145 1046.935 5631.425 1194.99 ;
      RECT 5630.585 1048.035 5630.865 1195.205 ;
      RECT 5630.025 1048.035 5630.305 1194.78 ;
      RECT 5629.465 1048.035 5629.745 1194.54 ;
      RECT 5628.905 1048.035 5629.185 1194.3 ;
      RECT 5628.345 1048.035 5628.625 1194.06 ;
      RECT 5627.785 1048.035 5628.065 1193.82 ;
      RECT 5627.225 1048.035 5627.505 1193.58 ;
      RECT 5626.665 1048.035 5626.945 1193.34 ;
      RECT 5626.105 1048.035 5626.385 1193.1 ;
      RECT 5625.545 1048.035 5625.825 1192.86 ;
      RECT 5624.985 1048.035 5625.265 1192.62 ;
      RECT 5622.465 1048.035 5622.745 1191.795 ;
      RECT 5621.905 1048.035 5622.185 1191.555 ;
      RECT 5621.345 1048.035 5621.625 1191.315 ;
      RECT 5620.785 1046.935 5621.065 1191.075 ;
      RECT 5620.225 1048.035 5620.505 1190.835 ;
      RECT 5619.665 1046.935 5619.945 1190.595 ;
      RECT 5619.105 1048.035 5619.385 1190.355 ;
      RECT 5618.545 1048.035 5618.825 1190.115 ;
      RECT 5591.945 1048.035 5592.225 1201.16 ;
      RECT 5591.385 1046.935 5591.665 1201.4 ;
      RECT 5590.825 1048.035 5591.105 1201.64 ;
      RECT 5590.265 1046.935 5590.545 1201.885 ;
      RECT 5589.705 1048.035 5589.985 1202.125 ;
      RECT 5589.145 1046.935 5589.425 1202.365 ;
      RECT 5588.585 1048.035 5588.865 1202.605 ;
      RECT 5588.025 1048.035 5588.305 1202.845 ;
      RECT 5587.465 1048.035 5587.745 1188.465 ;
      RECT 5586.905 1048.035 5587.185 1188.225 ;
      RECT 5586.345 1048.035 5586.625 1187.985 ;
      RECT 5585.785 1048.035 5586.065 1187.745 ;
      RECT 5585.225 1048.035 5585.505 1187.505 ;
      RECT 5584.665 1048.035 5584.945 1187.265 ;
      RECT 5584.105 1048.035 5584.385 1187.025 ;
      RECT 5583.545 1048.035 5583.825 1186.785 ;
      RECT 5582.985 1048.035 5583.265 1186.545 ;
      RECT 5582.425 1048.035 5582.705 1186.305 ;
      RECT 5581.865 1046.935 5582.145 1186.065 ;
      RECT 5581.305 1048.035 5581.585 1185.825 ;
      RECT 5580.745 1046.935 5581.025 1185.585 ;
      RECT 5580.185 1048.035 5580.465 1185.345 ;
      RECT 5566.185 1046.935 5566.465 1191.465 ;
      RECT 5565.625 1048.035 5565.905 1191.225 ;
      RECT 5565.065 1048.035 5565.345 1190.985 ;
      RECT 5564.505 1048.035 5564.785 1190.745 ;
      RECT 5563.945 1048.035 5564.225 1190.505 ;
      RECT 5563.385 1048.035 5563.665 1190.265 ;
      RECT 5562.825 1048.035 5563.105 1190.025 ;
      RECT 5562.265 1048.035 5562.545 1189.785 ;
      RECT 5561.705 1048.035 5561.985 1189.545 ;
      RECT 5561.145 1046.935 5561.425 1189.305 ;
      RECT 5560.585 1048.035 5560.865 1189.065 ;
      RECT 5560.025 1046.935 5560.305 1188.825 ;
      RECT 5559.465 1048.035 5559.745 1188.585 ;
      RECT 5558.905 1048.035 5559.185 1188.345 ;
      RECT 5558.345 1048.035 5558.625 1188.105 ;
      RECT 5557.785 1048.035 5558.065 1187.865 ;
      RECT 5557.225 1048.035 5557.505 1187.625 ;
      RECT 5556.665 1048.035 5556.945 1187.385 ;
      RECT 5556.105 1048.035 5556.385 1187.145 ;
      RECT 5555.545 1048.035 5555.825 1186.905 ;
      RECT 5554.985 1048.035 5555.265 1186.665 ;
      RECT 5554.425 1048.035 5554.705 1186.425 ;
      RECT 5553.865 1048.035 5554.145 1186.185 ;
      RECT 5514.665 1048.035 5514.945 1193.09 ;
      RECT 5514.105 1048.035 5514.385 1193.33 ;
      RECT 5513.545 1048.035 5513.825 1193.57 ;
      RECT 5512.985 1046.935 5513.265 1193.81 ;
      RECT 5512.425 1048.035 5512.705 1194.05 ;
      RECT 5511.865 1046.935 5512.145 1194.29 ;
      RECT 5511.305 1048.035 5511.585 1194.53 ;
      RECT 5510.745 1048.035 5511.025 1194.77 ;
      RECT 5510.185 1048.035 5510.465 1195.01 ;
      RECT 5509.625 1046.935 5509.905 1195.25 ;
      RECT 5509.065 1048.035 5509.345 1195.49 ;
      RECT 5508.505 1046.935 5508.785 1195.73 ;
      RECT 5507.945 1048.035 5508.225 1195.97 ;
      RECT 5507.385 1046.935 5507.665 1196.21 ;
      RECT 5506.825 1048.035 5507.105 1196.45 ;
      RECT 5506.265 1048.035 5506.545 1196.69 ;
      RECT 5505.705 1048.035 5505.985 1196.69 ;
      RECT 5505.145 1048.035 5505.425 1196.45 ;
      RECT 5504.585 1048.035 5504.865 1196.21 ;
      RECT 5504.025 1048.035 5504.305 1195.97 ;
      RECT 5503.465 1048.035 5503.745 1195.73 ;
      RECT 5502.905 1048.035 5503.185 1195.49 ;
      RECT 5502.345 1048.035 5502.625 1195.25 ;
      RECT 5501.785 1048.035 5502.065 1195.01 ;
      RECT 5501.225 1048.035 5501.505 1194.77 ;
      RECT 5492.265 1048.035 5492.545 1194.285 ;
      RECT 5491.705 1046.935 5491.985 1194.045 ;
      RECT 5491.145 1048.035 5491.425 1193.805 ;
      RECT 5490.585 1046.935 5490.865 1193.565 ;
      RECT 5490.025 1048.035 5490.305 1193.325 ;
      RECT 5489.465 1046.935 5489.745 1193.085 ;
      RECT 5488.905 1048.035 5489.185 1192.845 ;
      RECT 5488.345 1048.035 5488.625 1192.605 ;
      RECT 5487.785 1048.035 5488.065 1192.365 ;
      RECT 5487.225 1048.035 5487.505 1192.125 ;
      RECT 5486.665 1048.035 5486.945 1191.885 ;
      RECT 5486.105 1048.035 5486.385 1191.645 ;
      RECT 5485.545 1048.035 5485.825 1191.405 ;
      RECT 5484.985 1048.035 5485.265 1191.165 ;
      RECT 5482.465 1046.935 5482.745 1192.885 ;
      RECT 5481.905 1048.035 5482.185 1192.645 ;
      RECT 5481.345 1046.935 5481.625 1192.405 ;
      RECT 5480.785 1048.035 5481.065 1192.165 ;
      RECT 5480.225 1048.035 5480.505 1191.925 ;
      RECT 5479.665 1048.035 5479.945 1191.685 ;
      RECT 5479.105 1048.035 5479.385 1191.445 ;
      RECT 5478.545 1048.035 5478.825 1191.205 ;
      RECT 5452.505 1048.035 5452.785 1188.855 ;
      RECT 5451.945 1048.035 5452.225 1189.095 ;
      RECT 5451.385 1048.035 5451.665 1189.335 ;
      RECT 5450.825 1048.035 5451.105 1189.58 ;
      RECT 5450.265 1048.035 5450.545 1189.82 ;
      RECT 5449.705 1048.035 5449.985 1190.06 ;
      RECT 5449.145 1048.035 5449.425 1190.06 ;
      RECT 5448.585 1048.035 5448.865 1189.82 ;
      RECT 5448.025 1048.035 5448.305 1189.58 ;
      RECT 5447.465 1046.935 5447.745 1189.34 ;
      RECT 5446.905 1048.035 5447.185 1189.1 ;
      RECT 5446.345 1046.935 5446.625 1188.86 ;
      RECT 5445.785 1048.035 5446.065 1188.62 ;
      RECT 5445.225 1048.035 5445.505 1188.38 ;
      RECT 5444.665 1048.035 5444.945 1188.14 ;
      RECT 5444.105 1046.935 5444.385 1187.9 ;
      RECT 5443.545 1048.035 5443.825 1187.66 ;
      RECT 5442.985 1046.935 5443.265 1187.42 ;
      RECT 5442.425 1048.035 5442.705 1187.18 ;
      RECT 5441.865 1046.935 5442.145 1186.94 ;
      RECT 5441.305 1048.035 5441.585 1186.7 ;
      RECT 5440.745 1048.035 5441.025 1186.46 ;
      RECT 5440.185 1048.035 5440.465 1186.22 ;
      RECT 5439.625 1048.035 5439.905 1185.98 ;
      RECT 5426.185 1048.035 5426.465 1191.78 ;
      RECT 5425.625 1048.035 5425.905 1191.54 ;
      RECT 5425.065 1048.035 5425.345 1191.3 ;
      RECT 5424.505 1048.035 5424.785 1191.06 ;
      RECT 5423.945 1048.035 5424.225 1190.82 ;
      RECT 5423.385 1048.035 5423.665 1190.58 ;
      RECT 5422.825 1048.035 5423.105 1190.34 ;
      RECT 5422.265 1048.035 5422.545 1190.1 ;
      RECT 5421.705 1046.935 5421.985 1189.86 ;
      RECT 5421.145 1048.035 5421.425 1189.62 ;
      RECT 5420.585 1046.935 5420.865 1189.3 ;
      RECT 5420.025 1048.035 5420.305 1189.14 ;
      RECT 5419.465 1046.935 5419.745 1188.9 ;
      RECT 5418.905 1048.035 5419.185 1188.66 ;
      RECT 5418.345 1048.035 5418.625 1188.42 ;
      RECT 5417.785 1048.035 5418.065 1188.18 ;
      RECT 5417.225 1048.035 5417.505 1187.94 ;
      RECT 5416.665 1048.035 5416.945 1187.7 ;
      RECT 5416.105 1048.035 5416.385 1187.46 ;
      RECT 5415.545 1048.035 5415.825 1187.22 ;
      RECT 5414.985 1048.035 5415.265 1186.98 ;
      RECT 5414.425 1046.935 5414.705 1186.74 ;
      RECT 5413.865 1048.035 5414.145 1186.5 ;
      RECT 5413.305 1046.935 5413.585 1186.26 ;
      RECT 5374.105 1048.035 5374.385 1191.87 ;
      RECT 5373.545 1048.035 5373.825 1192.11 ;
      RECT 5372.985 1048.035 5373.265 1192.35 ;
      RECT 5372.425 1048.035 5372.705 1192.59 ;
      RECT 5371.865 1048.035 5372.145 1192.83 ;
      RECT 5371.305 1048.035 5371.585 1193.07 ;
      RECT 5370.745 1048.035 5371.025 1193.31 ;
      RECT 5370.185 1048.035 5370.465 1193.55 ;
      RECT 5369.625 1048.035 5369.905 1193.79 ;
      RECT 5369.065 1048.035 5369.345 1194.03 ;
      RECT 5368.505 1048.035 5368.785 1194.27 ;
      RECT 5367.945 1048.035 5368.225 1194.51 ;
      RECT 5367.385 1048.035 5367.665 1194.75 ;
      RECT 5366.825 1048.035 5367.105 1194.75 ;
      RECT 5366.265 1046.935 5366.545 1194.51 ;
      RECT 5365.705 1048.035 5365.985 1194.27 ;
      RECT 5365.145 1046.935 5365.425 1194.03 ;
      RECT 5364.585 1048.035 5364.865 1193.79 ;
      RECT 5364.025 1048.035 5364.305 1193.55 ;
      RECT 5363.465 1048.035 5363.745 1193.31 ;
      RECT 5362.905 1046.935 5363.185 1193.045 ;
      RECT 5362.345 1048.035 5362.625 1192.805 ;
      RECT 5361.785 1046.935 5362.065 1192.565 ;
      RECT 5361.225 1048.035 5361.505 1192.325 ;
      RECT 5352.265 1046.935 5352.545 1186.16 ;
      RECT 5351.705 1048.035 5351.985 1186.4 ;
      RECT 5351.145 1048.035 5351.425 1186.64 ;
      RECT 5350.585 1048.035 5350.865 1186.64 ;
      RECT 5350.025 1048.035 5350.305 1186.4 ;
      RECT 5349.465 1048.035 5349.745 1186.16 ;
      RECT 5348.905 1048.035 5349.185 1185.92 ;
      RECT 5348.345 1048.035 5348.625 1185.68 ;
      RECT 5347.785 1048.035 5348.065 1185.44 ;
      RECT 5347.225 1048.035 5347.505 1185.2 ;
      RECT 5346.665 1048.035 5346.945 1184.96 ;
      RECT 5346.105 1048.035 5346.385 1184.72 ;
      RECT 5345.545 1048.035 5345.825 1184.48 ;
      RECT 5344.985 1046.935 5345.265 1184.24 ;
      RECT 5342.465 1048.035 5342.745 1185.96 ;
      RECT 5341.905 1046.935 5342.185 1185.72 ;
      RECT 5341.345 1048.035 5341.625 1185.48 ;
      RECT 5340.785 1046.935 5341.065 1185.24 ;
      RECT 5340.225 1048.035 5340.505 1185 ;
      RECT 5339.665 1048.035 5339.945 1184.76 ;
      RECT 5339.105 1048.035 5339.385 1184.52 ;
      RECT 5313.065 1048.035 5313.345 1187.305 ;
      RECT 5312.505 1048.035 5312.785 1187.545 ;
      RECT 5311.945 1048.035 5312.225 1187.785 ;
      RECT 5311.385 1048.035 5311.665 1188.025 ;
      RECT 5310.825 1048.035 5311.105 1188.265 ;
      RECT 5310.265 1046.935 5310.545 1188.505 ;
      RECT 5309.705 1048.035 5309.985 1188.745 ;
      RECT 5309.145 1046.935 5309.425 1188.985 ;
      RECT 5308.585 1048.035 5308.865 1189.225 ;
      RECT 5308.025 1048.035 5308.305 1189.465 ;
      RECT 5307.465 1048.035 5307.745 1189.705 ;
      RECT 5306.905 1048.035 5307.185 1189.945 ;
      RECT 5306.345 1048.035 5306.625 1190.185 ;
      RECT 5305.785 1048.035 5306.065 1190.425 ;
      RECT 5305.225 1048.035 5305.505 1190.665 ;
      RECT 5304.665 1048.035 5304.945 1190.665 ;
      RECT 5304.105 1048.035 5304.385 1190.425 ;
      RECT 5303.545 1048.035 5303.825 1190.185 ;
      RECT 5302.985 1048.035 5303.265 1189.945 ;
      RECT 5302.425 1048.035 5302.705 1189.7 ;
      RECT 5301.865 1048.035 5302.145 1189.46 ;
      RECT 5301.305 1048.035 5301.585 1189.22 ;
      RECT 5300.745 1046.935 5301.025 1188.98 ;
      RECT 5300.185 1048.035 5300.465 1188.74 ;
      RECT 5286.745 1046.935 5287.025 1186.22 ;
      RECT 5286.185 1048.035 5286.465 1185.98 ;
      RECT 5285.625 1048.035 5285.905 1185.74 ;
      RECT 5285.065 1048.035 5285.345 1185.5 ;
      RECT 5284.505 1046.935 5284.785 1185.26 ;
      RECT 5283.945 1048.035 5284.225 1185.02 ;
      RECT 5283.385 1046.935 5283.665 1184.78 ;
      RECT 5282.825 1048.035 5283.105 1184.54 ;
      RECT 5282.265 1046.935 5282.545 1184.3 ;
      RECT 5281.705 1048.035 5281.985 1184.06 ;
      RECT 5281.145 1048.035 5281.425 1183.82 ;
      RECT 5280.585 1048.035 5280.865 1183.58 ;
      RECT 5280.025 1048.035 5280.305 1183.34 ;
      RECT 5279.465 1048.035 5279.745 1183.1 ;
      RECT 5278.905 1048.035 5279.185 1182.86 ;
      RECT 5278.345 1048.035 5278.625 1182.62 ;
      RECT 5277.785 1048.035 5278.065 1182.38 ;
      RECT 5277.225 1048.035 5277.505 1182.14 ;
      RECT 5276.665 1048.035 5276.945 1181.9 ;
      RECT 5276.105 1048.035 5276.385 1181.66 ;
      RECT 5275.545 1048.035 5275.825 1181.42 ;
      RECT 5274.985 1046.935 5275.265 1181.18 ;
      RECT 5274.425 1048.035 5274.705 1180.94 ;
      RECT 5273.865 1046.935 5274.145 1180.7 ;
      RECT 5234.105 1048.035 5234.385 1191.17 ;
      RECT 5233.545 1046.935 5233.825 1191.41 ;
      RECT 5232.985 1048.035 5233.265 1191.65 ;
      RECT 5232.425 1048.035 5232.705 1191.89 ;
      RECT 5231.865 1048.035 5232.145 1192.13 ;
      RECT 5231.305 1048.035 5231.585 1192.37 ;
      RECT 5230.745 1048.035 5231.025 1192.61 ;
      RECT 5230.185 1048.035 5230.465 1192.855 ;
      RECT 5229.625 1048.035 5229.905 1193.095 ;
      RECT 5229.065 1048.035 5229.345 1193.335 ;
      RECT 5228.505 1046.935 5228.785 1193.575 ;
      RECT 5227.945 1048.035 5228.225 1193.815 ;
      RECT 5227.385 1046.935 5227.665 1194.055 ;
      RECT 5226.825 1048.035 5227.105 1194.295 ;
      RECT 5226.265 1048.035 5226.545 1194.535 ;
      RECT 5225.705 1048.035 5225.985 1194.775 ;
      RECT 5225.145 1048.035 5225.425 1195.015 ;
      RECT 5224.585 1048.035 5224.865 1195.255 ;
      RECT 5224.025 1048.035 5224.305 1195.495 ;
      RECT 5223.465 1048.035 5223.745 1195.735 ;
      RECT 5222.905 1048.035 5223.185 1195.975 ;
      RECT 5222.345 1048.035 5222.625 1196.215 ;
      RECT 5221.785 1048.035 5222.065 1196.455 ;
      RECT 5221.225 1048.035 5221.505 1196.695 ;
      RECT 5212.265 1048.035 5212.545 1192.28 ;
      RECT 5211.705 1048.035 5211.985 1192.04 ;
      RECT 5211.145 1048.035 5211.425 1191.8 ;
      RECT 5210.585 1046.935 5210.865 1191.56 ;
      RECT 5210.025 1048.035 5210.305 1191.32 ;
      RECT 5209.465 1046.935 5209.745 1191.08 ;
      RECT 5208.905 1048.035 5209.185 1190.84 ;
      RECT 5208.345 1048.035 5208.625 1190.6 ;
      RECT 5207.785 1048.035 5208.065 1190.36 ;
      RECT 5207.225 1046.935 5207.505 1190.12 ;
      RECT 5206.665 1048.035 5206.945 1189.88 ;
      RECT 5206.105 1046.935 5206.385 1189.64 ;
      RECT 5205.545 1048.035 5205.825 1189.4 ;
      RECT 5204.985 1046.935 5205.265 1189.16 ;
      RECT 5202.465 1048.035 5202.745 1181.56 ;
      RECT 5201.905 1048.035 5202.185 1181.32 ;
      RECT 5201.345 1048.035 5201.625 1181.08 ;
      RECT 5200.785 1048.035 5201.065 1180.84 ;
      RECT 5200.225 1048.035 5200.505 1180.6 ;
      RECT 5199.665 1048.035 5199.945 1180.36 ;
      RECT 5199.105 1048.035 5199.385 1180.12 ;
      RECT 5173.065 1048.035 5173.345 1193.995 ;
      RECT 5172.505 1048.035 5172.785 1194.235 ;
      RECT 5171.945 1048.035 5172.225 1194.475 ;
      RECT 5171.385 1048.035 5171.665 1194.715 ;
      RECT 5170.825 1048.035 5171.105 1194.955 ;
      RECT 5170.265 1046.935 5170.545 1194.955 ;
      RECT 5169.705 1048.035 5169.985 1194.715 ;
      RECT 5169.145 1046.935 5169.425 1194.47 ;
      RECT 5168.585 1048.035 5168.865 1194.23 ;
      RECT 5168.025 1046.935 5168.305 1193.99 ;
      RECT 5167.465 1048.035 5167.745 1193.75 ;
      RECT 5166.905 1048.035 5167.185 1193.51 ;
      RECT 5166.345 1048.035 5166.625 1193.27 ;
      RECT 5165.785 1048.035 5166.065 1193.03 ;
      RECT 5165.225 1048.035 5165.505 1192.79 ;
      RECT 5164.665 1048.035 5164.945 1192.55 ;
      RECT 5164.105 1048.035 5164.385 1192.31 ;
      RECT 5163.545 1048.035 5163.825 1192.07 ;
      RECT 5162.985 1046.935 5163.265 1191.83 ;
      RECT 5162.425 1048.035 5162.705 1191.59 ;
      RECT 5161.865 1046.935 5162.145 1191.35 ;
      RECT 5161.305 1048.035 5161.585 1191.11 ;
      RECT 5160.745 1048.035 5161.025 1190.87 ;
      RECT 5160.185 1048.035 5160.465 1190.63 ;
      RECT 5146.745 1048.035 5147.025 1194.03 ;
      RECT 5146.185 1048.035 5146.465 1194.27 ;
      RECT 5145.625 1048.035 5145.905 1194.515 ;
      RECT 5145.065 1048.035 5145.345 1194.755 ;
      RECT 5144.505 1048.035 5144.785 1194.995 ;
      RECT 5143.945 1048.035 5144.225 1194.995 ;
      RECT 5143.385 1048.035 5143.665 1194.755 ;
      RECT 5142.825 1048.035 5143.105 1194.515 ;
      RECT 5142.265 1048.035 5142.545 1187.5 ;
      RECT 5141.705 1048.035 5141.985 1187.26 ;
      RECT 5141.145 1048.035 5141.425 1187.02 ;
      RECT 5140.585 1046.935 5140.865 1186.78 ;
      RECT 5140.025 1048.035 5140.305 1186.54 ;
      RECT 5139.465 1046.935 5139.745 1186.3 ;
      RECT 5138.905 1048.035 5139.185 1186.06 ;
      RECT 5138.345 1048.035 5138.625 1185.82 ;
      RECT 5137.785 1048.035 5138.065 1185.58 ;
      RECT 5137.225 1046.935 5137.505 1185.34 ;
      RECT 5136.665 1048.035 5136.945 1185.1 ;
      RECT 5136.105 1046.935 5136.385 1184.86 ;
      RECT 5135.545 1048.035 5135.825 1184.62 ;
      RECT 5134.985 1046.935 5135.265 1184.38 ;
      RECT 5134.425 1048.035 5134.705 1184.14 ;
      RECT 5133.865 1048.035 5134.145 1183.9 ;
      RECT 5093.545 1048.035 5093.825 1192.795 ;
      RECT 5092.985 1048.035 5093.265 1193.035 ;
      RECT 5092.425 1048.035 5092.705 1193.28 ;
      RECT 5091.865 1048.035 5092.145 1193.52 ;
      RECT 5091.305 1048.035 5091.585 1193.76 ;
      RECT 5090.745 1048.035 5091.025 1194 ;
      RECT 5090.185 1048.035 5090.465 1194.24 ;
      RECT 5089.625 1048.035 5089.905 1194.48 ;
      RECT 5089.065 1048.035 5089.345 1194.72 ;
      RECT 5088.505 1048.035 5088.785 1194.96 ;
      RECT 5087.945 1046.935 5088.225 1195.2 ;
      RECT 5087.385 1048.035 5087.665 1195.44 ;
      RECT 5086.825 1046.935 5087.105 1195.68 ;
      RECT 5086.265 1048.035 5086.545 1195.92 ;
      RECT 5085.705 1046.935 5085.985 1196.16 ;
      RECT 5085.145 1048.035 5085.425 1196.16 ;
      RECT 5084.585 1048.035 5084.865 1195.92 ;
      RECT 5084.025 1048.035 5084.305 1195.68 ;
      RECT 5083.465 1048.035 5083.745 1195.44 ;
      RECT 5082.905 1048.035 5083.185 1195.2 ;
      RECT 5082.345 1048.035 5082.625 1194.96 ;
      RECT 5081.785 1048.035 5082.065 1194.72 ;
      RECT 5081.225 1048.035 5081.505 1194.48 ;
      RECT 5072.265 1046.935 5072.545 1194.51 ;
      RECT 5071.705 1048.035 5071.985 1194.75 ;
      RECT 5071.145 1046.935 5071.425 1194.99 ;
      RECT 5070.585 1048.035 5070.865 1195.205 ;
      RECT 5070.025 1048.035 5070.305 1194.78 ;
      RECT 5069.465 1048.035 5069.745 1194.54 ;
      RECT 5068.905 1048.035 5069.185 1194.3 ;
      RECT 5068.345 1048.035 5068.625 1194.06 ;
      RECT 5067.785 1048.035 5068.065 1193.82 ;
      RECT 5067.225 1048.035 5067.505 1193.58 ;
      RECT 5066.665 1048.035 5066.945 1193.34 ;
      RECT 5066.105 1048.035 5066.385 1193.1 ;
      RECT 5065.545 1048.035 5065.825 1192.86 ;
      RECT 5064.985 1048.035 5065.265 1192.62 ;
      RECT 5062.465 1048.035 5062.745 1191.795 ;
      RECT 5061.905 1048.035 5062.185 1191.555 ;
      RECT 5061.345 1048.035 5061.625 1191.315 ;
      RECT 5060.785 1046.935 5061.065 1191.075 ;
      RECT 5060.225 1048.035 5060.505 1190.835 ;
      RECT 5059.665 1046.935 5059.945 1190.595 ;
      RECT 5059.105 1048.035 5059.385 1190.355 ;
      RECT 5058.545 1048.035 5058.825 1190.115 ;
      RECT 5031.945 1048.035 5032.225 1201.16 ;
      RECT 5031.385 1046.935 5031.665 1201.4 ;
      RECT 5030.825 1048.035 5031.105 1201.64 ;
      RECT 5030.265 1046.935 5030.545 1201.885 ;
      RECT 5029.705 1048.035 5029.985 1202.125 ;
      RECT 5029.145 1046.935 5029.425 1202.365 ;
      RECT 5028.585 1048.035 5028.865 1202.605 ;
      RECT 5028.025 1048.035 5028.305 1202.845 ;
      RECT 5027.465 1048.035 5027.745 1188.465 ;
      RECT 5026.905 1048.035 5027.185 1188.225 ;
      RECT 5026.345 1048.035 5026.625 1187.985 ;
      RECT 5025.785 1048.035 5026.065 1187.745 ;
      RECT 5025.225 1048.035 5025.505 1187.505 ;
      RECT 5024.665 1048.035 5024.945 1187.265 ;
      RECT 5024.105 1048.035 5024.385 1187.025 ;
      RECT 5023.545 1048.035 5023.825 1186.785 ;
      RECT 5022.985 1048.035 5023.265 1186.545 ;
      RECT 5022.425 1048.035 5022.705 1186.305 ;
      RECT 5021.865 1046.935 5022.145 1186.065 ;
      RECT 5021.305 1048.035 5021.585 1185.825 ;
      RECT 5020.745 1046.935 5021.025 1185.585 ;
      RECT 5020.185 1048.035 5020.465 1185.345 ;
      RECT 5006.185 1046.935 5006.465 1191.465 ;
      RECT 5005.625 1048.035 5005.905 1191.225 ;
      RECT 5005.065 1048.035 5005.345 1190.985 ;
      RECT 5004.505 1048.035 5004.785 1190.745 ;
      RECT 5003.945 1048.035 5004.225 1190.505 ;
      RECT 5003.385 1048.035 5003.665 1190.265 ;
      RECT 5002.825 1048.035 5003.105 1190.025 ;
      RECT 5002.265 1048.035 5002.545 1189.785 ;
      RECT 5001.705 1048.035 5001.985 1189.545 ;
      RECT 5001.145 1046.935 5001.425 1189.305 ;
      RECT 5000.585 1048.035 5000.865 1189.065 ;
      RECT 5000.025 1046.935 5000.305 1188.825 ;
      RECT 4999.465 1048.035 4999.745 1188.585 ;
      RECT 4998.905 1048.035 4999.185 1188.345 ;
      RECT 4998.345 1048.035 4998.625 1188.105 ;
      RECT 4997.785 1048.035 4998.065 1187.865 ;
      RECT 4997.225 1048.035 4997.505 1187.625 ;
      RECT 4996.665 1048.035 4996.945 1187.385 ;
      RECT 4996.105 1048.035 4996.385 1187.145 ;
      RECT 4995.545 1048.035 4995.825 1186.905 ;
      RECT 4994.985 1048.035 4995.265 1186.665 ;
      RECT 4994.425 1048.035 4994.705 1186.425 ;
      RECT 4993.865 1048.035 4994.145 1186.185 ;
      RECT 4954.665 1048.035 4954.945 1193.09 ;
      RECT 4954.105 1048.035 4954.385 1193.33 ;
      RECT 4953.545 1048.035 4953.825 1193.57 ;
      RECT 4952.985 1046.935 4953.265 1193.81 ;
      RECT 4952.425 1048.035 4952.705 1194.05 ;
      RECT 4951.865 1046.935 4952.145 1194.29 ;
      RECT 4951.305 1048.035 4951.585 1194.53 ;
      RECT 4950.745 1048.035 4951.025 1194.77 ;
      RECT 4950.185 1048.035 4950.465 1195.01 ;
      RECT 4949.625 1046.935 4949.905 1195.25 ;
      RECT 4949.065 1048.035 4949.345 1195.49 ;
      RECT 4948.505 1046.935 4948.785 1195.73 ;
      RECT 4947.945 1048.035 4948.225 1195.97 ;
      RECT 4947.385 1046.935 4947.665 1196.21 ;
      RECT 4946.825 1048.035 4947.105 1196.45 ;
      RECT 4946.265 1048.035 4946.545 1196.69 ;
      RECT 4945.705 1048.035 4945.985 1196.69 ;
      RECT 4945.145 1048.035 4945.425 1196.45 ;
      RECT 4944.585 1048.035 4944.865 1196.21 ;
      RECT 4944.025 1048.035 4944.305 1195.97 ;
      RECT 4943.465 1048.035 4943.745 1195.73 ;
      RECT 4942.905 1048.035 4943.185 1195.49 ;
      RECT 4942.345 1048.035 4942.625 1195.25 ;
      RECT 4941.785 1048.035 4942.065 1195.01 ;
      RECT 4941.225 1048.035 4941.505 1194.77 ;
      RECT 4932.265 1048.035 4932.545 1194.285 ;
      RECT 4931.705 1046.935 4931.985 1194.045 ;
      RECT 4931.145 1048.035 4931.425 1193.805 ;
      RECT 4930.585 1046.935 4930.865 1193.565 ;
      RECT 4930.025 1048.035 4930.305 1193.325 ;
      RECT 4929.465 1046.935 4929.745 1193.085 ;
      RECT 4928.905 1048.035 4929.185 1192.845 ;
      RECT 4928.345 1048.035 4928.625 1192.605 ;
      RECT 4927.785 1048.035 4928.065 1192.365 ;
      RECT 4927.225 1048.035 4927.505 1192.125 ;
      RECT 4926.665 1048.035 4926.945 1191.885 ;
      RECT 4926.105 1048.035 4926.385 1191.645 ;
      RECT 4925.545 1048.035 4925.825 1191.405 ;
      RECT 4924.985 1048.035 4925.265 1191.165 ;
      RECT 4922.465 1046.935 4922.745 1192.885 ;
      RECT 4921.905 1048.035 4922.185 1192.645 ;
      RECT 4921.345 1046.935 4921.625 1192.405 ;
      RECT 4920.785 1048.035 4921.065 1192.165 ;
      RECT 4920.225 1048.035 4920.505 1191.925 ;
      RECT 4919.665 1048.035 4919.945 1191.685 ;
      RECT 4919.105 1048.035 4919.385 1191.445 ;
      RECT 4918.545 1048.035 4918.825 1191.205 ;
      RECT 4892.505 1048.035 4892.785 1188.855 ;
      RECT 4891.945 1048.035 4892.225 1189.095 ;
      RECT 4891.385 1048.035 4891.665 1189.335 ;
      RECT 4890.825 1048.035 4891.105 1189.58 ;
      RECT 4890.265 1048.035 4890.545 1189.82 ;
      RECT 4889.705 1048.035 4889.985 1190.06 ;
      RECT 4889.145 1048.035 4889.425 1190.06 ;
      RECT 4888.585 1048.035 4888.865 1189.82 ;
      RECT 4888.025 1048.035 4888.305 1189.58 ;
      RECT 4887.465 1046.935 4887.745 1189.34 ;
      RECT 4886.905 1048.035 4887.185 1189.1 ;
      RECT 4886.345 1046.935 4886.625 1188.86 ;
      RECT 4885.785 1048.035 4886.065 1188.62 ;
      RECT 4885.225 1048.035 4885.505 1188.38 ;
      RECT 4884.665 1048.035 4884.945 1188.14 ;
      RECT 4884.105 1046.935 4884.385 1187.9 ;
      RECT 4883.545 1048.035 4883.825 1187.66 ;
      RECT 4882.985 1046.935 4883.265 1187.42 ;
      RECT 4882.425 1048.035 4882.705 1187.18 ;
      RECT 4881.865 1046.935 4882.145 1186.94 ;
      RECT 4881.305 1048.035 4881.585 1186.7 ;
      RECT 4880.745 1048.035 4881.025 1186.46 ;
      RECT 4880.185 1048.035 4880.465 1186.22 ;
      RECT 4879.625 1048.035 4879.905 1185.98 ;
      RECT 4866.185 1048.035 4866.465 1191.78 ;
      RECT 4865.625 1048.035 4865.905 1191.54 ;
      RECT 4865.065 1048.035 4865.345 1191.3 ;
      RECT 4864.505 1048.035 4864.785 1191.06 ;
      RECT 4863.945 1048.035 4864.225 1190.82 ;
      RECT 4863.385 1048.035 4863.665 1190.58 ;
      RECT 4862.825 1048.035 4863.105 1190.34 ;
      RECT 4862.265 1048.035 4862.545 1190.1 ;
      RECT 4861.705 1046.935 4861.985 1189.86 ;
      RECT 4861.145 1048.035 4861.425 1189.62 ;
      RECT 4860.585 1046.935 4860.865 1189.3 ;
      RECT 4860.025 1048.035 4860.305 1189.14 ;
      RECT 4859.465 1046.935 4859.745 1188.9 ;
      RECT 4858.905 1048.035 4859.185 1188.66 ;
      RECT 4858.345 1048.035 4858.625 1188.42 ;
      RECT 4857.785 1048.035 4858.065 1188.18 ;
      RECT 4857.225 1048.035 4857.505 1187.94 ;
      RECT 4856.665 1048.035 4856.945 1187.7 ;
      RECT 4856.105 1048.035 4856.385 1187.46 ;
      RECT 4855.545 1048.035 4855.825 1187.22 ;
      RECT 4854.985 1048.035 4855.265 1186.98 ;
      RECT 4854.425 1046.935 4854.705 1186.74 ;
      RECT 4853.865 1048.035 4854.145 1186.5 ;
      RECT 4853.305 1046.935 4853.585 1186.26 ;
      RECT 4814.105 1048.035 4814.385 1191.87 ;
      RECT 4813.545 1048.035 4813.825 1192.11 ;
      RECT 4812.985 1048.035 4813.265 1192.35 ;
      RECT 4812.425 1048.035 4812.705 1192.59 ;
      RECT 4811.865 1048.035 4812.145 1192.83 ;
      RECT 4811.305 1048.035 4811.585 1193.07 ;
      RECT 4810.745 1048.035 4811.025 1193.31 ;
      RECT 4810.185 1048.035 4810.465 1193.55 ;
      RECT 4809.625 1048.035 4809.905 1193.79 ;
      RECT 4809.065 1048.035 4809.345 1194.03 ;
      RECT 4808.505 1048.035 4808.785 1194.27 ;
      RECT 4807.945 1048.035 4808.225 1194.51 ;
      RECT 4807.385 1048.035 4807.665 1194.75 ;
      RECT 4806.825 1048.035 4807.105 1194.75 ;
      RECT 4806.265 1046.935 4806.545 1194.51 ;
      RECT 4805.705 1048.035 4805.985 1194.27 ;
      RECT 4805.145 1046.935 4805.425 1194.03 ;
      RECT 4804.585 1048.035 4804.865 1193.79 ;
      RECT 4804.025 1048.035 4804.305 1193.55 ;
      RECT 4803.465 1048.035 4803.745 1193.31 ;
      RECT 4802.905 1046.935 4803.185 1193.045 ;
      RECT 4802.345 1048.035 4802.625 1192.805 ;
      RECT 4801.785 1046.935 4802.065 1192.565 ;
      RECT 4801.225 1048.035 4801.505 1192.325 ;
      RECT 4792.265 1046.935 4792.545 1186.16 ;
      RECT 4791.705 1048.035 4791.985 1186.4 ;
      RECT 4791.145 1048.035 4791.425 1186.64 ;
      RECT 4790.585 1048.035 4790.865 1186.64 ;
      RECT 4790.025 1048.035 4790.305 1186.4 ;
      RECT 4789.465 1048.035 4789.745 1186.16 ;
      RECT 4788.905 1048.035 4789.185 1185.92 ;
      RECT 4788.345 1048.035 4788.625 1185.68 ;
      RECT 4787.785 1048.035 4788.065 1185.44 ;
      RECT 4787.225 1048.035 4787.505 1185.2 ;
      RECT 4786.665 1048.035 4786.945 1184.96 ;
      RECT 4786.105 1048.035 4786.385 1184.72 ;
      RECT 4785.545 1048.035 4785.825 1184.48 ;
      RECT 4784.985 1046.935 4785.265 1184.24 ;
      RECT 4782.465 1048.035 4782.745 1185.96 ;
      RECT 4781.905 1046.935 4782.185 1185.72 ;
      RECT 4781.345 1048.035 4781.625 1185.48 ;
      RECT 4780.785 1046.935 4781.065 1185.24 ;
      RECT 4780.225 1048.035 4780.505 1185 ;
      RECT 4779.665 1048.035 4779.945 1184.76 ;
      RECT 4779.105 1048.035 4779.385 1184.52 ;
      RECT 4753.065 1048.035 4753.345 1187.305 ;
      RECT 4752.505 1048.035 4752.785 1187.545 ;
      RECT 4751.945 1048.035 4752.225 1187.785 ;
      RECT 4751.385 1048.035 4751.665 1188.025 ;
      RECT 4750.825 1048.035 4751.105 1188.265 ;
      RECT 4750.265 1046.935 4750.545 1188.505 ;
      RECT 4749.705 1048.035 4749.985 1188.745 ;
      RECT 4749.145 1046.935 4749.425 1188.985 ;
      RECT 4748.585 1048.035 4748.865 1189.225 ;
      RECT 4748.025 1048.035 4748.305 1189.465 ;
      RECT 4747.465 1048.035 4747.745 1189.705 ;
      RECT 4746.905 1048.035 4747.185 1189.945 ;
      RECT 4746.345 1048.035 4746.625 1190.185 ;
      RECT 4745.785 1048.035 4746.065 1190.425 ;
      RECT 4745.225 1048.035 4745.505 1190.665 ;
      RECT 4744.665 1048.035 4744.945 1190.665 ;
      RECT 4744.105 1048.035 4744.385 1190.425 ;
      RECT 4743.545 1048.035 4743.825 1190.185 ;
      RECT 4742.985 1048.035 4743.265 1189.945 ;
      RECT 4742.425 1048.035 4742.705 1189.7 ;
      RECT 4741.865 1048.035 4742.145 1189.46 ;
      RECT 4741.305 1048.035 4741.585 1189.22 ;
      RECT 4740.745 1046.935 4741.025 1188.98 ;
      RECT 4740.185 1048.035 4740.465 1188.74 ;
      RECT 4726.745 1046.935 4727.025 1186.22 ;
      RECT 4726.185 1048.035 4726.465 1185.98 ;
      RECT 4725.625 1048.035 4725.905 1185.74 ;
      RECT 4725.065 1048.035 4725.345 1185.5 ;
      RECT 4724.505 1046.935 4724.785 1185.26 ;
      RECT 4723.945 1048.035 4724.225 1185.02 ;
      RECT 4723.385 1046.935 4723.665 1184.78 ;
      RECT 4722.825 1048.035 4723.105 1184.54 ;
      RECT 4722.265 1046.935 4722.545 1184.3 ;
      RECT 4721.705 1048.035 4721.985 1184.06 ;
      RECT 4721.145 1048.035 4721.425 1183.82 ;
      RECT 4720.585 1048.035 4720.865 1183.58 ;
      RECT 4720.025 1048.035 4720.305 1183.34 ;
      RECT 4719.465 1048.035 4719.745 1183.1 ;
      RECT 4718.905 1048.035 4719.185 1182.86 ;
      RECT 4718.345 1048.035 4718.625 1182.62 ;
      RECT 4717.785 1048.035 4718.065 1182.38 ;
      RECT 4717.225 1048.035 4717.505 1182.14 ;
      RECT 4716.665 1048.035 4716.945 1181.9 ;
      RECT 4716.105 1048.035 4716.385 1181.66 ;
      RECT 4715.545 1048.035 4715.825 1181.42 ;
      RECT 4714.985 1046.935 4715.265 1181.18 ;
      RECT 4714.425 1048.035 4714.705 1180.94 ;
      RECT 4713.865 1046.935 4714.145 1180.7 ;
      RECT 4674.105 1048.035 4674.385 1191.17 ;
      RECT 4673.545 1046.935 4673.825 1191.41 ;
      RECT 4672.985 1048.035 4673.265 1191.65 ;
      RECT 4672.425 1048.035 4672.705 1191.89 ;
      RECT 4671.865 1048.035 4672.145 1192.13 ;
      RECT 4671.305 1048.035 4671.585 1192.37 ;
      RECT 4670.745 1048.035 4671.025 1192.61 ;
      RECT 4670.185 1048.035 4670.465 1192.855 ;
      RECT 4669.625 1048.035 4669.905 1193.095 ;
      RECT 4669.065 1048.035 4669.345 1193.335 ;
      RECT 4668.505 1046.935 4668.785 1193.575 ;
      RECT 4667.945 1048.035 4668.225 1193.815 ;
      RECT 4667.385 1046.935 4667.665 1194.055 ;
      RECT 4666.825 1048.035 4667.105 1194.295 ;
      RECT 4666.265 1048.035 4666.545 1194.535 ;
      RECT 4665.705 1048.035 4665.985 1194.775 ;
      RECT 4665.145 1048.035 4665.425 1195.015 ;
      RECT 4664.585 1048.035 4664.865 1195.255 ;
      RECT 4664.025 1048.035 4664.305 1195.495 ;
      RECT 4663.465 1048.035 4663.745 1195.735 ;
      RECT 4662.905 1048.035 4663.185 1195.975 ;
      RECT 4662.345 1048.035 4662.625 1196.215 ;
      RECT 4661.785 1048.035 4662.065 1196.455 ;
      RECT 4661.225 1048.035 4661.505 1196.695 ;
      RECT 4652.265 1048.035 4652.545 1192.28 ;
      RECT 4651.705 1048.035 4651.985 1192.04 ;
      RECT 4651.145 1048.035 4651.425 1191.8 ;
      RECT 4650.585 1046.935 4650.865 1191.56 ;
      RECT 4650.025 1048.035 4650.305 1191.32 ;
      RECT 4649.465 1046.935 4649.745 1191.08 ;
      RECT 4648.905 1048.035 4649.185 1190.84 ;
      RECT 4648.345 1048.035 4648.625 1190.6 ;
      RECT 4647.785 1048.035 4648.065 1190.36 ;
      RECT 4647.225 1046.935 4647.505 1190.12 ;
      RECT 4646.665 1048.035 4646.945 1189.88 ;
      RECT 4646.105 1046.935 4646.385 1189.64 ;
      RECT 4645.545 1048.035 4645.825 1189.4 ;
      RECT 4644.985 1046.935 4645.265 1189.16 ;
      RECT 4642.465 1048.035 4642.745 1181.56 ;
      RECT 4641.905 1048.035 4642.185 1181.32 ;
      RECT 4641.345 1048.035 4641.625 1181.08 ;
      RECT 4640.785 1048.035 4641.065 1180.84 ;
      RECT 4640.225 1048.035 4640.505 1180.6 ;
      RECT 4639.665 1048.035 4639.945 1180.36 ;
      RECT 4639.105 1048.035 4639.385 1180.12 ;
      RECT 4613.065 1048.035 4613.345 1193.995 ;
      RECT 4612.505 1048.035 4612.785 1194.235 ;
      RECT 4611.945 1048.035 4612.225 1194.475 ;
      RECT 4611.385 1048.035 4611.665 1194.715 ;
      RECT 4610.825 1048.035 4611.105 1194.955 ;
      RECT 4610.265 1046.935 4610.545 1194.955 ;
      RECT 4609.705 1048.035 4609.985 1194.715 ;
      RECT 4609.145 1046.935 4609.425 1194.47 ;
      RECT 4608.585 1048.035 4608.865 1194.23 ;
      RECT 4608.025 1046.935 4608.305 1193.99 ;
      RECT 4607.465 1048.035 4607.745 1193.75 ;
      RECT 4606.905 1048.035 4607.185 1193.51 ;
      RECT 4606.345 1048.035 4606.625 1193.27 ;
      RECT 4605.785 1048.035 4606.065 1193.03 ;
      RECT 4605.225 1048.035 4605.505 1192.79 ;
      RECT 4604.665 1048.035 4604.945 1192.55 ;
      RECT 4604.105 1048.035 4604.385 1192.31 ;
      RECT 4603.545 1048.035 4603.825 1192.07 ;
      RECT 4602.985 1046.935 4603.265 1191.83 ;
      RECT 4602.425 1048.035 4602.705 1191.59 ;
      RECT 4601.865 1046.935 4602.145 1191.35 ;
      RECT 4601.305 1048.035 4601.585 1191.11 ;
      RECT 4600.745 1048.035 4601.025 1190.87 ;
      RECT 4600.185 1048.035 4600.465 1190.63 ;
      RECT 4586.745 1048.035 4587.025 1194.03 ;
      RECT 4586.185 1048.035 4586.465 1194.27 ;
      RECT 4585.625 1048.035 4585.905 1194.515 ;
      RECT 4585.065 1048.035 4585.345 1194.755 ;
      RECT 4584.505 1048.035 4584.785 1194.995 ;
      RECT 4583.945 1048.035 4584.225 1194.995 ;
      RECT 4583.385 1048.035 4583.665 1194.755 ;
      RECT 4582.825 1048.035 4583.105 1194.515 ;
      RECT 4582.265 1048.035 4582.545 1187.5 ;
      RECT 4581.705 1048.035 4581.985 1187.26 ;
      RECT 4581.145 1048.035 4581.425 1187.02 ;
      RECT 4580.585 1046.935 4580.865 1186.78 ;
      RECT 4580.025 1048.035 4580.305 1186.54 ;
      RECT 4579.465 1046.935 4579.745 1186.3 ;
      RECT 4578.905 1048.035 4579.185 1186.06 ;
      RECT 4578.345 1048.035 4578.625 1185.82 ;
      RECT 4577.785 1048.035 4578.065 1185.58 ;
      RECT 4577.225 1046.935 4577.505 1185.34 ;
      RECT 4576.665 1048.035 4576.945 1185.1 ;
      RECT 4576.105 1046.935 4576.385 1184.86 ;
      RECT 4575.545 1048.035 4575.825 1184.62 ;
      RECT 4574.985 1046.935 4575.265 1184.38 ;
      RECT 4574.425 1048.035 4574.705 1184.14 ;
      RECT 4573.865 1048.035 4574.145 1183.9 ;
      RECT 4533.545 1048.035 4533.825 1192.795 ;
      RECT 4532.985 1048.035 4533.265 1193.035 ;
      RECT 4532.425 1048.035 4532.705 1193.28 ;
      RECT 4531.865 1048.035 4532.145 1193.52 ;
      RECT 4531.305 1048.035 4531.585 1193.76 ;
      RECT 4530.745 1048.035 4531.025 1194 ;
      RECT 4530.185 1048.035 4530.465 1194.24 ;
      RECT 4529.625 1048.035 4529.905 1194.48 ;
      RECT 4529.065 1048.035 4529.345 1194.72 ;
      RECT 4528.505 1048.035 4528.785 1194.96 ;
      RECT 4527.945 1046.935 4528.225 1195.2 ;
      RECT 4527.385 1048.035 4527.665 1195.44 ;
      RECT 4526.825 1046.935 4527.105 1195.68 ;
      RECT 4526.265 1048.035 4526.545 1195.92 ;
      RECT 4525.705 1046.935 4525.985 1196.16 ;
      RECT 4525.145 1048.035 4525.425 1196.16 ;
      RECT 4524.585 1048.035 4524.865 1195.92 ;
      RECT 4524.025 1048.035 4524.305 1195.68 ;
      RECT 4523.465 1048.035 4523.745 1195.44 ;
      RECT 4522.905 1048.035 4523.185 1195.2 ;
      RECT 4522.345 1048.035 4522.625 1194.96 ;
      RECT 4521.785 1048.035 4522.065 1194.72 ;
      RECT 4521.225 1048.035 4521.505 1194.48 ;
      RECT 4512.265 1046.935 4512.545 1194.51 ;
      RECT 4511.705 1048.035 4511.985 1194.75 ;
      RECT 4511.145 1046.935 4511.425 1194.99 ;
      RECT 4510.585 1048.035 4510.865 1195.205 ;
      RECT 4510.025 1048.035 4510.305 1194.78 ;
      RECT 4509.465 1048.035 4509.745 1194.54 ;
      RECT 4508.905 1048.035 4509.185 1194.3 ;
      RECT 4508.345 1048.035 4508.625 1194.06 ;
      RECT 4507.785 1048.035 4508.065 1193.82 ;
      RECT 4507.225 1048.035 4507.505 1193.58 ;
      RECT 4506.665 1048.035 4506.945 1193.34 ;
      RECT 4506.105 1048.035 4506.385 1193.1 ;
      RECT 4505.545 1048.035 4505.825 1192.86 ;
      RECT 4504.985 1048.035 4505.265 1192.62 ;
      RECT 4502.465 1048.035 4502.745 1191.795 ;
      RECT 4501.905 1048.035 4502.185 1191.555 ;
      RECT 4501.345 1048.035 4501.625 1191.315 ;
      RECT 4500.785 1046.935 4501.065 1191.075 ;
      RECT 4500.225 1048.035 4500.505 1190.835 ;
      RECT 4499.665 1046.935 4499.945 1190.595 ;
      RECT 4499.105 1048.035 4499.385 1190.355 ;
      RECT 4498.545 1048.035 4498.825 1190.115 ;
      RECT 4471.945 1048.035 4472.225 1201.16 ;
      RECT 4471.385 1046.935 4471.665 1201.4 ;
      RECT 4470.825 1048.035 4471.105 1201.64 ;
      RECT 4470.265 1046.935 4470.545 1201.885 ;
      RECT 4469.705 1048.035 4469.985 1202.125 ;
      RECT 4469.145 1046.935 4469.425 1202.365 ;
      RECT 4468.585 1048.035 4468.865 1202.605 ;
      RECT 4468.025 1048.035 4468.305 1202.845 ;
      RECT 4467.465 1048.035 4467.745 1188.465 ;
      RECT 4466.905 1048.035 4467.185 1188.225 ;
      RECT 4466.345 1048.035 4466.625 1187.985 ;
      RECT 4465.785 1048.035 4466.065 1187.745 ;
      RECT 4465.225 1048.035 4465.505 1187.505 ;
      RECT 4464.665 1048.035 4464.945 1187.265 ;
      RECT 4464.105 1048.035 4464.385 1187.025 ;
      RECT 4463.545 1048.035 4463.825 1186.785 ;
      RECT 4462.985 1048.035 4463.265 1186.545 ;
      RECT 4462.425 1048.035 4462.705 1186.305 ;
      RECT 4461.865 1046.935 4462.145 1186.065 ;
      RECT 4461.305 1048.035 4461.585 1185.825 ;
      RECT 4460.745 1046.935 4461.025 1185.585 ;
      RECT 4460.185 1048.035 4460.465 1185.345 ;
      RECT 4446.185 1046.935 4446.465 1191.465 ;
      RECT 4445.625 1048.035 4445.905 1191.225 ;
      RECT 4445.065 1048.035 4445.345 1190.985 ;
      RECT 4444.505 1048.035 4444.785 1190.745 ;
      RECT 4443.945 1048.035 4444.225 1190.505 ;
      RECT 4443.385 1048.035 4443.665 1190.265 ;
      RECT 4442.825 1048.035 4443.105 1190.025 ;
      RECT 4442.265 1048.035 4442.545 1189.785 ;
      RECT 4441.705 1048.035 4441.985 1189.545 ;
      RECT 4441.145 1046.935 4441.425 1189.305 ;
      RECT 4440.585 1048.035 4440.865 1189.065 ;
      RECT 4440.025 1046.935 4440.305 1188.825 ;
      RECT 4439.465 1048.035 4439.745 1188.585 ;
      RECT 4438.905 1048.035 4439.185 1188.345 ;
      RECT 4438.345 1048.035 4438.625 1188.105 ;
      RECT 4437.785 1048.035 4438.065 1187.865 ;
      RECT 4437.225 1048.035 4437.505 1187.625 ;
      RECT 4436.665 1048.035 4436.945 1187.385 ;
      RECT 4436.105 1048.035 4436.385 1187.145 ;
      RECT 4435.545 1048.035 4435.825 1186.905 ;
      RECT 4434.985 1048.035 4435.265 1186.665 ;
      RECT 4434.425 1048.035 4434.705 1186.425 ;
      RECT 4433.865 1048.035 4434.145 1186.185 ;
      RECT 4394.665 1048.035 4394.945 1193.09 ;
      RECT 4394.105 1048.035 4394.385 1193.33 ;
      RECT 4393.545 1048.035 4393.825 1193.57 ;
      RECT 4392.985 1046.935 4393.265 1193.81 ;
      RECT 4392.425 1048.035 4392.705 1194.05 ;
      RECT 4391.865 1046.935 4392.145 1194.29 ;
      RECT 4391.305 1048.035 4391.585 1194.53 ;
      RECT 4390.745 1048.035 4391.025 1194.77 ;
      RECT 4390.185 1048.035 4390.465 1195.01 ;
      RECT 4389.625 1046.935 4389.905 1195.25 ;
      RECT 4389.065 1048.035 4389.345 1195.49 ;
      RECT 4388.505 1046.935 4388.785 1195.73 ;
      RECT 4387.945 1048.035 4388.225 1195.97 ;
      RECT 4387.385 1046.935 4387.665 1196.21 ;
      RECT 4386.825 1048.035 4387.105 1196.45 ;
      RECT 4386.265 1048.035 4386.545 1196.69 ;
      RECT 4385.705 1048.035 4385.985 1196.69 ;
      RECT 4385.145 1048.035 4385.425 1196.45 ;
      RECT 4384.585 1048.035 4384.865 1196.21 ;
      RECT 4384.025 1048.035 4384.305 1195.97 ;
      RECT 4383.465 1048.035 4383.745 1195.73 ;
      RECT 4382.905 1048.035 4383.185 1195.49 ;
      RECT 4382.345 1048.035 4382.625 1195.25 ;
      RECT 4381.785 1048.035 4382.065 1195.01 ;
      RECT 4381.225 1048.035 4381.505 1194.77 ;
      RECT 4372.265 1048.035 4372.545 1194.285 ;
      RECT 4371.705 1046.935 4371.985 1194.045 ;
      RECT 4371.145 1048.035 4371.425 1193.805 ;
      RECT 4370.585 1046.935 4370.865 1193.565 ;
      RECT 4370.025 1048.035 4370.305 1193.325 ;
      RECT 4369.465 1046.935 4369.745 1193.085 ;
      RECT 4368.905 1048.035 4369.185 1192.845 ;
      RECT 4368.345 1048.035 4368.625 1192.605 ;
      RECT 4367.785 1048.035 4368.065 1192.365 ;
      RECT 4367.225 1048.035 4367.505 1192.125 ;
      RECT 4366.665 1048.035 4366.945 1191.885 ;
      RECT 4366.105 1048.035 4366.385 1191.645 ;
      RECT 4365.545 1048.035 4365.825 1191.405 ;
      RECT 4364.985 1048.035 4365.265 1191.165 ;
      RECT 4362.465 1046.935 4362.745 1192.885 ;
      RECT 4361.905 1048.035 4362.185 1192.645 ;
      RECT 4361.345 1046.935 4361.625 1192.405 ;
      RECT 4360.785 1048.035 4361.065 1192.165 ;
      RECT 4360.225 1048.035 4360.505 1191.925 ;
      RECT 4359.665 1048.035 4359.945 1191.685 ;
      RECT 4359.105 1048.035 4359.385 1191.445 ;
      RECT 4358.545 1048.035 4358.825 1191.205 ;
      RECT 4332.505 1048.035 4332.785 1188.855 ;
      RECT 4331.945 1048.035 4332.225 1189.095 ;
      RECT 4331.385 1048.035 4331.665 1189.335 ;
      RECT 4330.825 1048.035 4331.105 1189.58 ;
      RECT 4330.265 1048.035 4330.545 1189.82 ;
      RECT 4329.705 1048.035 4329.985 1190.06 ;
      RECT 4329.145 1048.035 4329.425 1190.06 ;
      RECT 4328.585 1048.035 4328.865 1189.82 ;
      RECT 4328.025 1048.035 4328.305 1189.58 ;
      RECT 4327.465 1046.935 4327.745 1189.34 ;
      RECT 4326.905 1048.035 4327.185 1189.1 ;
      RECT 4326.345 1046.935 4326.625 1188.86 ;
      RECT 4325.785 1048.035 4326.065 1188.62 ;
      RECT 4325.225 1048.035 4325.505 1188.38 ;
      RECT 4324.665 1048.035 4324.945 1188.14 ;
      RECT 4324.105 1046.935 4324.385 1187.9 ;
      RECT 4323.545 1048.035 4323.825 1187.66 ;
      RECT 4322.985 1046.935 4323.265 1187.42 ;
      RECT 4322.425 1048.035 4322.705 1187.18 ;
      RECT 4321.865 1046.935 4322.145 1186.94 ;
      RECT 4321.305 1048.035 4321.585 1186.7 ;
      RECT 4320.745 1048.035 4321.025 1186.46 ;
      RECT 4320.185 1048.035 4320.465 1186.22 ;
      RECT 4319.625 1048.035 4319.905 1185.98 ;
      RECT 4306.185 1048.035 4306.465 1191.78 ;
      RECT 4305.625 1048.035 4305.905 1191.54 ;
      RECT 4305.065 1048.035 4305.345 1191.3 ;
      RECT 4304.505 1048.035 4304.785 1191.06 ;
      RECT 4303.945 1048.035 4304.225 1190.82 ;
      RECT 4303.385 1048.035 4303.665 1190.58 ;
      RECT 4302.825 1048.035 4303.105 1190.34 ;
      RECT 4302.265 1048.035 4302.545 1190.1 ;
      RECT 4301.705 1046.935 4301.985 1189.86 ;
      RECT 4301.145 1048.035 4301.425 1189.62 ;
      RECT 4300.585 1046.935 4300.865 1189.3 ;
      RECT 4300.025 1048.035 4300.305 1189.14 ;
      RECT 4299.465 1046.935 4299.745 1188.9 ;
      RECT 4298.905 1048.035 4299.185 1188.66 ;
      RECT 4298.345 1048.035 4298.625 1188.42 ;
      RECT 4297.785 1048.035 4298.065 1188.18 ;
      RECT 4297.225 1048.035 4297.505 1187.94 ;
      RECT 4296.665 1048.035 4296.945 1187.7 ;
      RECT 4296.105 1048.035 4296.385 1187.46 ;
      RECT 4295.545 1048.035 4295.825 1187.22 ;
      RECT 4294.985 1048.035 4295.265 1186.98 ;
      RECT 4294.425 1046.935 4294.705 1186.74 ;
      RECT 4293.865 1048.035 4294.145 1186.5 ;
      RECT 4293.305 1046.935 4293.585 1186.26 ;
      RECT 4254.105 1048.035 4254.385 1191.87 ;
      RECT 4253.545 1048.035 4253.825 1192.11 ;
      RECT 4252.985 1048.035 4253.265 1192.35 ;
      RECT 4252.425 1048.035 4252.705 1192.59 ;
      RECT 4251.865 1048.035 4252.145 1192.83 ;
      RECT 4251.305 1048.035 4251.585 1193.07 ;
      RECT 4250.745 1048.035 4251.025 1193.31 ;
      RECT 4250.185 1048.035 4250.465 1193.55 ;
      RECT 4249.625 1048.035 4249.905 1193.79 ;
      RECT 4249.065 1048.035 4249.345 1194.03 ;
      RECT 4248.505 1048.035 4248.785 1194.27 ;
      RECT 4247.945 1048.035 4248.225 1194.51 ;
      RECT 4247.385 1048.035 4247.665 1194.75 ;
      RECT 4246.825 1048.035 4247.105 1194.75 ;
      RECT 4246.265 1046.935 4246.545 1194.51 ;
      RECT 4245.705 1048.035 4245.985 1194.27 ;
      RECT 4245.145 1046.935 4245.425 1194.03 ;
      RECT 4244.585 1048.035 4244.865 1193.79 ;
      RECT 4244.025 1048.035 4244.305 1193.55 ;
      RECT 4243.465 1048.035 4243.745 1193.31 ;
      RECT 4242.905 1046.935 4243.185 1193.045 ;
      RECT 4242.345 1048.035 4242.625 1192.805 ;
      RECT 4241.785 1046.935 4242.065 1192.565 ;
      RECT 4241.225 1048.035 4241.505 1192.325 ;
      RECT 4232.265 1046.935 4232.545 1186.16 ;
      RECT 4231.705 1048.035 4231.985 1186.4 ;
      RECT 4231.145 1048.035 4231.425 1186.64 ;
      RECT 4230.585 1048.035 4230.865 1186.64 ;
      RECT 4230.025 1048.035 4230.305 1186.4 ;
      RECT 4229.465 1048.035 4229.745 1186.16 ;
      RECT 4228.905 1048.035 4229.185 1185.92 ;
      RECT 4228.345 1048.035 4228.625 1185.68 ;
      RECT 4227.785 1048.035 4228.065 1185.44 ;
      RECT 4227.225 1048.035 4227.505 1185.2 ;
      RECT 4226.665 1048.035 4226.945 1184.96 ;
      RECT 4226.105 1048.035 4226.385 1184.72 ;
      RECT 4225.545 1048.035 4225.825 1184.48 ;
      RECT 4224.985 1046.935 4225.265 1184.24 ;
      RECT 4222.465 1048.035 4222.745 1185.96 ;
      RECT 4221.905 1046.935 4222.185 1185.72 ;
      RECT 4221.345 1048.035 4221.625 1185.48 ;
      RECT 4220.785 1046.935 4221.065 1185.24 ;
      RECT 4220.225 1048.035 4220.505 1185 ;
      RECT 4219.665 1048.035 4219.945 1184.76 ;
      RECT 4219.105 1048.035 4219.385 1184.52 ;
      RECT 4193.065 1048.035 4193.345 1187.305 ;
      RECT 4192.505 1048.035 4192.785 1187.545 ;
      RECT 4191.945 1048.035 4192.225 1187.785 ;
      RECT 4191.385 1048.035 4191.665 1188.025 ;
      RECT 4190.825 1048.035 4191.105 1188.265 ;
      RECT 4190.265 1046.935 4190.545 1188.505 ;
      RECT 4189.705 1048.035 4189.985 1188.745 ;
      RECT 4189.145 1046.935 4189.425 1188.985 ;
      RECT 4188.585 1048.035 4188.865 1189.225 ;
      RECT 4188.025 1048.035 4188.305 1189.465 ;
      RECT 4187.465 1048.035 4187.745 1189.705 ;
      RECT 4186.905 1048.035 4187.185 1189.945 ;
      RECT 4186.345 1048.035 4186.625 1190.185 ;
      RECT 4185.785 1048.035 4186.065 1190.425 ;
      RECT 4185.225 1048.035 4185.505 1190.665 ;
      RECT 4184.665 1048.035 4184.945 1190.665 ;
      RECT 4184.105 1048.035 4184.385 1190.425 ;
      RECT 4183.545 1048.035 4183.825 1190.185 ;
      RECT 4182.985 1048.035 4183.265 1189.945 ;
      RECT 4182.425 1048.035 4182.705 1189.7 ;
      RECT 4181.865 1048.035 4182.145 1189.46 ;
      RECT 4181.305 1048.035 4181.585 1189.22 ;
      RECT 4180.745 1046.935 4181.025 1188.98 ;
      RECT 4180.185 1048.035 4180.465 1188.74 ;
      RECT 4166.745 1046.935 4167.025 1186.22 ;
      RECT 4166.185 1048.035 4166.465 1185.98 ;
      RECT 4165.625 1048.035 4165.905 1185.74 ;
      RECT 4165.065 1048.035 4165.345 1185.5 ;
      RECT 4164.505 1046.935 4164.785 1185.26 ;
      RECT 4163.945 1048.035 4164.225 1185.02 ;
      RECT 4163.385 1046.935 4163.665 1184.78 ;
      RECT 4162.825 1048.035 4163.105 1184.54 ;
      RECT 4162.265 1046.935 4162.545 1184.3 ;
      RECT 4161.705 1048.035 4161.985 1184.06 ;
      RECT 4161.145 1048.035 4161.425 1183.82 ;
      RECT 4160.585 1048.035 4160.865 1183.58 ;
      RECT 4160.025 1048.035 4160.305 1183.34 ;
      RECT 4159.465 1048.035 4159.745 1183.1 ;
      RECT 4158.905 1048.035 4159.185 1182.86 ;
      RECT 4158.345 1048.035 4158.625 1182.62 ;
      RECT 4157.785 1048.035 4158.065 1182.38 ;
      RECT 4157.225 1048.035 4157.505 1182.14 ;
      RECT 4156.665 1048.035 4156.945 1181.9 ;
      RECT 4156.105 1048.035 4156.385 1181.66 ;
      RECT 4155.545 1048.035 4155.825 1181.42 ;
      RECT 4154.985 1046.935 4155.265 1181.18 ;
      RECT 4154.425 1048.035 4154.705 1180.94 ;
      RECT 4153.865 1046.935 4154.145 1180.7 ;
      RECT 4114.105 1048.035 4114.385 1191.17 ;
      RECT 4113.545 1046.935 4113.825 1191.41 ;
      RECT 4112.985 1048.035 4113.265 1191.65 ;
      RECT 4112.425 1048.035 4112.705 1191.89 ;
      RECT 4111.865 1048.035 4112.145 1192.13 ;
      RECT 4111.305 1048.035 4111.585 1192.37 ;
      RECT 4110.745 1048.035 4111.025 1192.61 ;
      RECT 4110.185 1048.035 4110.465 1192.855 ;
      RECT 4109.625 1048.035 4109.905 1193.095 ;
      RECT 4109.065 1048.035 4109.345 1193.335 ;
      RECT 4108.505 1046.935 4108.785 1193.575 ;
      RECT 4107.945 1048.035 4108.225 1193.815 ;
      RECT 4107.385 1046.935 4107.665 1194.055 ;
      RECT 4106.825 1048.035 4107.105 1194.295 ;
      RECT 4106.265 1048.035 4106.545 1194.535 ;
      RECT 4105.705 1048.035 4105.985 1194.775 ;
      RECT 4105.145 1048.035 4105.425 1195.015 ;
      RECT 4104.585 1048.035 4104.865 1195.255 ;
      RECT 4104.025 1048.035 4104.305 1195.495 ;
      RECT 4103.465 1048.035 4103.745 1195.735 ;
      RECT 4102.905 1048.035 4103.185 1195.975 ;
      RECT 4102.345 1048.035 4102.625 1196.215 ;
      RECT 4101.785 1048.035 4102.065 1196.455 ;
      RECT 4101.225 1048.035 4101.505 1196.695 ;
      RECT 4092.265 1048.035 4092.545 1192.28 ;
      RECT 4091.705 1048.035 4091.985 1192.04 ;
      RECT 4091.145 1048.035 4091.425 1191.8 ;
      RECT 4090.585 1046.935 4090.865 1191.56 ;
      RECT 4090.025 1048.035 4090.305 1191.32 ;
      RECT 4089.465 1046.935 4089.745 1191.08 ;
      RECT 4088.905 1048.035 4089.185 1190.84 ;
      RECT 4088.345 1048.035 4088.625 1190.6 ;
      RECT 4087.785 1048.035 4088.065 1190.36 ;
      RECT 4087.225 1046.935 4087.505 1190.12 ;
      RECT 4086.665 1048.035 4086.945 1189.88 ;
      RECT 4086.105 1046.935 4086.385 1189.64 ;
      RECT 4085.545 1048.035 4085.825 1189.4 ;
      RECT 4084.985 1046.935 4085.265 1189.16 ;
      RECT 4082.465 1048.035 4082.745 1181.56 ;
      RECT 4081.905 1048.035 4082.185 1181.32 ;
      RECT 4081.345 1048.035 4081.625 1181.08 ;
      RECT 4080.785 1048.035 4081.065 1180.84 ;
      RECT 4080.225 1048.035 4080.505 1180.6 ;
      RECT 4079.665 1048.035 4079.945 1180.36 ;
      RECT 4079.105 1048.035 4079.385 1180.12 ;
      RECT 4053.065 1048.035 4053.345 1193.995 ;
      RECT 4052.505 1048.035 4052.785 1194.235 ;
      RECT 4051.945 1048.035 4052.225 1194.475 ;
      RECT 4051.385 1048.035 4051.665 1194.715 ;
      RECT 4050.825 1048.035 4051.105 1194.955 ;
      RECT 4050.265 1046.935 4050.545 1194.955 ;
      RECT 4049.705 1048.035 4049.985 1194.715 ;
      RECT 4049.145 1046.935 4049.425 1194.47 ;
      RECT 4048.585 1048.035 4048.865 1194.23 ;
      RECT 4048.025 1046.935 4048.305 1193.99 ;
      RECT 4047.465 1048.035 4047.745 1193.75 ;
      RECT 4046.905 1048.035 4047.185 1193.51 ;
      RECT 4046.345 1048.035 4046.625 1193.27 ;
      RECT 4045.785 1048.035 4046.065 1193.03 ;
      RECT 4045.225 1048.035 4045.505 1192.79 ;
      RECT 4044.665 1048.035 4044.945 1192.55 ;
      RECT 4044.105 1048.035 4044.385 1192.31 ;
      RECT 4043.545 1048.035 4043.825 1192.07 ;
      RECT 4042.985 1046.935 4043.265 1191.83 ;
      RECT 4042.425 1048.035 4042.705 1191.59 ;
      RECT 4041.865 1046.935 4042.145 1191.35 ;
      RECT 4041.305 1048.035 4041.585 1191.11 ;
      RECT 4040.745 1048.035 4041.025 1190.87 ;
      RECT 4040.185 1048.035 4040.465 1190.63 ;
      RECT 4026.745 1048.035 4027.025 1194.03 ;
      RECT 4026.185 1048.035 4026.465 1194.27 ;
      RECT 4025.625 1048.035 4025.905 1194.515 ;
      RECT 4025.065 1048.035 4025.345 1194.755 ;
      RECT 4024.505 1048.035 4024.785 1194.995 ;
      RECT 4023.945 1048.035 4024.225 1194.995 ;
      RECT 4023.385 1048.035 4023.665 1194.755 ;
      RECT 4022.825 1048.035 4023.105 1194.515 ;
      RECT 4022.265 1048.035 4022.545 1187.5 ;
      RECT 4021.705 1048.035 4021.985 1187.26 ;
      RECT 4021.145 1048.035 4021.425 1187.02 ;
      RECT 4020.585 1046.935 4020.865 1186.78 ;
      RECT 4020.025 1048.035 4020.305 1186.54 ;
      RECT 4019.465 1046.935 4019.745 1186.3 ;
      RECT 4018.905 1048.035 4019.185 1186.06 ;
      RECT 4018.345 1048.035 4018.625 1185.82 ;
      RECT 4017.785 1048.035 4018.065 1185.58 ;
      RECT 4017.225 1046.935 4017.505 1185.34 ;
      RECT 4016.665 1048.035 4016.945 1185.1 ;
      RECT 4016.105 1046.935 4016.385 1184.86 ;
      RECT 4015.545 1048.035 4015.825 1184.62 ;
      RECT 4014.985 1046.935 4015.265 1184.38 ;
      RECT 4014.425 1048.035 4014.705 1184.14 ;
      RECT 4013.865 1048.035 4014.145 1183.9 ;
      RECT 3973.545 1048.035 3973.825 1192.795 ;
      RECT 3972.985 1048.035 3973.265 1193.035 ;
      RECT 3972.425 1048.035 3972.705 1193.28 ;
      RECT 3971.865 1048.035 3972.145 1193.52 ;
      RECT 3971.305 1048.035 3971.585 1193.76 ;
      RECT 3970.745 1048.035 3971.025 1194 ;
      RECT 3970.185 1048.035 3970.465 1194.24 ;
      RECT 3969.625 1048.035 3969.905 1194.48 ;
      RECT 3969.065 1048.035 3969.345 1194.72 ;
      RECT 3968.505 1048.035 3968.785 1194.96 ;
      RECT 3967.945 1046.935 3968.225 1195.2 ;
      RECT 3967.385 1048.035 3967.665 1195.44 ;
      RECT 3966.825 1046.935 3967.105 1195.68 ;
      RECT 3966.265 1048.035 3966.545 1195.92 ;
      RECT 3965.705 1046.935 3965.985 1196.16 ;
      RECT 3965.145 1048.035 3965.425 1196.16 ;
      RECT 3964.585 1048.035 3964.865 1195.92 ;
      RECT 3964.025 1048.035 3964.305 1195.68 ;
      RECT 3963.465 1048.035 3963.745 1195.44 ;
      RECT 3962.905 1048.035 3963.185 1195.2 ;
      RECT 3962.345 1048.035 3962.625 1194.96 ;
      RECT 3961.785 1048.035 3962.065 1194.72 ;
      RECT 3961.225 1048.035 3961.505 1194.48 ;
      RECT 3952.265 1046.935 3952.545 1194.51 ;
      RECT 3951.705 1048.035 3951.985 1194.75 ;
      RECT 3951.145 1046.935 3951.425 1194.99 ;
      RECT 3950.585 1048.035 3950.865 1195.205 ;
      RECT 3950.025 1048.035 3950.305 1194.78 ;
      RECT 3949.465 1048.035 3949.745 1194.54 ;
      RECT 3948.905 1048.035 3949.185 1194.3 ;
      RECT 3948.345 1048.035 3948.625 1194.06 ;
      RECT 3947.785 1048.035 3948.065 1193.82 ;
      RECT 3947.225 1048.035 3947.505 1193.58 ;
      RECT 3946.665 1048.035 3946.945 1193.34 ;
      RECT 3946.105 1048.035 3946.385 1193.1 ;
      RECT 3945.545 1048.035 3945.825 1192.86 ;
      RECT 3944.985 1048.035 3945.265 1192.62 ;
      RECT 3942.465 1048.035 3942.745 1191.795 ;
      RECT 3941.905 1048.035 3942.185 1191.555 ;
      RECT 3941.345 1048.035 3941.625 1191.315 ;
      RECT 3940.785 1046.935 3941.065 1191.075 ;
      RECT 3940.225 1048.035 3940.505 1190.835 ;
      RECT 3939.665 1046.935 3939.945 1190.595 ;
      RECT 3939.105 1048.035 3939.385 1190.355 ;
      RECT 3938.545 1048.035 3938.825 1190.115 ;
      RECT 3911.945 1048.035 3912.225 1201.16 ;
      RECT 3911.385 1046.935 3911.665 1201.4 ;
      RECT 3910.825 1048.035 3911.105 1201.64 ;
      RECT 3910.265 1046.935 3910.545 1201.885 ;
      RECT 3909.705 1048.035 3909.985 1202.125 ;
      RECT 3909.145 1046.935 3909.425 1202.365 ;
      RECT 3908.585 1048.035 3908.865 1202.605 ;
      RECT 3908.025 1048.035 3908.305 1202.845 ;
      RECT 3907.465 1048.035 3907.745 1188.465 ;
      RECT 3906.905 1048.035 3907.185 1188.225 ;
      RECT 3906.345 1048.035 3906.625 1187.985 ;
      RECT 3905.785 1048.035 3906.065 1187.745 ;
      RECT 3905.225 1048.035 3905.505 1187.505 ;
      RECT 3904.665 1048.035 3904.945 1187.265 ;
      RECT 3904.105 1048.035 3904.385 1187.025 ;
      RECT 3903.545 1048.035 3903.825 1186.785 ;
      RECT 3902.985 1048.035 3903.265 1186.545 ;
      RECT 3902.425 1048.035 3902.705 1186.305 ;
      RECT 3901.865 1046.935 3902.145 1186.065 ;
      RECT 3901.305 1048.035 3901.585 1185.825 ;
      RECT 3900.745 1046.935 3901.025 1185.585 ;
      RECT 3900.185 1048.035 3900.465 1185.345 ;
      RECT 3886.185 1046.935 3886.465 1191.465 ;
      RECT 3885.625 1048.035 3885.905 1191.225 ;
      RECT 3885.065 1048.035 3885.345 1190.985 ;
      RECT 3884.505 1048.035 3884.785 1190.745 ;
      RECT 3883.945 1048.035 3884.225 1190.505 ;
      RECT 3883.385 1048.035 3883.665 1190.265 ;
      RECT 3882.825 1048.035 3883.105 1190.025 ;
      RECT 3882.265 1048.035 3882.545 1189.785 ;
      RECT 3881.705 1048.035 3881.985 1189.545 ;
      RECT 3881.145 1046.935 3881.425 1189.305 ;
      RECT 3880.585 1048.035 3880.865 1189.065 ;
      RECT 3880.025 1046.935 3880.305 1188.825 ;
      RECT 3879.465 1048.035 3879.745 1188.585 ;
      RECT 3878.905 1048.035 3879.185 1188.345 ;
      RECT 3878.345 1048.035 3878.625 1188.105 ;
      RECT 3877.785 1048.035 3878.065 1187.865 ;
      RECT 3877.225 1048.035 3877.505 1187.625 ;
      RECT 3876.665 1048.035 3876.945 1187.385 ;
      RECT 3876.105 1048.035 3876.385 1187.145 ;
      RECT 3875.545 1048.035 3875.825 1186.905 ;
      RECT 3874.985 1048.035 3875.265 1186.665 ;
      RECT 3874.425 1048.035 3874.705 1186.425 ;
      RECT 3873.865 1048.035 3874.145 1186.185 ;
      RECT 3834.665 1048.035 3834.945 1193.09 ;
      RECT 3834.105 1048.035 3834.385 1193.33 ;
      RECT 3833.545 1048.035 3833.825 1193.57 ;
      RECT 3832.985 1046.935 3833.265 1193.81 ;
      RECT 3832.425 1048.035 3832.705 1194.05 ;
      RECT 3831.865 1046.935 3832.145 1194.29 ;
      RECT 3831.305 1048.035 3831.585 1194.53 ;
      RECT 3830.745 1048.035 3831.025 1194.77 ;
      RECT 3830.185 1048.035 3830.465 1195.01 ;
      RECT 3829.625 1046.935 3829.905 1195.25 ;
      RECT 3829.065 1048.035 3829.345 1195.49 ;
      RECT 3828.505 1046.935 3828.785 1195.73 ;
      RECT 3827.945 1048.035 3828.225 1195.97 ;
      RECT 3827.385 1046.935 3827.665 1196.21 ;
      RECT 3826.825 1048.035 3827.105 1196.45 ;
      RECT 3826.265 1048.035 3826.545 1196.69 ;
      RECT 3825.705 1048.035 3825.985 1196.69 ;
      RECT 3825.145 1048.035 3825.425 1196.45 ;
      RECT 3824.585 1048.035 3824.865 1196.21 ;
      RECT 3824.025 1048.035 3824.305 1195.97 ;
      RECT 3823.465 1048.035 3823.745 1195.73 ;
      RECT 3822.905 1048.035 3823.185 1195.49 ;
      RECT 3822.345 1048.035 3822.625 1195.25 ;
      RECT 3821.785 1048.035 3822.065 1195.01 ;
      RECT 3821.225 1048.035 3821.505 1194.77 ;
      RECT 3812.265 1048.035 3812.545 1194.285 ;
      RECT 3811.705 1046.935 3811.985 1194.045 ;
      RECT 3811.145 1048.035 3811.425 1193.805 ;
      RECT 3810.585 1046.935 3810.865 1193.565 ;
      RECT 3810.025 1048.035 3810.305 1193.325 ;
      RECT 3809.465 1046.935 3809.745 1193.085 ;
      RECT 3808.905 1048.035 3809.185 1192.845 ;
      RECT 3808.345 1048.035 3808.625 1192.605 ;
      RECT 3807.785 1048.035 3808.065 1192.365 ;
      RECT 3807.225 1048.035 3807.505 1192.125 ;
      RECT 3806.665 1048.035 3806.945 1191.885 ;
      RECT 3806.105 1048.035 3806.385 1191.645 ;
      RECT 3805.545 1048.035 3805.825 1191.405 ;
      RECT 3804.985 1048.035 3805.265 1191.165 ;
      RECT 3802.465 1046.935 3802.745 1192.885 ;
      RECT 3801.905 1048.035 3802.185 1192.645 ;
      RECT 3801.345 1046.935 3801.625 1192.405 ;
      RECT 3800.785 1048.035 3801.065 1192.165 ;
      RECT 3800.225 1048.035 3800.505 1191.925 ;
      RECT 3799.665 1048.035 3799.945 1191.685 ;
      RECT 3799.105 1048.035 3799.385 1191.445 ;
      RECT 3798.545 1048.035 3798.825 1191.205 ;
      RECT 3772.505 1048.035 3772.785 1188.855 ;
      RECT 3771.945 1048.035 3772.225 1189.095 ;
      RECT 3771.385 1048.035 3771.665 1189.335 ;
      RECT 3770.825 1048.035 3771.105 1189.58 ;
      RECT 3770.265 1048.035 3770.545 1189.82 ;
      RECT 3769.705 1048.035 3769.985 1190.06 ;
      RECT 3769.145 1048.035 3769.425 1190.06 ;
      RECT 3768.585 1048.035 3768.865 1189.82 ;
      RECT 3768.025 1048.035 3768.305 1189.58 ;
      RECT 3767.465 1046.935 3767.745 1189.34 ;
      RECT 3766.905 1048.035 3767.185 1189.1 ;
      RECT 3766.345 1046.935 3766.625 1188.86 ;
      RECT 3765.785 1048.035 3766.065 1188.62 ;
      RECT 3765.225 1048.035 3765.505 1188.38 ;
      RECT 3764.665 1048.035 3764.945 1188.14 ;
      RECT 3764.105 1046.935 3764.385 1187.9 ;
      RECT 3763.545 1048.035 3763.825 1187.66 ;
      RECT 3762.985 1046.935 3763.265 1187.42 ;
      RECT 3762.425 1048.035 3762.705 1187.18 ;
      RECT 3761.865 1046.935 3762.145 1186.94 ;
      RECT 3761.305 1048.035 3761.585 1186.7 ;
      RECT 3760.745 1048.035 3761.025 1186.46 ;
      RECT 3760.185 1048.035 3760.465 1186.22 ;
      RECT 3759.625 1048.035 3759.905 1185.98 ;
      RECT 3746.185 1048.035 3746.465 1191.78 ;
      RECT 3745.625 1048.035 3745.905 1191.54 ;
      RECT 3745.065 1048.035 3745.345 1191.3 ;
      RECT 3744.505 1048.035 3744.785 1191.06 ;
      RECT 3743.945 1048.035 3744.225 1190.82 ;
      RECT 3743.385 1048.035 3743.665 1190.58 ;
      RECT 3742.825 1048.035 3743.105 1190.34 ;
      RECT 3742.265 1048.035 3742.545 1190.1 ;
      RECT 3741.705 1046.935 3741.985 1189.86 ;
      RECT 3741.145 1048.035 3741.425 1189.62 ;
      RECT 3740.585 1046.935 3740.865 1189.3 ;
      RECT 3740.025 1048.035 3740.305 1189.14 ;
      RECT 3739.465 1046.935 3739.745 1188.9 ;
      RECT 3738.905 1048.035 3739.185 1188.66 ;
      RECT 3738.345 1048.035 3738.625 1188.42 ;
      RECT 3737.785 1048.035 3738.065 1188.18 ;
      RECT 3737.225 1048.035 3737.505 1187.94 ;
      RECT 3736.665 1048.035 3736.945 1187.7 ;
      RECT 3736.105 1048.035 3736.385 1187.46 ;
      RECT 3735.545 1048.035 3735.825 1187.22 ;
      RECT 3734.985 1048.035 3735.265 1186.98 ;
      RECT 3734.425 1046.935 3734.705 1186.74 ;
      RECT 3733.865 1048.035 3734.145 1186.5 ;
      RECT 3733.305 1046.935 3733.585 1186.26 ;
      RECT 3694.105 1048.035 3694.385 1191.87 ;
      RECT 3693.545 1048.035 3693.825 1192.11 ;
      RECT 3692.985 1048.035 3693.265 1192.35 ;
      RECT 3692.425 1048.035 3692.705 1192.59 ;
      RECT 3691.865 1048.035 3692.145 1192.83 ;
      RECT 3691.305 1048.035 3691.585 1193.07 ;
      RECT 3690.745 1048.035 3691.025 1193.31 ;
      RECT 3690.185 1048.035 3690.465 1193.55 ;
      RECT 3689.625 1048.035 3689.905 1193.79 ;
      RECT 3689.065 1048.035 3689.345 1194.03 ;
      RECT 3688.505 1048.035 3688.785 1194.27 ;
      RECT 3687.945 1048.035 3688.225 1194.51 ;
      RECT 3687.385 1048.035 3687.665 1194.75 ;
      RECT 3686.825 1048.035 3687.105 1194.75 ;
      RECT 3686.265 1046.935 3686.545 1194.51 ;
      RECT 3685.705 1048.035 3685.985 1194.27 ;
      RECT 3685.145 1046.935 3685.425 1194.03 ;
      RECT 3684.585 1048.035 3684.865 1193.79 ;
      RECT 3684.025 1048.035 3684.305 1193.55 ;
      RECT 3683.465 1048.035 3683.745 1193.31 ;
      RECT 3682.905 1046.935 3683.185 1193.045 ;
      RECT 3682.345 1048.035 3682.625 1192.805 ;
      RECT 3681.785 1046.935 3682.065 1192.565 ;
      RECT 3681.225 1048.035 3681.505 1192.325 ;
      RECT 3672.265 1046.935 3672.545 1186.16 ;
      RECT 3671.705 1048.035 3671.985 1186.4 ;
      RECT 3671.145 1048.035 3671.425 1186.64 ;
      RECT 3670.585 1048.035 3670.865 1186.64 ;
      RECT 3670.025 1048.035 3670.305 1186.4 ;
      RECT 3669.465 1048.035 3669.745 1186.16 ;
      RECT 3668.905 1048.035 3669.185 1185.92 ;
      RECT 3668.345 1048.035 3668.625 1185.68 ;
      RECT 3667.785 1048.035 3668.065 1185.44 ;
      RECT 3667.225 1048.035 3667.505 1185.2 ;
      RECT 3666.665 1048.035 3666.945 1184.96 ;
      RECT 3666.105 1048.035 3666.385 1184.72 ;
      RECT 3665.545 1048.035 3665.825 1184.48 ;
      RECT 3664.985 1046.935 3665.265 1184.24 ;
      RECT 3662.465 1048.035 3662.745 1185.96 ;
      RECT 3661.905 1046.935 3662.185 1185.72 ;
      RECT 3661.345 1048.035 3661.625 1185.48 ;
      RECT 3660.785 1046.935 3661.065 1185.24 ;
      RECT 3660.225 1048.035 3660.505 1185 ;
      RECT 3659.665 1048.035 3659.945 1184.76 ;
      RECT 3659.105 1048.035 3659.385 1184.52 ;
      RECT 3633.065 1048.035 3633.345 1187.305 ;
      RECT 3632.505 1048.035 3632.785 1187.545 ;
      RECT 3631.945 1048.035 3632.225 1187.785 ;
      RECT 3631.385 1048.035 3631.665 1188.025 ;
      RECT 3630.825 1048.035 3631.105 1188.265 ;
      RECT 3630.265 1046.935 3630.545 1188.505 ;
      RECT 3629.705 1048.035 3629.985 1188.745 ;
      RECT 3629.145 1046.935 3629.425 1188.985 ;
      RECT 3628.585 1048.035 3628.865 1189.225 ;
      RECT 3628.025 1048.035 3628.305 1189.465 ;
      RECT 3627.465 1048.035 3627.745 1189.705 ;
      RECT 3626.905 1048.035 3627.185 1189.945 ;
      RECT 3626.345 1048.035 3626.625 1190.185 ;
      RECT 3625.785 1048.035 3626.065 1190.425 ;
      RECT 3625.225 1048.035 3625.505 1190.665 ;
      RECT 3624.665 1048.035 3624.945 1190.665 ;
      RECT 3624.105 1048.035 3624.385 1190.425 ;
      RECT 3623.545 1048.035 3623.825 1190.185 ;
      RECT 3622.985 1048.035 3623.265 1189.945 ;
      RECT 3622.425 1048.035 3622.705 1189.7 ;
      RECT 3621.865 1048.035 3622.145 1189.46 ;
      RECT 3621.305 1048.035 3621.585 1189.22 ;
      RECT 3620.745 1046.935 3621.025 1188.98 ;
      RECT 3620.185 1048.035 3620.465 1188.74 ;
      RECT 3606.745 1046.935 3607.025 1186.22 ;
      RECT 3606.185 1048.035 3606.465 1185.98 ;
      RECT 3605.625 1048.035 3605.905 1185.74 ;
      RECT 3605.065 1048.035 3605.345 1185.5 ;
      RECT 3604.505 1046.935 3604.785 1185.26 ;
      RECT 3603.945 1048.035 3604.225 1185.02 ;
      RECT 3603.385 1046.935 3603.665 1184.78 ;
      RECT 3602.825 1048.035 3603.105 1184.54 ;
      RECT 3602.265 1046.935 3602.545 1184.3 ;
      RECT 3601.705 1048.035 3601.985 1184.06 ;
      RECT 3601.145 1048.035 3601.425 1183.82 ;
      RECT 3600.585 1048.035 3600.865 1183.58 ;
      RECT 3600.025 1048.035 3600.305 1183.34 ;
      RECT 3599.465 1048.035 3599.745 1183.1 ;
      RECT 3598.905 1048.035 3599.185 1182.86 ;
      RECT 3598.345 1048.035 3598.625 1182.62 ;
      RECT 3597.785 1048.035 3598.065 1182.38 ;
      RECT 3597.225 1048.035 3597.505 1182.14 ;
      RECT 3596.665 1048.035 3596.945 1181.9 ;
      RECT 3596.105 1048.035 3596.385 1181.66 ;
      RECT 3595.545 1048.035 3595.825 1181.42 ;
      RECT 3594.985 1046.935 3595.265 1181.18 ;
      RECT 3594.425 1048.035 3594.705 1180.94 ;
      RECT 3593.865 1046.935 3594.145 1180.7 ;
      RECT 3554.105 1048.035 3554.385 1191.17 ;
      RECT 3553.545 1046.935 3553.825 1191.41 ;
      RECT 3552.985 1048.035 3553.265 1191.65 ;
      RECT 3552.425 1048.035 3552.705 1191.89 ;
      RECT 3551.865 1048.035 3552.145 1192.13 ;
      RECT 3551.305 1048.035 3551.585 1192.37 ;
      RECT 3550.745 1048.035 3551.025 1192.61 ;
      RECT 3550.185 1048.035 3550.465 1192.855 ;
      RECT 3549.625 1048.035 3549.905 1193.095 ;
      RECT 3549.065 1048.035 3549.345 1193.335 ;
      RECT 3548.505 1046.935 3548.785 1193.575 ;
      RECT 3547.945 1048.035 3548.225 1193.815 ;
      RECT 3547.385 1046.935 3547.665 1194.055 ;
      RECT 3546.825 1048.035 3547.105 1194.295 ;
      RECT 3546.265 1048.035 3546.545 1194.535 ;
      RECT 3545.705 1048.035 3545.985 1194.775 ;
      RECT 3545.145 1048.035 3545.425 1195.015 ;
      RECT 3544.585 1048.035 3544.865 1195.255 ;
      RECT 3544.025 1048.035 3544.305 1195.495 ;
      RECT 3543.465 1048.035 3543.745 1195.735 ;
      RECT 3542.905 1048.035 3543.185 1195.975 ;
      RECT 3542.345 1048.035 3542.625 1196.215 ;
      RECT 3541.785 1048.035 3542.065 1196.455 ;
      RECT 3541.225 1048.035 3541.505 1196.695 ;
      RECT 3532.265 1048.035 3532.545 1192.28 ;
      RECT 3531.705 1048.035 3531.985 1192.04 ;
      RECT 3531.145 1048.035 3531.425 1191.8 ;
      RECT 3530.585 1046.935 3530.865 1191.56 ;
      RECT 3530.025 1048.035 3530.305 1191.32 ;
      RECT 3529.465 1046.935 3529.745 1191.08 ;
      RECT 3528.905 1048.035 3529.185 1190.84 ;
      RECT 3528.345 1048.035 3528.625 1190.6 ;
      RECT 3527.785 1048.035 3528.065 1190.36 ;
      RECT 3527.225 1046.935 3527.505 1190.12 ;
      RECT 3526.665 1048.035 3526.945 1189.88 ;
      RECT 3526.105 1046.935 3526.385 1189.64 ;
      RECT 3525.545 1048.035 3525.825 1189.4 ;
      RECT 3524.985 1046.935 3525.265 1189.16 ;
      RECT 3522.465 1048.035 3522.745 1181.56 ;
      RECT 3521.905 1048.035 3522.185 1181.32 ;
      RECT 3521.345 1048.035 3521.625 1181.08 ;
      RECT 3520.785 1048.035 3521.065 1180.84 ;
      RECT 3520.225 1048.035 3520.505 1180.6 ;
      RECT 3519.665 1048.035 3519.945 1180.36 ;
      RECT 3519.105 1048.035 3519.385 1180.12 ;
      RECT 3493.065 1048.035 3493.345 1193.995 ;
      RECT 3492.505 1048.035 3492.785 1194.235 ;
      RECT 3491.945 1048.035 3492.225 1194.475 ;
      RECT 3491.385 1048.035 3491.665 1194.715 ;
      RECT 3490.825 1048.035 3491.105 1194.955 ;
      RECT 3490.265 1046.935 3490.545 1194.955 ;
      RECT 3489.705 1048.035 3489.985 1194.715 ;
      RECT 3489.145 1046.935 3489.425 1194.47 ;
      RECT 3488.585 1048.035 3488.865 1194.23 ;
      RECT 3488.025 1046.935 3488.305 1193.99 ;
      RECT 3487.465 1048.035 3487.745 1193.75 ;
      RECT 3486.905 1048.035 3487.185 1193.51 ;
      RECT 3486.345 1048.035 3486.625 1193.27 ;
      RECT 3485.785 1048.035 3486.065 1193.03 ;
      RECT 3485.225 1048.035 3485.505 1192.79 ;
      RECT 3484.665 1048.035 3484.945 1192.55 ;
      RECT 3484.105 1048.035 3484.385 1192.31 ;
      RECT 3483.545 1048.035 3483.825 1192.07 ;
      RECT 3482.985 1046.935 3483.265 1191.83 ;
      RECT 3482.425 1048.035 3482.705 1191.59 ;
      RECT 3481.865 1046.935 3482.145 1191.35 ;
      RECT 3481.305 1048.035 3481.585 1191.11 ;
      RECT 3480.745 1048.035 3481.025 1190.87 ;
      RECT 3480.185 1048.035 3480.465 1190.63 ;
      RECT 3466.745 1048.035 3467.025 1194.03 ;
      RECT 3466.185 1048.035 3466.465 1194.27 ;
      RECT 3465.625 1048.035 3465.905 1194.515 ;
      RECT 3465.065 1048.035 3465.345 1194.755 ;
      RECT 3464.505 1048.035 3464.785 1194.995 ;
      RECT 3463.945 1048.035 3464.225 1194.995 ;
      RECT 3463.385 1048.035 3463.665 1194.755 ;
      RECT 3462.825 1048.035 3463.105 1194.515 ;
      RECT 3462.265 1048.035 3462.545 1187.5 ;
      RECT 3461.705 1048.035 3461.985 1187.26 ;
      RECT 3461.145 1048.035 3461.425 1187.02 ;
      RECT 3460.585 1046.935 3460.865 1186.78 ;
      RECT 3460.025 1048.035 3460.305 1186.54 ;
      RECT 3459.465 1046.935 3459.745 1186.3 ;
      RECT 3458.905 1048.035 3459.185 1186.06 ;
      RECT 3458.345 1048.035 3458.625 1185.82 ;
      RECT 3457.785 1048.035 3458.065 1185.58 ;
      RECT 3457.225 1046.935 3457.505 1185.34 ;
      RECT 3456.665 1048.035 3456.945 1185.1 ;
      RECT 3456.105 1046.935 3456.385 1184.86 ;
      RECT 3455.545 1048.035 3455.825 1184.62 ;
      RECT 3454.985 1046.935 3455.265 1184.38 ;
      RECT 3454.425 1048.035 3454.705 1184.14 ;
      RECT 3453.865 1048.035 3454.145 1183.9 ;
      RECT 3413.545 1048.035 3413.825 1192.795 ;
      RECT 3412.985 1048.035 3413.265 1193.035 ;
      RECT 3412.425 1048.035 3412.705 1193.28 ;
      RECT 3411.865 1048.035 3412.145 1193.52 ;
      RECT 3411.305 1048.035 3411.585 1193.76 ;
      RECT 3410.745 1048.035 3411.025 1194 ;
      RECT 3410.185 1048.035 3410.465 1194.24 ;
      RECT 3409.625 1048.035 3409.905 1194.48 ;
      RECT 3409.065 1048.035 3409.345 1194.72 ;
      RECT 3408.505 1048.035 3408.785 1194.96 ;
      RECT 3407.945 1046.935 3408.225 1195.2 ;
      RECT 3407.385 1048.035 3407.665 1195.44 ;
      RECT 3406.825 1046.935 3407.105 1195.68 ;
      RECT 3406.265 1048.035 3406.545 1195.92 ;
      RECT 3405.705 1046.935 3405.985 1196.16 ;
      RECT 3405.145 1048.035 3405.425 1196.16 ;
      RECT 3404.585 1048.035 3404.865 1195.92 ;
      RECT 3404.025 1048.035 3404.305 1195.68 ;
      RECT 3403.465 1048.035 3403.745 1195.44 ;
      RECT 3402.905 1048.035 3403.185 1195.2 ;
      RECT 3402.345 1048.035 3402.625 1194.96 ;
      RECT 3401.785 1048.035 3402.065 1194.72 ;
      RECT 3401.225 1048.035 3401.505 1194.48 ;
      RECT 3392.265 1046.935 3392.545 1194.51 ;
      RECT 3391.705 1048.035 3391.985 1194.75 ;
      RECT 3391.145 1046.935 3391.425 1194.99 ;
      RECT 3390.585 1048.035 3390.865 1195.205 ;
      RECT 3390.025 1048.035 3390.305 1194.78 ;
      RECT 3389.465 1048.035 3389.745 1194.54 ;
      RECT 3388.905 1048.035 3389.185 1194.3 ;
      RECT 3388.345 1048.035 3388.625 1194.06 ;
      RECT 3387.785 1048.035 3388.065 1193.82 ;
      RECT 3387.225 1048.035 3387.505 1193.58 ;
      RECT 3386.665 1048.035 3386.945 1193.34 ;
      RECT 3386.105 1048.035 3386.385 1193.1 ;
      RECT 3385.545 1048.035 3385.825 1192.86 ;
      RECT 3384.985 1048.035 3385.265 1192.62 ;
      RECT 3382.465 1048.035 3382.745 1191.795 ;
      RECT 3381.905 1048.035 3382.185 1191.555 ;
      RECT 3381.345 1048.035 3381.625 1191.315 ;
      RECT 3380.785 1046.935 3381.065 1191.075 ;
      RECT 3380.225 1048.035 3380.505 1190.835 ;
      RECT 3379.665 1046.935 3379.945 1190.595 ;
      RECT 3379.105 1048.035 3379.385 1190.355 ;
      RECT 3378.545 1048.035 3378.825 1190.115 ;
      RECT 3351.945 1048.035 3352.225 1201.16 ;
      RECT 3351.385 1046.935 3351.665 1201.4 ;
      RECT 3350.825 1048.035 3351.105 1201.64 ;
      RECT 3350.265 1046.935 3350.545 1201.885 ;
      RECT 3349.705 1048.035 3349.985 1202.125 ;
      RECT 3349.145 1046.935 3349.425 1202.365 ;
      RECT 3348.585 1048.035 3348.865 1202.605 ;
      RECT 3348.025 1048.035 3348.305 1202.845 ;
      RECT 3347.465 1048.035 3347.745 1188.465 ;
      RECT 3346.905 1048.035 3347.185 1188.225 ;
      RECT 3346.345 1048.035 3346.625 1187.985 ;
      RECT 3345.785 1048.035 3346.065 1187.745 ;
      RECT 3345.225 1048.035 3345.505 1187.505 ;
      RECT 3344.665 1048.035 3344.945 1187.265 ;
      RECT 3344.105 1048.035 3344.385 1187.025 ;
      RECT 3343.545 1048.035 3343.825 1186.785 ;
      RECT 3342.985 1048.035 3343.265 1186.545 ;
      RECT 3342.425 1048.035 3342.705 1186.305 ;
      RECT 3341.865 1046.935 3342.145 1186.065 ;
      RECT 3341.305 1048.035 3341.585 1185.825 ;
      RECT 3340.745 1046.935 3341.025 1185.585 ;
      RECT 3340.185 1048.035 3340.465 1185.345 ;
      RECT 3326.185 1046.935 3326.465 1191.465 ;
      RECT 3325.625 1048.035 3325.905 1191.225 ;
      RECT 3325.065 1048.035 3325.345 1190.985 ;
      RECT 3324.505 1048.035 3324.785 1190.745 ;
      RECT 3323.945 1048.035 3324.225 1190.505 ;
      RECT 3323.385 1048.035 3323.665 1190.265 ;
      RECT 3322.825 1048.035 3323.105 1190.025 ;
      RECT 3322.265 1048.035 3322.545 1189.785 ;
      RECT 3321.705 1048.035 3321.985 1189.545 ;
      RECT 3321.145 1046.935 3321.425 1189.305 ;
      RECT 3320.585 1048.035 3320.865 1189.065 ;
      RECT 3320.025 1046.935 3320.305 1188.825 ;
      RECT 3319.465 1048.035 3319.745 1188.585 ;
      RECT 3318.905 1048.035 3319.185 1188.345 ;
      RECT 3318.345 1048.035 3318.625 1188.105 ;
      RECT 3317.785 1048.035 3318.065 1187.865 ;
      RECT 3317.225 1048.035 3317.505 1187.625 ;
      RECT 3316.665 1048.035 3316.945 1187.385 ;
      RECT 3316.105 1048.035 3316.385 1187.145 ;
      RECT 3315.545 1048.035 3315.825 1186.905 ;
      RECT 3314.985 1048.035 3315.265 1186.665 ;
      RECT 3314.425 1048.035 3314.705 1186.425 ;
      RECT 3313.865 1048.035 3314.145 1186.185 ;
      RECT 3274.665 1048.035 3274.945 1193.09 ;
      RECT 3274.105 1048.035 3274.385 1193.33 ;
      RECT 3273.545 1048.035 3273.825 1193.57 ;
      RECT 3272.985 1046.935 3273.265 1193.81 ;
      RECT 3272.425 1048.035 3272.705 1194.05 ;
      RECT 3271.865 1046.935 3272.145 1194.29 ;
      RECT 3271.305 1048.035 3271.585 1194.53 ;
      RECT 3270.745 1048.035 3271.025 1194.77 ;
      RECT 3270.185 1048.035 3270.465 1195.01 ;
      RECT 3269.625 1046.935 3269.905 1195.25 ;
      RECT 3269.065 1048.035 3269.345 1195.49 ;
      RECT 3268.505 1046.935 3268.785 1195.73 ;
      RECT 3267.945 1048.035 3268.225 1195.97 ;
      RECT 3267.385 1046.935 3267.665 1196.21 ;
      RECT 3266.825 1048.035 3267.105 1196.45 ;
      RECT 3266.265 1048.035 3266.545 1196.69 ;
      RECT 3265.705 1048.035 3265.985 1196.69 ;
      RECT 3265.145 1048.035 3265.425 1196.45 ;
      RECT 3264.585 1048.035 3264.865 1196.21 ;
      RECT 3264.025 1048.035 3264.305 1195.97 ;
      RECT 3263.465 1048.035 3263.745 1195.73 ;
      RECT 3262.905 1048.035 3263.185 1195.49 ;
      RECT 3262.345 1048.035 3262.625 1195.25 ;
      RECT 3261.785 1048.035 3262.065 1195.01 ;
      RECT 3261.225 1048.035 3261.505 1194.77 ;
      RECT 3252.265 1048.035 3252.545 1194.285 ;
      RECT 3251.705 1046.935 3251.985 1194.045 ;
      RECT 3251.145 1048.035 3251.425 1193.805 ;
      RECT 3250.585 1046.935 3250.865 1193.565 ;
      RECT 3250.025 1048.035 3250.305 1193.325 ;
      RECT 3249.465 1046.935 3249.745 1193.085 ;
      RECT 3248.905 1048.035 3249.185 1192.845 ;
      RECT 3248.345 1048.035 3248.625 1192.605 ;
      RECT 3247.785 1048.035 3248.065 1192.365 ;
      RECT 3247.225 1048.035 3247.505 1192.125 ;
      RECT 3246.665 1048.035 3246.945 1191.885 ;
      RECT 3246.105 1048.035 3246.385 1191.645 ;
      RECT 3245.545 1048.035 3245.825 1191.405 ;
      RECT 3244.985 1048.035 3245.265 1191.165 ;
      RECT 3242.465 1046.935 3242.745 1192.885 ;
      RECT 3241.905 1048.035 3242.185 1192.645 ;
      RECT 3241.345 1046.935 3241.625 1192.405 ;
      RECT 3240.785 1048.035 3241.065 1192.165 ;
      RECT 3240.225 1048.035 3240.505 1191.925 ;
      RECT 3239.665 1048.035 3239.945 1191.685 ;
      RECT 3239.105 1048.035 3239.385 1191.445 ;
      RECT 3238.545 1048.035 3238.825 1191.205 ;
      RECT 3212.505 1048.035 3212.785 1188.855 ;
      RECT 3211.945 1048.035 3212.225 1189.095 ;
      RECT 3211.385 1048.035 3211.665 1189.335 ;
      RECT 3210.825 1048.035 3211.105 1189.58 ;
      RECT 3210.265 1048.035 3210.545 1189.82 ;
      RECT 3209.705 1048.035 3209.985 1190.06 ;
      RECT 3209.145 1048.035 3209.425 1190.06 ;
      RECT 3208.585 1048.035 3208.865 1189.82 ;
      RECT 3208.025 1048.035 3208.305 1189.58 ;
      RECT 3207.465 1046.935 3207.745 1189.34 ;
      RECT 3206.905 1048.035 3207.185 1189.1 ;
      RECT 3206.345 1046.935 3206.625 1188.86 ;
      RECT 3205.785 1048.035 3206.065 1188.62 ;
      RECT 3205.225 1048.035 3205.505 1188.38 ;
      RECT 3204.665 1048.035 3204.945 1188.14 ;
      RECT 3204.105 1046.935 3204.385 1187.9 ;
      RECT 3203.545 1048.035 3203.825 1187.66 ;
      RECT 3202.985 1046.935 3203.265 1187.42 ;
      RECT 3202.425 1048.035 3202.705 1187.18 ;
      RECT 3201.865 1046.935 3202.145 1186.94 ;
      RECT 3201.305 1048.035 3201.585 1186.7 ;
      RECT 3200.745 1048.035 3201.025 1186.46 ;
      RECT 3200.185 1048.035 3200.465 1186.22 ;
      RECT 3199.625 1048.035 3199.905 1185.98 ;
      RECT 3186.185 1048.035 3186.465 1191.78 ;
      RECT 3185.625 1048.035 3185.905 1191.54 ;
      RECT 3185.065 1048.035 3185.345 1191.3 ;
      RECT 3184.505 1048.035 3184.785 1191.06 ;
      RECT 3183.945 1048.035 3184.225 1190.82 ;
      RECT 3183.385 1048.035 3183.665 1190.58 ;
      RECT 3182.825 1048.035 3183.105 1190.34 ;
      RECT 3182.265 1048.035 3182.545 1190.1 ;
      RECT 3181.705 1046.935 3181.985 1189.86 ;
      RECT 3181.145 1048.035 3181.425 1189.62 ;
      RECT 3180.585 1046.935 3180.865 1189.3 ;
      RECT 3180.025 1048.035 3180.305 1189.14 ;
      RECT 3179.465 1046.935 3179.745 1188.9 ;
      RECT 3178.905 1048.035 3179.185 1188.66 ;
      RECT 3178.345 1048.035 3178.625 1188.42 ;
      RECT 3177.785 1048.035 3178.065 1188.18 ;
      RECT 3177.225 1048.035 3177.505 1187.94 ;
      RECT 3176.665 1048.035 3176.945 1187.7 ;
      RECT 3176.105 1048.035 3176.385 1187.46 ;
      RECT 3175.545 1048.035 3175.825 1187.22 ;
      RECT 3174.985 1048.035 3175.265 1186.98 ;
      RECT 3174.425 1046.935 3174.705 1186.74 ;
      RECT 3173.865 1048.035 3174.145 1186.5 ;
      RECT 3173.305 1046.935 3173.585 1186.26 ;
      RECT 3134.105 1048.035 3134.385 1191.87 ;
      RECT 3133.545 1048.035 3133.825 1192.11 ;
      RECT 3132.985 1048.035 3133.265 1192.35 ;
      RECT 3132.425 1048.035 3132.705 1192.59 ;
      RECT 3131.865 1048.035 3132.145 1192.83 ;
      RECT 3131.305 1048.035 3131.585 1193.07 ;
      RECT 3130.745 1048.035 3131.025 1193.31 ;
      RECT 3130.185 1048.035 3130.465 1193.55 ;
      RECT 3129.625 1048.035 3129.905 1193.79 ;
      RECT 3129.065 1048.035 3129.345 1194.03 ;
      RECT 3128.505 1048.035 3128.785 1194.27 ;
      RECT 3127.945 1048.035 3128.225 1194.51 ;
      RECT 3127.385 1048.035 3127.665 1194.75 ;
      RECT 3126.825 1048.035 3127.105 1194.75 ;
      RECT 3126.265 1046.935 3126.545 1194.51 ;
      RECT 3125.705 1048.035 3125.985 1194.27 ;
      RECT 3125.145 1046.935 3125.425 1194.03 ;
      RECT 3124.585 1048.035 3124.865 1193.79 ;
      RECT 3124.025 1048.035 3124.305 1193.55 ;
      RECT 3123.465 1048.035 3123.745 1193.31 ;
      RECT 3122.905 1046.935 3123.185 1193.045 ;
      RECT 3122.345 1048.035 3122.625 1192.805 ;
      RECT 3121.785 1046.935 3122.065 1192.565 ;
      RECT 3121.225 1048.035 3121.505 1192.325 ;
      RECT 3112.265 1046.935 3112.545 1186.16 ;
      RECT 3111.705 1048.035 3111.985 1186.4 ;
      RECT 3111.145 1048.035 3111.425 1186.64 ;
      RECT 3110.585 1048.035 3110.865 1186.64 ;
      RECT 3110.025 1048.035 3110.305 1186.4 ;
      RECT 3109.465 1048.035 3109.745 1186.16 ;
      RECT 3108.905 1048.035 3109.185 1185.92 ;
      RECT 3108.345 1048.035 3108.625 1185.68 ;
      RECT 3107.785 1048.035 3108.065 1185.44 ;
      RECT 3107.225 1048.035 3107.505 1185.2 ;
      RECT 3106.665 1048.035 3106.945 1184.96 ;
      RECT 3106.105 1048.035 3106.385 1184.72 ;
      RECT 3105.545 1048.035 3105.825 1184.48 ;
      RECT 3104.985 1046.935 3105.265 1184.24 ;
      RECT 3102.465 1048.035 3102.745 1185.96 ;
      RECT 3101.905 1046.935 3102.185 1185.72 ;
      RECT 3101.345 1048.035 3101.625 1185.48 ;
      RECT 3100.785 1046.935 3101.065 1185.24 ;
      RECT 3100.225 1048.035 3100.505 1185 ;
      RECT 3099.665 1048.035 3099.945 1184.76 ;
      RECT 3099.105 1048.035 3099.385 1184.52 ;
      RECT 3073.065 1048.035 3073.345 1187.305 ;
      RECT 3072.505 1048.035 3072.785 1187.545 ;
      RECT 3071.945 1048.035 3072.225 1187.785 ;
      RECT 3071.385 1048.035 3071.665 1188.025 ;
      RECT 3070.825 1048.035 3071.105 1188.265 ;
      RECT 3070.265 1046.935 3070.545 1188.505 ;
      RECT 3069.705 1048.035 3069.985 1188.745 ;
      RECT 3069.145 1046.935 3069.425 1188.985 ;
      RECT 3068.585 1048.035 3068.865 1189.225 ;
      RECT 3068.025 1048.035 3068.305 1189.465 ;
      RECT 3067.465 1048.035 3067.745 1189.705 ;
      RECT 3066.905 1048.035 3067.185 1189.945 ;
      RECT 3066.345 1048.035 3066.625 1190.185 ;
      RECT 3065.785 1048.035 3066.065 1190.425 ;
      RECT 3065.225 1048.035 3065.505 1190.665 ;
      RECT 3064.665 1048.035 3064.945 1190.665 ;
      RECT 3064.105 1048.035 3064.385 1190.425 ;
      RECT 3063.545 1048.035 3063.825 1190.185 ;
      RECT 3062.985 1048.035 3063.265 1189.945 ;
      RECT 3062.425 1048.035 3062.705 1189.7 ;
      RECT 3061.865 1048.035 3062.145 1189.46 ;
      RECT 3061.305 1048.035 3061.585 1189.22 ;
      RECT 3060.745 1046.935 3061.025 1188.98 ;
      RECT 3060.185 1048.035 3060.465 1188.74 ;
      RECT 3046.745 1046.935 3047.025 1186.22 ;
      RECT 3046.185 1048.035 3046.465 1185.98 ;
      RECT 3045.625 1048.035 3045.905 1185.74 ;
      RECT 3045.065 1048.035 3045.345 1185.5 ;
      RECT 3044.505 1046.935 3044.785 1185.26 ;
      RECT 3043.945 1048.035 3044.225 1185.02 ;
      RECT 3043.385 1046.935 3043.665 1184.78 ;
      RECT 3042.825 1048.035 3043.105 1184.54 ;
      RECT 3042.265 1046.935 3042.545 1184.3 ;
      RECT 3041.705 1048.035 3041.985 1184.06 ;
      RECT 3041.145 1048.035 3041.425 1183.82 ;
      RECT 3040.585 1048.035 3040.865 1183.58 ;
      RECT 3040.025 1048.035 3040.305 1183.34 ;
      RECT 3039.465 1048.035 3039.745 1183.1 ;
      RECT 3038.905 1048.035 3039.185 1182.86 ;
      RECT 3038.345 1048.035 3038.625 1182.62 ;
      RECT 3037.785 1048.035 3038.065 1182.38 ;
      RECT 3037.225 1048.035 3037.505 1182.14 ;
      RECT 3036.665 1048.035 3036.945 1181.9 ;
      RECT 3036.105 1048.035 3036.385 1181.66 ;
      RECT 3035.545 1048.035 3035.825 1181.42 ;
      RECT 3034.985 1046.935 3035.265 1181.18 ;
      RECT 3034.425 1048.035 3034.705 1180.94 ;
      RECT 3033.865 1046.935 3034.145 1180.7 ;
      RECT 2994.105 1048.035 2994.385 1191.17 ;
      RECT 2993.545 1046.935 2993.825 1191.41 ;
      RECT 2992.985 1048.035 2993.265 1191.65 ;
      RECT 2992.425 1048.035 2992.705 1191.89 ;
      RECT 2991.865 1048.035 2992.145 1192.13 ;
      RECT 2991.305 1048.035 2991.585 1192.37 ;
      RECT 2990.745 1048.035 2991.025 1192.61 ;
      RECT 2990.185 1048.035 2990.465 1192.855 ;
      RECT 2989.625 1048.035 2989.905 1193.095 ;
      RECT 2989.065 1048.035 2989.345 1193.335 ;
      RECT 2988.505 1046.935 2988.785 1193.575 ;
      RECT 2987.945 1048.035 2988.225 1193.815 ;
      RECT 2987.385 1046.935 2987.665 1194.055 ;
      RECT 2986.825 1048.035 2987.105 1194.295 ;
      RECT 2986.265 1048.035 2986.545 1194.535 ;
      RECT 2985.705 1048.035 2985.985 1194.775 ;
      RECT 2985.145 1048.035 2985.425 1195.015 ;
      RECT 2984.585 1048.035 2984.865 1195.255 ;
      RECT 2984.025 1048.035 2984.305 1195.495 ;
      RECT 2983.465 1048.035 2983.745 1195.735 ;
      RECT 2982.905 1048.035 2983.185 1195.975 ;
      RECT 2982.345 1048.035 2982.625 1196.215 ;
      RECT 2981.785 1048.035 2982.065 1196.455 ;
      RECT 2981.225 1048.035 2981.505 1196.695 ;
      RECT 2972.265 1048.035 2972.545 1192.28 ;
      RECT 2971.705 1048.035 2971.985 1192.04 ;
      RECT 2971.145 1048.035 2971.425 1191.8 ;
      RECT 2970.585 1046.935 2970.865 1191.56 ;
      RECT 2970.025 1048.035 2970.305 1191.32 ;
      RECT 2969.465 1046.935 2969.745 1191.08 ;
      RECT 2968.905 1048.035 2969.185 1190.84 ;
      RECT 2968.345 1048.035 2968.625 1190.6 ;
      RECT 2967.785 1048.035 2968.065 1190.36 ;
      RECT 2967.225 1046.935 2967.505 1190.12 ;
      RECT 2966.665 1048.035 2966.945 1189.88 ;
      RECT 2966.105 1046.935 2966.385 1189.64 ;
      RECT 2965.545 1048.035 2965.825 1189.4 ;
      RECT 2964.985 1046.935 2965.265 1189.16 ;
      RECT 2962.465 1048.035 2962.745 1181.56 ;
      RECT 2961.905 1048.035 2962.185 1181.32 ;
      RECT 2961.345 1048.035 2961.625 1181.08 ;
      RECT 2960.785 1048.035 2961.065 1180.84 ;
      RECT 2960.225 1048.035 2960.505 1180.6 ;
      RECT 2959.665 1048.035 2959.945 1180.36 ;
      RECT 2959.105 1048.035 2959.385 1180.12 ;
      RECT 2933.065 1048.035 2933.345 1193.995 ;
      RECT 2932.505 1048.035 2932.785 1194.235 ;
      RECT 2931.945 1048.035 2932.225 1194.475 ;
      RECT 2931.385 1048.035 2931.665 1194.715 ;
      RECT 2930.825 1048.035 2931.105 1194.955 ;
      RECT 2930.265 1046.935 2930.545 1194.955 ;
      RECT 2929.705 1048.035 2929.985 1194.715 ;
      RECT 2929.145 1046.935 2929.425 1194.47 ;
      RECT 2928.585 1048.035 2928.865 1194.23 ;
      RECT 2928.025 1046.935 2928.305 1193.99 ;
      RECT 2927.465 1048.035 2927.745 1193.75 ;
      RECT 2926.905 1048.035 2927.185 1193.51 ;
      RECT 2926.345 1048.035 2926.625 1193.27 ;
      RECT 2925.785 1048.035 2926.065 1193.03 ;
      RECT 2925.225 1048.035 2925.505 1192.79 ;
      RECT 2924.665 1048.035 2924.945 1192.55 ;
      RECT 2924.105 1048.035 2924.385 1192.31 ;
      RECT 2923.545 1048.035 2923.825 1192.07 ;
      RECT 2922.985 1046.935 2923.265 1191.83 ;
      RECT 2922.425 1048.035 2922.705 1191.59 ;
      RECT 2921.865 1046.935 2922.145 1191.35 ;
      RECT 2921.305 1048.035 2921.585 1191.11 ;
      RECT 2920.745 1048.035 2921.025 1190.87 ;
      RECT 2920.185 1048.035 2920.465 1190.63 ;
      RECT 2906.745 1048.035 2907.025 1194.03 ;
      RECT 2906.185 1048.035 2906.465 1194.27 ;
      RECT 2905.625 1048.035 2905.905 1194.515 ;
      RECT 2905.065 1048.035 2905.345 1194.755 ;
      RECT 2904.505 1048.035 2904.785 1194.995 ;
      RECT 2903.945 1048.035 2904.225 1194.995 ;
      RECT 2903.385 1048.035 2903.665 1194.755 ;
      RECT 2902.825 1048.035 2903.105 1194.515 ;
      RECT 2902.265 1048.035 2902.545 1187.5 ;
      RECT 2901.705 1048.035 2901.985 1187.26 ;
      RECT 2901.145 1048.035 2901.425 1187.02 ;
      RECT 2900.585 1046.935 2900.865 1186.78 ;
      RECT 2900.025 1048.035 2900.305 1186.54 ;
      RECT 2899.465 1046.935 2899.745 1186.3 ;
      RECT 2898.905 1048.035 2899.185 1186.06 ;
      RECT 2898.345 1048.035 2898.625 1185.82 ;
      RECT 2897.785 1048.035 2898.065 1185.58 ;
      RECT 2897.225 1046.935 2897.505 1185.34 ;
      RECT 2896.665 1048.035 2896.945 1185.1 ;
      RECT 2896.105 1046.935 2896.385 1184.86 ;
      RECT 2895.545 1048.035 2895.825 1184.62 ;
      RECT 2894.985 1046.935 2895.265 1184.38 ;
      RECT 2894.425 1048.035 2894.705 1184.14 ;
      RECT 2893.865 1048.035 2894.145 1183.9 ;
      RECT 2853.545 1048.035 2853.825 1192.795 ;
      RECT 2852.985 1048.035 2853.265 1193.035 ;
      RECT 2852.425 1048.035 2852.705 1193.28 ;
      RECT 2851.865 1048.035 2852.145 1193.52 ;
      RECT 2851.305 1048.035 2851.585 1193.76 ;
      RECT 2850.745 1048.035 2851.025 1194 ;
      RECT 2850.185 1048.035 2850.465 1194.24 ;
      RECT 2849.625 1048.035 2849.905 1194.48 ;
      RECT 2849.065 1048.035 2849.345 1194.72 ;
      RECT 2848.505 1048.035 2848.785 1194.96 ;
      RECT 2847.945 1046.935 2848.225 1195.2 ;
      RECT 2847.385 1048.035 2847.665 1195.44 ;
      RECT 2846.825 1046.935 2847.105 1195.68 ;
      RECT 2846.265 1048.035 2846.545 1195.92 ;
      RECT 2845.705 1046.935 2845.985 1196.16 ;
      RECT 2845.145 1048.035 2845.425 1196.16 ;
      RECT 2844.585 1048.035 2844.865 1195.92 ;
      RECT 2844.025 1048.035 2844.305 1195.68 ;
      RECT 2843.465 1048.035 2843.745 1195.44 ;
      RECT 2842.905 1048.035 2843.185 1195.2 ;
      RECT 2842.345 1048.035 2842.625 1194.96 ;
      RECT 2841.785 1048.035 2842.065 1194.72 ;
      RECT 2841.225 1048.035 2841.505 1194.48 ;
      RECT 2832.265 1046.935 2832.545 1194.51 ;
      RECT 2831.705 1048.035 2831.985 1194.75 ;
      RECT 2831.145 1046.935 2831.425 1194.99 ;
      RECT 2830.585 1048.035 2830.865 1195.205 ;
      RECT 2830.025 1048.035 2830.305 1194.78 ;
      RECT 2829.465 1048.035 2829.745 1194.54 ;
      RECT 2828.905 1048.035 2829.185 1194.3 ;
      RECT 2828.345 1048.035 2828.625 1194.06 ;
      RECT 2827.785 1048.035 2828.065 1193.82 ;
      RECT 2827.225 1048.035 2827.505 1193.58 ;
      RECT 2826.665 1048.035 2826.945 1193.34 ;
      RECT 2826.105 1048.035 2826.385 1193.1 ;
      RECT 2825.545 1048.035 2825.825 1192.86 ;
      RECT 2824.985 1048.035 2825.265 1192.62 ;
      RECT 2822.465 1048.035 2822.745 1191.795 ;
      RECT 2821.905 1048.035 2822.185 1191.555 ;
      RECT 2821.345 1048.035 2821.625 1191.315 ;
      RECT 2820.785 1046.935 2821.065 1191.075 ;
      RECT 2820.225 1048.035 2820.505 1190.835 ;
      RECT 2819.665 1046.935 2819.945 1190.595 ;
      RECT 2819.105 1048.035 2819.385 1190.355 ;
      RECT 2818.545 1048.035 2818.825 1190.115 ;
      RECT 2791.945 1048.035 2792.225 1201.16 ;
      RECT 2791.385 1046.935 2791.665 1201.4 ;
      RECT 2790.825 1048.035 2791.105 1201.64 ;
      RECT 2790.265 1046.935 2790.545 1201.885 ;
      RECT 2789.705 1048.035 2789.985 1202.125 ;
      RECT 2789.145 1046.935 2789.425 1202.365 ;
      RECT 2788.585 1048.035 2788.865 1202.605 ;
      RECT 2788.025 1048.035 2788.305 1202.845 ;
      RECT 2787.465 1048.035 2787.745 1188.465 ;
      RECT 2786.905 1048.035 2787.185 1188.225 ;
      RECT 2786.345 1048.035 2786.625 1187.985 ;
      RECT 2785.785 1048.035 2786.065 1187.745 ;
      RECT 2785.225 1048.035 2785.505 1187.505 ;
      RECT 2784.665 1048.035 2784.945 1187.265 ;
      RECT 2784.105 1048.035 2784.385 1187.025 ;
      RECT 2783.545 1048.035 2783.825 1186.785 ;
      RECT 2782.985 1048.035 2783.265 1186.545 ;
      RECT 2782.425 1048.035 2782.705 1186.305 ;
      RECT 2781.865 1046.935 2782.145 1186.065 ;
      RECT 2781.305 1048.035 2781.585 1185.825 ;
      RECT 2780.745 1046.935 2781.025 1185.585 ;
      RECT 2780.185 1048.035 2780.465 1185.345 ;
      RECT 2766.185 1046.935 2766.465 1191.465 ;
      RECT 2765.625 1048.035 2765.905 1191.225 ;
      RECT 2765.065 1048.035 2765.345 1190.985 ;
      RECT 2764.505 1048.035 2764.785 1190.745 ;
      RECT 2763.945 1048.035 2764.225 1190.505 ;
      RECT 2763.385 1048.035 2763.665 1190.265 ;
      RECT 2762.825 1048.035 2763.105 1190.025 ;
      RECT 2762.265 1048.035 2762.545 1189.785 ;
      RECT 2761.705 1048.035 2761.985 1189.545 ;
      RECT 2761.145 1046.935 2761.425 1189.305 ;
      RECT 2760.585 1048.035 2760.865 1189.065 ;
      RECT 2760.025 1046.935 2760.305 1188.825 ;
      RECT 2759.465 1048.035 2759.745 1188.585 ;
      RECT 2758.905 1048.035 2759.185 1188.345 ;
      RECT 2758.345 1048.035 2758.625 1188.105 ;
      RECT 2757.785 1048.035 2758.065 1187.865 ;
      RECT 2757.225 1048.035 2757.505 1187.625 ;
      RECT 2756.665 1048.035 2756.945 1187.385 ;
      RECT 2756.105 1048.035 2756.385 1187.145 ;
      RECT 2755.545 1048.035 2755.825 1186.905 ;
      RECT 2754.985 1048.035 2755.265 1186.665 ;
      RECT 2754.425 1048.035 2754.705 1186.425 ;
      RECT 2753.865 1048.035 2754.145 1186.185 ;
      RECT 2714.665 1048.035 2714.945 1193.09 ;
      RECT 2714.105 1048.035 2714.385 1193.33 ;
      RECT 2713.545 1048.035 2713.825 1193.57 ;
      RECT 2712.985 1046.935 2713.265 1193.81 ;
      RECT 2712.425 1048.035 2712.705 1194.05 ;
      RECT 2711.865 1046.935 2712.145 1194.29 ;
      RECT 2711.305 1048.035 2711.585 1194.53 ;
      RECT 2710.745 1048.035 2711.025 1194.77 ;
      RECT 2710.185 1048.035 2710.465 1195.01 ;
      RECT 2709.625 1046.935 2709.905 1195.25 ;
      RECT 2709.065 1048.035 2709.345 1195.49 ;
      RECT 2708.505 1046.935 2708.785 1195.73 ;
      RECT 2707.945 1048.035 2708.225 1195.97 ;
      RECT 2707.385 1046.935 2707.665 1196.21 ;
      RECT 2706.825 1048.035 2707.105 1196.45 ;
      RECT 2706.265 1048.035 2706.545 1196.69 ;
      RECT 2705.705 1048.035 2705.985 1196.69 ;
      RECT 2705.145 1048.035 2705.425 1196.45 ;
      RECT 2704.585 1048.035 2704.865 1196.21 ;
      RECT 2704.025 1048.035 2704.305 1195.97 ;
      RECT 2703.465 1048.035 2703.745 1195.73 ;
      RECT 2702.905 1048.035 2703.185 1195.49 ;
      RECT 2702.345 1048.035 2702.625 1195.25 ;
      RECT 2701.785 1048.035 2702.065 1195.01 ;
      RECT 2701.225 1048.035 2701.505 1194.77 ;
      RECT 2692.265 1048.035 2692.545 1194.285 ;
      RECT 2691.705 1046.935 2691.985 1194.045 ;
      RECT 2691.145 1048.035 2691.425 1193.805 ;
      RECT 2690.585 1046.935 2690.865 1193.565 ;
      RECT 2690.025 1048.035 2690.305 1193.325 ;
      RECT 2689.465 1046.935 2689.745 1193.085 ;
      RECT 2688.905 1048.035 2689.185 1192.845 ;
      RECT 2688.345 1048.035 2688.625 1192.605 ;
      RECT 2687.785 1048.035 2688.065 1192.365 ;
      RECT 2687.225 1048.035 2687.505 1192.125 ;
      RECT 2686.665 1048.035 2686.945 1191.885 ;
      RECT 2686.105 1048.035 2686.385 1191.645 ;
      RECT 2685.545 1048.035 2685.825 1191.405 ;
      RECT 2684.985 1048.035 2685.265 1191.165 ;
      RECT 2682.465 1046.935 2682.745 1192.885 ;
      RECT 2681.905 1048.035 2682.185 1192.645 ;
      RECT 2681.345 1046.935 2681.625 1192.405 ;
      RECT 2680.785 1048.035 2681.065 1192.165 ;
      RECT 2680.225 1048.035 2680.505 1191.925 ;
      RECT 2679.665 1048.035 2679.945 1191.685 ;
      RECT 2679.105 1048.035 2679.385 1191.445 ;
      RECT 2678.545 1048.035 2678.825 1191.205 ;
      RECT 2652.505 1048.035 2652.785 1188.855 ;
      RECT 2651.945 1048.035 2652.225 1189.095 ;
      RECT 2651.385 1048.035 2651.665 1189.335 ;
      RECT 2650.825 1048.035 2651.105 1189.58 ;
      RECT 2650.265 1048.035 2650.545 1189.82 ;
      RECT 2649.705 1048.035 2649.985 1190.06 ;
      RECT 2649.145 1048.035 2649.425 1190.06 ;
      RECT 2648.585 1048.035 2648.865 1189.82 ;
      RECT 2648.025 1048.035 2648.305 1189.58 ;
      RECT 2647.465 1046.935 2647.745 1189.34 ;
      RECT 2646.905 1048.035 2647.185 1189.1 ;
      RECT 2646.345 1046.935 2646.625 1188.86 ;
      RECT 2645.785 1048.035 2646.065 1188.62 ;
      RECT 2645.225 1048.035 2645.505 1188.38 ;
      RECT 2644.665 1048.035 2644.945 1188.14 ;
      RECT 2644.105 1046.935 2644.385 1187.9 ;
      RECT 2643.545 1048.035 2643.825 1187.66 ;
      RECT 2642.985 1046.935 2643.265 1187.42 ;
      RECT 2642.425 1048.035 2642.705 1187.18 ;
      RECT 2641.865 1046.935 2642.145 1186.94 ;
      RECT 2641.305 1048.035 2641.585 1186.7 ;
      RECT 2640.745 1048.035 2641.025 1186.46 ;
      RECT 2640.185 1048.035 2640.465 1186.22 ;
      RECT 2639.625 1048.035 2639.905 1185.98 ;
      RECT 2626.185 1048.035 2626.465 1191.78 ;
      RECT 2625.625 1048.035 2625.905 1191.54 ;
      RECT 2625.065 1048.035 2625.345 1191.3 ;
      RECT 2624.505 1048.035 2624.785 1191.06 ;
      RECT 2623.945 1048.035 2624.225 1190.82 ;
      RECT 2623.385 1048.035 2623.665 1190.58 ;
      RECT 2622.825 1048.035 2623.105 1190.34 ;
      RECT 2622.265 1048.035 2622.545 1190.1 ;
      RECT 2621.705 1046.935 2621.985 1189.86 ;
      RECT 2621.145 1048.035 2621.425 1189.62 ;
      RECT 2620.585 1046.935 2620.865 1189.3 ;
      RECT 2620.025 1048.035 2620.305 1189.14 ;
      RECT 2619.465 1046.935 2619.745 1188.9 ;
      RECT 2618.905 1048.035 2619.185 1188.66 ;
      RECT 2618.345 1048.035 2618.625 1188.42 ;
      RECT 2617.785 1048.035 2618.065 1188.18 ;
      RECT 2617.225 1048.035 2617.505 1187.94 ;
      RECT 2616.665 1048.035 2616.945 1187.7 ;
      RECT 2616.105 1048.035 2616.385 1187.46 ;
      RECT 2615.545 1048.035 2615.825 1187.22 ;
      RECT 2614.985 1048.035 2615.265 1186.98 ;
      RECT 2614.425 1046.935 2614.705 1186.74 ;
      RECT 2613.865 1048.035 2614.145 1186.5 ;
      RECT 2613.305 1046.935 2613.585 1186.26 ;
      RECT 2574.105 1048.035 2574.385 1191.87 ;
      RECT 2573.545 1048.035 2573.825 1192.11 ;
      RECT 2572.985 1048.035 2573.265 1192.35 ;
      RECT 2572.425 1048.035 2572.705 1192.59 ;
      RECT 2571.865 1048.035 2572.145 1192.83 ;
      RECT 2571.305 1048.035 2571.585 1193.07 ;
      RECT 2570.745 1048.035 2571.025 1193.31 ;
      RECT 2570.185 1048.035 2570.465 1193.55 ;
      RECT 2569.625 1048.035 2569.905 1193.79 ;
      RECT 2569.065 1048.035 2569.345 1194.03 ;
      RECT 2568.505 1048.035 2568.785 1194.27 ;
      RECT 2567.945 1048.035 2568.225 1194.51 ;
      RECT 2567.385 1048.035 2567.665 1194.75 ;
      RECT 2566.825 1048.035 2567.105 1194.75 ;
      RECT 2566.265 1046.935 2566.545 1194.51 ;
      RECT 2565.705 1048.035 2565.985 1194.27 ;
      RECT 2565.145 1046.935 2565.425 1194.03 ;
      RECT 2564.585 1048.035 2564.865 1193.79 ;
      RECT 2564.025 1048.035 2564.305 1193.55 ;
      RECT 2563.465 1048.035 2563.745 1193.31 ;
      RECT 2562.905 1046.935 2563.185 1193.045 ;
      RECT 2562.345 1048.035 2562.625 1192.805 ;
      RECT 2561.785 1046.935 2562.065 1192.565 ;
      RECT 2561.225 1048.035 2561.505 1192.325 ;
      RECT 2552.265 1046.935 2552.545 1186.16 ;
      RECT 2551.705 1048.035 2551.985 1186.4 ;
      RECT 2551.145 1048.035 2551.425 1186.64 ;
      RECT 2550.585 1048.035 2550.865 1186.64 ;
      RECT 2550.025 1048.035 2550.305 1186.4 ;
      RECT 2549.465 1048.035 2549.745 1186.16 ;
      RECT 2548.905 1048.035 2549.185 1185.92 ;
      RECT 2548.345 1048.035 2548.625 1185.68 ;
      RECT 2547.785 1048.035 2548.065 1185.44 ;
      RECT 2547.225 1048.035 2547.505 1185.2 ;
      RECT 2546.665 1048.035 2546.945 1184.96 ;
      RECT 2546.105 1048.035 2546.385 1184.72 ;
      RECT 2545.545 1048.035 2545.825 1184.48 ;
      RECT 2544.985 1046.935 2545.265 1184.24 ;
      RECT 2542.465 1048.035 2542.745 1185.96 ;
      RECT 2541.905 1046.935 2542.185 1185.72 ;
      RECT 2541.345 1048.035 2541.625 1185.48 ;
      RECT 2540.785 1046.935 2541.065 1185.24 ;
      RECT 2540.225 1048.035 2540.505 1185 ;
      RECT 2539.665 1048.035 2539.945 1184.76 ;
      RECT 2539.105 1048.035 2539.385 1184.52 ;
      RECT 2513.065 1048.035 2513.345 1187.305 ;
      RECT 2512.505 1048.035 2512.785 1187.545 ;
      RECT 2511.945 1048.035 2512.225 1187.785 ;
      RECT 2511.385 1048.035 2511.665 1188.025 ;
      RECT 2510.825 1048.035 2511.105 1188.265 ;
      RECT 2510.265 1046.935 2510.545 1188.505 ;
      RECT 2509.705 1048.035 2509.985 1188.745 ;
      RECT 2509.145 1046.935 2509.425 1188.985 ;
      RECT 2508.585 1048.035 2508.865 1189.225 ;
      RECT 2508.025 1048.035 2508.305 1189.465 ;
      RECT 2507.465 1048.035 2507.745 1189.705 ;
      RECT 2506.905 1048.035 2507.185 1189.945 ;
      RECT 2506.345 1048.035 2506.625 1190.185 ;
      RECT 2505.785 1048.035 2506.065 1190.425 ;
      RECT 2505.225 1048.035 2505.505 1190.665 ;
      RECT 2504.665 1048.035 2504.945 1190.665 ;
      RECT 2504.105 1048.035 2504.385 1190.425 ;
      RECT 2503.545 1048.035 2503.825 1190.185 ;
      RECT 2502.985 1048.035 2503.265 1189.945 ;
      RECT 2502.425 1048.035 2502.705 1189.7 ;
      RECT 2501.865 1048.035 2502.145 1189.46 ;
      RECT 2501.305 1048.035 2501.585 1189.22 ;
      RECT 2500.745 1046.935 2501.025 1188.98 ;
      RECT 2500.185 1048.035 2500.465 1188.74 ;
      RECT 2486.745 1046.935 2487.025 1186.22 ;
      RECT 2486.185 1048.035 2486.465 1185.98 ;
      RECT 2485.625 1048.035 2485.905 1185.74 ;
      RECT 2485.065 1048.035 2485.345 1185.5 ;
      RECT 2484.505 1046.935 2484.785 1185.26 ;
      RECT 2483.945 1048.035 2484.225 1185.02 ;
      RECT 2483.385 1046.935 2483.665 1184.78 ;
      RECT 2482.825 1048.035 2483.105 1184.54 ;
      RECT 2482.265 1046.935 2482.545 1184.3 ;
      RECT 2481.705 1048.035 2481.985 1184.06 ;
      RECT 2481.145 1048.035 2481.425 1183.82 ;
      RECT 2480.585 1048.035 2480.865 1183.58 ;
      RECT 2480.025 1048.035 2480.305 1183.34 ;
      RECT 2479.465 1048.035 2479.745 1183.1 ;
      RECT 2478.905 1048.035 2479.185 1182.86 ;
      RECT 2478.345 1048.035 2478.625 1182.62 ;
      RECT 2477.785 1048.035 2478.065 1182.38 ;
      RECT 2477.225 1048.035 2477.505 1182.14 ;
      RECT 2476.665 1048.035 2476.945 1181.9 ;
      RECT 2476.105 1048.035 2476.385 1181.66 ;
      RECT 2475.545 1048.035 2475.825 1181.42 ;
      RECT 2474.985 1046.935 2475.265 1181.18 ;
      RECT 2474.425 1048.035 2474.705 1180.94 ;
      RECT 2473.865 1046.935 2474.145 1180.7 ;
      RECT 2434.105 1048.035 2434.385 1191.17 ;
      RECT 2433.545 1046.935 2433.825 1191.41 ;
      RECT 2432.985 1048.035 2433.265 1191.65 ;
      RECT 2432.425 1048.035 2432.705 1191.89 ;
      RECT 2431.865 1048.035 2432.145 1192.13 ;
      RECT 2431.305 1048.035 2431.585 1192.37 ;
      RECT 2430.745 1048.035 2431.025 1192.61 ;
      RECT 2430.185 1048.035 2430.465 1192.855 ;
      RECT 2429.625 1048.035 2429.905 1193.095 ;
      RECT 2429.065 1048.035 2429.345 1193.335 ;
      RECT 2428.505 1046.935 2428.785 1193.575 ;
      RECT 2427.945 1048.035 2428.225 1193.815 ;
      RECT 2427.385 1046.935 2427.665 1194.055 ;
      RECT 2426.825 1048.035 2427.105 1194.295 ;
      RECT 2426.265 1048.035 2426.545 1194.535 ;
      RECT 2425.705 1048.035 2425.985 1194.775 ;
      RECT 2425.145 1048.035 2425.425 1195.015 ;
      RECT 2424.585 1048.035 2424.865 1195.255 ;
      RECT 2424.025 1048.035 2424.305 1195.495 ;
      RECT 2423.465 1048.035 2423.745 1195.735 ;
      RECT 2422.905 1048.035 2423.185 1195.975 ;
      RECT 2422.345 1048.035 2422.625 1196.215 ;
      RECT 2421.785 1048.035 2422.065 1196.455 ;
      RECT 2421.225 1048.035 2421.505 1196.695 ;
      RECT 2412.265 1048.035 2412.545 1192.28 ;
      RECT 2411.705 1048.035 2411.985 1192.04 ;
      RECT 2411.145 1048.035 2411.425 1191.8 ;
      RECT 2410.585 1046.935 2410.865 1191.56 ;
      RECT 2410.025 1048.035 2410.305 1191.32 ;
      RECT 2409.465 1046.935 2409.745 1191.08 ;
      RECT 2408.905 1048.035 2409.185 1190.84 ;
      RECT 2408.345 1048.035 2408.625 1190.6 ;
      RECT 2407.785 1048.035 2408.065 1190.36 ;
      RECT 2407.225 1046.935 2407.505 1190.12 ;
      RECT 2406.665 1048.035 2406.945 1189.88 ;
      RECT 2406.105 1046.935 2406.385 1189.64 ;
      RECT 2405.545 1048.035 2405.825 1189.4 ;
      RECT 2404.985 1046.935 2405.265 1189.16 ;
      RECT 2402.465 1048.035 2402.745 1181.56 ;
      RECT 2401.905 1048.035 2402.185 1181.32 ;
      RECT 2401.345 1048.035 2401.625 1181.08 ;
      RECT 2400.785 1048.035 2401.065 1180.84 ;
      RECT 2400.225 1048.035 2400.505 1180.6 ;
      RECT 2399.665 1048.035 2399.945 1180.36 ;
      RECT 2399.105 1048.035 2399.385 1180.12 ;
      RECT 2373.065 1048.035 2373.345 1193.995 ;
      RECT 2372.505 1048.035 2372.785 1194.235 ;
      RECT 2371.945 1048.035 2372.225 1194.475 ;
      RECT 2371.385 1048.035 2371.665 1194.715 ;
      RECT 2370.825 1048.035 2371.105 1194.955 ;
      RECT 2370.265 1046.935 2370.545 1194.955 ;
      RECT 2369.705 1048.035 2369.985 1194.715 ;
      RECT 2369.145 1046.935 2369.425 1194.47 ;
      RECT 2368.585 1048.035 2368.865 1194.23 ;
      RECT 2368.025 1046.935 2368.305 1193.99 ;
      RECT 2367.465 1048.035 2367.745 1193.75 ;
      RECT 2366.905 1048.035 2367.185 1193.51 ;
      RECT 2366.345 1048.035 2366.625 1193.27 ;
      RECT 2365.785 1048.035 2366.065 1193.03 ;
      RECT 2365.225 1048.035 2365.505 1192.79 ;
      RECT 2364.665 1048.035 2364.945 1192.55 ;
      RECT 2364.105 1048.035 2364.385 1192.31 ;
      RECT 2363.545 1048.035 2363.825 1192.07 ;
      RECT 2362.985 1046.935 2363.265 1191.83 ;
      RECT 2362.425 1048.035 2362.705 1191.59 ;
      RECT 2361.865 1046.935 2362.145 1191.35 ;
      RECT 2361.305 1048.035 2361.585 1191.11 ;
      RECT 2360.745 1048.035 2361.025 1190.87 ;
      RECT 2360.185 1048.035 2360.465 1190.63 ;
      RECT 2346.745 1048.035 2347.025 1194.03 ;
      RECT 2346.185 1048.035 2346.465 1194.27 ;
      RECT 2345.625 1048.035 2345.905 1194.515 ;
      RECT 2345.065 1048.035 2345.345 1194.755 ;
      RECT 2344.505 1048.035 2344.785 1194.995 ;
      RECT 2343.945 1048.035 2344.225 1194.995 ;
      RECT 2343.385 1048.035 2343.665 1194.755 ;
      RECT 2342.825 1048.035 2343.105 1194.515 ;
      RECT 2342.265 1048.035 2342.545 1187.5 ;
      RECT 2341.705 1048.035 2341.985 1187.26 ;
      RECT 2341.145 1048.035 2341.425 1187.02 ;
      RECT 2340.585 1046.935 2340.865 1186.78 ;
      RECT 2340.025 1048.035 2340.305 1186.54 ;
      RECT 2339.465 1046.935 2339.745 1186.3 ;
      RECT 2338.905 1048.035 2339.185 1186.06 ;
      RECT 2338.345 1048.035 2338.625 1185.82 ;
      RECT 2337.785 1048.035 2338.065 1185.58 ;
      RECT 2337.225 1046.935 2337.505 1185.34 ;
      RECT 2336.665 1048.035 2336.945 1185.1 ;
      RECT 2336.105 1046.935 2336.385 1184.86 ;
      RECT 2335.545 1048.035 2335.825 1184.62 ;
      RECT 2334.985 1046.935 2335.265 1184.38 ;
      RECT 2334.425 1048.035 2334.705 1184.14 ;
      RECT 2333.865 1048.035 2334.145 1183.9 ;
      RECT 2293.545 1048.035 2293.825 1192.795 ;
      RECT 2292.985 1048.035 2293.265 1193.035 ;
      RECT 2292.425 1048.035 2292.705 1193.28 ;
      RECT 2291.865 1048.035 2292.145 1193.52 ;
      RECT 2291.305 1048.035 2291.585 1193.76 ;
      RECT 2290.745 1048.035 2291.025 1194 ;
      RECT 2290.185 1048.035 2290.465 1194.24 ;
      RECT 2289.625 1048.035 2289.905 1194.48 ;
      RECT 2289.065 1048.035 2289.345 1194.72 ;
      RECT 2288.505 1048.035 2288.785 1194.96 ;
      RECT 2287.945 1046.935 2288.225 1195.2 ;
      RECT 2287.385 1048.035 2287.665 1195.44 ;
      RECT 2286.825 1046.935 2287.105 1195.68 ;
      RECT 2286.265 1048.035 2286.545 1195.92 ;
      RECT 2285.705 1046.935 2285.985 1196.16 ;
      RECT 2285.145 1048.035 2285.425 1196.16 ;
      RECT 2284.585 1048.035 2284.865 1195.92 ;
      RECT 2284.025 1048.035 2284.305 1195.68 ;
      RECT 2283.465 1048.035 2283.745 1195.44 ;
      RECT 2282.905 1048.035 2283.185 1195.2 ;
      RECT 2282.345 1048.035 2282.625 1194.96 ;
      RECT 2281.785 1048.035 2282.065 1194.72 ;
      RECT 2281.225 1048.035 2281.505 1194.48 ;
      RECT 2272.265 1046.935 2272.545 1194.51 ;
      RECT 2271.705 1048.035 2271.985 1194.75 ;
      RECT 2271.145 1046.935 2271.425 1194.99 ;
      RECT 2270.585 1048.035 2270.865 1195.205 ;
      RECT 2270.025 1048.035 2270.305 1194.78 ;
      RECT 2269.465 1048.035 2269.745 1194.54 ;
      RECT 2268.905 1048.035 2269.185 1194.3 ;
      RECT 2268.345 1048.035 2268.625 1194.06 ;
      RECT 2267.785 1048.035 2268.065 1193.82 ;
      RECT 2267.225 1048.035 2267.505 1193.58 ;
      RECT 2266.665 1048.035 2266.945 1193.34 ;
      RECT 2266.105 1048.035 2266.385 1193.1 ;
      RECT 2265.545 1048.035 2265.825 1192.86 ;
      RECT 2264.985 1048.035 2265.265 1192.62 ;
      RECT 2262.465 1048.035 2262.745 1191.795 ;
      RECT 2261.905 1048.035 2262.185 1191.555 ;
      RECT 2261.345 1048.035 2261.625 1191.315 ;
      RECT 2260.785 1046.935 2261.065 1191.075 ;
      RECT 2260.225 1048.035 2260.505 1190.835 ;
      RECT 2259.665 1046.935 2259.945 1190.595 ;
      RECT 2259.105 1048.035 2259.385 1190.355 ;
      RECT 2258.545 1048.035 2258.825 1190.115 ;
      RECT 2231.945 1048.035 2232.225 1201.16 ;
      RECT 2231.385 1046.935 2231.665 1201.4 ;
      RECT 2230.825 1048.035 2231.105 1201.64 ;
      RECT 2230.265 1046.935 2230.545 1201.885 ;
      RECT 2229.705 1048.035 2229.985 1202.125 ;
      RECT 2229.145 1046.935 2229.425 1202.365 ;
      RECT 2228.585 1048.035 2228.865 1202.605 ;
      RECT 2228.025 1048.035 2228.305 1202.845 ;
      RECT 2227.465 1048.035 2227.745 1188.465 ;
      RECT 2226.905 1048.035 2227.185 1188.225 ;
      RECT 2226.345 1048.035 2226.625 1187.985 ;
      RECT 2225.785 1048.035 2226.065 1187.745 ;
      RECT 2225.225 1048.035 2225.505 1187.505 ;
      RECT 2224.665 1048.035 2224.945 1187.265 ;
      RECT 2224.105 1048.035 2224.385 1187.025 ;
      RECT 2223.545 1048.035 2223.825 1186.785 ;
      RECT 2222.985 1048.035 2223.265 1186.545 ;
      RECT 2222.425 1048.035 2222.705 1186.305 ;
      RECT 2221.865 1046.935 2222.145 1186.065 ;
      RECT 2221.305 1048.035 2221.585 1185.825 ;
      RECT 2220.745 1046.935 2221.025 1185.585 ;
      RECT 2220.185 1048.035 2220.465 1185.345 ;
      RECT 2206.185 1046.935 2206.465 1191.465 ;
      RECT 2205.625 1048.035 2205.905 1191.225 ;
      RECT 2205.065 1048.035 2205.345 1190.985 ;
      RECT 2204.505 1048.035 2204.785 1190.745 ;
      RECT 2203.945 1048.035 2204.225 1190.505 ;
      RECT 2203.385 1048.035 2203.665 1190.265 ;
      RECT 2202.825 1048.035 2203.105 1190.025 ;
      RECT 2202.265 1048.035 2202.545 1189.785 ;
      RECT 2201.705 1048.035 2201.985 1189.545 ;
      RECT 2201.145 1046.935 2201.425 1189.305 ;
      RECT 2200.585 1048.035 2200.865 1189.065 ;
      RECT 2200.025 1046.935 2200.305 1188.825 ;
      RECT 2199.465 1048.035 2199.745 1188.585 ;
      RECT 2198.905 1048.035 2199.185 1188.345 ;
      RECT 2198.345 1048.035 2198.625 1188.105 ;
      RECT 2197.785 1048.035 2198.065 1187.865 ;
      RECT 2197.225 1048.035 2197.505 1187.625 ;
      RECT 2196.665 1048.035 2196.945 1187.385 ;
      RECT 2196.105 1048.035 2196.385 1187.145 ;
      RECT 2195.545 1048.035 2195.825 1186.905 ;
      RECT 2194.985 1048.035 2195.265 1186.665 ;
      RECT 2194.425 1048.035 2194.705 1186.425 ;
      RECT 2193.865 1048.035 2194.145 1186.185 ;
      RECT 2154.665 1048.035 2154.945 1193.09 ;
      RECT 2154.105 1048.035 2154.385 1193.33 ;
      RECT 2153.545 1048.035 2153.825 1193.57 ;
      RECT 2152.985 1046.935 2153.265 1193.81 ;
      RECT 2152.425 1048.035 2152.705 1194.05 ;
      RECT 2151.865 1046.935 2152.145 1194.29 ;
      RECT 2151.305 1048.035 2151.585 1194.53 ;
      RECT 2150.745 1048.035 2151.025 1194.77 ;
      RECT 2150.185 1048.035 2150.465 1195.01 ;
      RECT 2149.625 1046.935 2149.905 1195.25 ;
      RECT 2149.065 1048.035 2149.345 1195.49 ;
      RECT 2148.505 1046.935 2148.785 1195.73 ;
      RECT 2147.945 1048.035 2148.225 1195.97 ;
      RECT 2147.385 1046.935 2147.665 1196.21 ;
      RECT 2146.825 1048.035 2147.105 1196.45 ;
      RECT 2146.265 1048.035 2146.545 1196.69 ;
      RECT 2145.705 1048.035 2145.985 1196.69 ;
      RECT 2145.145 1048.035 2145.425 1196.45 ;
      RECT 2144.585 1048.035 2144.865 1196.21 ;
      RECT 2144.025 1048.035 2144.305 1195.97 ;
      RECT 2143.465 1048.035 2143.745 1195.73 ;
      RECT 2142.905 1048.035 2143.185 1195.49 ;
      RECT 2142.345 1048.035 2142.625 1195.25 ;
      RECT 2141.785 1048.035 2142.065 1195.01 ;
      RECT 2141.225 1048.035 2141.505 1194.77 ;
      RECT 2132.265 1048.035 2132.545 1194.285 ;
      RECT 2131.705 1046.935 2131.985 1194.045 ;
      RECT 2131.145 1048.035 2131.425 1193.805 ;
      RECT 2130.585 1046.935 2130.865 1193.565 ;
      RECT 2130.025 1048.035 2130.305 1193.325 ;
      RECT 2129.465 1046.935 2129.745 1193.085 ;
      RECT 2128.905 1048.035 2129.185 1192.845 ;
      RECT 2128.345 1048.035 2128.625 1192.605 ;
      RECT 2127.785 1048.035 2128.065 1192.365 ;
      RECT 2127.225 1048.035 2127.505 1192.125 ;
      RECT 2126.665 1048.035 2126.945 1191.885 ;
      RECT 2126.105 1048.035 2126.385 1191.645 ;
      RECT 2125.545 1048.035 2125.825 1191.405 ;
      RECT 2124.985 1048.035 2125.265 1191.165 ;
      RECT 2122.465 1046.935 2122.745 1192.885 ;
      RECT 2121.905 1048.035 2122.185 1192.645 ;
      RECT 2121.345 1046.935 2121.625 1192.405 ;
      RECT 2120.785 1048.035 2121.065 1192.165 ;
      RECT 2120.225 1048.035 2120.505 1191.925 ;
      RECT 2119.665 1048.035 2119.945 1191.685 ;
      RECT 2119.105 1048.035 2119.385 1191.445 ;
      RECT 2118.545 1048.035 2118.825 1191.205 ;
      RECT 2092.505 1048.035 2092.785 1188.855 ;
      RECT 2091.945 1048.035 2092.225 1189.095 ;
      RECT 2091.385 1048.035 2091.665 1189.335 ;
      RECT 2090.825 1048.035 2091.105 1189.58 ;
      RECT 2090.265 1048.035 2090.545 1189.82 ;
      RECT 2089.705 1048.035 2089.985 1190.06 ;
      RECT 2089.145 1048.035 2089.425 1190.06 ;
      RECT 2088.585 1048.035 2088.865 1189.82 ;
      RECT 2088.025 1048.035 2088.305 1189.58 ;
      RECT 2087.465 1046.935 2087.745 1189.34 ;
      RECT 2086.905 1048.035 2087.185 1189.1 ;
      RECT 2086.345 1046.935 2086.625 1188.86 ;
      RECT 2085.785 1048.035 2086.065 1188.62 ;
      RECT 2085.225 1048.035 2085.505 1188.38 ;
      RECT 2084.665 1048.035 2084.945 1188.14 ;
      RECT 2084.105 1046.935 2084.385 1187.9 ;
      RECT 2083.545 1048.035 2083.825 1187.66 ;
      RECT 2082.985 1046.935 2083.265 1187.42 ;
      RECT 2082.425 1048.035 2082.705 1187.18 ;
      RECT 2081.865 1046.935 2082.145 1186.94 ;
      RECT 2081.305 1048.035 2081.585 1186.7 ;
      RECT 2080.745 1048.035 2081.025 1186.46 ;
      RECT 2080.185 1048.035 2080.465 1186.22 ;
      RECT 2079.625 1048.035 2079.905 1185.98 ;
      RECT 2066.185 1048.035 2066.465 1191.78 ;
      RECT 2065.625 1048.035 2065.905 1191.54 ;
      RECT 2065.065 1048.035 2065.345 1191.3 ;
      RECT 2064.505 1048.035 2064.785 1191.06 ;
      RECT 2063.945 1048.035 2064.225 1190.82 ;
      RECT 2063.385 1048.035 2063.665 1190.58 ;
      RECT 2062.825 1048.035 2063.105 1190.34 ;
      RECT 2062.265 1048.035 2062.545 1190.1 ;
      RECT 2061.705 1046.935 2061.985 1189.86 ;
      RECT 2061.145 1048.035 2061.425 1189.62 ;
      RECT 2060.585 1046.935 2060.865 1189.3 ;
      RECT 2060.025 1048.035 2060.305 1189.14 ;
      RECT 2059.465 1046.935 2059.745 1188.9 ;
      RECT 2058.905 1048.035 2059.185 1188.66 ;
      RECT 2058.345 1048.035 2058.625 1188.42 ;
      RECT 2057.785 1048.035 2058.065 1188.18 ;
      RECT 2057.225 1048.035 2057.505 1187.94 ;
      RECT 2056.665 1048.035 2056.945 1187.7 ;
      RECT 2056.105 1048.035 2056.385 1187.46 ;
      RECT 2055.545 1048.035 2055.825 1187.22 ;
      RECT 2054.985 1048.035 2055.265 1186.98 ;
      RECT 2054.425 1046.935 2054.705 1186.74 ;
      RECT 2053.865 1048.035 2054.145 1186.5 ;
      RECT 2053.305 1046.935 2053.585 1186.26 ;
      RECT 2014.105 1048.035 2014.385 1191.87 ;
      RECT 2013.545 1048.035 2013.825 1192.11 ;
      RECT 2012.985 1048.035 2013.265 1192.35 ;
      RECT 2012.425 1048.035 2012.705 1192.59 ;
      RECT 2011.865 1048.035 2012.145 1192.83 ;
      RECT 2011.305 1048.035 2011.585 1193.07 ;
      RECT 2010.745 1048.035 2011.025 1193.31 ;
      RECT 2010.185 1048.035 2010.465 1193.55 ;
      RECT 2009.625 1048.035 2009.905 1193.79 ;
      RECT 2009.065 1048.035 2009.345 1194.03 ;
      RECT 2008.505 1048.035 2008.785 1194.27 ;
      RECT 2007.945 1048.035 2008.225 1194.51 ;
      RECT 2007.385 1048.035 2007.665 1194.75 ;
      RECT 2006.825 1048.035 2007.105 1194.75 ;
      RECT 2006.265 1046.935 2006.545 1194.51 ;
      RECT 2005.705 1048.035 2005.985 1194.27 ;
      RECT 2005.145 1046.935 2005.425 1194.03 ;
      RECT 2004.585 1048.035 2004.865 1193.79 ;
      RECT 2004.025 1048.035 2004.305 1193.55 ;
      RECT 2003.465 1048.035 2003.745 1193.31 ;
      RECT 2002.905 1046.935 2003.185 1193.045 ;
      RECT 2002.345 1048.035 2002.625 1192.805 ;
      RECT 2001.785 1046.935 2002.065 1192.565 ;
      RECT 2001.225 1048.035 2001.505 1192.325 ;
      RECT 1992.265 1046.935 1992.545 1186.16 ;
      RECT 1991.705 1048.035 1991.985 1186.4 ;
      RECT 1991.145 1048.035 1991.425 1186.64 ;
      RECT 1990.585 1048.035 1990.865 1186.64 ;
      RECT 1990.025 1048.035 1990.305 1186.4 ;
      RECT 1989.465 1048.035 1989.745 1186.16 ;
      RECT 1988.905 1048.035 1989.185 1185.92 ;
      RECT 1988.345 1048.035 1988.625 1185.68 ;
      RECT 1987.785 1048.035 1988.065 1185.44 ;
      RECT 1987.225 1048.035 1987.505 1185.2 ;
      RECT 1986.665 1048.035 1986.945 1184.96 ;
      RECT 1986.105 1048.035 1986.385 1184.72 ;
      RECT 1985.545 1048.035 1985.825 1184.48 ;
      RECT 1984.985 1046.935 1985.265 1184.24 ;
      RECT 1982.465 1048.035 1982.745 1185.96 ;
      RECT 1981.905 1046.935 1982.185 1185.72 ;
      RECT 1981.345 1048.035 1981.625 1185.48 ;
      RECT 1980.785 1046.935 1981.065 1185.24 ;
      RECT 1980.225 1048.035 1980.505 1185 ;
      RECT 1979.665 1048.035 1979.945 1184.76 ;
      RECT 1979.105 1048.035 1979.385 1184.52 ;
      RECT 1953.065 1048.035 1953.345 1187.305 ;
      RECT 1952.505 1048.035 1952.785 1187.545 ;
      RECT 1951.945 1048.035 1952.225 1187.785 ;
      RECT 1951.385 1048.035 1951.665 1188.025 ;
      RECT 1950.825 1048.035 1951.105 1188.265 ;
      RECT 1950.265 1046.935 1950.545 1188.505 ;
      RECT 1949.705 1048.035 1949.985 1188.745 ;
      RECT 1949.145 1046.935 1949.425 1188.985 ;
      RECT 1948.585 1048.035 1948.865 1189.225 ;
      RECT 1948.025 1048.035 1948.305 1189.465 ;
      RECT 1947.465 1048.035 1947.745 1189.705 ;
      RECT 1946.905 1048.035 1947.185 1189.945 ;
      RECT 1946.345 1048.035 1946.625 1190.185 ;
      RECT 1945.785 1048.035 1946.065 1190.425 ;
      RECT 1945.225 1048.035 1945.505 1190.665 ;
      RECT 1944.665 1048.035 1944.945 1190.665 ;
      RECT 1944.105 1048.035 1944.385 1190.425 ;
      RECT 1943.545 1048.035 1943.825 1190.185 ;
      RECT 1942.985 1048.035 1943.265 1189.945 ;
      RECT 1942.425 1048.035 1942.705 1189.7 ;
      RECT 1941.865 1048.035 1942.145 1189.46 ;
      RECT 1941.305 1048.035 1941.585 1189.22 ;
      RECT 1940.745 1046.935 1941.025 1188.98 ;
      RECT 1940.185 1048.035 1940.465 1188.74 ;
      RECT 1926.745 1046.935 1927.025 1186.22 ;
      RECT 1926.185 1048.035 1926.465 1185.98 ;
      RECT 1925.625 1048.035 1925.905 1185.74 ;
      RECT 1925.065 1048.035 1925.345 1185.5 ;
      RECT 1924.505 1046.935 1924.785 1185.26 ;
      RECT 1923.945 1048.035 1924.225 1185.02 ;
      RECT 1923.385 1046.935 1923.665 1184.78 ;
      RECT 1922.825 1048.035 1923.105 1184.54 ;
      RECT 1922.265 1046.935 1922.545 1184.3 ;
      RECT 1921.705 1048.035 1921.985 1184.06 ;
      RECT 1921.145 1048.035 1921.425 1183.82 ;
      RECT 1920.585 1048.035 1920.865 1183.58 ;
      RECT 1920.025 1048.035 1920.305 1183.34 ;
      RECT 1919.465 1048.035 1919.745 1183.1 ;
      RECT 1918.905 1048.035 1919.185 1182.86 ;
      RECT 1918.345 1048.035 1918.625 1182.62 ;
      RECT 1917.785 1048.035 1918.065 1182.38 ;
      RECT 1917.225 1048.035 1917.505 1182.14 ;
      RECT 1916.665 1048.035 1916.945 1181.9 ;
      RECT 1916.105 1048.035 1916.385 1181.66 ;
      RECT 1915.545 1048.035 1915.825 1181.42 ;
      RECT 1914.985 1046.935 1915.265 1181.18 ;
      RECT 1914.425 1048.035 1914.705 1180.94 ;
      RECT 1913.865 1046.935 1914.145 1180.7 ;
      RECT 1874.105 1048.035 1874.385 1191.17 ;
      RECT 1873.545 1046.935 1873.825 1191.41 ;
      RECT 1872.985 1048.035 1873.265 1191.65 ;
      RECT 1872.425 1048.035 1872.705 1191.89 ;
      RECT 1871.865 1048.035 1872.145 1192.13 ;
      RECT 1871.305 1048.035 1871.585 1192.37 ;
      RECT 1870.745 1048.035 1871.025 1192.61 ;
      RECT 1870.185 1048.035 1870.465 1192.855 ;
      RECT 1869.625 1048.035 1869.905 1193.095 ;
      RECT 1869.065 1048.035 1869.345 1193.335 ;
      RECT 1868.505 1046.935 1868.785 1193.575 ;
      RECT 1867.945 1048.035 1868.225 1193.815 ;
      RECT 1867.385 1046.935 1867.665 1194.055 ;
      RECT 1866.825 1048.035 1867.105 1194.295 ;
      RECT 1866.265 1048.035 1866.545 1194.535 ;
      RECT 1865.705 1048.035 1865.985 1194.775 ;
      RECT 1865.145 1048.035 1865.425 1195.015 ;
      RECT 1864.585 1048.035 1864.865 1195.255 ;
      RECT 1864.025 1048.035 1864.305 1195.495 ;
      RECT 1863.465 1048.035 1863.745 1195.735 ;
      RECT 1862.905 1048.035 1863.185 1195.975 ;
      RECT 1862.345 1048.035 1862.625 1196.215 ;
      RECT 1861.785 1048.035 1862.065 1196.455 ;
      RECT 1861.225 1048.035 1861.505 1196.695 ;
      RECT 1852.265 1048.035 1852.545 1192.28 ;
      RECT 1851.705 1048.035 1851.985 1192.04 ;
      RECT 1851.145 1048.035 1851.425 1191.8 ;
      RECT 1850.585 1046.935 1850.865 1191.56 ;
      RECT 1850.025 1048.035 1850.305 1191.32 ;
      RECT 1849.465 1046.935 1849.745 1191.08 ;
      RECT 1848.905 1048.035 1849.185 1190.84 ;
      RECT 1848.345 1048.035 1848.625 1190.6 ;
      RECT 1847.785 1048.035 1848.065 1190.36 ;
      RECT 1847.225 1046.935 1847.505 1190.12 ;
      RECT 1846.665 1048.035 1846.945 1189.88 ;
      RECT 1846.105 1046.935 1846.385 1189.64 ;
      RECT 1845.545 1048.035 1845.825 1189.4 ;
      RECT 1844.985 1046.935 1845.265 1189.16 ;
      RECT 1842.465 1048.035 1842.745 1181.56 ;
      RECT 1841.905 1048.035 1842.185 1181.32 ;
      RECT 1841.345 1048.035 1841.625 1181.08 ;
      RECT 1840.785 1048.035 1841.065 1180.84 ;
      RECT 1840.225 1048.035 1840.505 1180.6 ;
      RECT 1839.665 1048.035 1839.945 1180.36 ;
      RECT 1839.105 1048.035 1839.385 1180.12 ;
      RECT 1813.065 1048.035 1813.345 1193.995 ;
      RECT 1812.505 1048.035 1812.785 1194.235 ;
      RECT 1811.945 1048.035 1812.225 1194.475 ;
      RECT 1811.385 1048.035 1811.665 1194.715 ;
      RECT 1810.825 1048.035 1811.105 1194.955 ;
      RECT 1810.265 1046.935 1810.545 1194.955 ;
      RECT 1809.705 1048.035 1809.985 1194.715 ;
      RECT 1809.145 1046.935 1809.425 1194.47 ;
      RECT 1808.585 1048.035 1808.865 1194.23 ;
      RECT 1808.025 1046.935 1808.305 1193.99 ;
      RECT 1807.465 1048.035 1807.745 1193.75 ;
      RECT 1806.905 1048.035 1807.185 1193.51 ;
      RECT 1806.345 1048.035 1806.625 1193.27 ;
      RECT 1805.785 1048.035 1806.065 1193.03 ;
      RECT 1805.225 1048.035 1805.505 1192.79 ;
      RECT 1804.665 1048.035 1804.945 1192.55 ;
      RECT 1804.105 1048.035 1804.385 1192.31 ;
      RECT 1803.545 1048.035 1803.825 1192.07 ;
      RECT 1802.985 1046.935 1803.265 1191.83 ;
      RECT 1802.425 1048.035 1802.705 1191.59 ;
      RECT 1801.865 1046.935 1802.145 1191.35 ;
      RECT 1801.305 1048.035 1801.585 1191.11 ;
      RECT 1800.745 1048.035 1801.025 1190.87 ;
      RECT 1800.185 1048.035 1800.465 1190.63 ;
      RECT 1786.745 1048.035 1787.025 1194.03 ;
      RECT 1786.185 1048.035 1786.465 1194.27 ;
      RECT 1785.625 1048.035 1785.905 1194.515 ;
      RECT 1785.065 1048.035 1785.345 1194.755 ;
      RECT 1784.505 1048.035 1784.785 1194.995 ;
      RECT 1783.945 1048.035 1784.225 1194.995 ;
      RECT 1783.385 1048.035 1783.665 1194.755 ;
      RECT 1782.825 1048.035 1783.105 1194.515 ;
      RECT 1782.265 1048.035 1782.545 1187.5 ;
      RECT 1781.705 1048.035 1781.985 1187.26 ;
      RECT 1781.145 1048.035 1781.425 1187.02 ;
      RECT 1780.585 1046.935 1780.865 1186.78 ;
      RECT 1780.025 1048.035 1780.305 1186.54 ;
      RECT 1779.465 1046.935 1779.745 1186.3 ;
      RECT 1778.905 1048.035 1779.185 1186.06 ;
      RECT 1778.345 1048.035 1778.625 1185.82 ;
      RECT 1777.785 1048.035 1778.065 1185.58 ;
      RECT 1777.225 1046.935 1777.505 1185.34 ;
      RECT 1776.665 1048.035 1776.945 1185.1 ;
      RECT 1776.105 1046.935 1776.385 1184.86 ;
      RECT 1775.545 1048.035 1775.825 1184.62 ;
      RECT 1774.985 1046.935 1775.265 1184.38 ;
      RECT 1774.425 1048.035 1774.705 1184.14 ;
      RECT 1773.865 1048.035 1774.145 1183.9 ;
      RECT 1733.545 1048.035 1733.825 1192.795 ;
      RECT 1732.985 1048.035 1733.265 1193.035 ;
      RECT 1732.425 1048.035 1732.705 1193.28 ;
      RECT 1731.865 1048.035 1732.145 1193.52 ;
      RECT 1731.305 1048.035 1731.585 1193.76 ;
      RECT 1730.745 1048.035 1731.025 1194 ;
      RECT 1730.185 1048.035 1730.465 1194.24 ;
      RECT 1729.625 1048.035 1729.905 1194.48 ;
      RECT 1729.065 1048.035 1729.345 1194.72 ;
      RECT 1728.505 1048.035 1728.785 1194.96 ;
      RECT 1727.945 1046.935 1728.225 1195.2 ;
      RECT 1727.385 1048.035 1727.665 1195.44 ;
      RECT 1726.825 1046.935 1727.105 1195.68 ;
      RECT 1726.265 1048.035 1726.545 1195.92 ;
      RECT 1725.705 1046.935 1725.985 1196.16 ;
      RECT 1725.145 1048.035 1725.425 1196.16 ;
      RECT 1724.585 1048.035 1724.865 1195.92 ;
      RECT 1724.025 1048.035 1724.305 1195.68 ;
      RECT 1723.465 1048.035 1723.745 1195.44 ;
      RECT 1722.905 1048.035 1723.185 1195.2 ;
      RECT 1722.345 1048.035 1722.625 1194.96 ;
      RECT 1721.785 1048.035 1722.065 1194.72 ;
      RECT 1721.225 1048.035 1721.505 1194.48 ;
      RECT 1712.265 1046.935 1712.545 1194.51 ;
      RECT 1711.705 1048.035 1711.985 1194.75 ;
      RECT 1711.145 1046.935 1711.425 1194.99 ;
      RECT 1710.585 1048.035 1710.865 1195.205 ;
      RECT 1710.025 1048.035 1710.305 1194.78 ;
      RECT 1709.465 1048.035 1709.745 1194.54 ;
      RECT 1708.905 1048.035 1709.185 1194.3 ;
      RECT 1708.345 1048.035 1708.625 1194.06 ;
      RECT 1707.785 1048.035 1708.065 1193.82 ;
      RECT 1707.225 1048.035 1707.505 1193.58 ;
      RECT 1706.665 1048.035 1706.945 1193.34 ;
      RECT 1706.105 1048.035 1706.385 1193.1 ;
      RECT 1705.545 1048.035 1705.825 1192.86 ;
      RECT 1704.985 1048.035 1705.265 1192.62 ;
      RECT 1702.465 1048.035 1702.745 1191.795 ;
      RECT 1701.905 1048.035 1702.185 1191.555 ;
      RECT 1701.345 1048.035 1701.625 1191.315 ;
      RECT 1700.785 1046.935 1701.065 1191.075 ;
      RECT 1700.225 1048.035 1700.505 1190.835 ;
      RECT 1699.665 1046.935 1699.945 1190.595 ;
      RECT 1699.105 1048.035 1699.385 1190.355 ;
      RECT 1698.545 1048.035 1698.825 1190.115 ;
      RECT 1671.945 1048.035 1672.225 1201.16 ;
      RECT 1671.385 1046.935 1671.665 1201.4 ;
      RECT 1670.825 1048.035 1671.105 1201.64 ;
      RECT 1670.265 1046.935 1670.545 1201.885 ;
      RECT 1669.705 1048.035 1669.985 1202.125 ;
      RECT 1669.145 1046.935 1669.425 1202.365 ;
      RECT 1668.585 1048.035 1668.865 1202.605 ;
      RECT 1668.025 1048.035 1668.305 1202.845 ;
      RECT 1667.465 1048.035 1667.745 1188.465 ;
      RECT 1666.905 1048.035 1667.185 1188.225 ;
      RECT 1666.345 1048.035 1666.625 1187.985 ;
      RECT 1665.785 1048.035 1666.065 1187.745 ;
      RECT 1665.225 1048.035 1665.505 1187.505 ;
      RECT 1664.665 1048.035 1664.945 1187.265 ;
      RECT 1664.105 1048.035 1664.385 1187.025 ;
      RECT 1663.545 1048.035 1663.825 1186.785 ;
      RECT 1662.985 1048.035 1663.265 1186.545 ;
      RECT 1662.425 1048.035 1662.705 1186.305 ;
      RECT 1661.865 1046.935 1662.145 1186.065 ;
      RECT 1661.305 1048.035 1661.585 1185.825 ;
      RECT 1660.745 1046.935 1661.025 1185.585 ;
      RECT 1660.185 1048.035 1660.465 1185.345 ;
      RECT 1646.185 1046.935 1646.465 1191.465 ;
      RECT 1645.625 1048.035 1645.905 1191.225 ;
      RECT 1645.065 1048.035 1645.345 1190.985 ;
      RECT 1644.505 1048.035 1644.785 1190.745 ;
      RECT 1643.945 1048.035 1644.225 1190.505 ;
      RECT 1643.385 1048.035 1643.665 1190.265 ;
      RECT 1642.825 1048.035 1643.105 1190.025 ;
      RECT 1642.265 1048.035 1642.545 1189.785 ;
      RECT 1641.705 1048.035 1641.985 1189.545 ;
      RECT 1641.145 1046.935 1641.425 1189.305 ;
      RECT 1640.585 1048.035 1640.865 1189.065 ;
      RECT 1640.025 1046.935 1640.305 1188.825 ;
      RECT 1639.465 1048.035 1639.745 1188.585 ;
      RECT 1638.905 1048.035 1639.185 1188.345 ;
      RECT 1638.345 1048.035 1638.625 1188.105 ;
      RECT 1637.785 1048.035 1638.065 1187.865 ;
      RECT 1637.225 1048.035 1637.505 1187.625 ;
      RECT 1636.665 1048.035 1636.945 1187.385 ;
      RECT 1636.105 1048.035 1636.385 1187.145 ;
      RECT 1635.545 1048.035 1635.825 1186.905 ;
      RECT 1634.985 1048.035 1635.265 1186.665 ;
      RECT 1634.425 1048.035 1634.705 1186.425 ;
      RECT 1633.865 1048.035 1634.145 1186.185 ;
      RECT 1594.665 1048.035 1594.945 1193.09 ;
      RECT 1594.105 1048.035 1594.385 1193.33 ;
      RECT 1593.545 1048.035 1593.825 1193.57 ;
      RECT 1592.985 1046.935 1593.265 1193.81 ;
      RECT 1592.425 1048.035 1592.705 1194.05 ;
      RECT 1591.865 1046.935 1592.145 1194.29 ;
      RECT 1591.305 1048.035 1591.585 1194.53 ;
      RECT 1590.745 1048.035 1591.025 1194.77 ;
      RECT 1590.185 1048.035 1590.465 1195.01 ;
      RECT 1589.625 1046.935 1589.905 1195.25 ;
      RECT 1589.065 1048.035 1589.345 1195.49 ;
      RECT 1588.505 1046.935 1588.785 1195.73 ;
      RECT 1587.945 1048.035 1588.225 1195.97 ;
      RECT 1587.385 1046.935 1587.665 1196.21 ;
      RECT 1586.825 1048.035 1587.105 1196.45 ;
      RECT 1586.265 1048.035 1586.545 1196.69 ;
      RECT 1585.705 1048.035 1585.985 1196.69 ;
      RECT 1585.145 1048.035 1585.425 1196.45 ;
      RECT 1584.585 1048.035 1584.865 1196.21 ;
      RECT 1584.025 1048.035 1584.305 1195.97 ;
      RECT 1583.465 1048.035 1583.745 1195.73 ;
      RECT 1582.905 1048.035 1583.185 1195.49 ;
      RECT 1582.345 1048.035 1582.625 1195.25 ;
      RECT 1581.785 1048.035 1582.065 1195.01 ;
      RECT 1581.225 1048.035 1581.505 1194.77 ;
      RECT 1572.265 1048.035 1572.545 1194.285 ;
      RECT 1571.705 1046.935 1571.985 1194.045 ;
      RECT 1571.145 1048.035 1571.425 1193.805 ;
      RECT 1570.585 1046.935 1570.865 1193.565 ;
      RECT 1570.025 1048.035 1570.305 1193.325 ;
      RECT 1569.465 1046.935 1569.745 1193.085 ;
      RECT 1568.905 1048.035 1569.185 1192.845 ;
      RECT 1568.345 1048.035 1568.625 1192.605 ;
      RECT 1567.785 1048.035 1568.065 1192.365 ;
      RECT 1567.225 1048.035 1567.505 1192.125 ;
      RECT 1566.665 1048.035 1566.945 1191.885 ;
      RECT 1566.105 1048.035 1566.385 1191.645 ;
      RECT 1565.545 1048.035 1565.825 1191.405 ;
      RECT 1564.985 1048.035 1565.265 1191.165 ;
      RECT 1562.465 1046.935 1562.745 1192.885 ;
      RECT 1561.905 1048.035 1562.185 1192.645 ;
      RECT 1561.345 1046.935 1561.625 1192.405 ;
      RECT 1560.785 1048.035 1561.065 1192.165 ;
      RECT 1560.225 1048.035 1560.505 1191.925 ;
      RECT 1559.665 1048.035 1559.945 1191.685 ;
      RECT 1559.105 1048.035 1559.385 1191.445 ;
      RECT 1558.545 1048.035 1558.825 1191.205 ;
      RECT 1532.505 1048.035 1532.785 1188.855 ;
      RECT 1531.945 1048.035 1532.225 1189.095 ;
      RECT 1531.385 1048.035 1531.665 1189.335 ;
      RECT 1530.825 1048.035 1531.105 1189.58 ;
      RECT 1530.265 1048.035 1530.545 1189.82 ;
      RECT 1529.705 1048.035 1529.985 1190.06 ;
      RECT 1529.145 1048.035 1529.425 1190.06 ;
      RECT 1528.585 1048.035 1528.865 1189.82 ;
      RECT 1528.025 1048.035 1528.305 1189.58 ;
      RECT 1527.465 1046.935 1527.745 1189.34 ;
      RECT 1526.905 1048.035 1527.185 1189.1 ;
      RECT 1526.345 1046.935 1526.625 1188.86 ;
      RECT 1525.785 1048.035 1526.065 1188.62 ;
      RECT 1525.225 1048.035 1525.505 1188.38 ;
      RECT 1524.665 1048.035 1524.945 1188.14 ;
      RECT 1524.105 1046.935 1524.385 1187.9 ;
      RECT 1523.545 1048.035 1523.825 1187.66 ;
      RECT 1522.985 1046.935 1523.265 1187.42 ;
      RECT 1522.425 1048.035 1522.705 1187.18 ;
      RECT 1521.865 1046.935 1522.145 1186.94 ;
      RECT 1521.305 1048.035 1521.585 1186.7 ;
      RECT 1520.745 1048.035 1521.025 1186.46 ;
      RECT 1520.185 1048.035 1520.465 1186.22 ;
      RECT 1519.625 1048.035 1519.905 1185.98 ;
      RECT 1506.185 1048.035 1506.465 1191.78 ;
      RECT 1505.625 1048.035 1505.905 1191.54 ;
      RECT 1505.065 1048.035 1505.345 1191.3 ;
      RECT 1504.505 1048.035 1504.785 1191.06 ;
      RECT 1503.945 1048.035 1504.225 1190.82 ;
      RECT 1503.385 1048.035 1503.665 1190.58 ;
      RECT 1502.825 1048.035 1503.105 1190.34 ;
      RECT 1502.265 1048.035 1502.545 1190.1 ;
      RECT 1501.705 1046.935 1501.985 1189.86 ;
      RECT 1501.145 1048.035 1501.425 1189.62 ;
      RECT 1500.585 1046.935 1500.865 1189.3 ;
      RECT 1500.025 1048.035 1500.305 1189.14 ;
      RECT 1499.465 1046.935 1499.745 1188.9 ;
      RECT 1498.905 1048.035 1499.185 1188.66 ;
      RECT 1498.345 1048.035 1498.625 1188.42 ;
      RECT 1497.785 1048.035 1498.065 1188.18 ;
      RECT 1497.225 1048.035 1497.505 1187.94 ;
      RECT 1496.665 1048.035 1496.945 1187.7 ;
      RECT 1496.105 1048.035 1496.385 1187.46 ;
      RECT 1495.545 1048.035 1495.825 1187.22 ;
      RECT 1494.985 1048.035 1495.265 1186.98 ;
      RECT 1494.425 1046.935 1494.705 1186.74 ;
      RECT 1493.865 1048.035 1494.145 1186.5 ;
      RECT 1493.305 1046.935 1493.585 1186.26 ;
      RECT 1454.105 1048.035 1454.385 1191.87 ;
      RECT 1453.545 1048.035 1453.825 1192.11 ;
      RECT 1452.985 1048.035 1453.265 1192.35 ;
      RECT 1452.425 1048.035 1452.705 1192.59 ;
      RECT 1451.865 1048.035 1452.145 1192.83 ;
      RECT 1451.305 1048.035 1451.585 1193.07 ;
      RECT 1450.745 1048.035 1451.025 1193.31 ;
      RECT 1450.185 1048.035 1450.465 1193.55 ;
      RECT 1449.625 1048.035 1449.905 1193.79 ;
      RECT 1449.065 1048.035 1449.345 1194.03 ;
      RECT 1448.505 1048.035 1448.785 1194.27 ;
      RECT 1447.945 1048.035 1448.225 1194.51 ;
      RECT 1447.385 1048.035 1447.665 1194.75 ;
      RECT 1446.825 1048.035 1447.105 1194.75 ;
      RECT 1446.265 1046.935 1446.545 1194.51 ;
      RECT 1445.705 1048.035 1445.985 1194.27 ;
      RECT 1445.145 1046.935 1445.425 1194.03 ;
      RECT 1444.585 1048.035 1444.865 1193.79 ;
      RECT 1444.025 1048.035 1444.305 1193.55 ;
      RECT 1443.465 1048.035 1443.745 1193.31 ;
      RECT 1442.905 1046.935 1443.185 1193.045 ;
      RECT 1442.345 1048.035 1442.625 1192.805 ;
      RECT 1441.785 1046.935 1442.065 1192.565 ;
      RECT 1441.225 1048.035 1441.505 1192.325 ;
      RECT 1432.265 1046.935 1432.545 1186.16 ;
      RECT 1431.705 1048.035 1431.985 1186.4 ;
      RECT 1431.145 1048.035 1431.425 1186.64 ;
      RECT 1430.585 1048.035 1430.865 1186.64 ;
      RECT 1430.025 1048.035 1430.305 1186.4 ;
      RECT 1429.465 1048.035 1429.745 1186.16 ;
      RECT 1428.905 1048.035 1429.185 1185.92 ;
      RECT 1428.345 1048.035 1428.625 1185.68 ;
      RECT 1427.785 1048.035 1428.065 1185.44 ;
      RECT 1427.225 1048.035 1427.505 1185.2 ;
      RECT 1426.665 1048.035 1426.945 1184.96 ;
      RECT 1426.105 1048.035 1426.385 1184.72 ;
      RECT 1425.545 1048.035 1425.825 1184.48 ;
      RECT 1424.985 1046.935 1425.265 1184.24 ;
      RECT 1422.465 1048.035 1422.745 1185.96 ;
      RECT 1421.905 1046.935 1422.185 1185.72 ;
      RECT 1421.345 1048.035 1421.625 1185.48 ;
      RECT 1420.785 1046.935 1421.065 1185.24 ;
      RECT 1420.225 1048.035 1420.505 1185 ;
      RECT 1419.665 1048.035 1419.945 1184.76 ;
      RECT 1419.105 1048.035 1419.385 1184.52 ;
      RECT 1393.065 1048.035 1393.345 1187.305 ;
      RECT 1392.505 1048.035 1392.785 1187.545 ;
      RECT 1391.945 1048.035 1392.225 1187.785 ;
      RECT 1391.385 1048.035 1391.665 1188.025 ;
      RECT 1390.825 1048.035 1391.105 1188.265 ;
      RECT 1390.265 1046.935 1390.545 1188.505 ;
      RECT 1389.705 1048.035 1389.985 1188.745 ;
      RECT 1389.145 1046.935 1389.425 1188.985 ;
      RECT 1388.585 1048.035 1388.865 1189.225 ;
      RECT 1388.025 1048.035 1388.305 1189.465 ;
      RECT 1387.465 1048.035 1387.745 1189.705 ;
      RECT 1386.905 1048.035 1387.185 1189.945 ;
      RECT 1386.345 1048.035 1386.625 1190.185 ;
      RECT 1385.785 1048.035 1386.065 1190.425 ;
      RECT 1385.225 1048.035 1385.505 1190.665 ;
      RECT 1384.665 1048.035 1384.945 1190.665 ;
      RECT 1384.105 1048.035 1384.385 1190.425 ;
      RECT 1383.545 1048.035 1383.825 1190.185 ;
      RECT 1382.985 1048.035 1383.265 1189.945 ;
      RECT 1382.425 1048.035 1382.705 1189.7 ;
      RECT 1381.865 1048.035 1382.145 1189.46 ;
      RECT 1381.305 1048.035 1381.585 1189.22 ;
      RECT 1380.745 1046.935 1381.025 1188.98 ;
      RECT 1380.185 1048.035 1380.465 1188.74 ;
      RECT 1366.745 1046.935 1367.025 1186.22 ;
      RECT 1366.185 1048.035 1366.465 1185.98 ;
      RECT 1365.625 1048.035 1365.905 1185.74 ;
      RECT 1365.065 1048.035 1365.345 1185.5 ;
      RECT 1364.505 1046.935 1364.785 1185.26 ;
      RECT 1363.945 1048.035 1364.225 1185.02 ;
      RECT 1363.385 1046.935 1363.665 1184.78 ;
      RECT 1362.825 1048.035 1363.105 1184.54 ;
      RECT 1362.265 1046.935 1362.545 1184.3 ;
      RECT 1361.705 1048.035 1361.985 1184.06 ;
      RECT 1361.145 1048.035 1361.425 1183.82 ;
      RECT 1360.585 1048.035 1360.865 1183.58 ;
      RECT 1360.025 1048.035 1360.305 1183.34 ;
      RECT 1359.465 1048.035 1359.745 1183.1 ;
      RECT 1358.905 1048.035 1359.185 1182.86 ;
      RECT 1358.345 1048.035 1358.625 1182.62 ;
      RECT 1357.785 1048.035 1358.065 1182.38 ;
      RECT 1357.225 1048.035 1357.505 1182.14 ;
      RECT 1356.665 1048.035 1356.945 1181.9 ;
      RECT 1356.105 1048.035 1356.385 1181.66 ;
      RECT 1355.545 1048.035 1355.825 1181.42 ;
      RECT 1354.985 1046.935 1355.265 1181.18 ;
      RECT 1354.425 1048.035 1354.705 1180.94 ;
      RECT 1353.865 1046.935 1354.145 1180.7 ;
      RECT 1314.105 1048.035 1314.385 1191.17 ;
      RECT 1313.545 1046.935 1313.825 1191.41 ;
      RECT 1312.985 1048.035 1313.265 1191.65 ;
      RECT 1312.425 1048.035 1312.705 1191.89 ;
      RECT 1311.865 1048.035 1312.145 1192.13 ;
      RECT 1311.305 1048.035 1311.585 1192.37 ;
      RECT 1310.745 1048.035 1311.025 1192.61 ;
      RECT 1310.185 1048.035 1310.465 1192.855 ;
      RECT 1309.625 1048.035 1309.905 1193.095 ;
      RECT 1309.065 1048.035 1309.345 1193.335 ;
      RECT 1308.505 1046.935 1308.785 1193.575 ;
      RECT 1307.945 1048.035 1308.225 1193.815 ;
      RECT 1307.385 1046.935 1307.665 1194.055 ;
      RECT 1306.825 1048.035 1307.105 1194.295 ;
      RECT 1306.265 1048.035 1306.545 1194.535 ;
      RECT 1305.705 1048.035 1305.985 1194.775 ;
      RECT 1305.145 1048.035 1305.425 1195.015 ;
      RECT 1304.585 1048.035 1304.865 1195.255 ;
      RECT 1304.025 1048.035 1304.305 1195.495 ;
      RECT 1303.465 1048.035 1303.745 1195.735 ;
      RECT 1302.905 1048.035 1303.185 1195.975 ;
      RECT 1302.345 1048.035 1302.625 1196.215 ;
      RECT 1301.785 1048.035 1302.065 1196.455 ;
      RECT 1301.225 1048.035 1301.505 1196.695 ;
      RECT 1292.265 1048.035 1292.545 1192.28 ;
      RECT 1291.705 1048.035 1291.985 1192.04 ;
      RECT 1291.145 1048.035 1291.425 1191.8 ;
      RECT 1290.585 1046.935 1290.865 1191.56 ;
      RECT 1290.025 1048.035 1290.305 1191.32 ;
      RECT 1289.465 1046.935 1289.745 1191.08 ;
      RECT 1288.905 1048.035 1289.185 1190.84 ;
      RECT 1288.345 1048.035 1288.625 1190.6 ;
      RECT 1287.785 1048.035 1288.065 1190.36 ;
      RECT 1287.225 1046.935 1287.505 1190.12 ;
      RECT 1286.665 1048.035 1286.945 1189.88 ;
      RECT 1286.105 1046.935 1286.385 1189.64 ;
      RECT 1285.545 1048.035 1285.825 1189.4 ;
      RECT 1284.985 1046.935 1285.265 1189.16 ;
      RECT 1282.465 1048.035 1282.745 1181.56 ;
      RECT 1281.905 1048.035 1282.185 1181.32 ;
      RECT 1281.345 1048.035 1281.625 1181.08 ;
      RECT 1280.785 1048.035 1281.065 1180.84 ;
      RECT 1280.225 1048.035 1280.505 1180.6 ;
      RECT 1279.665 1048.035 1279.945 1180.36 ;
      RECT 1279.105 1048.035 1279.385 1180.12 ;
      RECT 1253.065 1048.035 1253.345 1193.995 ;
      RECT 1252.505 1048.035 1252.785 1194.235 ;
      RECT 1251.945 1048.035 1252.225 1194.475 ;
      RECT 1251.385 1048.035 1251.665 1194.715 ;
      RECT 1250.825 1048.035 1251.105 1194.955 ;
      RECT 1250.265 1046.935 1250.545 1194.955 ;
      RECT 1249.705 1048.035 1249.985 1194.715 ;
      RECT 1249.145 1046.935 1249.425 1194.47 ;
      RECT 1248.585 1048.035 1248.865 1194.23 ;
      RECT 1248.025 1046.935 1248.305 1193.99 ;
      RECT 1247.465 1048.035 1247.745 1193.75 ;
      RECT 1246.905 1048.035 1247.185 1193.51 ;
      RECT 1246.345 1048.035 1246.625 1193.27 ;
      RECT 1245.785 1048.035 1246.065 1193.03 ;
      RECT 1245.225 1048.035 1245.505 1192.79 ;
      RECT 1244.665 1048.035 1244.945 1192.55 ;
      RECT 1244.105 1048.035 1244.385 1192.31 ;
      RECT 1243.545 1048.035 1243.825 1192.07 ;
      RECT 1242.985 1046.935 1243.265 1191.83 ;
      RECT 1242.425 1048.035 1242.705 1191.59 ;
      RECT 1241.865 1046.935 1242.145 1191.35 ;
      RECT 1241.305 1048.035 1241.585 1191.11 ;
      RECT 1240.745 1048.035 1241.025 1190.87 ;
      RECT 1240.185 1048.035 1240.465 1190.63 ;
      RECT 1226.745 1048.035 1227.025 1194.03 ;
      RECT 1226.185 1048.035 1226.465 1194.27 ;
      RECT 1225.625 1048.035 1225.905 1194.515 ;
      RECT 1225.065 1048.035 1225.345 1194.755 ;
      RECT 1224.505 1048.035 1224.785 1194.995 ;
      RECT 1223.945 1048.035 1224.225 1194.995 ;
      RECT 1223.385 1048.035 1223.665 1194.755 ;
      RECT 1222.825 1048.035 1223.105 1194.515 ;
      RECT 1222.265 1048.035 1222.545 1187.5 ;
      RECT 1221.705 1048.035 1221.985 1187.26 ;
      RECT 1221.145 1048.035 1221.425 1187.02 ;
      RECT 1220.585 1046.935 1220.865 1186.78 ;
      RECT 1220.025 1048.035 1220.305 1186.54 ;
      RECT 1219.465 1046.935 1219.745 1186.3 ;
      RECT 1218.905 1048.035 1219.185 1186.06 ;
      RECT 1218.345 1048.035 1218.625 1185.82 ;
      RECT 1217.785 1048.035 1218.065 1185.58 ;
      RECT 1217.225 1046.935 1217.505 1185.34 ;
      RECT 1216.665 1048.035 1216.945 1185.1 ;
      RECT 1216.105 1046.935 1216.385 1184.86 ;
      RECT 1215.545 1048.035 1215.825 1184.62 ;
      RECT 1214.985 1046.935 1215.265 1184.38 ;
      RECT 1214.425 1048.035 1214.705 1184.14 ;
      RECT 1213.865 1048.035 1214.145 1183.9 ;
      RECT 1173.545 1048.035 1173.825 1192.795 ;
      RECT 1172.985 1048.035 1173.265 1193.035 ;
      RECT 1172.425 1048.035 1172.705 1193.28 ;
      RECT 1171.865 1048.035 1172.145 1193.52 ;
      RECT 1171.305 1048.035 1171.585 1193.76 ;
      RECT 1170.745 1048.035 1171.025 1194 ;
      RECT 1170.185 1048.035 1170.465 1194.24 ;
      RECT 1169.625 1048.035 1169.905 1194.48 ;
      RECT 1169.065 1048.035 1169.345 1194.72 ;
      RECT 1168.505 1048.035 1168.785 1194.96 ;
      RECT 1167.945 1046.935 1168.225 1195.2 ;
      RECT 1167.385 1048.035 1167.665 1195.44 ;
      RECT 1166.825 1046.935 1167.105 1195.68 ;
      RECT 1166.265 1048.035 1166.545 1195.92 ;
      RECT 1165.705 1046.935 1165.985 1196.16 ;
      RECT 1165.145 1048.035 1165.425 1196.16 ;
      RECT 1164.585 1048.035 1164.865 1195.92 ;
      RECT 1164.025 1048.035 1164.305 1195.68 ;
      RECT 1163.465 1048.035 1163.745 1195.44 ;
      RECT 1162.905 1048.035 1163.185 1195.2 ;
      RECT 1162.345 1048.035 1162.625 1194.96 ;
      RECT 1161.785 1048.035 1162.065 1194.72 ;
      RECT 1161.225 1048.035 1161.505 1194.48 ;
      RECT 1152.265 1046.935 1152.545 1194.51 ;
      RECT 1151.705 1048.035 1151.985 1194.75 ;
      RECT 1151.145 1046.935 1151.425 1194.99 ;
      RECT 1150.585 1048.035 1150.865 1195.205 ;
      RECT 1150.025 1048.035 1150.305 1194.78 ;
      RECT 1149.465 1048.035 1149.745 1194.54 ;
      RECT 1148.905 1048.035 1149.185 1194.3 ;
      RECT 1148.345 1048.035 1148.625 1194.06 ;
      RECT 1147.785 1048.035 1148.065 1193.82 ;
      RECT 1147.225 1048.035 1147.505 1193.58 ;
      RECT 1146.665 1048.035 1146.945 1193.34 ;
      RECT 1146.105 1048.035 1146.385 1193.1 ;
      RECT 1145.545 1048.035 1145.825 1192.86 ;
      RECT 1144.985 1048.035 1145.265 1192.62 ;
      RECT 1142.465 1048.035 1142.745 1191.795 ;
      RECT 1141.905 1048.035 1142.185 1191.555 ;
      RECT 1141.345 1048.035 1141.625 1191.315 ;
      RECT 1140.785 1046.935 1141.065 1191.075 ;
      RECT 1140.225 1048.035 1140.505 1190.835 ;
      RECT 1139.665 1046.935 1139.945 1190.595 ;
      RECT 1139.105 1048.035 1139.385 1190.355 ;
      RECT 1138.545 1048.035 1138.825 1190.115 ;
      RECT 1137.985 1048.035 1138.265 1154.13 ;
      RECT 990 9497.56 1010 9527.56 ;
      RECT 990 9529.56 1010 9559.56 ;
      RECT 990 9617.56 1010 9647.56 ;
      RECT 990 9649.56 1010 9679.56 ;
      RECT 990 9737.56 1010 9767.56 ;
      RECT 990 9769.56 1010 9799.56 ;
      RECT 990 9857.56 1010 9887.56 ;
      RECT 990 9889.56 1010 9919.56 ;
      RECT 992.1 1057.81 1001.84 1058.61 ;
      RECT 992.1 1087.58 1001.84 1088.38 ;
      RECT 992.1 1090.38 1001.84 1091.18 ;
      RECT 992.1 1116.79 1001.84 1117.59 ;
      RECT 992.1 1119.19 1001.84 1119.99 ;
      RECT 992.1 1121.59 1001.84 1122.39 ;
      RECT 992.1 1123.99 1001.84 1124.79 ;
      RECT 992.1 1126.39 1001.84 1127.19 ;
    LAYER M4 SPACING 0.28 ;
      RECT 14234.005 1047.855 19161.9 10000 ;
      RECT 19033.205 1046.435 19161.9 10000 ;
      RECT 19031.385 1046.935 19031.665 10000 ;
      RECT 19030.265 1046.935 19030.545 10000 ;
      RECT 19029.145 1046.935 19029.425 10000 ;
      RECT 19021.865 1046.935 19022.145 10000 ;
      RECT 19020.745 1046.935 19021.025 10000 ;
      RECT 19006.185 1046.935 19019.765 10000 ;
      RECT 19006.325 1046.435 19019.765 10000 ;
      RECT 19001.145 1046.935 19001.425 10000 ;
      RECT 19000.025 1046.935 19000.305 10000 ;
      RECT 18955.365 1046.435 18993.445 10000 ;
      RECT 18952.985 1046.935 18953.265 10000 ;
      RECT 18951.865 1046.935 18952.145 10000 ;
      RECT 18949.625 1046.935 18949.905 10000 ;
      RECT 18948.505 1046.935 18948.785 10000 ;
      RECT 18947.385 1046.935 18947.665 10000 ;
      RECT 18932.965 1046.435 18940.805 10000 ;
      RECT 18931.705 1046.935 18931.985 10000 ;
      RECT 18930.585 1046.935 18930.865 10000 ;
      RECT 18929.465 1046.935 18929.745 10000 ;
      RECT 18922.465 1046.935 18924.565 10000 ;
      RECT 18922.605 1046.435 18924.565 10000 ;
      RECT 18921.345 1046.935 18921.625 10000 ;
      RECT 18893.205 1046.435 18918.125 10000 ;
      RECT 18887.465 1046.935 18887.745 10000 ;
      RECT 18886.345 1046.935 18886.625 10000 ;
      RECT 18884.105 1046.935 18884.385 10000 ;
      RECT 18882.985 1046.935 18883.265 10000 ;
      RECT 18881.865 1046.935 18882.145 10000 ;
      RECT 18866.885 1046.435 18879.205 10000 ;
      RECT 18861.705 1046.935 18861.985 10000 ;
      RECT 18860.585 1046.935 18860.865 10000 ;
      RECT 18859.465 1046.935 18859.745 10000 ;
      RECT 18854.425 1046.935 18854.705 10000 ;
      RECT 18814.805 1046.935 18853.585 10000 ;
      RECT 18806.265 1046.935 18806.545 10000 ;
      RECT 18805.145 1046.935 18805.425 10000 ;
      RECT 18802.905 1046.935 18803.185 10000 ;
      RECT 18801.785 1046.935 18802.065 10000 ;
      RECT 18792.265 1046.935 18800.805 10000 ;
      RECT 18792.405 1046.435 18800.805 10000 ;
      RECT 18783.165 1046.935 18785.265 10000 ;
      RECT 18781.905 1046.935 18782.185 10000 ;
      RECT 18780.785 1046.935 18781.065 10000 ;
      RECT 18753.765 1046.435 18778.685 10000 ;
      RECT 18750.265 1046.935 18750.545 10000 ;
      RECT 18749.145 1046.935 18749.425 10000 ;
      RECT 18740.745 1046.935 18741.025 10000 ;
      RECT 18726.745 1046.935 18739.765 10000 ;
      RECT 18726.885 1046.435 18739.765 10000 ;
      RECT 18724.505 1046.935 18724.785 10000 ;
      RECT 18723.385 1046.935 18723.665 10000 ;
      RECT 18722.265 1046.935 18722.545 10000 ;
      RECT 18714.985 1046.935 18715.265 10000 ;
      RECT 18674.805 1046.935 18714.145 10000 ;
      RECT 18673.545 1046.935 18673.825 10000 ;
      RECT 18668.505 1046.935 18668.785 10000 ;
      RECT 18667.385 1046.935 18667.665 10000 ;
      RECT 18652.965 1046.435 18660.805 10000 ;
      RECT 18650.585 1046.935 18650.865 10000 ;
      RECT 18649.465 1046.935 18649.745 10000 ;
      RECT 18647.225 1046.935 18647.505 10000 ;
      RECT 18646.105 1046.935 18646.385 10000 ;
      RECT 18643.165 1046.935 18645.265 10000 ;
      RECT 18613.765 1046.435 18638.685 10000 ;
      RECT 18610.265 1046.935 18610.545 10000 ;
      RECT 18609.145 1046.935 18609.425 10000 ;
      RECT 18608.025 1046.935 18608.305 10000 ;
      RECT 18602.985 1046.935 18603.265 10000 ;
      RECT 18601.865 1046.935 18602.145 10000 ;
      RECT 18587.445 1046.435 18599.765 10000 ;
      RECT 18580.585 1046.935 18580.865 10000 ;
      RECT 18579.465 1046.935 18579.745 10000 ;
      RECT 18577.225 1046.935 18577.505 10000 ;
      RECT 18576.105 1046.935 18576.385 10000 ;
      RECT 18574.985 1046.935 18575.265 10000 ;
      RECT 18534.245 1046.435 18573.445 10000 ;
      RECT 18527.945 1046.935 18528.225 10000 ;
      RECT 18526.825 1046.935 18527.105 10000 ;
      RECT 18525.705 1046.935 18525.985 10000 ;
      RECT 18512.265 1046.935 18520.805 10000 ;
      RECT 18512.405 1046.435 18520.805 10000 ;
      RECT 18511.145 1046.935 18511.425 10000 ;
      RECT 18503.165 1046.435 18504.565 10000 ;
      RECT 18500.785 1046.935 18501.065 10000 ;
      RECT 18499.665 1046.935 18499.945 10000 ;
      RECT 18472.645 1046.435 18498.125 10000 ;
      RECT 18471.385 1046.935 18471.665 10000 ;
      RECT 18470.265 1046.935 18470.545 10000 ;
      RECT 18469.145 1046.935 18469.425 10000 ;
      RECT 18461.865 1046.935 18462.145 10000 ;
      RECT 18460.745 1046.935 18461.025 10000 ;
      RECT 18446.185 1046.935 18459.765 10000 ;
      RECT 18446.325 1046.435 18459.765 10000 ;
      RECT 18441.145 1046.935 18441.425 10000 ;
      RECT 18440.025 1046.935 18440.305 10000 ;
      RECT 18395.365 1046.435 18433.445 10000 ;
      RECT 18392.985 1046.935 18393.265 10000 ;
      RECT 18391.865 1046.935 18392.145 10000 ;
      RECT 18389.625 1046.935 18389.905 10000 ;
      RECT 18388.505 1046.935 18388.785 10000 ;
      RECT 18387.385 1046.935 18387.665 10000 ;
      RECT 18372.965 1046.435 18380.805 10000 ;
      RECT 18371.705 1046.935 18371.985 10000 ;
      RECT 18370.585 1046.935 18370.865 10000 ;
      RECT 18369.465 1046.935 18369.745 10000 ;
      RECT 18362.465 1046.935 18364.565 10000 ;
      RECT 18362.605 1046.435 18364.565 10000 ;
      RECT 18361.345 1046.935 18361.625 10000 ;
      RECT 18333.205 1046.435 18358.125 10000 ;
      RECT 18327.465 1046.935 18327.745 10000 ;
      RECT 18326.345 1046.935 18326.625 10000 ;
      RECT 18324.105 1046.935 18324.385 10000 ;
      RECT 18322.985 1046.935 18323.265 10000 ;
      RECT 18321.865 1046.935 18322.145 10000 ;
      RECT 18306.885 1046.435 18319.205 10000 ;
      RECT 18301.705 1046.935 18301.985 10000 ;
      RECT 18300.585 1046.935 18300.865 10000 ;
      RECT 18299.465 1046.935 18299.745 10000 ;
      RECT 18294.425 1046.935 18294.705 10000 ;
      RECT 18254.805 1046.935 18293.585 10000 ;
      RECT 18246.265 1046.935 18246.545 10000 ;
      RECT 18245.145 1046.935 18245.425 10000 ;
      RECT 18242.905 1046.935 18243.185 10000 ;
      RECT 18241.785 1046.935 18242.065 10000 ;
      RECT 18232.265 1046.935 18240.805 10000 ;
      RECT 18232.405 1046.435 18240.805 10000 ;
      RECT 18223.165 1046.935 18225.265 10000 ;
      RECT 18221.905 1046.935 18222.185 10000 ;
      RECT 18220.785 1046.935 18221.065 10000 ;
      RECT 18193.765 1046.435 18218.685 10000 ;
      RECT 18190.265 1046.935 18190.545 10000 ;
      RECT 18189.145 1046.935 18189.425 10000 ;
      RECT 18180.745 1046.935 18181.025 10000 ;
      RECT 18166.745 1046.935 18179.765 10000 ;
      RECT 18166.885 1046.435 18179.765 10000 ;
      RECT 18164.505 1046.935 18164.785 10000 ;
      RECT 18163.385 1046.935 18163.665 10000 ;
      RECT 18162.265 1046.935 18162.545 10000 ;
      RECT 18154.985 1046.935 18155.265 10000 ;
      RECT 18114.805 1046.935 18154.145 10000 ;
      RECT 18113.545 1046.935 18113.825 10000 ;
      RECT 18108.505 1046.935 18108.785 10000 ;
      RECT 18107.385 1046.935 18107.665 10000 ;
      RECT 18092.965 1046.435 18100.805 10000 ;
      RECT 18090.585 1046.935 18090.865 10000 ;
      RECT 18089.465 1046.935 18089.745 10000 ;
      RECT 18087.225 1046.935 18087.505 10000 ;
      RECT 18086.105 1046.935 18086.385 10000 ;
      RECT 18083.165 1046.935 18085.265 10000 ;
      RECT 18053.765 1046.435 18078.685 10000 ;
      RECT 18050.265 1046.935 18050.545 10000 ;
      RECT 18049.145 1046.935 18049.425 10000 ;
      RECT 18048.025 1046.935 18048.305 10000 ;
      RECT 18042.985 1046.935 18043.265 10000 ;
      RECT 18041.865 1046.935 18042.145 10000 ;
      RECT 18027.445 1046.435 18039.765 10000 ;
      RECT 18020.585 1046.935 18020.865 10000 ;
      RECT 18019.465 1046.935 18019.745 10000 ;
      RECT 18017.225 1046.935 18017.505 10000 ;
      RECT 18016.105 1046.935 18016.385 10000 ;
      RECT 18014.985 1046.935 18015.265 10000 ;
      RECT 17974.245 1046.435 18013.445 10000 ;
      RECT 17967.945 1046.935 17968.225 10000 ;
      RECT 17966.825 1046.935 17967.105 10000 ;
      RECT 17965.705 1046.935 17965.985 10000 ;
      RECT 17952.265 1046.935 17960.805 10000 ;
      RECT 17952.405 1046.435 17960.805 10000 ;
      RECT 17951.145 1046.935 17951.425 10000 ;
      RECT 17943.165 1046.435 17944.565 10000 ;
      RECT 17940.785 1046.935 17941.065 10000 ;
      RECT 17939.665 1046.935 17939.945 10000 ;
      RECT 17912.645 1046.435 17938.125 10000 ;
      RECT 17911.385 1046.935 17911.665 10000 ;
      RECT 17910.265 1046.935 17910.545 10000 ;
      RECT 17909.145 1046.935 17909.425 10000 ;
      RECT 17901.865 1046.935 17902.145 10000 ;
      RECT 17900.745 1046.935 17901.025 10000 ;
      RECT 17886.185 1046.935 17899.765 10000 ;
      RECT 17886.325 1046.435 17899.765 10000 ;
      RECT 17881.145 1046.935 17881.425 10000 ;
      RECT 17880.025 1046.935 17880.305 10000 ;
      RECT 17835.365 1046.435 17873.445 10000 ;
      RECT 17832.985 1046.935 17833.265 10000 ;
      RECT 17831.865 1046.935 17832.145 10000 ;
      RECT 17829.625 1046.935 17829.905 10000 ;
      RECT 17828.505 1046.935 17828.785 10000 ;
      RECT 17827.385 1046.935 17827.665 10000 ;
      RECT 17812.965 1046.435 17820.805 10000 ;
      RECT 17811.705 1046.935 17811.985 10000 ;
      RECT 17810.585 1046.935 17810.865 10000 ;
      RECT 17809.465 1046.935 17809.745 10000 ;
      RECT 17802.465 1046.935 17804.565 10000 ;
      RECT 17802.605 1046.435 17804.565 10000 ;
      RECT 17801.345 1046.935 17801.625 10000 ;
      RECT 17773.205 1046.435 17798.125 10000 ;
      RECT 17767.465 1046.935 17767.745 10000 ;
      RECT 17766.345 1046.935 17766.625 10000 ;
      RECT 17764.105 1046.935 17764.385 10000 ;
      RECT 17762.985 1046.935 17763.265 10000 ;
      RECT 17761.865 1046.935 17762.145 10000 ;
      RECT 17746.885 1046.435 17759.205 10000 ;
      RECT 17741.705 1046.935 17741.985 10000 ;
      RECT 17740.585 1046.935 17740.865 10000 ;
      RECT 17739.465 1046.935 17739.745 10000 ;
      RECT 17734.425 1046.935 17734.705 10000 ;
      RECT 17694.805 1046.935 17733.585 10000 ;
      RECT 17686.265 1046.935 17686.545 10000 ;
      RECT 17685.145 1046.935 17685.425 10000 ;
      RECT 17682.905 1046.935 17683.185 10000 ;
      RECT 17681.785 1046.935 17682.065 10000 ;
      RECT 17672.265 1046.935 17680.805 10000 ;
      RECT 17672.405 1046.435 17680.805 10000 ;
      RECT 17663.165 1046.935 17665.265 10000 ;
      RECT 17661.905 1046.935 17662.185 10000 ;
      RECT 17660.785 1046.935 17661.065 10000 ;
      RECT 17633.765 1046.435 17658.685 10000 ;
      RECT 17630.265 1046.935 17630.545 10000 ;
      RECT 17629.145 1046.935 17629.425 10000 ;
      RECT 17620.745 1046.935 17621.025 10000 ;
      RECT 17606.745 1046.935 17619.765 10000 ;
      RECT 17606.885 1046.435 17619.765 10000 ;
      RECT 17604.505 1046.935 17604.785 10000 ;
      RECT 17603.385 1046.935 17603.665 10000 ;
      RECT 17602.265 1046.935 17602.545 10000 ;
      RECT 17594.985 1046.935 17595.265 10000 ;
      RECT 17554.805 1046.935 17594.145 10000 ;
      RECT 17553.545 1046.935 17553.825 10000 ;
      RECT 17548.505 1046.935 17548.785 10000 ;
      RECT 17547.385 1046.935 17547.665 10000 ;
      RECT 17532.965 1046.435 17540.805 10000 ;
      RECT 17530.585 1046.935 17530.865 10000 ;
      RECT 17529.465 1046.935 17529.745 10000 ;
      RECT 17527.225 1046.935 17527.505 10000 ;
      RECT 17526.105 1046.935 17526.385 10000 ;
      RECT 17523.165 1046.935 17525.265 10000 ;
      RECT 17493.765 1046.435 17518.685 10000 ;
      RECT 17490.265 1046.935 17490.545 10000 ;
      RECT 17489.145 1046.935 17489.425 10000 ;
      RECT 17488.025 1046.935 17488.305 10000 ;
      RECT 17482.985 1046.935 17483.265 10000 ;
      RECT 17481.865 1046.935 17482.145 10000 ;
      RECT 17467.445 1046.435 17479.765 10000 ;
      RECT 17460.585 1046.935 17460.865 10000 ;
      RECT 17459.465 1046.935 17459.745 10000 ;
      RECT 17457.225 1046.935 17457.505 10000 ;
      RECT 17456.105 1046.935 17456.385 10000 ;
      RECT 17454.985 1046.935 17455.265 10000 ;
      RECT 17414.245 1046.435 17453.445 10000 ;
      RECT 17407.945 1046.935 17408.225 10000 ;
      RECT 17406.825 1046.935 17407.105 10000 ;
      RECT 17405.705 1046.935 17405.985 10000 ;
      RECT 17392.265 1046.935 17400.805 10000 ;
      RECT 17392.405 1046.435 17400.805 10000 ;
      RECT 17391.145 1046.935 17391.425 10000 ;
      RECT 17383.165 1046.435 17384.565 10000 ;
      RECT 17380.785 1046.935 17381.065 10000 ;
      RECT 17379.665 1046.935 17379.945 10000 ;
      RECT 17352.645 1046.435 17378.125 10000 ;
      RECT 17351.385 1046.935 17351.665 10000 ;
      RECT 17350.265 1046.935 17350.545 10000 ;
      RECT 17349.145 1046.935 17349.425 10000 ;
      RECT 17341.865 1046.935 17342.145 10000 ;
      RECT 17340.745 1046.935 17341.025 10000 ;
      RECT 17326.185 1046.935 17339.765 10000 ;
      RECT 17326.325 1046.435 17339.765 10000 ;
      RECT 17321.145 1046.935 17321.425 10000 ;
      RECT 17320.025 1046.935 17320.305 10000 ;
      RECT 17275.365 1046.435 17313.445 10000 ;
      RECT 17272.985 1046.935 17273.265 10000 ;
      RECT 17271.865 1046.935 17272.145 10000 ;
      RECT 17269.625 1046.935 17269.905 10000 ;
      RECT 17268.505 1046.935 17268.785 10000 ;
      RECT 17267.385 1046.935 17267.665 10000 ;
      RECT 17252.965 1046.435 17260.805 10000 ;
      RECT 17251.705 1046.935 17251.985 10000 ;
      RECT 17250.585 1046.935 17250.865 10000 ;
      RECT 17249.465 1046.935 17249.745 10000 ;
      RECT 17242.465 1046.935 17244.565 10000 ;
      RECT 17242.605 1046.435 17244.565 10000 ;
      RECT 17241.345 1046.935 17241.625 10000 ;
      RECT 17213.205 1046.435 17238.125 10000 ;
      RECT 17207.465 1046.935 17207.745 10000 ;
      RECT 17206.345 1046.935 17206.625 10000 ;
      RECT 17204.105 1046.935 17204.385 10000 ;
      RECT 17202.985 1046.935 17203.265 10000 ;
      RECT 17201.865 1046.935 17202.145 10000 ;
      RECT 17186.885 1046.435 17199.205 10000 ;
      RECT 17181.705 1046.935 17181.985 10000 ;
      RECT 17180.585 1046.935 17180.865 10000 ;
      RECT 17179.465 1046.935 17179.745 10000 ;
      RECT 17174.425 1046.935 17174.705 10000 ;
      RECT 17134.805 1046.935 17173.585 10000 ;
      RECT 17126.265 1046.935 17126.545 10000 ;
      RECT 17125.145 1046.935 17125.425 10000 ;
      RECT 17122.905 1046.935 17123.185 10000 ;
      RECT 17121.785 1046.935 17122.065 10000 ;
      RECT 17112.265 1046.935 17120.805 10000 ;
      RECT 17112.405 1046.435 17120.805 10000 ;
      RECT 17103.165 1046.935 17105.265 10000 ;
      RECT 17101.905 1046.935 17102.185 10000 ;
      RECT 17100.785 1046.935 17101.065 10000 ;
      RECT 17073.765 1046.435 17098.685 10000 ;
      RECT 17070.265 1046.935 17070.545 10000 ;
      RECT 17069.145 1046.935 17069.425 10000 ;
      RECT 17060.745 1046.935 17061.025 10000 ;
      RECT 17046.745 1046.935 17059.765 10000 ;
      RECT 17046.885 1046.435 17059.765 10000 ;
      RECT 17044.505 1046.935 17044.785 10000 ;
      RECT 17043.385 1046.935 17043.665 10000 ;
      RECT 17042.265 1046.935 17042.545 10000 ;
      RECT 17034.985 1046.935 17035.265 10000 ;
      RECT 16994.805 1046.935 17034.145 10000 ;
      RECT 16993.545 1046.935 16993.825 10000 ;
      RECT 16988.505 1046.935 16988.785 10000 ;
      RECT 16987.385 1046.935 16987.665 10000 ;
      RECT 16972.965 1046.435 16980.805 10000 ;
      RECT 16970.585 1046.935 16970.865 10000 ;
      RECT 16969.465 1046.935 16969.745 10000 ;
      RECT 16967.225 1046.935 16967.505 10000 ;
      RECT 16966.105 1046.935 16966.385 10000 ;
      RECT 16963.165 1046.935 16965.265 10000 ;
      RECT 16933.765 1046.435 16958.685 10000 ;
      RECT 16930.265 1046.935 16930.545 10000 ;
      RECT 16929.145 1046.935 16929.425 10000 ;
      RECT 16928.025 1046.935 16928.305 10000 ;
      RECT 16922.985 1046.935 16923.265 10000 ;
      RECT 16921.865 1046.935 16922.145 10000 ;
      RECT 16907.445 1046.435 16919.765 10000 ;
      RECT 16900.585 1046.935 16900.865 10000 ;
      RECT 16899.465 1046.935 16899.745 10000 ;
      RECT 16897.225 1046.935 16897.505 10000 ;
      RECT 16896.105 1046.935 16896.385 10000 ;
      RECT 16894.985 1046.935 16895.265 10000 ;
      RECT 16854.245 1046.435 16893.445 10000 ;
      RECT 16847.945 1046.935 16848.225 10000 ;
      RECT 16846.825 1046.935 16847.105 10000 ;
      RECT 16845.705 1046.935 16845.985 10000 ;
      RECT 16832.265 1046.935 16840.805 10000 ;
      RECT 16832.405 1046.435 16840.805 10000 ;
      RECT 16831.145 1046.935 16831.425 10000 ;
      RECT 16823.165 1046.435 16824.565 10000 ;
      RECT 16820.785 1046.935 16821.065 10000 ;
      RECT 16819.665 1046.935 16819.945 10000 ;
      RECT 16792.645 1046.435 16818.125 10000 ;
      RECT 16791.385 1046.935 16791.665 10000 ;
      RECT 16790.265 1046.935 16790.545 10000 ;
      RECT 16789.145 1046.935 16789.425 10000 ;
      RECT 16781.865 1046.935 16782.145 10000 ;
      RECT 16780.745 1046.935 16781.025 10000 ;
      RECT 16766.185 1046.935 16779.765 10000 ;
      RECT 16766.325 1046.435 16779.765 10000 ;
      RECT 16761.145 1046.935 16761.425 10000 ;
      RECT 16760.025 1046.935 16760.305 10000 ;
      RECT 16715.365 1046.435 16753.445 10000 ;
      RECT 16712.985 1046.935 16713.265 10000 ;
      RECT 16711.865 1046.935 16712.145 10000 ;
      RECT 16709.625 1046.935 16709.905 10000 ;
      RECT 16708.505 1046.935 16708.785 10000 ;
      RECT 16707.385 1046.935 16707.665 10000 ;
      RECT 16692.965 1046.435 16700.805 10000 ;
      RECT 16691.705 1046.935 16691.985 10000 ;
      RECT 16690.585 1046.935 16690.865 10000 ;
      RECT 16689.465 1046.935 16689.745 10000 ;
      RECT 16682.465 1046.935 16684.565 10000 ;
      RECT 16682.605 1046.435 16684.565 10000 ;
      RECT 16681.345 1046.935 16681.625 10000 ;
      RECT 16653.205 1046.435 16678.125 10000 ;
      RECT 16647.465 1046.935 16647.745 10000 ;
      RECT 16646.345 1046.935 16646.625 10000 ;
      RECT 16644.105 1046.935 16644.385 10000 ;
      RECT 16642.985 1046.935 16643.265 10000 ;
      RECT 16641.865 1046.935 16642.145 10000 ;
      RECT 16626.885 1046.435 16639.205 10000 ;
      RECT 16621.705 1046.935 16621.985 10000 ;
      RECT 16620.585 1046.935 16620.865 10000 ;
      RECT 16619.465 1046.935 16619.745 10000 ;
      RECT 16614.425 1046.935 16614.705 10000 ;
      RECT 16574.805 1046.935 16613.585 10000 ;
      RECT 16566.265 1046.935 16566.545 10000 ;
      RECT 16565.145 1046.935 16565.425 10000 ;
      RECT 16562.905 1046.935 16563.185 10000 ;
      RECT 16561.785 1046.935 16562.065 10000 ;
      RECT 16552.265 1046.935 16560.805 10000 ;
      RECT 16552.405 1046.435 16560.805 10000 ;
      RECT 16543.165 1046.935 16545.265 10000 ;
      RECT 16541.905 1046.935 16542.185 10000 ;
      RECT 16540.785 1046.935 16541.065 10000 ;
      RECT 16513.765 1046.435 16538.685 10000 ;
      RECT 16510.265 1046.935 16510.545 10000 ;
      RECT 16509.145 1046.935 16509.425 10000 ;
      RECT 16500.745 1046.935 16501.025 10000 ;
      RECT 16486.745 1046.935 16499.765 10000 ;
      RECT 16486.885 1046.435 16499.765 10000 ;
      RECT 16484.505 1046.935 16484.785 10000 ;
      RECT 16483.385 1046.935 16483.665 10000 ;
      RECT 16482.265 1046.935 16482.545 10000 ;
      RECT 16474.985 1046.935 16475.265 10000 ;
      RECT 16434.805 1046.935 16474.145 10000 ;
      RECT 16433.545 1046.935 16433.825 10000 ;
      RECT 16428.505 1046.935 16428.785 10000 ;
      RECT 16427.385 1046.935 16427.665 10000 ;
      RECT 16412.965 1046.435 16420.805 10000 ;
      RECT 16410.585 1046.935 16410.865 10000 ;
      RECT 16409.465 1046.935 16409.745 10000 ;
      RECT 16407.225 1046.935 16407.505 10000 ;
      RECT 16406.105 1046.935 16406.385 10000 ;
      RECT 16403.165 1046.935 16405.265 10000 ;
      RECT 16373.765 1046.435 16398.685 10000 ;
      RECT 16370.265 1046.935 16370.545 10000 ;
      RECT 16369.145 1046.935 16369.425 10000 ;
      RECT 16368.025 1046.935 16368.305 10000 ;
      RECT 16362.985 1046.935 16363.265 10000 ;
      RECT 16361.865 1046.935 16362.145 10000 ;
      RECT 16347.445 1046.435 16359.765 10000 ;
      RECT 16340.585 1046.935 16340.865 10000 ;
      RECT 16339.465 1046.935 16339.745 10000 ;
      RECT 16337.225 1046.935 16337.505 10000 ;
      RECT 16336.105 1046.935 16336.385 10000 ;
      RECT 16334.985 1046.935 16335.265 10000 ;
      RECT 16294.245 1046.435 16333.445 10000 ;
      RECT 16287.945 1046.935 16288.225 10000 ;
      RECT 16286.825 1046.935 16287.105 10000 ;
      RECT 16285.705 1046.935 16285.985 10000 ;
      RECT 16272.265 1046.935 16280.805 10000 ;
      RECT 16272.405 1046.435 16280.805 10000 ;
      RECT 16271.145 1046.935 16271.425 10000 ;
      RECT 16263.165 1046.435 16264.565 10000 ;
      RECT 16260.785 1046.935 16261.065 10000 ;
      RECT 16259.665 1046.935 16259.945 10000 ;
      RECT 16232.645 1046.435 16258.125 10000 ;
      RECT 16231.385 1046.935 16231.665 10000 ;
      RECT 16230.265 1046.935 16230.545 10000 ;
      RECT 16229.145 1046.935 16229.425 10000 ;
      RECT 16221.865 1046.935 16222.145 10000 ;
      RECT 16220.745 1046.935 16221.025 10000 ;
      RECT 16206.185 1046.935 16219.765 10000 ;
      RECT 16206.325 1046.435 16219.765 10000 ;
      RECT 16201.145 1046.935 16201.425 10000 ;
      RECT 16200.025 1046.935 16200.305 10000 ;
      RECT 16155.365 1046.435 16193.445 10000 ;
      RECT 16152.985 1046.935 16153.265 10000 ;
      RECT 16151.865 1046.935 16152.145 10000 ;
      RECT 16149.625 1046.935 16149.905 10000 ;
      RECT 16148.505 1046.935 16148.785 10000 ;
      RECT 16147.385 1046.935 16147.665 10000 ;
      RECT 16132.965 1046.435 16140.805 10000 ;
      RECT 16131.705 1046.935 16131.985 10000 ;
      RECT 16130.585 1046.935 16130.865 10000 ;
      RECT 16129.465 1046.935 16129.745 10000 ;
      RECT 16122.465 1046.935 16124.565 10000 ;
      RECT 16122.605 1046.435 16124.565 10000 ;
      RECT 16121.345 1046.935 16121.625 10000 ;
      RECT 16093.205 1046.435 16118.125 10000 ;
      RECT 16087.465 1046.935 16087.745 10000 ;
      RECT 16086.345 1046.935 16086.625 10000 ;
      RECT 16084.105 1046.935 16084.385 10000 ;
      RECT 16082.985 1046.935 16083.265 10000 ;
      RECT 16081.865 1046.935 16082.145 10000 ;
      RECT 16066.885 1046.435 16079.205 10000 ;
      RECT 16061.705 1046.935 16061.985 10000 ;
      RECT 16060.585 1046.935 16060.865 10000 ;
      RECT 16059.465 1046.935 16059.745 10000 ;
      RECT 16054.425 1046.935 16054.705 10000 ;
      RECT 16014.805 1046.935 16053.585 10000 ;
      RECT 16006.265 1046.935 16006.545 10000 ;
      RECT 16005.145 1046.935 16005.425 10000 ;
      RECT 16002.905 1046.935 16003.185 10000 ;
      RECT 16001.785 1046.935 16002.065 10000 ;
      RECT 15992.265 1046.935 16000.805 10000 ;
      RECT 15992.405 1046.435 16000.805 10000 ;
      RECT 15983.165 1046.935 15985.265 10000 ;
      RECT 15981.905 1046.935 15982.185 10000 ;
      RECT 15980.785 1046.935 15981.065 10000 ;
      RECT 15953.765 1046.435 15978.685 10000 ;
      RECT 15950.265 1046.935 15950.545 10000 ;
      RECT 15949.145 1046.935 15949.425 10000 ;
      RECT 15940.745 1046.935 15941.025 10000 ;
      RECT 15926.745 1046.935 15939.765 10000 ;
      RECT 15926.885 1046.435 15939.765 10000 ;
      RECT 15924.505 1046.935 15924.785 10000 ;
      RECT 15923.385 1046.935 15923.665 10000 ;
      RECT 15922.265 1046.935 15922.545 10000 ;
      RECT 15914.985 1046.935 15915.265 10000 ;
      RECT 15874.805 1046.935 15914.145 10000 ;
      RECT 15873.545 1046.935 15873.825 10000 ;
      RECT 15868.505 1046.935 15868.785 10000 ;
      RECT 15867.385 1046.935 15867.665 10000 ;
      RECT 15852.965 1046.435 15860.805 10000 ;
      RECT 15850.585 1046.935 15850.865 10000 ;
      RECT 15849.465 1046.935 15849.745 10000 ;
      RECT 15847.225 1046.935 15847.505 10000 ;
      RECT 15846.105 1046.935 15846.385 10000 ;
      RECT 15843.165 1046.935 15845.265 10000 ;
      RECT 15813.765 1046.435 15838.685 10000 ;
      RECT 15810.265 1046.935 15810.545 10000 ;
      RECT 15809.145 1046.935 15809.425 10000 ;
      RECT 15808.025 1046.935 15808.305 10000 ;
      RECT 15802.985 1046.935 15803.265 10000 ;
      RECT 15801.865 1046.935 15802.145 10000 ;
      RECT 15787.445 1046.435 15799.765 10000 ;
      RECT 15780.585 1046.935 15780.865 10000 ;
      RECT 15779.465 1046.935 15779.745 10000 ;
      RECT 15777.225 1046.935 15777.505 10000 ;
      RECT 15776.105 1046.935 15776.385 10000 ;
      RECT 15774.985 1046.935 15775.265 10000 ;
      RECT 15734.245 1046.435 15773.445 10000 ;
      RECT 15727.945 1046.935 15728.225 10000 ;
      RECT 15726.825 1046.935 15727.105 10000 ;
      RECT 15725.705 1046.935 15725.985 10000 ;
      RECT 15712.265 1046.935 15720.805 10000 ;
      RECT 15712.405 1046.435 15720.805 10000 ;
      RECT 15711.145 1046.935 15711.425 10000 ;
      RECT 15703.165 1046.435 15704.565 10000 ;
      RECT 15700.785 1046.935 15701.065 10000 ;
      RECT 15699.665 1046.935 15699.945 10000 ;
      RECT 15672.645 1046.435 15698.125 10000 ;
      RECT 15671.385 1046.935 15671.665 10000 ;
      RECT 15670.265 1046.935 15670.545 10000 ;
      RECT 15669.145 1046.935 15669.425 10000 ;
      RECT 15661.865 1046.935 15662.145 10000 ;
      RECT 15660.745 1046.935 15661.025 10000 ;
      RECT 15646.185 1046.935 15659.765 10000 ;
      RECT 15646.325 1046.435 15659.765 10000 ;
      RECT 15641.145 1046.935 15641.425 10000 ;
      RECT 15640.025 1046.935 15640.305 10000 ;
      RECT 15595.365 1046.435 15633.445 10000 ;
      RECT 15592.985 1046.935 15593.265 10000 ;
      RECT 15591.865 1046.935 15592.145 10000 ;
      RECT 15589.625 1046.935 15589.905 10000 ;
      RECT 15588.505 1046.935 15588.785 10000 ;
      RECT 15587.385 1046.935 15587.665 10000 ;
      RECT 15572.965 1046.435 15580.805 10000 ;
      RECT 15571.705 1046.935 15571.985 10000 ;
      RECT 15570.585 1046.935 15570.865 10000 ;
      RECT 15569.465 1046.935 15569.745 10000 ;
      RECT 15562.465 1046.935 15564.565 10000 ;
      RECT 15562.605 1046.435 15564.565 10000 ;
      RECT 15561.345 1046.935 15561.625 10000 ;
      RECT 15533.205 1046.435 15558.125 10000 ;
      RECT 15527.465 1046.935 15527.745 10000 ;
      RECT 15526.345 1046.935 15526.625 10000 ;
      RECT 15524.105 1046.935 15524.385 10000 ;
      RECT 15522.985 1046.935 15523.265 10000 ;
      RECT 15521.865 1046.935 15522.145 10000 ;
      RECT 15506.885 1046.435 15519.205 10000 ;
      RECT 15501.705 1046.935 15501.985 10000 ;
      RECT 15500.585 1046.935 15500.865 10000 ;
      RECT 15499.465 1046.935 15499.745 10000 ;
      RECT 15494.425 1046.935 15494.705 10000 ;
      RECT 15454.805 1046.935 15493.585 10000 ;
      RECT 15446.265 1046.935 15446.545 10000 ;
      RECT 15445.145 1046.935 15445.425 10000 ;
      RECT 15442.905 1046.935 15443.185 10000 ;
      RECT 15441.785 1046.935 15442.065 10000 ;
      RECT 15432.265 1046.935 15440.805 10000 ;
      RECT 15432.405 1046.435 15440.805 10000 ;
      RECT 15423.165 1046.935 15425.265 10000 ;
      RECT 15421.905 1046.935 15422.185 10000 ;
      RECT 15420.785 1046.935 15421.065 10000 ;
      RECT 15393.765 1046.435 15418.685 10000 ;
      RECT 15390.265 1046.935 15390.545 10000 ;
      RECT 15389.145 1046.935 15389.425 10000 ;
      RECT 15380.745 1046.935 15381.025 10000 ;
      RECT 15366.745 1046.935 15379.765 10000 ;
      RECT 15366.885 1046.435 15379.765 10000 ;
      RECT 15364.505 1046.935 15364.785 10000 ;
      RECT 15363.385 1046.935 15363.665 10000 ;
      RECT 15362.265 1046.935 15362.545 10000 ;
      RECT 15354.985 1046.935 15355.265 10000 ;
      RECT 15314.805 1046.935 15354.145 10000 ;
      RECT 15313.545 1046.935 15313.825 10000 ;
      RECT 15308.505 1046.935 15308.785 10000 ;
      RECT 15307.385 1046.935 15307.665 10000 ;
      RECT 15292.965 1046.435 15300.805 10000 ;
      RECT 15290.585 1046.935 15290.865 10000 ;
      RECT 15289.465 1046.935 15289.745 10000 ;
      RECT 15287.225 1046.935 15287.505 10000 ;
      RECT 15286.105 1046.935 15286.385 10000 ;
      RECT 15283.165 1046.935 15285.265 10000 ;
      RECT 15253.765 1046.435 15278.685 10000 ;
      RECT 15250.265 1046.935 15250.545 10000 ;
      RECT 15249.145 1046.935 15249.425 10000 ;
      RECT 15248.025 1046.935 15248.305 10000 ;
      RECT 15242.985 1046.935 15243.265 10000 ;
      RECT 15241.865 1046.935 15242.145 10000 ;
      RECT 15227.445 1046.435 15239.765 10000 ;
      RECT 15220.585 1046.935 15220.865 10000 ;
      RECT 15219.465 1046.935 15219.745 10000 ;
      RECT 15217.225 1046.935 15217.505 10000 ;
      RECT 15216.105 1046.935 15216.385 10000 ;
      RECT 15214.985 1046.935 15215.265 10000 ;
      RECT 15174.245 1046.435 15213.445 10000 ;
      RECT 15167.945 1046.935 15168.225 10000 ;
      RECT 15166.825 1046.935 15167.105 10000 ;
      RECT 15165.705 1046.935 15165.985 10000 ;
      RECT 15152.265 1046.935 15160.805 10000 ;
      RECT 15152.405 1046.435 15160.805 10000 ;
      RECT 15151.145 1046.935 15151.425 10000 ;
      RECT 15143.165 1046.435 15144.565 10000 ;
      RECT 15140.785 1046.935 15141.065 10000 ;
      RECT 15139.665 1046.935 15139.945 10000 ;
      RECT 15112.645 1046.435 15138.125 10000 ;
      RECT 15111.385 1046.935 15111.665 10000 ;
      RECT 15110.265 1046.935 15110.545 10000 ;
      RECT 15109.145 1046.935 15109.425 10000 ;
      RECT 15101.865 1046.935 15102.145 10000 ;
      RECT 15100.745 1046.935 15101.025 10000 ;
      RECT 15086.185 1046.935 15099.765 10000 ;
      RECT 15086.325 1046.435 15099.765 10000 ;
      RECT 15081.145 1046.935 15081.425 10000 ;
      RECT 15080.025 1046.935 15080.305 10000 ;
      RECT 15035.365 1046.435 15073.445 10000 ;
      RECT 15032.985 1046.935 15033.265 10000 ;
      RECT 15031.865 1046.935 15032.145 10000 ;
      RECT 15029.625 1046.935 15029.905 10000 ;
      RECT 15028.505 1046.935 15028.785 10000 ;
      RECT 15027.385 1046.935 15027.665 10000 ;
      RECT 15012.965 1046.435 15020.805 10000 ;
      RECT 15011.705 1046.935 15011.985 10000 ;
      RECT 15010.585 1046.935 15010.865 10000 ;
      RECT 15009.465 1046.935 15009.745 10000 ;
      RECT 15002.465 1046.935 15004.565 10000 ;
      RECT 15002.605 1046.435 15004.565 10000 ;
      RECT 15001.345 1046.935 15001.625 10000 ;
      RECT 14973.205 1046.435 14998.125 10000 ;
      RECT 14967.465 1046.935 14967.745 10000 ;
      RECT 14966.345 1046.935 14966.625 10000 ;
      RECT 14964.105 1046.935 14964.385 10000 ;
      RECT 14962.985 1046.935 14963.265 10000 ;
      RECT 14961.865 1046.935 14962.145 10000 ;
      RECT 14946.885 1046.435 14959.205 10000 ;
      RECT 14941.705 1046.935 14941.985 10000 ;
      RECT 14940.585 1046.935 14940.865 10000 ;
      RECT 14939.465 1046.935 14939.745 10000 ;
      RECT 14934.425 1046.935 14934.705 10000 ;
      RECT 14894.805 1046.935 14933.585 10000 ;
      RECT 14886.265 1046.935 14886.545 10000 ;
      RECT 14885.145 1046.935 14885.425 10000 ;
      RECT 14882.905 1046.935 14883.185 10000 ;
      RECT 14881.785 1046.935 14882.065 10000 ;
      RECT 14872.265 1046.935 14880.805 10000 ;
      RECT 14872.405 1046.435 14880.805 10000 ;
      RECT 14863.165 1046.935 14865.265 10000 ;
      RECT 14861.905 1046.935 14862.185 10000 ;
      RECT 14860.785 1046.935 14861.065 10000 ;
      RECT 14833.765 1046.435 14858.685 10000 ;
      RECT 14830.265 1046.935 14830.545 10000 ;
      RECT 14829.145 1046.935 14829.425 10000 ;
      RECT 14820.745 1046.935 14821.025 10000 ;
      RECT 14806.745 1046.935 14819.765 10000 ;
      RECT 14806.885 1046.435 14819.765 10000 ;
      RECT 14804.505 1046.935 14804.785 10000 ;
      RECT 14803.385 1046.935 14803.665 10000 ;
      RECT 14802.265 1046.935 14802.545 10000 ;
      RECT 14794.985 1046.935 14795.265 10000 ;
      RECT 14754.805 1046.935 14794.145 10000 ;
      RECT 14753.545 1046.935 14753.825 10000 ;
      RECT 14748.505 1046.935 14748.785 10000 ;
      RECT 14747.385 1046.935 14747.665 10000 ;
      RECT 14732.965 1046.435 14740.805 10000 ;
      RECT 14730.585 1046.935 14730.865 10000 ;
      RECT 14729.465 1046.935 14729.745 10000 ;
      RECT 14727.225 1046.935 14727.505 10000 ;
      RECT 14726.105 1046.935 14726.385 10000 ;
      RECT 14723.165 1046.935 14725.265 10000 ;
      RECT 14693.765 1046.435 14718.685 10000 ;
      RECT 14690.265 1046.935 14690.545 10000 ;
      RECT 14689.145 1046.935 14689.425 10000 ;
      RECT 14688.025 1046.935 14688.305 10000 ;
      RECT 14682.985 1046.935 14683.265 10000 ;
      RECT 14681.865 1046.935 14682.145 10000 ;
      RECT 14667.445 1046.435 14679.765 10000 ;
      RECT 14660.585 1046.935 14660.865 10000 ;
      RECT 14659.465 1046.935 14659.745 10000 ;
      RECT 14657.225 1046.935 14657.505 10000 ;
      RECT 14656.105 1046.935 14656.385 10000 ;
      RECT 14654.985 1046.935 14655.265 10000 ;
      RECT 14614.245 1046.435 14653.445 10000 ;
      RECT 14607.945 1046.935 14608.225 10000 ;
      RECT 14606.825 1046.935 14607.105 10000 ;
      RECT 14605.705 1046.935 14605.985 10000 ;
      RECT 14592.265 1046.935 14600.805 10000 ;
      RECT 14592.405 1046.435 14600.805 10000 ;
      RECT 14591.145 1046.935 14591.425 10000 ;
      RECT 14583.165 1046.435 14584.565 10000 ;
      RECT 14580.785 1046.935 14581.065 10000 ;
      RECT 14579.665 1046.935 14579.945 10000 ;
      RECT 14552.645 1046.435 14578.125 10000 ;
      RECT 14551.385 1046.935 14551.665 10000 ;
      RECT 14550.265 1046.935 14550.545 10000 ;
      RECT 14549.145 1046.935 14549.425 10000 ;
      RECT 14541.865 1046.935 14542.145 10000 ;
      RECT 14540.745 1046.935 14541.025 10000 ;
      RECT 14526.185 1046.935 14539.765 10000 ;
      RECT 14526.325 1046.435 14539.765 10000 ;
      RECT 14521.145 1046.935 14521.425 10000 ;
      RECT 14520.025 1046.935 14520.305 10000 ;
      RECT 14475.365 1046.435 14513.445 10000 ;
      RECT 14472.985 1046.935 14473.265 10000 ;
      RECT 14471.865 1046.935 14472.145 10000 ;
      RECT 14469.625 1046.935 14469.905 10000 ;
      RECT 14468.505 1046.935 14468.785 10000 ;
      RECT 14467.385 1046.935 14467.665 10000 ;
      RECT 14452.965 1046.435 14460.805 10000 ;
      RECT 14451.705 1046.935 14451.985 10000 ;
      RECT 14450.585 1046.935 14450.865 10000 ;
      RECT 14449.465 1046.935 14449.745 10000 ;
      RECT 14442.465 1046.935 14444.565 10000 ;
      RECT 14442.605 1046.435 14444.565 10000 ;
      RECT 14441.345 1046.935 14441.625 10000 ;
      RECT 14413.205 1046.435 14438.125 10000 ;
      RECT 14407.465 1046.935 14407.745 10000 ;
      RECT 14406.345 1046.935 14406.625 10000 ;
      RECT 14404.105 1046.935 14404.385 10000 ;
      RECT 14402.985 1046.935 14403.265 10000 ;
      RECT 14401.865 1046.935 14402.145 10000 ;
      RECT 14386.885 1046.435 14399.205 10000 ;
      RECT 14381.705 1046.935 14381.985 10000 ;
      RECT 14380.585 1046.935 14380.865 10000 ;
      RECT 14379.465 1046.935 14379.745 10000 ;
      RECT 14374.425 1046.935 14374.705 10000 ;
      RECT 14334.805 1046.935 14373.585 10000 ;
      RECT 14326.265 1046.935 14326.545 10000 ;
      RECT 14325.145 1046.935 14325.425 10000 ;
      RECT 14322.905 1046.935 14323.185 10000 ;
      RECT 14321.785 1046.935 14322.065 10000 ;
      RECT 14312.265 1046.935 14320.805 10000 ;
      RECT 14312.405 1046.435 14320.805 10000 ;
      RECT 14303.165 1046.935 14305.265 10000 ;
      RECT 14301.905 1046.935 14302.185 10000 ;
      RECT 14300.785 1046.935 14301.065 10000 ;
      RECT 14273.765 1046.435 14298.685 10000 ;
      RECT 14270.265 1046.935 14270.545 10000 ;
      RECT 14269.145 1046.935 14269.425 10000 ;
      RECT 14260.745 1046.935 14261.025 10000 ;
      RECT 14246.745 1046.935 14259.765 10000 ;
      RECT 14246.885 1046.435 14259.765 10000 ;
      RECT 14244.505 1046.935 14244.785 10000 ;
      RECT 14243.385 1046.935 14243.665 10000 ;
      RECT 14242.265 1046.935 14242.545 10000 ;
      RECT 14234.985 1046.935 14235.265 10000 ;
      RECT 14234.005 1046.935 14234.145 10000 ;
      RECT 18814.805 1046.435 18853.445 10000 ;
      RECT 18783.165 1046.435 18785.125 10000 ;
      RECT 18674.805 1046.435 18714.005 10000 ;
      RECT 18643.165 1046.435 18645.125 10000 ;
      RECT 18254.805 1046.435 18293.445 10000 ;
      RECT 18223.165 1046.435 18225.125 10000 ;
      RECT 18114.805 1046.435 18154.005 10000 ;
      RECT 18083.165 1046.435 18085.125 10000 ;
      RECT 17694.805 1046.435 17733.445 10000 ;
      RECT 17663.165 1046.435 17665.125 10000 ;
      RECT 17554.805 1046.435 17594.005 10000 ;
      RECT 17523.165 1046.435 17525.125 10000 ;
      RECT 17134.805 1046.435 17173.445 10000 ;
      RECT 17103.165 1046.435 17105.125 10000 ;
      RECT 16994.805 1046.435 17034.005 10000 ;
      RECT 16963.165 1046.435 16965.125 10000 ;
      RECT 16574.805 1046.435 16613.445 10000 ;
      RECT 16543.165 1046.435 16545.125 10000 ;
      RECT 16434.805 1046.435 16474.005 10000 ;
      RECT 16403.165 1046.435 16405.125 10000 ;
      RECT 16014.805 1046.435 16053.445 10000 ;
      RECT 15983.165 1046.435 15985.125 10000 ;
      RECT 15874.805 1046.435 15914.005 10000 ;
      RECT 15843.165 1046.435 15845.125 10000 ;
      RECT 15454.805 1046.435 15493.445 10000 ;
      RECT 15423.165 1046.435 15425.125 10000 ;
      RECT 15314.805 1046.435 15354.005 10000 ;
      RECT 15283.165 1046.435 15285.125 10000 ;
      RECT 14894.805 1046.435 14933.445 10000 ;
      RECT 14863.165 1046.435 14865.125 10000 ;
      RECT 14754.805 1046.435 14794.005 10000 ;
      RECT 14723.165 1046.435 14725.125 10000 ;
      RECT 14334.805 1046.435 14373.445 10000 ;
      RECT 14303.165 1046.435 14305.125 10000 ;
      RECT 7682.145 1047.855 14234.005 10000 ;
      RECT 14194.805 1046.435 14234.005 10000 ;
      RECT 14193.545 1046.935 14193.825 10000 ;
      RECT 14188.505 1046.935 14188.785 10000 ;
      RECT 14187.385 1046.935 14187.665 10000 ;
      RECT 14172.965 1046.435 14180.805 10000 ;
      RECT 14170.585 1046.935 14170.865 10000 ;
      RECT 14169.465 1046.935 14169.745 10000 ;
      RECT 14167.225 1046.935 14167.505 10000 ;
      RECT 14166.105 1046.935 14166.385 10000 ;
      RECT 14163.165 1046.935 14165.265 10000 ;
      RECT 14133.765 1046.435 14158.685 10000 ;
      RECT 14130.265 1046.935 14130.545 10000 ;
      RECT 14129.145 1046.935 14129.425 10000 ;
      RECT 14128.025 1046.935 14128.305 10000 ;
      RECT 14122.985 1046.935 14123.265 10000 ;
      RECT 14121.865 1046.935 14122.145 10000 ;
      RECT 14107.445 1046.435 14119.765 10000 ;
      RECT 14100.585 1046.935 14100.865 10000 ;
      RECT 14099.465 1046.935 14099.745 10000 ;
      RECT 14097.225 1046.935 14097.505 10000 ;
      RECT 14096.105 1046.935 14096.385 10000 ;
      RECT 14094.985 1046.935 14095.265 10000 ;
      RECT 14054.245 1046.435 14093.445 10000 ;
      RECT 14047.945 1046.935 14048.225 10000 ;
      RECT 14046.825 1046.935 14047.105 10000 ;
      RECT 14045.705 1046.935 14045.985 10000 ;
      RECT 14032.265 1046.935 14040.805 10000 ;
      RECT 14032.405 1046.435 14040.805 10000 ;
      RECT 14031.145 1046.935 14031.425 10000 ;
      RECT 14023.165 1046.435 14024.565 10000 ;
      RECT 14020.785 1046.935 14021.065 10000 ;
      RECT 14019.665 1046.935 14019.945 10000 ;
      RECT 13992.645 1046.435 14018.125 10000 ;
      RECT 13991.385 1046.935 13991.665 10000 ;
      RECT 13990.265 1046.935 13990.545 10000 ;
      RECT 13989.145 1046.935 13989.425 10000 ;
      RECT 13981.865 1046.935 13982.145 10000 ;
      RECT 13980.745 1046.935 13981.025 10000 ;
      RECT 13966.185 1046.935 13979.765 10000 ;
      RECT 13966.325 1046.435 13979.765 10000 ;
      RECT 13961.145 1046.935 13961.425 10000 ;
      RECT 13960.025 1046.935 13960.305 10000 ;
      RECT 13915.365 1046.435 13953.445 10000 ;
      RECT 13912.985 1046.935 13913.265 10000 ;
      RECT 13911.865 1046.935 13912.145 10000 ;
      RECT 13909.625 1046.935 13909.905 10000 ;
      RECT 13908.505 1046.935 13908.785 10000 ;
      RECT 13907.385 1046.935 13907.665 10000 ;
      RECT 13892.965 1046.435 13900.805 10000 ;
      RECT 13891.705 1046.935 13891.985 10000 ;
      RECT 13890.585 1046.935 13890.865 10000 ;
      RECT 13889.465 1046.935 13889.745 10000 ;
      RECT 13882.465 1046.935 13884.565 10000 ;
      RECT 13882.605 1046.435 13884.565 10000 ;
      RECT 13881.345 1046.935 13881.625 10000 ;
      RECT 13853.205 1046.435 13878.125 10000 ;
      RECT 13847.465 1046.935 13847.745 10000 ;
      RECT 13846.345 1046.935 13846.625 10000 ;
      RECT 13844.105 1046.935 13844.385 10000 ;
      RECT 13842.985 1046.935 13843.265 10000 ;
      RECT 13841.865 1046.935 13842.145 10000 ;
      RECT 13826.885 1046.435 13839.205 10000 ;
      RECT 13821.705 1046.935 13821.985 10000 ;
      RECT 13820.585 1046.935 13820.865 10000 ;
      RECT 13819.465 1046.935 13819.745 10000 ;
      RECT 13814.425 1046.935 13814.705 10000 ;
      RECT 13774.805 1046.935 13813.585 10000 ;
      RECT 13766.265 1046.935 13766.545 10000 ;
      RECT 13765.145 1046.935 13765.425 10000 ;
      RECT 13762.905 1046.935 13763.185 10000 ;
      RECT 13761.785 1046.935 13762.065 10000 ;
      RECT 13752.265 1046.935 13760.805 10000 ;
      RECT 13752.405 1046.435 13760.805 10000 ;
      RECT 13743.165 1046.935 13745.265 10000 ;
      RECT 13741.905 1046.935 13742.185 10000 ;
      RECT 13740.785 1046.935 13741.065 10000 ;
      RECT 13713.765 1046.435 13738.685 10000 ;
      RECT 13710.265 1046.935 13710.545 10000 ;
      RECT 13709.145 1046.935 13709.425 10000 ;
      RECT 13700.745 1046.935 13701.025 10000 ;
      RECT 13686.745 1046.935 13699.765 10000 ;
      RECT 13686.885 1046.435 13699.765 10000 ;
      RECT 13684.505 1046.935 13684.785 10000 ;
      RECT 13683.385 1046.935 13683.665 10000 ;
      RECT 13682.265 1046.935 13682.545 10000 ;
      RECT 13674.985 1046.935 13675.265 10000 ;
      RECT 13634.805 1046.935 13674.145 10000 ;
      RECT 13633.545 1046.935 13633.825 10000 ;
      RECT 13628.505 1046.935 13628.785 10000 ;
      RECT 13627.385 1046.935 13627.665 10000 ;
      RECT 13612.965 1046.435 13620.805 10000 ;
      RECT 13610.585 1046.935 13610.865 10000 ;
      RECT 13609.465 1046.935 13609.745 10000 ;
      RECT 13607.225 1046.935 13607.505 10000 ;
      RECT 13606.105 1046.935 13606.385 10000 ;
      RECT 13603.165 1046.935 13605.265 10000 ;
      RECT 13573.765 1046.435 13598.685 10000 ;
      RECT 13570.265 1046.935 13570.545 10000 ;
      RECT 13569.145 1046.935 13569.425 10000 ;
      RECT 13568.025 1046.935 13568.305 10000 ;
      RECT 13562.985 1046.935 13563.265 10000 ;
      RECT 13561.865 1046.935 13562.145 10000 ;
      RECT 13547.445 1046.435 13559.765 10000 ;
      RECT 13540.585 1046.935 13540.865 10000 ;
      RECT 13539.465 1046.935 13539.745 10000 ;
      RECT 13537.225 1046.935 13537.505 10000 ;
      RECT 13536.105 1046.935 13536.385 10000 ;
      RECT 13534.985 1046.935 13535.265 10000 ;
      RECT 13494.245 1046.435 13533.445 10000 ;
      RECT 13487.945 1046.935 13488.225 10000 ;
      RECT 13486.825 1046.935 13487.105 10000 ;
      RECT 13485.705 1046.935 13485.985 10000 ;
      RECT 13472.265 1046.935 13480.805 10000 ;
      RECT 13472.405 1046.435 13480.805 10000 ;
      RECT 13471.145 1046.935 13471.425 10000 ;
      RECT 13463.165 1046.435 13464.565 10000 ;
      RECT 13460.785 1046.935 13461.065 10000 ;
      RECT 13459.665 1046.935 13459.945 10000 ;
      RECT 13432.645 1046.435 13458.125 10000 ;
      RECT 13431.385 1046.935 13431.665 10000 ;
      RECT 13430.265 1046.935 13430.545 10000 ;
      RECT 13429.145 1046.935 13429.425 10000 ;
      RECT 13421.865 1046.935 13422.145 10000 ;
      RECT 13420.745 1046.935 13421.025 10000 ;
      RECT 13406.185 1046.935 13419.765 10000 ;
      RECT 13406.325 1046.435 13419.765 10000 ;
      RECT 13401.145 1046.935 13401.425 10000 ;
      RECT 13400.025 1046.935 13400.305 10000 ;
      RECT 13355.365 1046.435 13393.445 10000 ;
      RECT 13352.985 1046.935 13353.265 10000 ;
      RECT 13351.865 1046.935 13352.145 10000 ;
      RECT 13349.625 1046.935 13349.905 10000 ;
      RECT 13348.505 1046.935 13348.785 10000 ;
      RECT 13347.385 1046.935 13347.665 10000 ;
      RECT 13332.965 1046.435 13340.805 10000 ;
      RECT 13331.705 1046.935 13331.985 10000 ;
      RECT 13330.585 1046.935 13330.865 10000 ;
      RECT 13329.465 1046.935 13329.745 10000 ;
      RECT 13322.465 1046.935 13324.565 10000 ;
      RECT 13322.605 1046.435 13324.565 10000 ;
      RECT 13321.345 1046.935 13321.625 10000 ;
      RECT 13293.205 1046.435 13318.125 10000 ;
      RECT 13287.465 1046.935 13287.745 10000 ;
      RECT 13286.345 1046.935 13286.625 10000 ;
      RECT 13284.105 1046.935 13284.385 10000 ;
      RECT 13282.985 1046.935 13283.265 10000 ;
      RECT 13281.865 1046.935 13282.145 10000 ;
      RECT 13266.885 1046.435 13279.205 10000 ;
      RECT 13261.705 1046.935 13261.985 10000 ;
      RECT 13260.585 1046.935 13260.865 10000 ;
      RECT 13259.465 1046.935 13259.745 10000 ;
      RECT 13254.425 1046.935 13254.705 10000 ;
      RECT 13214.805 1046.935 13253.585 10000 ;
      RECT 13206.265 1046.935 13206.545 10000 ;
      RECT 13205.145 1046.935 13205.425 10000 ;
      RECT 13202.905 1046.935 13203.185 10000 ;
      RECT 13201.785 1046.935 13202.065 10000 ;
      RECT 13192.265 1046.935 13200.805 10000 ;
      RECT 13192.405 1046.435 13200.805 10000 ;
      RECT 13183.165 1046.935 13185.265 10000 ;
      RECT 13181.905 1046.935 13182.185 10000 ;
      RECT 13180.785 1046.935 13181.065 10000 ;
      RECT 13153.765 1046.435 13178.685 10000 ;
      RECT 13150.265 1046.935 13150.545 10000 ;
      RECT 13149.145 1046.935 13149.425 10000 ;
      RECT 13140.745 1046.935 13141.025 10000 ;
      RECT 13126.745 1046.935 13139.765 10000 ;
      RECT 13126.885 1046.435 13139.765 10000 ;
      RECT 13124.505 1046.935 13124.785 10000 ;
      RECT 13123.385 1046.935 13123.665 10000 ;
      RECT 13122.265 1046.935 13122.545 10000 ;
      RECT 13114.985 1046.935 13115.265 10000 ;
      RECT 13074.805 1046.935 13114.145 10000 ;
      RECT 13073.545 1046.935 13073.825 10000 ;
      RECT 13068.505 1046.935 13068.785 10000 ;
      RECT 13067.385 1046.935 13067.665 10000 ;
      RECT 13052.965 1046.435 13060.805 10000 ;
      RECT 13050.585 1046.935 13050.865 10000 ;
      RECT 13049.465 1046.935 13049.745 10000 ;
      RECT 13047.225 1046.935 13047.505 10000 ;
      RECT 13046.105 1046.935 13046.385 10000 ;
      RECT 13043.165 1046.935 13045.265 10000 ;
      RECT 13013.765 1046.435 13038.685 10000 ;
      RECT 13010.265 1046.935 13010.545 10000 ;
      RECT 13009.145 1046.935 13009.425 10000 ;
      RECT 13008.025 1046.935 13008.305 10000 ;
      RECT 13002.985 1046.935 13003.265 10000 ;
      RECT 13001.865 1046.935 13002.145 10000 ;
      RECT 12987.445 1046.435 12999.765 10000 ;
      RECT 12980.585 1046.935 12980.865 10000 ;
      RECT 12979.465 1046.935 12979.745 10000 ;
      RECT 12977.225 1046.935 12977.505 10000 ;
      RECT 12976.105 1046.935 12976.385 10000 ;
      RECT 12974.985 1046.935 12975.265 10000 ;
      RECT 12934.245 1046.435 12973.445 10000 ;
      RECT 12927.945 1046.935 12928.225 10000 ;
      RECT 12926.825 1046.935 12927.105 10000 ;
      RECT 12925.705 1046.935 12925.985 10000 ;
      RECT 12912.265 1046.935 12920.805 10000 ;
      RECT 12912.405 1046.435 12920.805 10000 ;
      RECT 12911.145 1046.935 12911.425 10000 ;
      RECT 12903.165 1046.435 12904.565 10000 ;
      RECT 12900.785 1046.935 12901.065 10000 ;
      RECT 12899.665 1046.935 12899.945 10000 ;
      RECT 12872.645 1046.435 12898.125 10000 ;
      RECT 12871.385 1046.935 12871.665 10000 ;
      RECT 12870.265 1046.935 12870.545 10000 ;
      RECT 12869.145 1046.935 12869.425 10000 ;
      RECT 12861.865 1046.935 12862.145 10000 ;
      RECT 12860.745 1046.935 12861.025 10000 ;
      RECT 12846.185 1046.935 12859.765 10000 ;
      RECT 12846.325 1046.435 12859.765 10000 ;
      RECT 12841.145 1046.935 12841.425 10000 ;
      RECT 12840.025 1046.935 12840.305 10000 ;
      RECT 12795.365 1046.435 12833.445 10000 ;
      RECT 12792.985 1046.935 12793.265 10000 ;
      RECT 12791.865 1046.935 12792.145 10000 ;
      RECT 12789.625 1046.935 12789.905 10000 ;
      RECT 12788.505 1046.935 12788.785 10000 ;
      RECT 12787.385 1046.935 12787.665 10000 ;
      RECT 12772.965 1046.435 12780.805 10000 ;
      RECT 12771.705 1046.935 12771.985 10000 ;
      RECT 12770.585 1046.935 12770.865 10000 ;
      RECT 12769.465 1046.935 12769.745 10000 ;
      RECT 12762.465 1046.935 12764.565 10000 ;
      RECT 12762.605 1046.435 12764.565 10000 ;
      RECT 12761.345 1046.935 12761.625 10000 ;
      RECT 12733.205 1046.435 12758.125 10000 ;
      RECT 12727.465 1046.935 12727.745 10000 ;
      RECT 12726.345 1046.935 12726.625 10000 ;
      RECT 12724.105 1046.935 12724.385 10000 ;
      RECT 12722.985 1046.935 12723.265 10000 ;
      RECT 12721.865 1046.935 12722.145 10000 ;
      RECT 12706.885 1046.435 12719.205 10000 ;
      RECT 12701.705 1046.935 12701.985 10000 ;
      RECT 12700.585 1046.935 12700.865 10000 ;
      RECT 12699.465 1046.935 12699.745 10000 ;
      RECT 12694.425 1046.935 12694.705 10000 ;
      RECT 12654.805 1046.935 12693.585 10000 ;
      RECT 12646.265 1046.935 12646.545 10000 ;
      RECT 12645.145 1046.935 12645.425 10000 ;
      RECT 12642.905 1046.935 12643.185 10000 ;
      RECT 12641.785 1046.935 12642.065 10000 ;
      RECT 12632.265 1046.935 12640.805 10000 ;
      RECT 12632.405 1046.435 12640.805 10000 ;
      RECT 12623.165 1046.935 12625.265 10000 ;
      RECT 12621.905 1046.935 12622.185 10000 ;
      RECT 12620.785 1046.935 12621.065 10000 ;
      RECT 12593.765 1046.435 12618.685 10000 ;
      RECT 12590.265 1046.935 12590.545 10000 ;
      RECT 12589.145 1046.935 12589.425 10000 ;
      RECT 12580.745 1046.935 12581.025 10000 ;
      RECT 12566.745 1046.935 12579.765 10000 ;
      RECT 12566.885 1046.435 12579.765 10000 ;
      RECT 12564.505 1046.935 12564.785 10000 ;
      RECT 12563.385 1046.935 12563.665 10000 ;
      RECT 12562.265 1046.935 12562.545 10000 ;
      RECT 12554.985 1046.935 12555.265 10000 ;
      RECT 12514.805 1046.935 12554.145 10000 ;
      RECT 12513.545 1046.935 12513.825 10000 ;
      RECT 12508.505 1046.935 12508.785 10000 ;
      RECT 12507.385 1046.935 12507.665 10000 ;
      RECT 12492.965 1046.435 12500.805 10000 ;
      RECT 12490.585 1046.935 12490.865 10000 ;
      RECT 12489.465 1046.935 12489.745 10000 ;
      RECT 12487.225 1046.935 12487.505 10000 ;
      RECT 12486.105 1046.935 12486.385 10000 ;
      RECT 12483.165 1046.935 12485.265 10000 ;
      RECT 12453.765 1046.435 12478.685 10000 ;
      RECT 12450.265 1046.935 12450.545 10000 ;
      RECT 12449.145 1046.935 12449.425 10000 ;
      RECT 12448.025 1046.935 12448.305 10000 ;
      RECT 12442.985 1046.935 12443.265 10000 ;
      RECT 12441.865 1046.935 12442.145 10000 ;
      RECT 12427.445 1046.435 12439.765 10000 ;
      RECT 12420.585 1046.935 12420.865 10000 ;
      RECT 12419.465 1046.935 12419.745 10000 ;
      RECT 12417.225 1046.935 12417.505 10000 ;
      RECT 12416.105 1046.935 12416.385 10000 ;
      RECT 12414.985 1046.935 12415.265 10000 ;
      RECT 12374.245 1046.435 12413.445 10000 ;
      RECT 12367.945 1046.935 12368.225 10000 ;
      RECT 12366.825 1046.935 12367.105 10000 ;
      RECT 12365.705 1046.935 12365.985 10000 ;
      RECT 12352.265 1046.935 12360.805 10000 ;
      RECT 12352.405 1046.435 12360.805 10000 ;
      RECT 12351.145 1046.935 12351.425 10000 ;
      RECT 12343.165 1046.435 12344.565 10000 ;
      RECT 12340.785 1046.935 12341.065 10000 ;
      RECT 12339.665 1046.935 12339.945 10000 ;
      RECT 12312.645 1046.435 12338.125 10000 ;
      RECT 12311.385 1046.935 12311.665 10000 ;
      RECT 12310.265 1046.935 12310.545 10000 ;
      RECT 12309.145 1046.935 12309.425 10000 ;
      RECT 12301.865 1046.935 12302.145 10000 ;
      RECT 12300.745 1046.935 12301.025 10000 ;
      RECT 12286.185 1046.935 12299.765 10000 ;
      RECT 12286.325 1046.435 12299.765 10000 ;
      RECT 12281.145 1046.935 12281.425 10000 ;
      RECT 12280.025 1046.935 12280.305 10000 ;
      RECT 12235.365 1046.435 12273.445 10000 ;
      RECT 12232.985 1046.935 12233.265 10000 ;
      RECT 12231.865 1046.935 12232.145 10000 ;
      RECT 12229.625 1046.935 12229.905 10000 ;
      RECT 12228.505 1046.935 12228.785 10000 ;
      RECT 12227.385 1046.935 12227.665 10000 ;
      RECT 12212.965 1046.435 12220.805 10000 ;
      RECT 12211.705 1046.935 12211.985 10000 ;
      RECT 12210.585 1046.935 12210.865 10000 ;
      RECT 12209.465 1046.935 12209.745 10000 ;
      RECT 12202.465 1046.935 12204.565 10000 ;
      RECT 12202.605 1046.435 12204.565 10000 ;
      RECT 12201.345 1046.935 12201.625 10000 ;
      RECT 12173.205 1046.435 12198.125 10000 ;
      RECT 12167.465 1046.935 12167.745 10000 ;
      RECT 12166.345 1046.935 12166.625 10000 ;
      RECT 12164.105 1046.935 12164.385 10000 ;
      RECT 12162.985 1046.935 12163.265 10000 ;
      RECT 12161.865 1046.935 12162.145 10000 ;
      RECT 12146.885 1046.435 12159.205 10000 ;
      RECT 12141.705 1046.935 12141.985 10000 ;
      RECT 12140.585 1046.935 12140.865 10000 ;
      RECT 12139.465 1046.935 12139.745 10000 ;
      RECT 12134.425 1046.935 12134.705 10000 ;
      RECT 12094.805 1046.935 12133.585 10000 ;
      RECT 12086.265 1046.935 12086.545 10000 ;
      RECT 12085.145 1046.935 12085.425 10000 ;
      RECT 12082.905 1046.935 12083.185 10000 ;
      RECT 12081.785 1046.935 12082.065 10000 ;
      RECT 12072.265 1046.935 12080.805 10000 ;
      RECT 12072.405 1046.435 12080.805 10000 ;
      RECT 12063.165 1046.935 12065.265 10000 ;
      RECT 12061.905 1046.935 12062.185 10000 ;
      RECT 12060.785 1046.935 12061.065 10000 ;
      RECT 12033.765 1046.435 12058.685 10000 ;
      RECT 12030.265 1046.935 12030.545 10000 ;
      RECT 12029.145 1046.935 12029.425 10000 ;
      RECT 12020.745 1046.935 12021.025 10000 ;
      RECT 12006.745 1046.935 12019.765 10000 ;
      RECT 12006.885 1046.435 12019.765 10000 ;
      RECT 12004.505 1046.935 12004.785 10000 ;
      RECT 12003.385 1046.935 12003.665 10000 ;
      RECT 12002.265 1046.935 12002.545 10000 ;
      RECT 11994.985 1046.935 11995.265 10000 ;
      RECT 11954.805 1046.935 11994.145 10000 ;
      RECT 11953.545 1046.935 11953.825 10000 ;
      RECT 11948.505 1046.935 11948.785 10000 ;
      RECT 11947.385 1046.935 11947.665 10000 ;
      RECT 11932.965 1046.435 11940.805 10000 ;
      RECT 11930.585 1046.935 11930.865 10000 ;
      RECT 11929.465 1046.935 11929.745 10000 ;
      RECT 11927.225 1046.935 11927.505 10000 ;
      RECT 11926.105 1046.935 11926.385 10000 ;
      RECT 11923.165 1046.935 11925.265 10000 ;
      RECT 11893.765 1046.435 11918.685 10000 ;
      RECT 11890.265 1046.935 11890.545 10000 ;
      RECT 11889.145 1046.935 11889.425 10000 ;
      RECT 11888.025 1046.935 11888.305 10000 ;
      RECT 11882.985 1046.935 11883.265 10000 ;
      RECT 11881.865 1046.935 11882.145 10000 ;
      RECT 11867.445 1046.435 11879.765 10000 ;
      RECT 11860.585 1046.935 11860.865 10000 ;
      RECT 11859.465 1046.935 11859.745 10000 ;
      RECT 11857.225 1046.935 11857.505 10000 ;
      RECT 11856.105 1046.935 11856.385 10000 ;
      RECT 11854.985 1046.935 11855.265 10000 ;
      RECT 11814.245 1046.435 11853.445 10000 ;
      RECT 11807.945 1046.935 11808.225 10000 ;
      RECT 11806.825 1046.935 11807.105 10000 ;
      RECT 11805.705 1046.935 11805.985 10000 ;
      RECT 11792.265 1046.935 11800.805 10000 ;
      RECT 11792.405 1046.435 11800.805 10000 ;
      RECT 11791.145 1046.935 11791.425 10000 ;
      RECT 11783.165 1046.435 11784.565 10000 ;
      RECT 11780.785 1046.935 11781.065 10000 ;
      RECT 11779.665 1046.935 11779.945 10000 ;
      RECT 11752.645 1046.435 11778.125 10000 ;
      RECT 11751.385 1046.935 11751.665 10000 ;
      RECT 11750.265 1046.935 11750.545 10000 ;
      RECT 11749.145 1046.935 11749.425 10000 ;
      RECT 11741.865 1046.935 11742.145 10000 ;
      RECT 11740.745 1046.935 11741.025 10000 ;
      RECT 11726.185 1046.935 11739.765 10000 ;
      RECT 11726.325 1046.435 11739.765 10000 ;
      RECT 11721.145 1046.935 11721.425 10000 ;
      RECT 11720.025 1046.935 11720.305 10000 ;
      RECT 11675.365 1046.435 11713.445 10000 ;
      RECT 11672.985 1046.935 11673.265 10000 ;
      RECT 11671.865 1046.935 11672.145 10000 ;
      RECT 11669.625 1046.935 11669.905 10000 ;
      RECT 11668.505 1046.935 11668.785 10000 ;
      RECT 11667.385 1046.935 11667.665 10000 ;
      RECT 11652.965 1046.435 11660.805 10000 ;
      RECT 11651.705 1046.935 11651.985 10000 ;
      RECT 11650.585 1046.935 11650.865 10000 ;
      RECT 11649.465 1046.935 11649.745 10000 ;
      RECT 11642.465 1046.935 11644.565 10000 ;
      RECT 11642.605 1046.435 11644.565 10000 ;
      RECT 11641.345 1046.935 11641.625 10000 ;
      RECT 11613.205 1046.435 11638.125 10000 ;
      RECT 11607.465 1046.935 11607.745 10000 ;
      RECT 11606.345 1046.935 11606.625 10000 ;
      RECT 11604.105 1046.935 11604.385 10000 ;
      RECT 11602.985 1046.935 11603.265 10000 ;
      RECT 11601.865 1046.935 11602.145 10000 ;
      RECT 11586.885 1046.435 11599.205 10000 ;
      RECT 11581.705 1046.935 11581.985 10000 ;
      RECT 11580.585 1046.935 11580.865 10000 ;
      RECT 11579.465 1046.935 11579.745 10000 ;
      RECT 11574.425 1046.935 11574.705 10000 ;
      RECT 11534.805 1046.935 11573.585 10000 ;
      RECT 11526.265 1046.935 11526.545 10000 ;
      RECT 11525.145 1046.935 11525.425 10000 ;
      RECT 11522.905 1046.935 11523.185 10000 ;
      RECT 11521.785 1046.935 11522.065 10000 ;
      RECT 11512.265 1046.935 11520.805 10000 ;
      RECT 11512.405 1046.435 11520.805 10000 ;
      RECT 11503.165 1046.935 11505.265 10000 ;
      RECT 11501.905 1046.935 11502.185 10000 ;
      RECT 11500.785 1046.935 11501.065 10000 ;
      RECT 11473.765 1046.435 11498.685 10000 ;
      RECT 11470.265 1046.935 11470.545 10000 ;
      RECT 11469.145 1046.935 11469.425 10000 ;
      RECT 11460.745 1046.935 11461.025 10000 ;
      RECT 11446.745 1046.935 11459.765 10000 ;
      RECT 11446.885 1046.435 11459.765 10000 ;
      RECT 11444.505 1046.935 11444.785 10000 ;
      RECT 11443.385 1046.935 11443.665 10000 ;
      RECT 11442.265 1046.935 11442.545 10000 ;
      RECT 11434.985 1046.935 11435.265 10000 ;
      RECT 11394.805 1046.935 11434.145 10000 ;
      RECT 11393.545 1046.935 11393.825 10000 ;
      RECT 11388.505 1046.935 11388.785 10000 ;
      RECT 11387.385 1046.935 11387.665 10000 ;
      RECT 11372.965 1046.435 11380.805 10000 ;
      RECT 11370.585 1046.935 11370.865 10000 ;
      RECT 11369.465 1046.935 11369.745 10000 ;
      RECT 11367.225 1046.935 11367.505 10000 ;
      RECT 11366.105 1046.935 11366.385 10000 ;
      RECT 11363.165 1046.935 11365.265 10000 ;
      RECT 11333.765 1046.435 11358.685 10000 ;
      RECT 11330.265 1046.935 11330.545 10000 ;
      RECT 11329.145 1046.935 11329.425 10000 ;
      RECT 11328.025 1046.935 11328.305 10000 ;
      RECT 11322.985 1046.935 11323.265 10000 ;
      RECT 11321.865 1046.935 11322.145 10000 ;
      RECT 11307.445 1046.435 11319.765 10000 ;
      RECT 11300.585 1046.935 11300.865 10000 ;
      RECT 11299.465 1046.935 11299.745 10000 ;
      RECT 11297.225 1046.935 11297.505 10000 ;
      RECT 11296.105 1046.935 11296.385 10000 ;
      RECT 11294.985 1046.935 11295.265 10000 ;
      RECT 11254.245 1046.435 11293.445 10000 ;
      RECT 11247.945 1046.935 11248.225 10000 ;
      RECT 11246.825 1046.935 11247.105 10000 ;
      RECT 11245.705 1046.935 11245.985 10000 ;
      RECT 11232.265 1046.935 11240.805 10000 ;
      RECT 11232.405 1046.435 11240.805 10000 ;
      RECT 11231.145 1046.935 11231.425 10000 ;
      RECT 11223.165 1046.435 11224.565 10000 ;
      RECT 11220.785 1046.935 11221.065 10000 ;
      RECT 11219.665 1046.935 11219.945 10000 ;
      RECT 11192.645 1046.435 11218.125 10000 ;
      RECT 11191.385 1046.935 11191.665 10000 ;
      RECT 11190.265 1046.935 11190.545 10000 ;
      RECT 11189.145 1046.935 11189.425 10000 ;
      RECT 11181.865 1046.935 11182.145 10000 ;
      RECT 11180.745 1046.935 11181.025 10000 ;
      RECT 11166.185 1046.935 11179.765 10000 ;
      RECT 11166.325 1046.435 11179.765 10000 ;
      RECT 11161.145 1046.935 11161.425 10000 ;
      RECT 11160.025 1046.935 11160.305 10000 ;
      RECT 11115.365 1046.435 11153.445 10000 ;
      RECT 11112.985 1046.935 11113.265 10000 ;
      RECT 11111.865 1046.935 11112.145 10000 ;
      RECT 11109.625 1046.935 11109.905 10000 ;
      RECT 11108.505 1046.935 11108.785 10000 ;
      RECT 11107.385 1046.935 11107.665 10000 ;
      RECT 11092.965 1046.435 11100.805 10000 ;
      RECT 11091.705 1046.935 11091.985 10000 ;
      RECT 11090.585 1046.935 11090.865 10000 ;
      RECT 11089.465 1046.935 11089.745 10000 ;
      RECT 11082.465 1046.935 11084.565 10000 ;
      RECT 11082.605 1046.435 11084.565 10000 ;
      RECT 11081.345 1046.935 11081.625 10000 ;
      RECT 11053.205 1046.435 11078.125 10000 ;
      RECT 11047.465 1046.935 11047.745 10000 ;
      RECT 11046.345 1046.935 11046.625 10000 ;
      RECT 11044.105 1046.935 11044.385 10000 ;
      RECT 11042.985 1046.935 11043.265 10000 ;
      RECT 11041.865 1046.935 11042.145 10000 ;
      RECT 11026.885 1046.435 11039.205 10000 ;
      RECT 11021.705 1046.935 11021.985 10000 ;
      RECT 11020.585 1046.935 11020.865 10000 ;
      RECT 11019.465 1046.935 11019.745 10000 ;
      RECT 11014.425 1046.935 11014.705 10000 ;
      RECT 10974.805 1046.935 11013.585 10000 ;
      RECT 10966.265 1046.935 10966.545 10000 ;
      RECT 10965.145 1046.935 10965.425 10000 ;
      RECT 10962.905 1046.935 10963.185 10000 ;
      RECT 10961.785 1046.935 10962.065 10000 ;
      RECT 10952.265 1046.935 10960.805 10000 ;
      RECT 10952.405 1046.435 10960.805 10000 ;
      RECT 10943.165 1046.935 10945.265 10000 ;
      RECT 10941.905 1046.935 10942.185 10000 ;
      RECT 10940.785 1046.935 10941.065 10000 ;
      RECT 10913.765 1046.435 10938.685 10000 ;
      RECT 10910.265 1046.935 10910.545 10000 ;
      RECT 10909.145 1046.935 10909.425 10000 ;
      RECT 10900.745 1046.935 10901.025 10000 ;
      RECT 10886.745 1046.935 10899.765 10000 ;
      RECT 10886.885 1046.435 10899.765 10000 ;
      RECT 10884.505 1046.935 10884.785 10000 ;
      RECT 10883.385 1046.935 10883.665 10000 ;
      RECT 10882.265 1046.935 10882.545 10000 ;
      RECT 10874.985 1046.935 10875.265 10000 ;
      RECT 10834.805 1046.935 10874.145 10000 ;
      RECT 10833.545 1046.935 10833.825 10000 ;
      RECT 10828.505 1046.935 10828.785 10000 ;
      RECT 10827.385 1046.935 10827.665 10000 ;
      RECT 10812.965 1046.435 10820.805 10000 ;
      RECT 10810.585 1046.935 10810.865 10000 ;
      RECT 10809.465 1046.935 10809.745 10000 ;
      RECT 10807.225 1046.935 10807.505 10000 ;
      RECT 10806.105 1046.935 10806.385 10000 ;
      RECT 10803.165 1046.935 10805.265 10000 ;
      RECT 10773.765 1046.435 10798.685 10000 ;
      RECT 10770.265 1046.935 10770.545 10000 ;
      RECT 10769.145 1046.935 10769.425 10000 ;
      RECT 10768.025 1046.935 10768.305 10000 ;
      RECT 10762.985 1046.935 10763.265 10000 ;
      RECT 10761.865 1046.935 10762.145 10000 ;
      RECT 10747.445 1046.435 10759.765 10000 ;
      RECT 10740.585 1046.935 10740.865 10000 ;
      RECT 10739.465 1046.935 10739.745 10000 ;
      RECT 10737.225 1046.935 10737.505 10000 ;
      RECT 10736.105 1046.935 10736.385 10000 ;
      RECT 10734.985 1046.935 10735.265 10000 ;
      RECT 10694.245 1046.435 10733.445 10000 ;
      RECT 10687.945 1046.935 10688.225 10000 ;
      RECT 10686.825 1046.935 10687.105 10000 ;
      RECT 10685.705 1046.935 10685.985 10000 ;
      RECT 10672.265 1046.935 10680.805 10000 ;
      RECT 10672.405 1046.435 10680.805 10000 ;
      RECT 10671.145 1046.935 10671.425 10000 ;
      RECT 10663.165 1046.435 10664.565 10000 ;
      RECT 10660.785 1046.935 10661.065 10000 ;
      RECT 10659.665 1046.935 10659.945 10000 ;
      RECT 10632.645 1046.435 10658.125 10000 ;
      RECT 10631.385 1046.935 10631.665 10000 ;
      RECT 10630.265 1046.935 10630.545 10000 ;
      RECT 10629.145 1046.935 10629.425 10000 ;
      RECT 10621.865 1046.935 10622.145 10000 ;
      RECT 10620.745 1046.935 10621.025 10000 ;
      RECT 10606.185 1046.935 10619.765 10000 ;
      RECT 10606.325 1046.435 10619.765 10000 ;
      RECT 10601.145 1046.935 10601.425 10000 ;
      RECT 10600.025 1046.935 10600.305 10000 ;
      RECT 10555.365 1046.435 10593.445 10000 ;
      RECT 10552.985 1046.935 10553.265 10000 ;
      RECT 10551.865 1046.935 10552.145 10000 ;
      RECT 10549.625 1046.935 10549.905 10000 ;
      RECT 10548.505 1046.935 10548.785 10000 ;
      RECT 10547.385 1046.935 10547.665 10000 ;
      RECT 10532.965 1046.435 10540.805 10000 ;
      RECT 10531.705 1046.935 10531.985 10000 ;
      RECT 10530.585 1046.935 10530.865 10000 ;
      RECT 10529.465 1046.935 10529.745 10000 ;
      RECT 10522.465 1046.935 10524.565 10000 ;
      RECT 10522.605 1046.435 10524.565 10000 ;
      RECT 10521.345 1046.935 10521.625 10000 ;
      RECT 10493.205 1046.435 10518.125 10000 ;
      RECT 10487.465 1046.935 10487.745 10000 ;
      RECT 10486.345 1046.935 10486.625 10000 ;
      RECT 10484.105 1046.935 10484.385 10000 ;
      RECT 10482.985 1046.935 10483.265 10000 ;
      RECT 10481.865 1046.935 10482.145 10000 ;
      RECT 10466.885 1046.435 10479.205 10000 ;
      RECT 10461.705 1046.935 10461.985 10000 ;
      RECT 10460.585 1046.935 10460.865 10000 ;
      RECT 10459.465 1046.935 10459.745 10000 ;
      RECT 10454.425 1046.935 10454.705 10000 ;
      RECT 10414.805 1046.935 10453.585 10000 ;
      RECT 10406.265 1046.935 10406.545 10000 ;
      RECT 10405.145 1046.935 10405.425 10000 ;
      RECT 10402.905 1046.935 10403.185 10000 ;
      RECT 10401.785 1046.935 10402.065 10000 ;
      RECT 10392.265 1046.935 10400.805 10000 ;
      RECT 10392.405 1046.435 10400.805 10000 ;
      RECT 10383.165 1046.935 10385.265 10000 ;
      RECT 10381.905 1046.935 10382.185 10000 ;
      RECT 10380.785 1046.935 10381.065 10000 ;
      RECT 10353.765 1046.435 10378.685 10000 ;
      RECT 10350.265 1046.935 10350.545 10000 ;
      RECT 10349.145 1046.935 10349.425 10000 ;
      RECT 10340.745 1046.935 10341.025 10000 ;
      RECT 10326.745 1046.935 10339.765 10000 ;
      RECT 10326.885 1046.435 10339.765 10000 ;
      RECT 10324.505 1046.935 10324.785 10000 ;
      RECT 10323.385 1046.935 10323.665 10000 ;
      RECT 10322.265 1046.935 10322.545 10000 ;
      RECT 10314.985 1046.935 10315.265 10000 ;
      RECT 10274.805 1046.935 10314.145 10000 ;
      RECT 10273.545 1046.935 10273.825 10000 ;
      RECT 10268.505 1046.935 10268.785 10000 ;
      RECT 10267.385 1046.935 10267.665 10000 ;
      RECT 10252.965 1046.435 10260.805 10000 ;
      RECT 10250.585 1046.935 10250.865 10000 ;
      RECT 10249.465 1046.935 10249.745 10000 ;
      RECT 10247.225 1046.935 10247.505 10000 ;
      RECT 10246.105 1046.935 10246.385 10000 ;
      RECT 10243.165 1046.935 10245.265 10000 ;
      RECT 10213.765 1046.435 10238.685 10000 ;
      RECT 10210.265 1046.935 10210.545 10000 ;
      RECT 10209.145 1046.935 10209.425 10000 ;
      RECT 10208.025 1046.935 10208.305 10000 ;
      RECT 10202.985 1046.935 10203.265 10000 ;
      RECT 10201.865 1046.935 10202.145 10000 ;
      RECT 10187.445 1046.435 10199.765 10000 ;
      RECT 10180.585 1046.935 10180.865 10000 ;
      RECT 10179.465 1046.935 10179.745 10000 ;
      RECT 10177.225 1046.935 10177.505 10000 ;
      RECT 10176.105 1046.935 10176.385 10000 ;
      RECT 10174.985 1046.935 10175.265 10000 ;
      RECT 10134.245 1046.435 10173.445 10000 ;
      RECT 10127.945 1046.935 10128.225 10000 ;
      RECT 10126.825 1046.935 10127.105 10000 ;
      RECT 10125.705 1046.935 10125.985 10000 ;
      RECT 10112.265 1046.935 10120.805 10000 ;
      RECT 10112.405 1046.435 10120.805 10000 ;
      RECT 10111.145 1046.935 10111.425 10000 ;
      RECT 10103.165 1046.435 10104.565 10000 ;
      RECT 10100.785 1046.935 10101.065 10000 ;
      RECT 10099.665 1046.935 10099.945 10000 ;
      RECT 10072.645 1046.435 10098.125 10000 ;
      RECT 10071.385 1046.935 10071.665 10000 ;
      RECT 10070.265 1046.935 10070.545 10000 ;
      RECT 10069.145 1046.935 10069.425 10000 ;
      RECT 10061.865 1046.935 10062.145 10000 ;
      RECT 10060.745 1046.935 10061.025 10000 ;
      RECT 10046.185 1046.935 10059.765 10000 ;
      RECT 10046.325 1046.435 10059.765 10000 ;
      RECT 10041.145 1046.935 10041.425 10000 ;
      RECT 10040.025 1046.935 10040.305 10000 ;
      RECT 9995.365 1046.435 10033.445 10000 ;
      RECT 9992.985 1046.935 9993.265 10000 ;
      RECT 9991.865 1046.935 9992.145 10000 ;
      RECT 9989.625 1046.935 9989.905 10000 ;
      RECT 9988.505 1046.935 9988.785 10000 ;
      RECT 9987.385 1046.935 9987.665 10000 ;
      RECT 9972.965 1046.435 9980.805 10000 ;
      RECT 9971.705 1046.935 9971.985 10000 ;
      RECT 9970.585 1046.935 9970.865 10000 ;
      RECT 9969.465 1046.935 9969.745 10000 ;
      RECT 9962.465 1046.935 9964.565 10000 ;
      RECT 9962.605 1046.435 9964.565 10000 ;
      RECT 9961.345 1046.935 9961.625 10000 ;
      RECT 9933.205 1046.435 9958.125 10000 ;
      RECT 9927.465 1046.935 9927.745 10000 ;
      RECT 9926.345 1046.935 9926.625 10000 ;
      RECT 9924.105 1046.935 9924.385 10000 ;
      RECT 9922.985 1046.935 9923.265 10000 ;
      RECT 9921.865 1046.935 9922.145 10000 ;
      RECT 9906.885 1046.435 9919.205 10000 ;
      RECT 9901.705 1046.935 9901.985 10000 ;
      RECT 9900.585 1046.935 9900.865 10000 ;
      RECT 9899.465 1046.935 9899.745 10000 ;
      RECT 9894.425 1046.935 9894.705 10000 ;
      RECT 9854.805 1046.935 9893.585 10000 ;
      RECT 9846.265 1046.935 9846.545 10000 ;
      RECT 9845.145 1046.935 9845.425 10000 ;
      RECT 9842.905 1046.935 9843.185 10000 ;
      RECT 9841.785 1046.935 9842.065 10000 ;
      RECT 9832.265 1046.935 9840.805 10000 ;
      RECT 9832.405 1046.435 9840.805 10000 ;
      RECT 9823.165 1046.935 9825.265 10000 ;
      RECT 9821.905 1046.935 9822.185 10000 ;
      RECT 9820.785 1046.935 9821.065 10000 ;
      RECT 9793.765 1046.435 9818.685 10000 ;
      RECT 9790.265 1046.935 9790.545 10000 ;
      RECT 9789.145 1046.935 9789.425 10000 ;
      RECT 9780.745 1046.935 9781.025 10000 ;
      RECT 9766.745 1046.935 9779.765 10000 ;
      RECT 9766.885 1046.435 9779.765 10000 ;
      RECT 9764.505 1046.935 9764.785 10000 ;
      RECT 9763.385 1046.935 9763.665 10000 ;
      RECT 9762.265 1046.935 9762.545 10000 ;
      RECT 9754.985 1046.935 9755.265 10000 ;
      RECT 9714.805 1046.935 9754.145 10000 ;
      RECT 9713.545 1046.935 9713.825 10000 ;
      RECT 9708.505 1046.935 9708.785 10000 ;
      RECT 9707.385 1046.935 9707.665 10000 ;
      RECT 9692.965 1046.435 9700.805 10000 ;
      RECT 9690.585 1046.935 9690.865 10000 ;
      RECT 9689.465 1046.935 9689.745 10000 ;
      RECT 9687.225 1046.935 9687.505 10000 ;
      RECT 9686.105 1046.935 9686.385 10000 ;
      RECT 9683.165 1046.935 9685.265 10000 ;
      RECT 9653.765 1046.435 9678.685 10000 ;
      RECT 9650.265 1046.935 9650.545 10000 ;
      RECT 9649.145 1046.935 9649.425 10000 ;
      RECT 9648.025 1046.935 9648.305 10000 ;
      RECT 9642.985 1046.935 9643.265 10000 ;
      RECT 9641.865 1046.935 9642.145 10000 ;
      RECT 9627.445 1046.435 9639.765 10000 ;
      RECT 9620.585 1046.935 9620.865 10000 ;
      RECT 9619.465 1046.935 9619.745 10000 ;
      RECT 9617.225 1046.935 9617.505 10000 ;
      RECT 9616.105 1046.935 9616.385 10000 ;
      RECT 9614.985 1046.935 9615.265 10000 ;
      RECT 9574.245 1046.435 9613.445 10000 ;
      RECT 9567.945 1046.935 9568.225 10000 ;
      RECT 9566.825 1046.935 9567.105 10000 ;
      RECT 9565.705 1046.935 9565.985 10000 ;
      RECT 9552.265 1046.935 9560.805 10000 ;
      RECT 9552.405 1046.435 9560.805 10000 ;
      RECT 9551.145 1046.935 9551.425 10000 ;
      RECT 9543.165 1046.435 9544.565 10000 ;
      RECT 9540.785 1046.935 9541.065 10000 ;
      RECT 9539.665 1046.935 9539.945 10000 ;
      RECT 9512.645 1046.435 9538.125 10000 ;
      RECT 9511.385 1046.935 9511.665 10000 ;
      RECT 9510.265 1046.935 9510.545 10000 ;
      RECT 9509.145 1046.935 9509.425 10000 ;
      RECT 9501.865 1046.935 9502.145 10000 ;
      RECT 9500.745 1046.935 9501.025 10000 ;
      RECT 9486.185 1046.935 9499.765 10000 ;
      RECT 9486.325 1046.435 9499.765 10000 ;
      RECT 9481.145 1046.935 9481.425 10000 ;
      RECT 9480.025 1046.935 9480.305 10000 ;
      RECT 9435.365 1046.435 9473.445 10000 ;
      RECT 9432.985 1046.935 9433.265 10000 ;
      RECT 9431.865 1046.935 9432.145 10000 ;
      RECT 9429.625 1046.935 9429.905 10000 ;
      RECT 9428.505 1046.935 9428.785 10000 ;
      RECT 9427.385 1046.935 9427.665 10000 ;
      RECT 9412.965 1046.435 9420.805 10000 ;
      RECT 9411.705 1046.935 9411.985 10000 ;
      RECT 9410.585 1046.935 9410.865 10000 ;
      RECT 9409.465 1046.935 9409.745 10000 ;
      RECT 9402.465 1046.935 9404.565 10000 ;
      RECT 9402.605 1046.435 9404.565 10000 ;
      RECT 9401.345 1046.935 9401.625 10000 ;
      RECT 9373.205 1046.435 9398.125 10000 ;
      RECT 9367.465 1046.935 9367.745 10000 ;
      RECT 9366.345 1046.935 9366.625 10000 ;
      RECT 9364.105 1046.935 9364.385 10000 ;
      RECT 9362.985 1046.935 9363.265 10000 ;
      RECT 9361.865 1046.935 9362.145 10000 ;
      RECT 9346.885 1046.435 9359.205 10000 ;
      RECT 9341.705 1046.935 9341.985 10000 ;
      RECT 9340.585 1046.935 9340.865 10000 ;
      RECT 9339.465 1046.935 9339.745 10000 ;
      RECT 9334.425 1046.935 9334.705 10000 ;
      RECT 9294.805 1046.935 9333.585 10000 ;
      RECT 9286.265 1046.935 9286.545 10000 ;
      RECT 9285.145 1046.935 9285.425 10000 ;
      RECT 9282.905 1046.935 9283.185 10000 ;
      RECT 9281.785 1046.935 9282.065 10000 ;
      RECT 9272.265 1046.935 9280.805 10000 ;
      RECT 9272.405 1046.435 9280.805 10000 ;
      RECT 9263.165 1046.935 9265.265 10000 ;
      RECT 9261.905 1046.935 9262.185 10000 ;
      RECT 9260.785 1046.935 9261.065 10000 ;
      RECT 9233.765 1046.435 9258.685 10000 ;
      RECT 9230.265 1046.935 9230.545 10000 ;
      RECT 9229.145 1046.935 9229.425 10000 ;
      RECT 9220.745 1046.935 9221.025 10000 ;
      RECT 9206.745 1046.935 9219.765 10000 ;
      RECT 9206.885 1046.435 9219.765 10000 ;
      RECT 9204.505 1046.935 9204.785 10000 ;
      RECT 9203.385 1046.935 9203.665 10000 ;
      RECT 9202.265 1046.935 9202.545 10000 ;
      RECT 9194.985 1046.935 9195.265 10000 ;
      RECT 9154.805 1046.935 9194.145 10000 ;
      RECT 9153.545 1046.935 9153.825 10000 ;
      RECT 9148.505 1046.935 9148.785 10000 ;
      RECT 9147.385 1046.935 9147.665 10000 ;
      RECT 9132.965 1046.435 9140.805 10000 ;
      RECT 9130.585 1046.935 9130.865 10000 ;
      RECT 9129.465 1046.935 9129.745 10000 ;
      RECT 9127.225 1046.935 9127.505 10000 ;
      RECT 9126.105 1046.935 9126.385 10000 ;
      RECT 9123.165 1046.935 9125.265 10000 ;
      RECT 9093.765 1046.435 9118.685 10000 ;
      RECT 9090.265 1046.935 9090.545 10000 ;
      RECT 9089.145 1046.935 9089.425 10000 ;
      RECT 9088.025 1046.935 9088.305 10000 ;
      RECT 9082.985 1046.935 9083.265 10000 ;
      RECT 9081.865 1046.935 9082.145 10000 ;
      RECT 9067.445 1046.435 9079.765 10000 ;
      RECT 9060.585 1046.935 9060.865 10000 ;
      RECT 9059.465 1046.935 9059.745 10000 ;
      RECT 9057.225 1046.935 9057.505 10000 ;
      RECT 9056.105 1046.935 9056.385 10000 ;
      RECT 9054.985 1046.935 9055.265 10000 ;
      RECT 9014.245 1046.435 9053.445 10000 ;
      RECT 9007.945 1046.935 9008.225 10000 ;
      RECT 9006.825 1046.935 9007.105 10000 ;
      RECT 9005.705 1046.935 9005.985 10000 ;
      RECT 8992.265 1046.935 9000.805 10000 ;
      RECT 8992.405 1046.435 9000.805 10000 ;
      RECT 8991.145 1046.935 8991.425 10000 ;
      RECT 8983.165 1046.435 8984.565 10000 ;
      RECT 8980.785 1046.935 8981.065 10000 ;
      RECT 8979.665 1046.935 8979.945 10000 ;
      RECT 8952.645 1046.435 8978.125 10000 ;
      RECT 8951.385 1046.935 8951.665 10000 ;
      RECT 8950.265 1046.935 8950.545 10000 ;
      RECT 8949.145 1046.935 8949.425 10000 ;
      RECT 8941.865 1046.935 8942.145 10000 ;
      RECT 8940.745 1046.935 8941.025 10000 ;
      RECT 8926.185 1046.935 8939.765 10000 ;
      RECT 8926.325 1046.435 8939.765 10000 ;
      RECT 8921.145 1046.935 8921.425 10000 ;
      RECT 8920.025 1046.935 8920.305 10000 ;
      RECT 8875.365 1046.435 8913.445 10000 ;
      RECT 8872.985 1046.935 8873.265 10000 ;
      RECT 8871.865 1046.935 8872.145 10000 ;
      RECT 8869.625 1046.935 8869.905 10000 ;
      RECT 8868.505 1046.935 8868.785 10000 ;
      RECT 8867.385 1046.935 8867.665 10000 ;
      RECT 8852.965 1046.435 8860.805 10000 ;
      RECT 8851.705 1046.935 8851.985 10000 ;
      RECT 8850.585 1046.935 8850.865 10000 ;
      RECT 8849.465 1046.935 8849.745 10000 ;
      RECT 8842.465 1046.935 8844.565 10000 ;
      RECT 8842.605 1046.435 8844.565 10000 ;
      RECT 8841.345 1046.935 8841.625 10000 ;
      RECT 8813.205 1046.435 8838.125 10000 ;
      RECT 8807.465 1046.935 8807.745 10000 ;
      RECT 8806.345 1046.935 8806.625 10000 ;
      RECT 8804.105 1046.935 8804.385 10000 ;
      RECT 8802.985 1046.935 8803.265 10000 ;
      RECT 8801.865 1046.935 8802.145 10000 ;
      RECT 8786.885 1046.435 8799.205 10000 ;
      RECT 8781.705 1046.935 8781.985 10000 ;
      RECT 8780.585 1046.935 8780.865 10000 ;
      RECT 8779.465 1046.935 8779.745 10000 ;
      RECT 8774.425 1046.935 8774.705 10000 ;
      RECT 8734.805 1046.935 8773.585 10000 ;
      RECT 8726.265 1046.935 8726.545 10000 ;
      RECT 8725.145 1046.935 8725.425 10000 ;
      RECT 8722.905 1046.935 8723.185 10000 ;
      RECT 8721.785 1046.935 8722.065 10000 ;
      RECT 8712.265 1046.935 8720.805 10000 ;
      RECT 8712.405 1046.435 8720.805 10000 ;
      RECT 8703.165 1046.935 8705.265 10000 ;
      RECT 8701.905 1046.935 8702.185 10000 ;
      RECT 8700.785 1046.935 8701.065 10000 ;
      RECT 8673.765 1046.435 8698.685 10000 ;
      RECT 8670.265 1046.935 8670.545 10000 ;
      RECT 8669.145 1046.935 8669.425 10000 ;
      RECT 8660.745 1046.935 8661.025 10000 ;
      RECT 8646.745 1046.935 8659.765 10000 ;
      RECT 8646.885 1046.435 8659.765 10000 ;
      RECT 8644.505 1046.935 8644.785 10000 ;
      RECT 8643.385 1046.935 8643.665 10000 ;
      RECT 8642.265 1046.935 8642.545 10000 ;
      RECT 8634.985 1046.935 8635.265 10000 ;
      RECT 8594.805 1046.935 8634.145 10000 ;
      RECT 8593.545 1046.935 8593.825 10000 ;
      RECT 8588.505 1046.935 8588.785 10000 ;
      RECT 8587.385 1046.935 8587.665 10000 ;
      RECT 8572.965 1046.435 8580.805 10000 ;
      RECT 8570.585 1046.935 8570.865 10000 ;
      RECT 8569.465 1046.935 8569.745 10000 ;
      RECT 8567.225 1046.935 8567.505 10000 ;
      RECT 8566.105 1046.935 8566.385 10000 ;
      RECT 8563.165 1046.935 8565.265 10000 ;
      RECT 8533.765 1046.435 8558.685 10000 ;
      RECT 8530.265 1046.935 8530.545 10000 ;
      RECT 8529.145 1046.935 8529.425 10000 ;
      RECT 8528.025 1046.935 8528.305 10000 ;
      RECT 8522.985 1046.935 8523.265 10000 ;
      RECT 8521.865 1046.935 8522.145 10000 ;
      RECT 8507.445 1046.435 8519.765 10000 ;
      RECT 8500.585 1046.935 8500.865 10000 ;
      RECT 8499.465 1046.935 8499.745 10000 ;
      RECT 8497.225 1046.935 8497.505 10000 ;
      RECT 8496.105 1046.935 8496.385 10000 ;
      RECT 8494.985 1046.935 8495.265 10000 ;
      RECT 8454.245 1046.435 8493.445 10000 ;
      RECT 8447.945 1046.935 8448.225 10000 ;
      RECT 8446.825 1046.935 8447.105 10000 ;
      RECT 8445.705 1046.935 8445.985 10000 ;
      RECT 8432.265 1046.935 8440.805 10000 ;
      RECT 8432.405 1046.435 8440.805 10000 ;
      RECT 8431.145 1046.935 8431.425 10000 ;
      RECT 8423.165 1046.435 8424.565 10000 ;
      RECT 8420.785 1046.935 8421.065 10000 ;
      RECT 8419.665 1046.935 8419.945 10000 ;
      RECT 8392.645 1046.435 8418.125 10000 ;
      RECT 8391.385 1046.935 8391.665 10000 ;
      RECT 8390.265 1046.935 8390.545 10000 ;
      RECT 8389.145 1046.935 8389.425 10000 ;
      RECT 8381.865 1046.935 8382.145 10000 ;
      RECT 8380.745 1046.935 8381.025 10000 ;
      RECT 8366.185 1046.935 8379.765 10000 ;
      RECT 8366.325 1046.435 8379.765 10000 ;
      RECT 8361.145 1046.935 8361.425 10000 ;
      RECT 8360.025 1046.935 8360.305 10000 ;
      RECT 8315.365 1046.435 8353.445 10000 ;
      RECT 8312.985 1046.935 8313.265 10000 ;
      RECT 8311.865 1046.935 8312.145 10000 ;
      RECT 8309.625 1046.935 8309.905 10000 ;
      RECT 8308.505 1046.935 8308.785 10000 ;
      RECT 8307.385 1046.935 8307.665 10000 ;
      RECT 8292.965 1046.435 8300.805 10000 ;
      RECT 8291.705 1046.935 8291.985 10000 ;
      RECT 8290.585 1046.935 8290.865 10000 ;
      RECT 8289.465 1046.935 8289.745 10000 ;
      RECT 8282.465 1046.935 8284.565 10000 ;
      RECT 8282.605 1046.435 8284.565 10000 ;
      RECT 8281.345 1046.935 8281.625 10000 ;
      RECT 8253.205 1046.435 8278.125 10000 ;
      RECT 8247.465 1046.935 8247.745 10000 ;
      RECT 8246.345 1046.935 8246.625 10000 ;
      RECT 8244.105 1046.935 8244.385 10000 ;
      RECT 8242.985 1046.935 8243.265 10000 ;
      RECT 8241.865 1046.935 8242.145 10000 ;
      RECT 8226.885 1046.435 8239.205 10000 ;
      RECT 8221.705 1046.935 8221.985 10000 ;
      RECT 8220.585 1046.935 8220.865 10000 ;
      RECT 8219.465 1046.935 8219.745 10000 ;
      RECT 8214.425 1046.935 8214.705 10000 ;
      RECT 8174.805 1046.935 8213.585 10000 ;
      RECT 8166.265 1046.935 8166.545 10000 ;
      RECT 8165.145 1046.935 8165.425 10000 ;
      RECT 8162.905 1046.935 8163.185 10000 ;
      RECT 8161.785 1046.935 8162.065 10000 ;
      RECT 8152.265 1046.935 8160.805 10000 ;
      RECT 8152.405 1046.435 8160.805 10000 ;
      RECT 8143.165 1046.935 8145.265 10000 ;
      RECT 8141.905 1046.935 8142.185 10000 ;
      RECT 8140.785 1046.935 8141.065 10000 ;
      RECT 8113.765 1046.435 8138.685 10000 ;
      RECT 8110.265 1046.935 8110.545 10000 ;
      RECT 8109.145 1046.935 8109.425 10000 ;
      RECT 8100.745 1046.935 8101.025 10000 ;
      RECT 8086.745 1046.935 8099.765 10000 ;
      RECT 8086.885 1046.435 8099.765 10000 ;
      RECT 8084.505 1046.935 8084.785 10000 ;
      RECT 8083.385 1046.935 8083.665 10000 ;
      RECT 8082.265 1046.935 8082.545 10000 ;
      RECT 8074.985 1046.935 8075.265 10000 ;
      RECT 8034.805 1046.935 8074.145 10000 ;
      RECT 8033.545 1046.935 8033.825 10000 ;
      RECT 8028.505 1046.935 8028.785 10000 ;
      RECT 8027.385 1046.935 8027.665 10000 ;
      RECT 8012.965 1046.435 8020.805 10000 ;
      RECT 8010.585 1046.935 8010.865 10000 ;
      RECT 8009.465 1046.935 8009.745 10000 ;
      RECT 8007.225 1046.935 8007.505 10000 ;
      RECT 8006.105 1046.935 8006.385 10000 ;
      RECT 8003.165 1046.935 8005.265 10000 ;
      RECT 7973.765 1046.435 7998.685 10000 ;
      RECT 7970.265 1046.935 7970.545 10000 ;
      RECT 7969.145 1046.935 7969.425 10000 ;
      RECT 7968.025 1046.935 7968.305 10000 ;
      RECT 7962.985 1046.935 7963.265 10000 ;
      RECT 7961.865 1046.935 7962.145 10000 ;
      RECT 7947.445 1046.435 7959.765 10000 ;
      RECT 7940.585 1046.935 7940.865 10000 ;
      RECT 7939.465 1046.935 7939.745 10000 ;
      RECT 7937.225 1046.935 7937.505 10000 ;
      RECT 7936.105 1046.935 7936.385 10000 ;
      RECT 7934.985 1046.935 7935.265 10000 ;
      RECT 7894.245 1046.435 7933.445 10000 ;
      RECT 7887.945 1046.935 7888.225 10000 ;
      RECT 7886.825 1046.935 7887.105 10000 ;
      RECT 7885.705 1046.935 7885.985 10000 ;
      RECT 7872.265 1046.935 7880.805 10000 ;
      RECT 7872.405 1046.435 7880.805 10000 ;
      RECT 7871.145 1046.935 7871.425 10000 ;
      RECT 7863.165 1046.435 7864.565 10000 ;
      RECT 7860.785 1046.935 7861.065 10000 ;
      RECT 7859.665 1046.935 7859.945 10000 ;
      RECT 7832.645 1046.435 7858.125 10000 ;
      RECT 7831.385 1046.935 7831.665 10000 ;
      RECT 7830.265 1046.935 7830.545 10000 ;
      RECT 7829.145 1046.935 7829.425 10000 ;
      RECT 7821.865 1046.935 7822.145 10000 ;
      RECT 7820.745 1046.935 7821.025 10000 ;
      RECT 7806.185 1046.935 7819.765 10000 ;
      RECT 7806.325 1046.435 7819.765 10000 ;
      RECT 7801.145 1046.935 7801.425 10000 ;
      RECT 7800.025 1046.935 7800.305 10000 ;
      RECT 7755.365 1046.435 7793.445 10000 ;
      RECT 7752.985 1046.935 7753.265 10000 ;
      RECT 7751.865 1046.935 7752.145 10000 ;
      RECT 7749.625 1046.935 7749.905 10000 ;
      RECT 7748.505 1046.935 7748.785 10000 ;
      RECT 7747.385 1046.935 7747.665 10000 ;
      RECT 7732.965 1046.435 7740.805 10000 ;
      RECT 7731.705 1046.935 7731.985 10000 ;
      RECT 7730.585 1046.935 7730.865 10000 ;
      RECT 7729.465 1046.935 7729.745 10000 ;
      RECT 7722.465 1046.935 7724.565 10000 ;
      RECT 7722.605 1046.435 7724.565 10000 ;
      RECT 7721.345 1046.935 7721.625 10000 ;
      RECT 7693.205 1046.435 7718.125 10000 ;
      RECT 7687.465 1046.935 7687.745 10000 ;
      RECT 7686.345 1046.935 7686.625 10000 ;
      RECT 7684.105 1046.935 7684.385 10000 ;
      RECT 7682.985 1046.935 7683.265 10000 ;
      RECT 14163.165 1046.435 14165.125 10000 ;
      RECT 13774.805 1046.435 13813.445 10000 ;
      RECT 13743.165 1046.435 13745.125 10000 ;
      RECT 13634.805 1046.435 13674.005 10000 ;
      RECT 13603.165 1046.435 13605.125 10000 ;
      RECT 13214.805 1046.435 13253.445 10000 ;
      RECT 13183.165 1046.435 13185.125 10000 ;
      RECT 13074.805 1046.435 13114.005 10000 ;
      RECT 13043.165 1046.435 13045.125 10000 ;
      RECT 12654.805 1046.435 12693.445 10000 ;
      RECT 12623.165 1046.435 12625.125 10000 ;
      RECT 12514.805 1046.435 12554.005 10000 ;
      RECT 12483.165 1046.435 12485.125 10000 ;
      RECT 12094.805 1046.435 12133.445 10000 ;
      RECT 12063.165 1046.435 12065.125 10000 ;
      RECT 11954.805 1046.435 11994.005 10000 ;
      RECT 11923.165 1046.435 11925.125 10000 ;
      RECT 11534.805 1046.435 11573.445 10000 ;
      RECT 11503.165 1046.435 11505.125 10000 ;
      RECT 11394.805 1046.435 11434.005 10000 ;
      RECT 11363.165 1046.435 11365.125 10000 ;
      RECT 10974.805 1046.435 11013.445 10000 ;
      RECT 10943.165 1046.435 10945.125 10000 ;
      RECT 10834.805 1046.435 10874.005 10000 ;
      RECT 10803.165 1046.435 10805.125 10000 ;
      RECT 10414.805 1046.435 10453.445 10000 ;
      RECT 10383.165 1046.435 10385.125 10000 ;
      RECT 10274.805 1046.435 10314.005 10000 ;
      RECT 10243.165 1046.435 10245.125 10000 ;
      RECT 9854.805 1046.435 9893.445 10000 ;
      RECT 9823.165 1046.435 9825.125 10000 ;
      RECT 9714.805 1046.435 9754.005 10000 ;
      RECT 9683.165 1046.435 9685.125 10000 ;
      RECT 9294.805 1046.435 9333.445 10000 ;
      RECT 9263.165 1046.435 9265.125 10000 ;
      RECT 9154.805 1046.435 9194.005 10000 ;
      RECT 9123.165 1046.435 9125.125 10000 ;
      RECT 8734.805 1046.435 8773.445 10000 ;
      RECT 8703.165 1046.435 8705.125 10000 ;
      RECT 8594.805 1046.435 8634.005 10000 ;
      RECT 8563.165 1046.435 8565.125 10000 ;
      RECT 8174.805 1046.435 8213.445 10000 ;
      RECT 8143.165 1046.435 8145.125 10000 ;
      RECT 8034.805 1046.435 8074.005 10000 ;
      RECT 8003.165 1046.435 8005.125 10000 ;
      RECT 998.1 1047.855 7682.145 10000 ;
      RECT 7681.865 1046.935 7682.145 10000 ;
      RECT 7666.885 1046.435 7679.205 10000 ;
      RECT 7661.705 1046.935 7661.985 10000 ;
      RECT 7660.585 1046.935 7660.865 10000 ;
      RECT 7659.465 1046.935 7659.745 10000 ;
      RECT 7654.425 1046.935 7654.705 10000 ;
      RECT 7614.805 1046.935 7653.585 10000 ;
      RECT 7606.265 1046.935 7606.545 10000 ;
      RECT 7605.145 1046.935 7605.425 10000 ;
      RECT 7602.905 1046.935 7603.185 10000 ;
      RECT 7601.785 1046.935 7602.065 10000 ;
      RECT 7592.265 1046.935 7600.805 10000 ;
      RECT 7592.405 1046.435 7600.805 10000 ;
      RECT 7583.165 1046.935 7585.265 10000 ;
      RECT 7581.905 1046.935 7582.185 10000 ;
      RECT 7580.785 1046.935 7581.065 10000 ;
      RECT 7553.765 1046.435 7578.685 10000 ;
      RECT 7550.265 1046.935 7550.545 10000 ;
      RECT 7549.145 1046.935 7549.425 10000 ;
      RECT 7540.745 1046.935 7541.025 10000 ;
      RECT 7526.745 1046.935 7539.765 10000 ;
      RECT 7526.885 1046.435 7539.765 10000 ;
      RECT 7524.505 1046.935 7524.785 10000 ;
      RECT 7523.385 1046.935 7523.665 10000 ;
      RECT 7522.265 1046.935 7522.545 10000 ;
      RECT 7514.985 1046.935 7515.265 10000 ;
      RECT 7474.805 1046.935 7514.145 10000 ;
      RECT 7473.545 1046.935 7473.825 10000 ;
      RECT 7468.505 1046.935 7468.785 10000 ;
      RECT 7467.385 1046.935 7467.665 10000 ;
      RECT 7452.965 1046.435 7460.805 10000 ;
      RECT 7450.585 1046.935 7450.865 10000 ;
      RECT 7449.465 1046.935 7449.745 10000 ;
      RECT 7447.225 1046.935 7447.505 10000 ;
      RECT 7446.105 1046.935 7446.385 10000 ;
      RECT 7443.165 1046.935 7445.265 10000 ;
      RECT 7413.765 1046.435 7438.685 10000 ;
      RECT 7410.265 1046.935 7410.545 10000 ;
      RECT 7409.145 1046.935 7409.425 10000 ;
      RECT 7408.025 1046.935 7408.305 10000 ;
      RECT 7402.985 1046.935 7403.265 10000 ;
      RECT 7401.865 1046.935 7402.145 10000 ;
      RECT 7387.445 1046.435 7399.765 10000 ;
      RECT 7380.585 1046.935 7380.865 10000 ;
      RECT 7379.465 1046.935 7379.745 10000 ;
      RECT 7377.225 1046.935 7377.505 10000 ;
      RECT 7376.105 1046.935 7376.385 10000 ;
      RECT 7374.985 1046.935 7375.265 10000 ;
      RECT 7334.245 1046.435 7373.445 10000 ;
      RECT 7327.945 1046.935 7328.225 10000 ;
      RECT 7326.825 1046.935 7327.105 10000 ;
      RECT 7325.705 1046.935 7325.985 10000 ;
      RECT 7312.265 1046.935 7320.805 10000 ;
      RECT 7312.405 1046.435 7320.805 10000 ;
      RECT 7311.145 1046.935 7311.425 10000 ;
      RECT 7303.165 1046.435 7304.565 10000 ;
      RECT 7300.785 1046.935 7301.065 10000 ;
      RECT 7299.665 1046.935 7299.945 10000 ;
      RECT 7272.645 1046.435 7298.125 10000 ;
      RECT 7271.385 1046.935 7271.665 10000 ;
      RECT 7270.265 1046.935 7270.545 10000 ;
      RECT 7269.145 1046.935 7269.425 10000 ;
      RECT 7261.865 1046.935 7262.145 10000 ;
      RECT 7260.745 1046.935 7261.025 10000 ;
      RECT 7246.185 1046.935 7259.765 10000 ;
      RECT 7246.325 1046.435 7259.765 10000 ;
      RECT 7241.145 1046.935 7241.425 10000 ;
      RECT 7240.025 1046.935 7240.305 10000 ;
      RECT 7195.365 1046.435 7233.445 10000 ;
      RECT 7192.985 1046.935 7193.265 10000 ;
      RECT 7191.865 1046.935 7192.145 10000 ;
      RECT 7189.625 1046.935 7189.905 10000 ;
      RECT 7188.505 1046.935 7188.785 10000 ;
      RECT 7187.385 1046.935 7187.665 10000 ;
      RECT 7172.965 1046.435 7180.805 10000 ;
      RECT 7171.705 1046.935 7171.985 10000 ;
      RECT 7170.585 1046.935 7170.865 10000 ;
      RECT 7169.465 1046.935 7169.745 10000 ;
      RECT 7162.465 1046.935 7164.565 10000 ;
      RECT 7162.605 1046.435 7164.565 10000 ;
      RECT 7161.345 1046.935 7161.625 10000 ;
      RECT 7133.205 1046.435 7158.125 10000 ;
      RECT 7127.465 1046.935 7127.745 10000 ;
      RECT 7126.345 1046.935 7126.625 10000 ;
      RECT 7124.105 1046.935 7124.385 10000 ;
      RECT 7122.985 1046.935 7123.265 10000 ;
      RECT 7121.865 1046.935 7122.145 10000 ;
      RECT 7106.885 1046.435 7119.205 10000 ;
      RECT 7101.705 1046.935 7101.985 10000 ;
      RECT 7100.585 1046.935 7100.865 10000 ;
      RECT 7099.465 1046.935 7099.745 10000 ;
      RECT 7094.425 1046.935 7094.705 10000 ;
      RECT 7054.805 1046.935 7093.585 10000 ;
      RECT 7046.265 1046.935 7046.545 10000 ;
      RECT 7045.145 1046.935 7045.425 10000 ;
      RECT 7042.905 1046.935 7043.185 10000 ;
      RECT 7041.785 1046.935 7042.065 10000 ;
      RECT 7032.265 1046.935 7040.805 10000 ;
      RECT 7032.405 1046.435 7040.805 10000 ;
      RECT 7023.165 1046.935 7025.265 10000 ;
      RECT 7021.905 1046.935 7022.185 10000 ;
      RECT 7020.785 1046.935 7021.065 10000 ;
      RECT 6993.765 1046.435 7018.685 10000 ;
      RECT 6990.265 1046.935 6990.545 10000 ;
      RECT 6989.145 1046.935 6989.425 10000 ;
      RECT 6980.745 1046.935 6981.025 10000 ;
      RECT 6966.745 1046.935 6979.765 10000 ;
      RECT 6966.885 1046.435 6979.765 10000 ;
      RECT 6964.505 1046.935 6964.785 10000 ;
      RECT 6963.385 1046.935 6963.665 10000 ;
      RECT 6962.265 1046.935 6962.545 10000 ;
      RECT 6954.985 1046.935 6955.265 10000 ;
      RECT 6914.805 1046.935 6954.145 10000 ;
      RECT 6913.545 1046.935 6913.825 10000 ;
      RECT 6908.505 1046.935 6908.785 10000 ;
      RECT 6907.385 1046.935 6907.665 10000 ;
      RECT 6892.965 1046.435 6900.805 10000 ;
      RECT 6890.585 1046.935 6890.865 10000 ;
      RECT 6889.465 1046.935 6889.745 10000 ;
      RECT 6887.225 1046.935 6887.505 10000 ;
      RECT 6886.105 1046.935 6886.385 10000 ;
      RECT 6883.165 1046.935 6885.265 10000 ;
      RECT 6853.765 1046.435 6878.685 10000 ;
      RECT 6850.265 1046.935 6850.545 10000 ;
      RECT 6849.145 1046.935 6849.425 10000 ;
      RECT 6848.025 1046.935 6848.305 10000 ;
      RECT 6842.985 1046.935 6843.265 10000 ;
      RECT 6841.865 1046.935 6842.145 10000 ;
      RECT 6827.445 1046.435 6839.765 10000 ;
      RECT 6820.585 1046.935 6820.865 10000 ;
      RECT 6819.465 1046.935 6819.745 10000 ;
      RECT 6817.225 1046.935 6817.505 10000 ;
      RECT 6816.105 1046.935 6816.385 10000 ;
      RECT 6814.985 1046.935 6815.265 10000 ;
      RECT 6774.245 1046.435 6813.445 10000 ;
      RECT 6767.945 1046.935 6768.225 10000 ;
      RECT 6766.825 1046.935 6767.105 10000 ;
      RECT 6765.705 1046.935 6765.985 10000 ;
      RECT 6752.265 1046.935 6760.805 10000 ;
      RECT 6752.405 1046.435 6760.805 10000 ;
      RECT 6751.145 1046.935 6751.425 10000 ;
      RECT 6743.165 1046.435 6744.565 10000 ;
      RECT 6740.785 1046.935 6741.065 10000 ;
      RECT 6739.665 1046.935 6739.945 10000 ;
      RECT 6712.645 1046.435 6738.125 10000 ;
      RECT 6711.385 1046.935 6711.665 10000 ;
      RECT 6710.265 1046.935 6710.545 10000 ;
      RECT 6709.145 1046.935 6709.425 10000 ;
      RECT 6701.865 1046.935 6702.145 10000 ;
      RECT 6700.745 1046.935 6701.025 10000 ;
      RECT 6686.185 1046.935 6699.765 10000 ;
      RECT 6686.325 1046.435 6699.765 10000 ;
      RECT 6681.145 1046.935 6681.425 10000 ;
      RECT 6680.025 1046.935 6680.305 10000 ;
      RECT 6635.365 1046.435 6673.445 10000 ;
      RECT 6632.985 1046.935 6633.265 10000 ;
      RECT 6631.865 1046.935 6632.145 10000 ;
      RECT 6629.625 1046.935 6629.905 10000 ;
      RECT 6628.505 1046.935 6628.785 10000 ;
      RECT 6627.385 1046.935 6627.665 10000 ;
      RECT 6612.965 1046.435 6620.805 10000 ;
      RECT 6611.705 1046.935 6611.985 10000 ;
      RECT 6610.585 1046.935 6610.865 10000 ;
      RECT 6609.465 1046.935 6609.745 10000 ;
      RECT 6602.465 1046.935 6604.565 10000 ;
      RECT 6602.605 1046.435 6604.565 10000 ;
      RECT 6601.345 1046.935 6601.625 10000 ;
      RECT 6573.205 1046.435 6598.125 10000 ;
      RECT 6567.465 1046.935 6567.745 10000 ;
      RECT 6566.345 1046.935 6566.625 10000 ;
      RECT 6564.105 1046.935 6564.385 10000 ;
      RECT 6562.985 1046.935 6563.265 10000 ;
      RECT 6561.865 1046.935 6562.145 10000 ;
      RECT 6546.885 1046.435 6559.205 10000 ;
      RECT 6541.705 1046.935 6541.985 10000 ;
      RECT 6540.585 1046.935 6540.865 10000 ;
      RECT 6539.465 1046.935 6539.745 10000 ;
      RECT 6534.425 1046.935 6534.705 10000 ;
      RECT 6494.805 1046.935 6533.585 10000 ;
      RECT 6486.265 1046.935 6486.545 10000 ;
      RECT 6485.145 1046.935 6485.425 10000 ;
      RECT 6482.905 1046.935 6483.185 10000 ;
      RECT 6481.785 1046.935 6482.065 10000 ;
      RECT 6472.265 1046.935 6480.805 10000 ;
      RECT 6472.405 1046.435 6480.805 10000 ;
      RECT 6463.165 1046.935 6465.265 10000 ;
      RECT 6461.905 1046.935 6462.185 10000 ;
      RECT 6460.785 1046.935 6461.065 10000 ;
      RECT 6433.765 1046.435 6458.685 10000 ;
      RECT 6430.265 1046.935 6430.545 10000 ;
      RECT 6429.145 1046.935 6429.425 10000 ;
      RECT 6420.745 1046.935 6421.025 10000 ;
      RECT 6406.745 1046.935 6419.765 10000 ;
      RECT 6406.885 1046.435 6419.765 10000 ;
      RECT 6404.505 1046.935 6404.785 10000 ;
      RECT 6403.385 1046.935 6403.665 10000 ;
      RECT 6402.265 1046.935 6402.545 10000 ;
      RECT 6394.985 1046.935 6395.265 10000 ;
      RECT 6354.805 1046.935 6394.145 10000 ;
      RECT 6353.545 1046.935 6353.825 10000 ;
      RECT 6348.505 1046.935 6348.785 10000 ;
      RECT 6347.385 1046.935 6347.665 10000 ;
      RECT 6332.965 1046.435 6340.805 10000 ;
      RECT 6330.585 1046.935 6330.865 10000 ;
      RECT 6329.465 1046.935 6329.745 10000 ;
      RECT 6327.225 1046.935 6327.505 10000 ;
      RECT 6326.105 1046.935 6326.385 10000 ;
      RECT 6323.165 1046.935 6325.265 10000 ;
      RECT 6293.765 1046.435 6318.685 10000 ;
      RECT 6290.265 1046.935 6290.545 10000 ;
      RECT 6289.145 1046.935 6289.425 10000 ;
      RECT 6288.025 1046.935 6288.305 10000 ;
      RECT 6282.985 1046.935 6283.265 10000 ;
      RECT 6281.865 1046.935 6282.145 10000 ;
      RECT 6267.445 1046.435 6279.765 10000 ;
      RECT 6260.585 1046.935 6260.865 10000 ;
      RECT 6259.465 1046.935 6259.745 10000 ;
      RECT 6257.225 1046.935 6257.505 10000 ;
      RECT 6256.105 1046.935 6256.385 10000 ;
      RECT 6254.985 1046.935 6255.265 10000 ;
      RECT 6214.245 1046.435 6253.445 10000 ;
      RECT 6207.945 1046.935 6208.225 10000 ;
      RECT 6206.825 1046.935 6207.105 10000 ;
      RECT 6205.705 1046.935 6205.985 10000 ;
      RECT 6192.265 1046.935 6200.805 10000 ;
      RECT 6192.405 1046.435 6200.805 10000 ;
      RECT 6191.145 1046.935 6191.425 10000 ;
      RECT 6183.165 1046.435 6184.565 10000 ;
      RECT 6180.785 1046.935 6181.065 10000 ;
      RECT 6179.665 1046.935 6179.945 10000 ;
      RECT 6152.645 1046.435 6178.125 10000 ;
      RECT 6151.385 1046.935 6151.665 10000 ;
      RECT 6150.265 1046.935 6150.545 10000 ;
      RECT 6149.145 1046.935 6149.425 10000 ;
      RECT 6141.865 1046.935 6142.145 10000 ;
      RECT 6140.745 1046.935 6141.025 10000 ;
      RECT 6126.185 1046.935 6139.765 10000 ;
      RECT 6126.325 1046.435 6139.765 10000 ;
      RECT 6121.145 1046.935 6121.425 10000 ;
      RECT 6120.025 1046.935 6120.305 10000 ;
      RECT 6075.365 1046.435 6113.445 10000 ;
      RECT 6072.985 1046.935 6073.265 10000 ;
      RECT 6071.865 1046.935 6072.145 10000 ;
      RECT 6069.625 1046.935 6069.905 10000 ;
      RECT 6068.505 1046.935 6068.785 10000 ;
      RECT 6067.385 1046.935 6067.665 10000 ;
      RECT 6052.965 1046.435 6060.805 10000 ;
      RECT 6051.705 1046.935 6051.985 10000 ;
      RECT 6050.585 1046.935 6050.865 10000 ;
      RECT 6049.465 1046.935 6049.745 10000 ;
      RECT 6042.465 1046.935 6044.565 10000 ;
      RECT 6042.605 1046.435 6044.565 10000 ;
      RECT 6041.345 1046.935 6041.625 10000 ;
      RECT 6013.205 1046.435 6038.125 10000 ;
      RECT 6007.465 1046.935 6007.745 10000 ;
      RECT 6006.345 1046.935 6006.625 10000 ;
      RECT 6004.105 1046.935 6004.385 10000 ;
      RECT 6002.985 1046.935 6003.265 10000 ;
      RECT 6001.865 1046.935 6002.145 10000 ;
      RECT 5986.885 1046.435 5999.205 10000 ;
      RECT 5981.705 1046.935 5981.985 10000 ;
      RECT 5980.585 1046.935 5980.865 10000 ;
      RECT 5979.465 1046.935 5979.745 10000 ;
      RECT 5974.425 1046.935 5974.705 10000 ;
      RECT 5934.805 1046.935 5973.585 10000 ;
      RECT 5926.265 1046.935 5926.545 10000 ;
      RECT 5925.145 1046.935 5925.425 10000 ;
      RECT 5922.905 1046.935 5923.185 10000 ;
      RECT 5921.785 1046.935 5922.065 10000 ;
      RECT 5912.265 1046.935 5920.805 10000 ;
      RECT 5912.405 1046.435 5920.805 10000 ;
      RECT 5903.165 1046.935 5905.265 10000 ;
      RECT 5901.905 1046.935 5902.185 10000 ;
      RECT 5900.785 1046.935 5901.065 10000 ;
      RECT 5873.765 1046.435 5898.685 10000 ;
      RECT 5870.265 1046.935 5870.545 10000 ;
      RECT 5869.145 1046.935 5869.425 10000 ;
      RECT 5860.745 1046.935 5861.025 10000 ;
      RECT 5846.745 1046.935 5859.765 10000 ;
      RECT 5846.885 1046.435 5859.765 10000 ;
      RECT 5844.505 1046.935 5844.785 10000 ;
      RECT 5843.385 1046.935 5843.665 10000 ;
      RECT 5842.265 1046.935 5842.545 10000 ;
      RECT 5834.985 1046.935 5835.265 10000 ;
      RECT 5794.805 1046.935 5834.145 10000 ;
      RECT 5793.545 1046.935 5793.825 10000 ;
      RECT 5788.505 1046.935 5788.785 10000 ;
      RECT 5787.385 1046.935 5787.665 10000 ;
      RECT 5772.965 1046.435 5780.805 10000 ;
      RECT 5770.585 1046.935 5770.865 10000 ;
      RECT 5769.465 1046.935 5769.745 10000 ;
      RECT 5767.225 1046.935 5767.505 10000 ;
      RECT 5766.105 1046.935 5766.385 10000 ;
      RECT 5763.165 1046.935 5765.265 10000 ;
      RECT 5733.765 1046.435 5758.685 10000 ;
      RECT 5730.265 1046.935 5730.545 10000 ;
      RECT 5729.145 1046.935 5729.425 10000 ;
      RECT 5728.025 1046.935 5728.305 10000 ;
      RECT 5722.985 1046.935 5723.265 10000 ;
      RECT 5721.865 1046.935 5722.145 10000 ;
      RECT 5707.445 1046.435 5719.765 10000 ;
      RECT 5700.585 1046.935 5700.865 10000 ;
      RECT 5699.465 1046.935 5699.745 10000 ;
      RECT 5697.225 1046.935 5697.505 10000 ;
      RECT 5696.105 1046.935 5696.385 10000 ;
      RECT 5694.985 1046.935 5695.265 10000 ;
      RECT 5654.245 1046.435 5693.445 10000 ;
      RECT 5647.945 1046.935 5648.225 10000 ;
      RECT 5646.825 1046.935 5647.105 10000 ;
      RECT 5645.705 1046.935 5645.985 10000 ;
      RECT 5632.265 1046.935 5640.805 10000 ;
      RECT 5632.405 1046.435 5640.805 10000 ;
      RECT 5631.145 1046.935 5631.425 10000 ;
      RECT 5623.165 1046.435 5624.565 10000 ;
      RECT 5620.785 1046.935 5621.065 10000 ;
      RECT 5619.665 1046.935 5619.945 10000 ;
      RECT 5592.645 1046.435 5618.125 10000 ;
      RECT 5591.385 1046.935 5591.665 10000 ;
      RECT 5590.265 1046.935 5590.545 10000 ;
      RECT 5589.145 1046.935 5589.425 10000 ;
      RECT 5581.865 1046.935 5582.145 10000 ;
      RECT 5580.745 1046.935 5581.025 10000 ;
      RECT 5566.185 1046.935 5579.765 10000 ;
      RECT 5566.325 1046.435 5579.765 10000 ;
      RECT 5561.145 1046.935 5561.425 10000 ;
      RECT 5560.025 1046.935 5560.305 10000 ;
      RECT 5515.365 1046.435 5553.445 10000 ;
      RECT 5512.985 1046.935 5513.265 10000 ;
      RECT 5511.865 1046.935 5512.145 10000 ;
      RECT 5509.625 1046.935 5509.905 10000 ;
      RECT 5508.505 1046.935 5508.785 10000 ;
      RECT 5507.385 1046.935 5507.665 10000 ;
      RECT 5492.965 1046.435 5500.805 10000 ;
      RECT 5491.705 1046.935 5491.985 10000 ;
      RECT 5490.585 1046.935 5490.865 10000 ;
      RECT 5489.465 1046.935 5489.745 10000 ;
      RECT 5482.465 1046.935 5484.565 10000 ;
      RECT 5482.605 1046.435 5484.565 10000 ;
      RECT 5481.345 1046.935 5481.625 10000 ;
      RECT 5453.205 1046.435 5478.125 10000 ;
      RECT 5447.465 1046.935 5447.745 10000 ;
      RECT 5446.345 1046.935 5446.625 10000 ;
      RECT 5444.105 1046.935 5444.385 10000 ;
      RECT 5442.985 1046.935 5443.265 10000 ;
      RECT 5441.865 1046.935 5442.145 10000 ;
      RECT 5426.885 1046.435 5439.205 10000 ;
      RECT 5421.705 1046.935 5421.985 10000 ;
      RECT 5420.585 1046.935 5420.865 10000 ;
      RECT 5419.465 1046.935 5419.745 10000 ;
      RECT 5414.425 1046.935 5414.705 10000 ;
      RECT 5374.805 1046.935 5413.585 10000 ;
      RECT 5366.265 1046.935 5366.545 10000 ;
      RECT 5365.145 1046.935 5365.425 10000 ;
      RECT 5362.905 1046.935 5363.185 10000 ;
      RECT 5361.785 1046.935 5362.065 10000 ;
      RECT 5352.265 1046.935 5360.805 10000 ;
      RECT 5352.405 1046.435 5360.805 10000 ;
      RECT 5343.165 1046.935 5345.265 10000 ;
      RECT 5341.905 1046.935 5342.185 10000 ;
      RECT 5340.785 1046.935 5341.065 10000 ;
      RECT 5313.765 1046.435 5338.685 10000 ;
      RECT 5310.265 1046.935 5310.545 10000 ;
      RECT 5309.145 1046.935 5309.425 10000 ;
      RECT 5300.745 1046.935 5301.025 10000 ;
      RECT 5286.745 1046.935 5299.765 10000 ;
      RECT 5286.885 1046.435 5299.765 10000 ;
      RECT 5284.505 1046.935 5284.785 10000 ;
      RECT 5283.385 1046.935 5283.665 10000 ;
      RECT 5282.265 1046.935 5282.545 10000 ;
      RECT 5274.985 1046.935 5275.265 10000 ;
      RECT 5234.805 1046.935 5274.145 10000 ;
      RECT 5233.545 1046.935 5233.825 10000 ;
      RECT 5228.505 1046.935 5228.785 10000 ;
      RECT 5227.385 1046.935 5227.665 10000 ;
      RECT 5212.965 1046.435 5220.805 10000 ;
      RECT 5210.585 1046.935 5210.865 10000 ;
      RECT 5209.465 1046.935 5209.745 10000 ;
      RECT 5207.225 1046.935 5207.505 10000 ;
      RECT 5206.105 1046.935 5206.385 10000 ;
      RECT 5203.165 1046.935 5205.265 10000 ;
      RECT 5173.765 1046.435 5198.685 10000 ;
      RECT 5170.265 1046.935 5170.545 10000 ;
      RECT 5169.145 1046.935 5169.425 10000 ;
      RECT 5168.025 1046.935 5168.305 10000 ;
      RECT 5162.985 1046.935 5163.265 10000 ;
      RECT 5161.865 1046.935 5162.145 10000 ;
      RECT 5147.445 1046.435 5159.765 10000 ;
      RECT 5140.585 1046.935 5140.865 10000 ;
      RECT 5139.465 1046.935 5139.745 10000 ;
      RECT 5137.225 1046.935 5137.505 10000 ;
      RECT 5136.105 1046.935 5136.385 10000 ;
      RECT 5134.985 1046.935 5135.265 10000 ;
      RECT 5094.245 1046.435 5133.445 10000 ;
      RECT 5087.945 1046.935 5088.225 10000 ;
      RECT 5086.825 1046.935 5087.105 10000 ;
      RECT 5085.705 1046.935 5085.985 10000 ;
      RECT 5072.265 1046.935 5080.805 10000 ;
      RECT 5072.405 1046.435 5080.805 10000 ;
      RECT 5071.145 1046.935 5071.425 10000 ;
      RECT 5063.165 1046.435 5064.565 10000 ;
      RECT 5060.785 1046.935 5061.065 10000 ;
      RECT 5059.665 1046.935 5059.945 10000 ;
      RECT 5032.645 1046.435 5058.125 10000 ;
      RECT 5031.385 1046.935 5031.665 10000 ;
      RECT 5030.265 1046.935 5030.545 10000 ;
      RECT 5029.145 1046.935 5029.425 10000 ;
      RECT 5021.865 1046.935 5022.145 10000 ;
      RECT 5020.745 1046.935 5021.025 10000 ;
      RECT 5006.185 1046.935 5019.765 10000 ;
      RECT 5006.325 1046.435 5019.765 10000 ;
      RECT 5001.145 1046.935 5001.425 10000 ;
      RECT 5000.025 1046.935 5000.305 10000 ;
      RECT 4955.365 1046.435 4993.445 10000 ;
      RECT 4952.985 1046.935 4953.265 10000 ;
      RECT 4951.865 1046.935 4952.145 10000 ;
      RECT 4949.625 1046.935 4949.905 10000 ;
      RECT 4948.505 1046.935 4948.785 10000 ;
      RECT 4947.385 1046.935 4947.665 10000 ;
      RECT 4932.965 1046.435 4940.805 10000 ;
      RECT 4931.705 1046.935 4931.985 10000 ;
      RECT 4930.585 1046.935 4930.865 10000 ;
      RECT 4929.465 1046.935 4929.745 10000 ;
      RECT 4922.465 1046.935 4924.565 10000 ;
      RECT 4922.605 1046.435 4924.565 10000 ;
      RECT 4921.345 1046.935 4921.625 10000 ;
      RECT 4893.205 1046.435 4918.125 10000 ;
      RECT 4887.465 1046.935 4887.745 10000 ;
      RECT 4886.345 1046.935 4886.625 10000 ;
      RECT 4884.105 1046.935 4884.385 10000 ;
      RECT 4882.985 1046.935 4883.265 10000 ;
      RECT 4881.865 1046.935 4882.145 10000 ;
      RECT 4866.885 1046.435 4879.205 10000 ;
      RECT 4861.705 1046.935 4861.985 10000 ;
      RECT 4860.585 1046.935 4860.865 10000 ;
      RECT 4859.465 1046.935 4859.745 10000 ;
      RECT 4854.425 1046.935 4854.705 10000 ;
      RECT 4814.805 1046.935 4853.585 10000 ;
      RECT 4806.265 1046.935 4806.545 10000 ;
      RECT 4805.145 1046.935 4805.425 10000 ;
      RECT 4802.905 1046.935 4803.185 10000 ;
      RECT 4801.785 1046.935 4802.065 10000 ;
      RECT 4792.265 1046.935 4800.805 10000 ;
      RECT 4792.405 1046.435 4800.805 10000 ;
      RECT 4783.165 1046.935 4785.265 10000 ;
      RECT 4781.905 1046.935 4782.185 10000 ;
      RECT 4780.785 1046.935 4781.065 10000 ;
      RECT 4753.765 1046.435 4778.685 10000 ;
      RECT 4750.265 1046.935 4750.545 10000 ;
      RECT 4749.145 1046.935 4749.425 10000 ;
      RECT 4740.745 1046.935 4741.025 10000 ;
      RECT 4726.745 1046.935 4739.765 10000 ;
      RECT 4726.885 1046.435 4739.765 10000 ;
      RECT 4724.505 1046.935 4724.785 10000 ;
      RECT 4723.385 1046.935 4723.665 10000 ;
      RECT 4722.265 1046.935 4722.545 10000 ;
      RECT 4714.985 1046.935 4715.265 10000 ;
      RECT 4674.805 1046.935 4714.145 10000 ;
      RECT 4673.545 1046.935 4673.825 10000 ;
      RECT 4668.505 1046.935 4668.785 10000 ;
      RECT 4667.385 1046.935 4667.665 10000 ;
      RECT 4652.965 1046.435 4660.805 10000 ;
      RECT 4650.585 1046.935 4650.865 10000 ;
      RECT 4649.465 1046.935 4649.745 10000 ;
      RECT 4647.225 1046.935 4647.505 10000 ;
      RECT 4646.105 1046.935 4646.385 10000 ;
      RECT 4643.165 1046.935 4645.265 10000 ;
      RECT 4613.765 1046.435 4638.685 10000 ;
      RECT 4610.265 1046.935 4610.545 10000 ;
      RECT 4609.145 1046.935 4609.425 10000 ;
      RECT 4608.025 1046.935 4608.305 10000 ;
      RECT 4602.985 1046.935 4603.265 10000 ;
      RECT 4601.865 1046.935 4602.145 10000 ;
      RECT 4587.445 1046.435 4599.765 10000 ;
      RECT 4580.585 1046.935 4580.865 10000 ;
      RECT 4579.465 1046.935 4579.745 10000 ;
      RECT 4577.225 1046.935 4577.505 10000 ;
      RECT 4576.105 1046.935 4576.385 10000 ;
      RECT 4574.985 1046.935 4575.265 10000 ;
      RECT 4534.245 1046.435 4573.445 10000 ;
      RECT 4527.945 1046.935 4528.225 10000 ;
      RECT 4526.825 1046.935 4527.105 10000 ;
      RECT 4525.705 1046.935 4525.985 10000 ;
      RECT 4512.265 1046.935 4520.805 10000 ;
      RECT 4512.405 1046.435 4520.805 10000 ;
      RECT 4511.145 1046.935 4511.425 10000 ;
      RECT 4503.165 1046.435 4504.565 10000 ;
      RECT 4500.785 1046.935 4501.065 10000 ;
      RECT 4499.665 1046.935 4499.945 10000 ;
      RECT 4472.645 1046.435 4498.125 10000 ;
      RECT 4471.385 1046.935 4471.665 10000 ;
      RECT 4470.265 1046.935 4470.545 10000 ;
      RECT 4469.145 1046.935 4469.425 10000 ;
      RECT 4461.865 1046.935 4462.145 10000 ;
      RECT 4460.745 1046.935 4461.025 10000 ;
      RECT 4446.185 1046.935 4459.765 10000 ;
      RECT 4446.325 1046.435 4459.765 10000 ;
      RECT 4441.145 1046.935 4441.425 10000 ;
      RECT 4440.025 1046.935 4440.305 10000 ;
      RECT 4395.365 1046.435 4433.445 10000 ;
      RECT 4392.985 1046.935 4393.265 10000 ;
      RECT 4391.865 1046.935 4392.145 10000 ;
      RECT 4389.625 1046.935 4389.905 10000 ;
      RECT 4388.505 1046.935 4388.785 10000 ;
      RECT 4387.385 1046.935 4387.665 10000 ;
      RECT 4372.965 1046.435 4380.805 10000 ;
      RECT 4371.705 1046.935 4371.985 10000 ;
      RECT 4370.585 1046.935 4370.865 10000 ;
      RECT 4369.465 1046.935 4369.745 10000 ;
      RECT 4362.465 1046.935 4364.565 10000 ;
      RECT 4362.605 1046.435 4364.565 10000 ;
      RECT 4361.345 1046.935 4361.625 10000 ;
      RECT 4333.205 1046.435 4358.125 10000 ;
      RECT 4327.465 1046.935 4327.745 10000 ;
      RECT 4326.345 1046.935 4326.625 10000 ;
      RECT 4324.105 1046.935 4324.385 10000 ;
      RECT 4322.985 1046.935 4323.265 10000 ;
      RECT 4321.865 1046.935 4322.145 10000 ;
      RECT 4306.885 1046.435 4319.205 10000 ;
      RECT 4301.705 1046.935 4301.985 10000 ;
      RECT 4300.585 1046.935 4300.865 10000 ;
      RECT 4299.465 1046.935 4299.745 10000 ;
      RECT 4294.425 1046.935 4294.705 10000 ;
      RECT 4254.805 1046.935 4293.585 10000 ;
      RECT 4246.265 1046.935 4246.545 10000 ;
      RECT 4245.145 1046.935 4245.425 10000 ;
      RECT 4242.905 1046.935 4243.185 10000 ;
      RECT 4241.785 1046.935 4242.065 10000 ;
      RECT 4232.265 1046.935 4240.805 10000 ;
      RECT 4232.405 1046.435 4240.805 10000 ;
      RECT 4223.165 1046.935 4225.265 10000 ;
      RECT 4221.905 1046.935 4222.185 10000 ;
      RECT 4220.785 1046.935 4221.065 10000 ;
      RECT 4193.765 1046.435 4218.685 10000 ;
      RECT 4190.265 1046.935 4190.545 10000 ;
      RECT 4189.145 1046.935 4189.425 10000 ;
      RECT 4180.745 1046.935 4181.025 10000 ;
      RECT 4166.745 1046.935 4179.765 10000 ;
      RECT 4166.885 1046.435 4179.765 10000 ;
      RECT 4164.505 1046.935 4164.785 10000 ;
      RECT 4163.385 1046.935 4163.665 10000 ;
      RECT 4162.265 1046.935 4162.545 10000 ;
      RECT 4154.985 1046.935 4155.265 10000 ;
      RECT 4114.805 1046.935 4154.145 10000 ;
      RECT 4113.545 1046.935 4113.825 10000 ;
      RECT 4108.505 1046.935 4108.785 10000 ;
      RECT 4107.385 1046.935 4107.665 10000 ;
      RECT 4092.965 1046.435 4100.805 10000 ;
      RECT 4090.585 1046.935 4090.865 10000 ;
      RECT 4089.465 1046.935 4089.745 10000 ;
      RECT 4087.225 1046.935 4087.505 10000 ;
      RECT 4086.105 1046.935 4086.385 10000 ;
      RECT 4083.165 1046.935 4085.265 10000 ;
      RECT 4053.765 1046.435 4078.685 10000 ;
      RECT 4050.265 1046.935 4050.545 10000 ;
      RECT 4049.145 1046.935 4049.425 10000 ;
      RECT 4048.025 1046.935 4048.305 10000 ;
      RECT 4042.985 1046.935 4043.265 10000 ;
      RECT 4041.865 1046.935 4042.145 10000 ;
      RECT 4027.445 1046.435 4039.765 10000 ;
      RECT 4020.585 1046.935 4020.865 10000 ;
      RECT 4019.465 1046.935 4019.745 10000 ;
      RECT 4017.225 1046.935 4017.505 10000 ;
      RECT 4016.105 1046.935 4016.385 10000 ;
      RECT 4014.985 1046.935 4015.265 10000 ;
      RECT 3974.245 1046.435 4013.445 10000 ;
      RECT 3967.945 1046.935 3968.225 10000 ;
      RECT 3966.825 1046.935 3967.105 10000 ;
      RECT 3965.705 1046.935 3965.985 10000 ;
      RECT 3952.265 1046.935 3960.805 10000 ;
      RECT 3952.405 1046.435 3960.805 10000 ;
      RECT 3951.145 1046.935 3951.425 10000 ;
      RECT 3943.165 1046.435 3944.565 10000 ;
      RECT 3940.785 1046.935 3941.065 10000 ;
      RECT 3939.665 1046.935 3939.945 10000 ;
      RECT 3912.645 1046.435 3938.125 10000 ;
      RECT 3911.385 1046.935 3911.665 10000 ;
      RECT 3910.265 1046.935 3910.545 10000 ;
      RECT 3909.145 1046.935 3909.425 10000 ;
      RECT 3901.865 1046.935 3902.145 10000 ;
      RECT 3900.745 1046.935 3901.025 10000 ;
      RECT 3886.185 1046.935 3899.765 10000 ;
      RECT 3886.325 1046.435 3899.765 10000 ;
      RECT 3881.145 1046.935 3881.425 10000 ;
      RECT 3880.025 1046.935 3880.305 10000 ;
      RECT 3835.365 1046.435 3873.445 10000 ;
      RECT 3832.985 1046.935 3833.265 10000 ;
      RECT 3831.865 1046.935 3832.145 10000 ;
      RECT 3829.625 1046.935 3829.905 10000 ;
      RECT 3828.505 1046.935 3828.785 10000 ;
      RECT 3827.385 1046.935 3827.665 10000 ;
      RECT 3812.965 1046.435 3820.805 10000 ;
      RECT 3811.705 1046.935 3811.985 10000 ;
      RECT 3810.585 1046.935 3810.865 10000 ;
      RECT 3809.465 1046.935 3809.745 10000 ;
      RECT 3802.465 1046.935 3804.565 10000 ;
      RECT 3802.605 1046.435 3804.565 10000 ;
      RECT 3801.345 1046.935 3801.625 10000 ;
      RECT 3773.205 1046.435 3798.125 10000 ;
      RECT 3767.465 1046.935 3767.745 10000 ;
      RECT 3766.345 1046.935 3766.625 10000 ;
      RECT 3764.105 1046.935 3764.385 10000 ;
      RECT 3762.985 1046.935 3763.265 10000 ;
      RECT 3761.865 1046.935 3762.145 10000 ;
      RECT 3746.885 1046.435 3759.205 10000 ;
      RECT 3741.705 1046.935 3741.985 10000 ;
      RECT 3740.585 1046.935 3740.865 10000 ;
      RECT 3739.465 1046.935 3739.745 10000 ;
      RECT 3734.425 1046.935 3734.705 10000 ;
      RECT 3694.805 1046.935 3733.585 10000 ;
      RECT 3686.265 1046.935 3686.545 10000 ;
      RECT 3685.145 1046.935 3685.425 10000 ;
      RECT 3682.905 1046.935 3683.185 10000 ;
      RECT 3681.785 1046.935 3682.065 10000 ;
      RECT 3672.265 1046.935 3680.805 10000 ;
      RECT 3672.405 1046.435 3680.805 10000 ;
      RECT 3663.165 1046.935 3665.265 10000 ;
      RECT 3661.905 1046.935 3662.185 10000 ;
      RECT 3660.785 1046.935 3661.065 10000 ;
      RECT 3633.765 1046.435 3658.685 10000 ;
      RECT 3630.265 1046.935 3630.545 10000 ;
      RECT 3629.145 1046.935 3629.425 10000 ;
      RECT 3620.745 1046.935 3621.025 10000 ;
      RECT 3606.745 1046.935 3619.765 10000 ;
      RECT 3606.885 1046.435 3619.765 10000 ;
      RECT 3604.505 1046.935 3604.785 10000 ;
      RECT 3603.385 1046.935 3603.665 10000 ;
      RECT 3602.265 1046.935 3602.545 10000 ;
      RECT 3594.985 1046.935 3595.265 10000 ;
      RECT 3554.805 1046.935 3594.145 10000 ;
      RECT 3553.545 1046.935 3553.825 10000 ;
      RECT 3548.505 1046.935 3548.785 10000 ;
      RECT 3547.385 1046.935 3547.665 10000 ;
      RECT 3532.965 1046.435 3540.805 10000 ;
      RECT 3530.585 1046.935 3530.865 10000 ;
      RECT 3529.465 1046.935 3529.745 10000 ;
      RECT 3527.225 1046.935 3527.505 10000 ;
      RECT 3526.105 1046.935 3526.385 10000 ;
      RECT 3523.165 1046.935 3525.265 10000 ;
      RECT 3493.765 1046.435 3518.685 10000 ;
      RECT 3490.265 1046.935 3490.545 10000 ;
      RECT 3489.145 1046.935 3489.425 10000 ;
      RECT 3488.025 1046.935 3488.305 10000 ;
      RECT 3482.985 1046.935 3483.265 10000 ;
      RECT 3481.865 1046.935 3482.145 10000 ;
      RECT 3467.445 1046.435 3479.765 10000 ;
      RECT 3460.585 1046.935 3460.865 10000 ;
      RECT 3459.465 1046.935 3459.745 10000 ;
      RECT 3457.225 1046.935 3457.505 10000 ;
      RECT 3456.105 1046.935 3456.385 10000 ;
      RECT 3454.985 1046.935 3455.265 10000 ;
      RECT 3414.245 1046.435 3453.445 10000 ;
      RECT 3407.945 1046.935 3408.225 10000 ;
      RECT 3406.825 1046.935 3407.105 10000 ;
      RECT 3405.705 1046.935 3405.985 10000 ;
      RECT 3392.265 1046.935 3400.805 10000 ;
      RECT 3392.405 1046.435 3400.805 10000 ;
      RECT 3391.145 1046.935 3391.425 10000 ;
      RECT 3383.165 1046.435 3384.565 10000 ;
      RECT 3380.785 1046.935 3381.065 10000 ;
      RECT 3379.665 1046.935 3379.945 10000 ;
      RECT 3352.645 1046.435 3378.125 10000 ;
      RECT 3351.385 1046.935 3351.665 10000 ;
      RECT 3350.265 1046.935 3350.545 10000 ;
      RECT 3349.145 1046.935 3349.425 10000 ;
      RECT 3341.865 1046.935 3342.145 10000 ;
      RECT 3340.745 1046.935 3341.025 10000 ;
      RECT 3326.185 1046.935 3339.765 10000 ;
      RECT 3326.325 1046.435 3339.765 10000 ;
      RECT 3321.145 1046.935 3321.425 10000 ;
      RECT 3320.025 1046.935 3320.305 10000 ;
      RECT 3275.365 1046.435 3313.445 10000 ;
      RECT 3272.985 1046.935 3273.265 10000 ;
      RECT 3271.865 1046.935 3272.145 10000 ;
      RECT 3269.625 1046.935 3269.905 10000 ;
      RECT 3268.505 1046.935 3268.785 10000 ;
      RECT 3267.385 1046.935 3267.665 10000 ;
      RECT 3252.965 1046.435 3260.805 10000 ;
      RECT 3251.705 1046.935 3251.985 10000 ;
      RECT 3250.585 1046.935 3250.865 10000 ;
      RECT 3249.465 1046.935 3249.745 10000 ;
      RECT 3242.465 1046.935 3244.565 10000 ;
      RECT 3242.605 1046.435 3244.565 10000 ;
      RECT 3241.345 1046.935 3241.625 10000 ;
      RECT 3213.205 1046.435 3238.125 10000 ;
      RECT 3207.465 1046.935 3207.745 10000 ;
      RECT 3206.345 1046.935 3206.625 10000 ;
      RECT 3204.105 1046.935 3204.385 10000 ;
      RECT 3202.985 1046.935 3203.265 10000 ;
      RECT 3201.865 1046.935 3202.145 10000 ;
      RECT 3186.885 1046.435 3199.205 10000 ;
      RECT 3181.705 1046.935 3181.985 10000 ;
      RECT 3180.585 1046.935 3180.865 10000 ;
      RECT 3179.465 1046.935 3179.745 10000 ;
      RECT 3174.425 1046.935 3174.705 10000 ;
      RECT 3134.805 1046.935 3173.585 10000 ;
      RECT 3126.265 1046.935 3126.545 10000 ;
      RECT 3125.145 1046.935 3125.425 10000 ;
      RECT 3122.905 1046.935 3123.185 10000 ;
      RECT 3121.785 1046.935 3122.065 10000 ;
      RECT 3112.265 1046.935 3120.805 10000 ;
      RECT 3112.405 1046.435 3120.805 10000 ;
      RECT 3103.165 1046.935 3105.265 10000 ;
      RECT 3101.905 1046.935 3102.185 10000 ;
      RECT 3100.785 1046.935 3101.065 10000 ;
      RECT 3073.765 1046.435 3098.685 10000 ;
      RECT 3070.265 1046.935 3070.545 10000 ;
      RECT 3069.145 1046.935 3069.425 10000 ;
      RECT 3060.745 1046.935 3061.025 10000 ;
      RECT 3046.745 1046.935 3059.765 10000 ;
      RECT 3046.885 1046.435 3059.765 10000 ;
      RECT 3044.505 1046.935 3044.785 10000 ;
      RECT 3043.385 1046.935 3043.665 10000 ;
      RECT 3042.265 1046.935 3042.545 10000 ;
      RECT 3034.985 1046.935 3035.265 10000 ;
      RECT 2994.805 1046.935 3034.145 10000 ;
      RECT 2993.545 1046.935 2993.825 10000 ;
      RECT 2988.505 1046.935 2988.785 10000 ;
      RECT 2987.385 1046.935 2987.665 10000 ;
      RECT 2972.965 1046.435 2980.805 10000 ;
      RECT 2970.585 1046.935 2970.865 10000 ;
      RECT 2969.465 1046.935 2969.745 10000 ;
      RECT 2967.225 1046.935 2967.505 10000 ;
      RECT 2966.105 1046.935 2966.385 10000 ;
      RECT 2963.165 1046.935 2965.265 10000 ;
      RECT 2933.765 1046.435 2958.685 10000 ;
      RECT 2930.265 1046.935 2930.545 10000 ;
      RECT 2929.145 1046.935 2929.425 10000 ;
      RECT 2928.025 1046.935 2928.305 10000 ;
      RECT 2922.985 1046.935 2923.265 10000 ;
      RECT 2921.865 1046.935 2922.145 10000 ;
      RECT 2907.445 1046.435 2919.765 10000 ;
      RECT 2900.585 1046.935 2900.865 10000 ;
      RECT 2899.465 1046.935 2899.745 10000 ;
      RECT 2897.225 1046.935 2897.505 10000 ;
      RECT 2896.105 1046.935 2896.385 10000 ;
      RECT 2894.985 1046.935 2895.265 10000 ;
      RECT 2854.245 1046.435 2893.445 10000 ;
      RECT 2847.945 1046.935 2848.225 10000 ;
      RECT 2846.825 1046.935 2847.105 10000 ;
      RECT 2845.705 1046.935 2845.985 10000 ;
      RECT 2832.265 1046.935 2840.805 10000 ;
      RECT 2832.405 1046.435 2840.805 10000 ;
      RECT 2831.145 1046.935 2831.425 10000 ;
      RECT 2823.165 1046.435 2824.565 10000 ;
      RECT 2820.785 1046.935 2821.065 10000 ;
      RECT 2819.665 1046.935 2819.945 10000 ;
      RECT 2792.645 1046.435 2818.125 10000 ;
      RECT 2791.385 1046.935 2791.665 10000 ;
      RECT 2790.265 1046.935 2790.545 10000 ;
      RECT 2789.145 1046.935 2789.425 10000 ;
      RECT 2781.865 1046.935 2782.145 10000 ;
      RECT 2780.745 1046.935 2781.025 10000 ;
      RECT 2766.185 1046.935 2779.765 10000 ;
      RECT 2766.325 1046.435 2779.765 10000 ;
      RECT 2761.145 1046.935 2761.425 10000 ;
      RECT 2760.025 1046.935 2760.305 10000 ;
      RECT 2715.365 1046.435 2753.445 10000 ;
      RECT 2712.985 1046.935 2713.265 10000 ;
      RECT 2711.865 1046.935 2712.145 10000 ;
      RECT 2709.625 1046.935 2709.905 10000 ;
      RECT 2708.505 1046.935 2708.785 10000 ;
      RECT 2707.385 1046.935 2707.665 10000 ;
      RECT 2692.965 1046.435 2700.805 10000 ;
      RECT 2691.705 1046.935 2691.985 10000 ;
      RECT 2690.585 1046.935 2690.865 10000 ;
      RECT 2689.465 1046.935 2689.745 10000 ;
      RECT 2682.465 1046.935 2684.565 10000 ;
      RECT 2682.605 1046.435 2684.565 10000 ;
      RECT 2681.345 1046.935 2681.625 10000 ;
      RECT 2653.205 1046.435 2678.125 10000 ;
      RECT 2647.465 1046.935 2647.745 10000 ;
      RECT 2646.345 1046.935 2646.625 10000 ;
      RECT 2644.105 1046.935 2644.385 10000 ;
      RECT 2642.985 1046.935 2643.265 10000 ;
      RECT 2641.865 1046.935 2642.145 10000 ;
      RECT 2626.885 1046.435 2639.205 10000 ;
      RECT 2621.705 1046.935 2621.985 10000 ;
      RECT 2620.585 1046.935 2620.865 10000 ;
      RECT 2619.465 1046.935 2619.745 10000 ;
      RECT 2614.425 1046.935 2614.705 10000 ;
      RECT 2574.805 1046.935 2613.585 10000 ;
      RECT 2566.265 1046.935 2566.545 10000 ;
      RECT 2565.145 1046.935 2565.425 10000 ;
      RECT 2562.905 1046.935 2563.185 10000 ;
      RECT 2561.785 1046.935 2562.065 10000 ;
      RECT 2552.265 1046.935 2560.805 10000 ;
      RECT 2552.405 1046.435 2560.805 10000 ;
      RECT 2543.165 1046.935 2545.265 10000 ;
      RECT 2541.905 1046.935 2542.185 10000 ;
      RECT 2540.785 1046.935 2541.065 10000 ;
      RECT 2513.765 1046.435 2538.685 10000 ;
      RECT 2510.265 1046.935 2510.545 10000 ;
      RECT 2509.145 1046.935 2509.425 10000 ;
      RECT 2500.745 1046.935 2501.025 10000 ;
      RECT 2486.745 1046.935 2499.765 10000 ;
      RECT 2486.885 1046.435 2499.765 10000 ;
      RECT 2484.505 1046.935 2484.785 10000 ;
      RECT 2483.385 1046.935 2483.665 10000 ;
      RECT 2482.265 1046.935 2482.545 10000 ;
      RECT 2474.985 1046.935 2475.265 10000 ;
      RECT 2434.805 1046.935 2474.145 10000 ;
      RECT 2433.545 1046.935 2433.825 10000 ;
      RECT 2428.505 1046.935 2428.785 10000 ;
      RECT 2427.385 1046.935 2427.665 10000 ;
      RECT 2412.965 1046.435 2420.805 10000 ;
      RECT 2410.585 1046.935 2410.865 10000 ;
      RECT 2409.465 1046.935 2409.745 10000 ;
      RECT 2407.225 1046.935 2407.505 10000 ;
      RECT 2406.105 1046.935 2406.385 10000 ;
      RECT 2403.165 1046.935 2405.265 10000 ;
      RECT 2373.765 1046.435 2398.685 10000 ;
      RECT 2370.265 1046.935 2370.545 10000 ;
      RECT 2369.145 1046.935 2369.425 10000 ;
      RECT 2368.025 1046.935 2368.305 10000 ;
      RECT 2362.985 1046.935 2363.265 10000 ;
      RECT 2361.865 1046.935 2362.145 10000 ;
      RECT 2347.445 1046.435 2359.765 10000 ;
      RECT 2340.585 1046.935 2340.865 10000 ;
      RECT 2339.465 1046.935 2339.745 10000 ;
      RECT 2337.225 1046.935 2337.505 10000 ;
      RECT 2336.105 1046.935 2336.385 10000 ;
      RECT 2334.985 1046.935 2335.265 10000 ;
      RECT 2294.245 1046.435 2333.445 10000 ;
      RECT 2287.945 1046.935 2288.225 10000 ;
      RECT 2286.825 1046.935 2287.105 10000 ;
      RECT 2285.705 1046.935 2285.985 10000 ;
      RECT 2272.265 1046.935 2280.805 10000 ;
      RECT 2272.405 1046.435 2280.805 10000 ;
      RECT 2271.145 1046.935 2271.425 10000 ;
      RECT 2263.165 1046.435 2264.565 10000 ;
      RECT 2260.785 1046.935 2261.065 10000 ;
      RECT 2259.665 1046.935 2259.945 10000 ;
      RECT 2232.645 1046.435 2258.125 10000 ;
      RECT 2231.385 1046.935 2231.665 10000 ;
      RECT 2230.265 1046.935 2230.545 10000 ;
      RECT 2229.145 1046.935 2229.425 10000 ;
      RECT 2221.865 1046.935 2222.145 10000 ;
      RECT 2220.745 1046.935 2221.025 10000 ;
      RECT 2206.185 1046.935 2219.765 10000 ;
      RECT 2206.325 1046.435 2219.765 10000 ;
      RECT 2201.145 1046.935 2201.425 10000 ;
      RECT 2200.025 1046.935 2200.305 10000 ;
      RECT 2155.365 1046.435 2193.445 10000 ;
      RECT 2152.985 1046.935 2153.265 10000 ;
      RECT 2151.865 1046.935 2152.145 10000 ;
      RECT 2149.625 1046.935 2149.905 10000 ;
      RECT 2148.505 1046.935 2148.785 10000 ;
      RECT 2147.385 1046.935 2147.665 10000 ;
      RECT 2132.965 1046.435 2140.805 10000 ;
      RECT 2131.705 1046.935 2131.985 10000 ;
      RECT 2130.585 1046.935 2130.865 10000 ;
      RECT 2129.465 1046.935 2129.745 10000 ;
      RECT 2122.465 1046.935 2124.565 10000 ;
      RECT 2122.605 1046.435 2124.565 10000 ;
      RECT 2121.345 1046.935 2121.625 10000 ;
      RECT 2093.205 1046.435 2118.125 10000 ;
      RECT 2087.465 1046.935 2087.745 10000 ;
      RECT 2086.345 1046.935 2086.625 10000 ;
      RECT 2084.105 1046.935 2084.385 10000 ;
      RECT 2082.985 1046.935 2083.265 10000 ;
      RECT 2081.865 1046.935 2082.145 10000 ;
      RECT 2066.885 1046.435 2079.205 10000 ;
      RECT 2061.705 1046.935 2061.985 10000 ;
      RECT 2060.585 1046.935 2060.865 10000 ;
      RECT 2059.465 1046.935 2059.745 10000 ;
      RECT 2054.425 1046.935 2054.705 10000 ;
      RECT 2014.805 1046.935 2053.585 10000 ;
      RECT 2006.265 1046.935 2006.545 10000 ;
      RECT 2005.145 1046.935 2005.425 10000 ;
      RECT 2002.905 1046.935 2003.185 10000 ;
      RECT 2001.785 1046.935 2002.065 10000 ;
      RECT 1992.265 1046.935 2000.805 10000 ;
      RECT 1992.405 1046.435 2000.805 10000 ;
      RECT 1983.165 1046.935 1985.265 10000 ;
      RECT 1981.905 1046.935 1982.185 10000 ;
      RECT 1980.785 1046.935 1981.065 10000 ;
      RECT 1953.765 1046.435 1978.685 10000 ;
      RECT 1950.265 1046.935 1950.545 10000 ;
      RECT 1949.145 1046.935 1949.425 10000 ;
      RECT 1940.745 1046.935 1941.025 10000 ;
      RECT 1926.745 1046.935 1939.765 10000 ;
      RECT 1926.885 1046.435 1939.765 10000 ;
      RECT 1924.505 1046.935 1924.785 10000 ;
      RECT 1923.385 1046.935 1923.665 10000 ;
      RECT 1922.265 1046.935 1922.545 10000 ;
      RECT 1914.985 1046.935 1915.265 10000 ;
      RECT 1874.805 1046.935 1914.145 10000 ;
      RECT 1873.545 1046.935 1873.825 10000 ;
      RECT 1868.505 1046.935 1868.785 10000 ;
      RECT 1867.385 1046.935 1867.665 10000 ;
      RECT 1852.965 1046.435 1860.805 10000 ;
      RECT 1850.585 1046.935 1850.865 10000 ;
      RECT 1849.465 1046.935 1849.745 10000 ;
      RECT 1847.225 1046.935 1847.505 10000 ;
      RECT 1846.105 1046.935 1846.385 10000 ;
      RECT 1843.165 1046.935 1845.265 10000 ;
      RECT 1813.765 1046.435 1838.685 10000 ;
      RECT 1810.265 1046.935 1810.545 10000 ;
      RECT 1809.145 1046.935 1809.425 10000 ;
      RECT 1808.025 1046.935 1808.305 10000 ;
      RECT 1802.985 1046.935 1803.265 10000 ;
      RECT 1801.865 1046.935 1802.145 10000 ;
      RECT 1787.445 1046.435 1799.765 10000 ;
      RECT 1780.585 1046.935 1780.865 10000 ;
      RECT 1779.465 1046.935 1779.745 10000 ;
      RECT 1777.225 1046.935 1777.505 10000 ;
      RECT 1776.105 1046.935 1776.385 10000 ;
      RECT 1774.985 1046.935 1775.265 10000 ;
      RECT 1734.245 1046.435 1773.445 10000 ;
      RECT 1727.945 1046.935 1728.225 10000 ;
      RECT 1726.825 1046.935 1727.105 10000 ;
      RECT 1725.705 1046.935 1725.985 10000 ;
      RECT 1712.265 1046.935 1720.805 10000 ;
      RECT 1712.405 1046.435 1720.805 10000 ;
      RECT 1711.145 1046.935 1711.425 10000 ;
      RECT 1703.165 1046.435 1704.565 10000 ;
      RECT 1700.785 1046.935 1701.065 10000 ;
      RECT 1699.665 1046.935 1699.945 10000 ;
      RECT 1672.645 1046.435 1698.125 10000 ;
      RECT 1671.385 1046.935 1671.665 10000 ;
      RECT 1670.265 1046.935 1670.545 10000 ;
      RECT 1669.145 1046.935 1669.425 10000 ;
      RECT 1661.865 1046.935 1662.145 10000 ;
      RECT 1660.745 1046.935 1661.025 10000 ;
      RECT 1646.185 1046.935 1659.765 10000 ;
      RECT 1646.325 1046.435 1659.765 10000 ;
      RECT 1641.145 1046.935 1641.425 10000 ;
      RECT 1640.025 1046.935 1640.305 10000 ;
      RECT 1595.365 1046.435 1633.445 10000 ;
      RECT 1592.985 1046.935 1593.265 10000 ;
      RECT 1591.865 1046.935 1592.145 10000 ;
      RECT 1589.625 1046.935 1589.905 10000 ;
      RECT 1588.505 1046.935 1588.785 10000 ;
      RECT 1587.385 1046.935 1587.665 10000 ;
      RECT 1572.965 1046.435 1580.805 10000 ;
      RECT 1571.705 1046.935 1571.985 10000 ;
      RECT 1570.585 1046.935 1570.865 10000 ;
      RECT 1569.465 1046.935 1569.745 10000 ;
      RECT 1562.465 1046.935 1564.565 10000 ;
      RECT 1562.605 1046.435 1564.565 10000 ;
      RECT 1561.345 1046.935 1561.625 10000 ;
      RECT 1533.205 1046.435 1558.125 10000 ;
      RECT 1527.465 1046.935 1527.745 10000 ;
      RECT 1526.345 1046.935 1526.625 10000 ;
      RECT 1524.105 1046.935 1524.385 10000 ;
      RECT 1522.985 1046.935 1523.265 10000 ;
      RECT 1521.865 1046.935 1522.145 10000 ;
      RECT 1506.885 1046.435 1519.205 10000 ;
      RECT 1501.705 1046.935 1501.985 10000 ;
      RECT 1500.585 1046.935 1500.865 10000 ;
      RECT 1499.465 1046.935 1499.745 10000 ;
      RECT 1494.425 1046.935 1494.705 10000 ;
      RECT 1454.805 1046.935 1493.585 10000 ;
      RECT 1446.265 1046.935 1446.545 10000 ;
      RECT 1445.145 1046.935 1445.425 10000 ;
      RECT 1442.905 1046.935 1443.185 10000 ;
      RECT 1441.785 1046.935 1442.065 10000 ;
      RECT 1432.265 1046.935 1440.805 10000 ;
      RECT 1432.405 1046.435 1440.805 10000 ;
      RECT 1423.165 1046.935 1425.265 10000 ;
      RECT 1421.905 1046.935 1422.185 10000 ;
      RECT 1420.785 1046.935 1421.065 10000 ;
      RECT 1393.765 1046.435 1418.685 10000 ;
      RECT 1390.265 1046.935 1390.545 10000 ;
      RECT 1389.145 1046.935 1389.425 10000 ;
      RECT 1380.745 1046.935 1381.025 10000 ;
      RECT 1366.745 1046.935 1379.765 10000 ;
      RECT 1366.885 1046.435 1379.765 10000 ;
      RECT 1364.505 1046.935 1364.785 10000 ;
      RECT 1363.385 1046.935 1363.665 10000 ;
      RECT 1362.265 1046.935 1362.545 10000 ;
      RECT 1354.985 1046.935 1355.265 10000 ;
      RECT 1314.805 1046.935 1354.145 10000 ;
      RECT 1313.545 1046.935 1313.825 10000 ;
      RECT 1308.505 1046.935 1308.785 10000 ;
      RECT 1307.385 1046.935 1307.665 10000 ;
      RECT 1292.965 1046.435 1300.805 10000 ;
      RECT 1290.585 1046.935 1290.865 10000 ;
      RECT 1289.465 1046.935 1289.745 10000 ;
      RECT 1287.225 1046.935 1287.505 10000 ;
      RECT 1286.105 1046.935 1286.385 10000 ;
      RECT 1283.165 1046.935 1285.265 10000 ;
      RECT 1253.765 1046.435 1278.685 10000 ;
      RECT 1250.265 1046.935 1250.545 10000 ;
      RECT 1249.145 1046.935 1249.425 10000 ;
      RECT 1248.025 1046.935 1248.305 10000 ;
      RECT 1242.985 1046.935 1243.265 10000 ;
      RECT 1241.865 1046.935 1242.145 10000 ;
      RECT 1227.445 1046.435 1239.765 10000 ;
      RECT 1220.585 1046.935 1220.865 10000 ;
      RECT 1219.465 1046.935 1219.745 10000 ;
      RECT 1217.225 1046.935 1217.505 10000 ;
      RECT 1216.105 1046.935 1216.385 10000 ;
      RECT 1214.985 1046.935 1215.265 10000 ;
      RECT 1174.245 1046.435 1213.445 10000 ;
      RECT 1167.945 1046.935 1168.225 10000 ;
      RECT 1166.825 1046.935 1167.105 10000 ;
      RECT 1165.705 1046.935 1165.985 10000 ;
      RECT 1152.265 1046.935 1160.805 10000 ;
      RECT 1152.405 1046.435 1160.805 10000 ;
      RECT 1151.145 1046.935 1151.425 10000 ;
      RECT 1143.165 1046.435 1144.565 10000 ;
      RECT 1140.785 1046.935 1141.065 10000 ;
      RECT 1139.665 1046.935 1139.945 10000 ;
      RECT 998.1 1046.435 1137.565 10000 ;
      RECT 7614.805 1046.435 7653.445 10000 ;
      RECT 7583.165 1046.435 7585.125 10000 ;
      RECT 7474.805 1046.435 7514.005 10000 ;
      RECT 7443.165 1046.435 7445.125 10000 ;
      RECT 7054.805 1046.435 7093.445 10000 ;
      RECT 7023.165 1046.435 7025.125 10000 ;
      RECT 6914.805 1046.435 6954.005 10000 ;
      RECT 6883.165 1046.435 6885.125 10000 ;
      RECT 6494.805 1046.435 6533.445 10000 ;
      RECT 6463.165 1046.435 6465.125 10000 ;
      RECT 6354.805 1046.435 6394.005 10000 ;
      RECT 6323.165 1046.435 6325.125 10000 ;
      RECT 5934.805 1046.435 5973.445 10000 ;
      RECT 5903.165 1046.435 5905.125 10000 ;
      RECT 5794.805 1046.435 5834.005 10000 ;
      RECT 5763.165 1046.435 5765.125 10000 ;
      RECT 5374.805 1046.435 5413.445 10000 ;
      RECT 5343.165 1046.435 5345.125 10000 ;
      RECT 5234.805 1046.435 5274.005 10000 ;
      RECT 5203.165 1046.435 5205.125 10000 ;
      RECT 4814.805 1046.435 4853.445 10000 ;
      RECT 4783.165 1046.435 4785.125 10000 ;
      RECT 4674.805 1046.435 4714.005 10000 ;
      RECT 4643.165 1046.435 4645.125 10000 ;
      RECT 4254.805 1046.435 4293.445 10000 ;
      RECT 4223.165 1046.435 4225.125 10000 ;
      RECT 4114.805 1046.435 4154.005 10000 ;
      RECT 4083.165 1046.435 4085.125 10000 ;
      RECT 3694.805 1046.435 3733.445 10000 ;
      RECT 3663.165 1046.435 3665.125 10000 ;
      RECT 3554.805 1046.435 3594.005 10000 ;
      RECT 3523.165 1046.435 3525.125 10000 ;
      RECT 3134.805 1046.435 3173.445 10000 ;
      RECT 3103.165 1046.435 3105.125 10000 ;
      RECT 2994.805 1046.435 3034.005 10000 ;
      RECT 2963.165 1046.435 2965.125 10000 ;
      RECT 2574.805 1046.435 2613.445 10000 ;
      RECT 2543.165 1046.435 2545.125 10000 ;
      RECT 2434.805 1046.435 2474.005 10000 ;
      RECT 2403.165 1046.435 2405.125 10000 ;
      RECT 2014.805 1046.435 2053.445 10000 ;
      RECT 1983.165 1046.435 1985.125 10000 ;
      RECT 1874.805 1046.435 1914.005 10000 ;
      RECT 1843.165 1046.435 1845.125 10000 ;
      RECT 1454.805 1046.435 1493.445 10000 ;
      RECT 1423.165 1046.435 1425.125 10000 ;
      RECT 1314.805 1046.435 1354.005 10000 ;
      RECT 1283.165 1046.435 1285.125 10000 ;
    LAYER M5 ;
      RECT 4.1 9990 20195.9 9995.9 ;
      RECT 20190 4.1 20195.9 9995.9 ;
      RECT 4.1 4.1 10 9995.9 ;
      RECT 4.1 4.1 20195.9 10 ;
      RECT 19160.9 1118.985 19167.9 1120.185 ;
      RECT 19158.16 1119.19 19167.9 1119.99 ;
      RECT 19160.9 1121.385 19167.9 1122.585 ;
      RECT 19158.16 1121.59 19167.9 1122.39 ;
      RECT 19160.9 1123.785 19167.9 1124.985 ;
      RECT 19158.16 1123.99 19167.9 1124.79 ;
      RECT 19160.9 1126.185 19167.9 1127.385 ;
      RECT 19158.16 1126.39 19167.9 1127.19 ;
      RECT 19033.5 1166.44 19040.475 1188.44 ;
      RECT 19040.475 1127.265 19046.5 1180.44 ;
      RECT 19033.5 1048.035 19035.565 1188.44 ;
      RECT 19033.5 1127.265 19046.5 1150.07 ;
      RECT 19033.5 1087.44 19039.865 1150.07 ;
      RECT 19033.5 1087.44 19046.5 1094.78 ;
      RECT 19042.56 1048.035 19046.5 1094.78 ;
      RECT 19040.475 1053.41 19046.5 1094.78 ;
      RECT 19033.5 1053.41 19046.5 1071.07 ;
      RECT 19033.5 1048.035 19039.07 1071.07 ;
      RECT 19033.5 1048.035 19046.5 1049.11 ;
      RECT 19016.52 1166.44 19029.52 1209.16 ;
      RECT 19018.145 1048.035 19029.52 1209.16 ;
      RECT 19016.52 1087.44 19029.52 1150.07 ;
      RECT 19016.52 1048.035 19029.52 1071.07 ;
      RECT 18986 1183.44 19014 1209.16 ;
      RECT 18992.145 1048.035 19008.565 1209.16 ;
      RECT 18986 1070.44 18987.235 1209.16 ;
      RECT 18986 1070.44 19013.235 1167.07 ;
      RECT 18986 1087.44 19014 1150.07 ;
      RECT 18988.365 1048.035 19008.565 1167.07 ;
      RECT 18986 1048.035 19014 1054.07 ;
      RECT 18970.48 1087.44 18983.48 1209.16 ;
      RECT 18970.48 1048.035 18976.835 1209.16 ;
      RECT 18970.48 1048.035 18983.48 1071.07 ;
      RECT 18953.5 1149.44 18966.5 1189.16 ;
      RECT 18964.63 1048.035 18966.5 1189.16 ;
      RECT 18962.865 1053.42 18966.5 1189.16 ;
      RECT 18953.5 1048.035 18955.115 1189.16 ;
      RECT 18953.5 1053.42 18966.5 1118.87 ;
      RECT 18953.5 1048.035 18961.85 1118.87 ;
      RECT 18953.5 1048.035 18966.5 1049.12 ;
      RECT 18936.52 1070.44 18949.52 1209.16 ;
      RECT 18936.865 1048.035 18949.52 1209.16 ;
      RECT 18936.52 1048.035 18949.52 1054.07 ;
      RECT 18906 1118.44 18934 1209.16 ;
      RECT 18918.375 1070.44 18934 1209.16 ;
      RECT 18906 1048.035 18910.625 1209.16 ;
      RECT 18906 1048.035 18931.955 1087.87 ;
      RECT 18906 1048.035 18934 1054.07 ;
      RECT 18890.48 1166.44 18903.48 1209.16 ;
      RECT 18900.475 1053.365 18903.48 1209.16 ;
      RECT 18890.48 1048.035 18895.565 1209.16 ;
      RECT 18890.48 1087.44 18903.48 1150.07 ;
      RECT 18890.48 1053.365 18903.48 1071.07 ;
      RECT 18890.48 1048.035 18898.81 1071.07 ;
      RECT 18890.48 1048.035 18903.48 1049.165 ;
      RECT 18873.5 1166.44 18886.5 1189.16 ;
      RECT 18878.145 1048.035 18886.5 1189.16 ;
      RECT 18877.98 1087.44 18886.5 1189.16 ;
      RECT 18873.5 1087.44 18886.5 1150.07 ;
      RECT 18873.5 1048.035 18886.5 1071.07 ;
      RECT 18856.52 1183.44 18869.52 1209.16 ;
      RECT 18856.52 1048.035 18868.565 1209.16 ;
      RECT 18856.52 1070.44 18869.52 1167.07 ;
      RECT 18856.52 1048.035 18869.52 1054.07 ;
      RECT 18826 1183.44 18854 1209.16 ;
      RECT 18852.145 1048.035 18854 1209.16 ;
      RECT 18826 1087.44 18847.235 1209.16 ;
      RECT 18849.555 1048.035 18854 1167.07 ;
      RECT 18832.55 1070.44 18854 1167.07 ;
      RECT 18826 1048.035 18844.645 1071.07 ;
      RECT 18826 1048.035 18854 1054.07 ;
      RECT 18810.48 1149.44 18823.48 1209.16 ;
      RECT 18822.865 1053.415 18823.48 1209.16 ;
      RECT 18810.48 1048.035 18815.115 1209.16 ;
      RECT 18810.48 1053.415 18823.48 1118.87 ;
      RECT 18810.48 1048.035 18821.85 1118.87 ;
      RECT 18810.48 1048.035 18823.48 1049.12 ;
      RECT 18793.5 1070.44 18806.5 1189.16 ;
      RECT 18796.865 1048.035 18806.5 1189.16 ;
      RECT 18793.5 1048.035 18806.5 1054.07 ;
      RECT 18776.52 1118.44 18789.52 1209.16 ;
      RECT 18778.375 1048.035 18789.52 1209.16 ;
      RECT 18776.52 1048.035 18789.52 1087.87 ;
      RECT 18746 1166.44 18774 1209.16 ;
      RECT 18760.475 1118.44 18774 1209.16 ;
      RECT 18746 1048.035 18755.565 1209.16 ;
      RECT 18746 1087.44 18770.625 1150.07 ;
      RECT 18764.53 1048.035 18774 1087.87 ;
      RECT 18760.475 1053.365 18774 1087.87 ;
      RECT 18746 1053.365 18774 1071.07 ;
      RECT 18746 1048.035 18758.81 1071.07 ;
      RECT 18746 1048.035 18774 1049.165 ;
      RECT 18730.48 1183.44 18743.48 1209.16 ;
      RECT 18738.145 1048.035 18743.48 1209.16 ;
      RECT 18733.475 1166.44 18743.48 1209.16 ;
      RECT 18730.48 1166.44 18743.48 1167.07 ;
      RECT 18730.48 1070.44 18733.235 1167.07 ;
      RECT 18730.48 1087.44 18743.48 1150.07 ;
      RECT 18730.48 1070.44 18743.48 1071.07 ;
      RECT 18733.475 1048.035 18743.48 1071.07 ;
      RECT 18730.48 1048.035 18743.48 1054.07 ;
      RECT 18696.52 1183.44 18709.52 1209.16 ;
      RECT 18696.52 1087.44 18707.235 1209.16 ;
      RECT 18701.75 1070.44 18709.52 1167.07 ;
      RECT 18696.52 1048.035 18704.565 1071.07 ;
      RECT 18696.52 1048.035 18709.52 1054.07 ;
      RECT 18666 1149.44 18694 1209.16 ;
      RECT 18684.63 1048.035 18694 1209.16 ;
      RECT 18682.865 1053.42 18694 1209.16 ;
      RECT 18666 1048.035 18675.115 1209.16 ;
      RECT 18666 1053.42 18694 1118.87 ;
      RECT 18666 1048.035 18681.85 1118.87 ;
      RECT 18666 1048.035 18694 1049.12 ;
      RECT 18650.48 1070.44 18663.48 1209.16 ;
      RECT 18656.865 1048.035 18663.48 1209.16 ;
      RECT 18650.48 1048.035 18651.955 1209.16 ;
      RECT 18650.48 1048.035 18663.48 1054.07 ;
      RECT 18633.5 1118.44 18646.5 1189.16 ;
      RECT 18638.375 1048.035 18646.5 1189.16 ;
      RECT 18633.5 1048.035 18646.5 1087.87 ;
      RECT 18616.52 1166.44 18629.52 1209.16 ;
      RECT 18624.53 1048.035 18629.52 1209.16 ;
      RECT 18620.475 1053.365 18629.52 1209.16 ;
      RECT 18616.52 1087.44 18629.52 1150.07 ;
      RECT 18616.52 1053.365 18629.52 1071.07 ;
      RECT 18616.52 1048.035 18618.81 1071.07 ;
      RECT 18616.52 1048.035 18629.52 1049.375 ;
      RECT 18586 1183.44 18614 1209.16 ;
      RECT 18598.145 1048.035 18614 1209.16 ;
      RECT 18593.475 1166.44 18614 1209.16 ;
      RECT 18586 1048.035 18588.565 1209.16 ;
      RECT 18586 1166.44 18614 1167.07 ;
      RECT 18586 1070.44 18593.235 1167.07 ;
      RECT 18586 1087.44 18614 1150.07 ;
      RECT 18586 1070.44 18614 1071.07 ;
      RECT 18593.475 1048.035 18614 1071.07 ;
      RECT 18586 1048.035 18614 1054.07 ;
      RECT 18570.48 1183.44 18583.48 1209.16 ;
      RECT 18572.145 1048.035 18583.48 1209.16 ;
      RECT 18570.48 1048.035 18583.48 1167.07 ;
      RECT 18553.5 1087.44 18566.5 1189.16 ;
      RECT 18560.13 1070.44 18566.5 1189.16 ;
      RECT 18553.5 1048.035 18563.455 1071.07 ;
      RECT 18553.5 1048.035 18566.5 1054.07 ;
      RECT 18536.52 1149.44 18549.52 1209.16 ;
      RECT 18544.63 1048.035 18549.52 1209.16 ;
      RECT 18542.865 1053.42 18549.52 1209.16 ;
      RECT 18536.52 1053.42 18549.52 1118.87 ;
      RECT 18536.52 1048.035 18541.85 1118.87 ;
      RECT 18536.52 1048.035 18549.52 1049.12 ;
      RECT 18506 1070.44 18534 1209.16 ;
      RECT 18516.865 1048.035 18534 1209.16 ;
      RECT 18506 1048.035 18511.955 1209.16 ;
      RECT 18506 1048.035 18534 1054.07 ;
      RECT 18490.48 1118.44 18503.48 1209.16 ;
      RECT 18498.375 1048.035 18503.48 1209.16 ;
      RECT 18490.48 1048.035 18503.48 1087.87 ;
      RECT 18473.5 1166.44 18486.5 1189.16 ;
      RECT 18484.43 1048.035 18486.5 1189.16 ;
      RECT 18480.475 1053.365 18486.5 1189.16 ;
      RECT 18473.5 1048.035 18475.565 1189.16 ;
      RECT 18473.5 1087.44 18486.5 1150.07 ;
      RECT 18473.5 1053.365 18486.5 1071.07 ;
      RECT 18473.5 1048.035 18478.81 1071.07 ;
      RECT 18473.5 1048.035 18486.5 1049.165 ;
      RECT 18456.52 1166.44 18469.52 1209.16 ;
      RECT 18458.145 1048.035 18469.52 1209.16 ;
      RECT 18456.52 1087.44 18469.52 1150.07 ;
      RECT 18456.52 1048.035 18469.52 1071.07 ;
      RECT 18426 1183.44 18454 1209.16 ;
      RECT 18432.145 1048.035 18448.565 1209.16 ;
      RECT 18426 1070.44 18427.235 1209.16 ;
      RECT 18426 1070.44 18453.235 1167.07 ;
      RECT 18426 1087.44 18454 1150.07 ;
      RECT 18428.365 1048.035 18448.565 1167.07 ;
      RECT 18426 1048.035 18454 1054.07 ;
      RECT 18410.48 1087.44 18423.48 1209.16 ;
      RECT 18410.48 1048.035 18416.835 1209.16 ;
      RECT 18410.48 1048.035 18423.48 1071.07 ;
      RECT 18393.5 1149.44 18406.5 1189.16 ;
      RECT 18404.63 1048.035 18406.5 1189.16 ;
      RECT 18402.865 1053.42 18406.5 1189.16 ;
      RECT 18393.5 1048.035 18395.115 1189.16 ;
      RECT 18393.5 1053.42 18406.5 1118.87 ;
      RECT 18393.5 1048.035 18401.85 1118.87 ;
      RECT 18393.5 1048.035 18406.5 1049.12 ;
      RECT 18376.52 1070.44 18389.52 1209.16 ;
      RECT 18376.865 1048.035 18389.52 1209.16 ;
      RECT 18376.52 1048.035 18389.52 1054.07 ;
      RECT 18346 1118.44 18374 1209.16 ;
      RECT 18358.375 1070.44 18374 1209.16 ;
      RECT 18346 1048.035 18350.625 1209.16 ;
      RECT 18346 1048.035 18371.955 1087.87 ;
      RECT 18346 1048.035 18374 1054.07 ;
      RECT 18330.48 1166.44 18343.48 1209.16 ;
      RECT 18340.475 1053.365 18343.48 1209.16 ;
      RECT 18330.48 1048.035 18335.565 1209.16 ;
      RECT 18330.48 1087.44 18343.48 1150.07 ;
      RECT 18330.48 1053.365 18343.48 1071.07 ;
      RECT 18330.48 1048.035 18338.81 1071.07 ;
      RECT 18330.48 1048.035 18343.48 1049.165 ;
      RECT 18313.5 1166.44 18326.5 1189.16 ;
      RECT 18318.145 1048.035 18326.5 1189.16 ;
      RECT 18317.98 1087.44 18326.5 1189.16 ;
      RECT 18313.5 1087.44 18326.5 1150.07 ;
      RECT 18313.5 1048.035 18326.5 1071.07 ;
      RECT 18296.52 1183.44 18309.52 1209.16 ;
      RECT 18296.52 1048.035 18308.565 1209.16 ;
      RECT 18296.52 1070.44 18309.52 1167.07 ;
      RECT 18296.52 1048.035 18309.52 1054.07 ;
      RECT 18266 1183.44 18294 1209.16 ;
      RECT 18292.145 1048.035 18294 1209.16 ;
      RECT 18266 1087.44 18287.235 1209.16 ;
      RECT 18289.555 1048.035 18294 1167.07 ;
      RECT 18272.55 1070.44 18294 1167.07 ;
      RECT 18266 1048.035 18284.645 1071.07 ;
      RECT 18266 1048.035 18294 1054.07 ;
      RECT 18250.48 1149.44 18263.48 1209.16 ;
      RECT 18262.865 1053.415 18263.48 1209.16 ;
      RECT 18250.48 1048.035 18255.115 1209.16 ;
      RECT 18250.48 1053.415 18263.48 1118.87 ;
      RECT 18250.48 1048.035 18261.85 1118.87 ;
      RECT 18250.48 1048.035 18263.48 1049.12 ;
      RECT 18233.5 1070.44 18246.5 1189.16 ;
      RECT 18236.865 1048.035 18246.5 1189.16 ;
      RECT 18233.5 1048.035 18246.5 1054.07 ;
      RECT 18216.52 1118.44 18229.52 1209.16 ;
      RECT 18218.375 1048.035 18229.52 1209.16 ;
      RECT 18216.52 1048.035 18229.52 1087.87 ;
      RECT 18186 1166.44 18214 1209.16 ;
      RECT 18200.475 1118.44 18214 1209.16 ;
      RECT 18186 1048.035 18195.565 1209.16 ;
      RECT 18186 1087.44 18210.625 1150.07 ;
      RECT 18204.53 1048.035 18214 1087.87 ;
      RECT 18200.475 1053.365 18214 1087.87 ;
      RECT 18186 1053.365 18214 1071.07 ;
      RECT 18186 1048.035 18198.81 1071.07 ;
      RECT 18186 1048.035 18214 1049.165 ;
      RECT 18170.48 1183.44 18183.48 1209.16 ;
      RECT 18178.145 1048.035 18183.48 1209.16 ;
      RECT 18173.475 1166.44 18183.48 1209.16 ;
      RECT 18170.48 1166.44 18183.48 1167.07 ;
      RECT 18170.48 1070.44 18173.235 1167.07 ;
      RECT 18170.48 1087.44 18183.48 1150.07 ;
      RECT 18170.48 1070.44 18183.48 1071.07 ;
      RECT 18173.475 1048.035 18183.48 1071.07 ;
      RECT 18170.48 1048.035 18183.48 1054.07 ;
      RECT 18136.52 1183.44 18149.52 1209.16 ;
      RECT 18136.52 1087.44 18147.235 1209.16 ;
      RECT 18141.75 1070.44 18149.52 1167.07 ;
      RECT 18136.52 1048.035 18144.565 1071.07 ;
      RECT 18136.52 1048.035 18149.52 1054.07 ;
      RECT 18106 1149.44 18134 1209.16 ;
      RECT 18124.63 1048.035 18134 1209.16 ;
      RECT 18122.865 1053.42 18134 1209.16 ;
      RECT 18106 1048.035 18115.115 1209.16 ;
      RECT 18106 1053.42 18134 1118.87 ;
      RECT 18106 1048.035 18121.85 1118.87 ;
      RECT 18106 1048.035 18134 1049.12 ;
      RECT 18090.48 1070.44 18103.48 1209.16 ;
      RECT 18096.865 1048.035 18103.48 1209.16 ;
      RECT 18090.48 1048.035 18091.955 1209.16 ;
      RECT 18090.48 1048.035 18103.48 1054.07 ;
      RECT 18073.5 1118.44 18086.5 1189.16 ;
      RECT 18078.375 1048.035 18086.5 1189.16 ;
      RECT 18073.5 1048.035 18086.5 1087.87 ;
      RECT 18056.52 1166.44 18069.52 1209.16 ;
      RECT 18064.53 1048.035 18069.52 1209.16 ;
      RECT 18060.475 1053.365 18069.52 1209.16 ;
      RECT 18056.52 1087.44 18069.52 1150.07 ;
      RECT 18056.52 1053.365 18069.52 1071.07 ;
      RECT 18056.52 1048.035 18058.81 1071.07 ;
      RECT 18056.52 1048.035 18069.52 1049.375 ;
      RECT 18026 1183.44 18054 1209.16 ;
      RECT 18038.145 1048.035 18054 1209.16 ;
      RECT 18033.475 1166.44 18054 1209.16 ;
      RECT 18026 1048.035 18028.565 1209.16 ;
      RECT 18026 1166.44 18054 1167.07 ;
      RECT 18026 1070.44 18033.235 1167.07 ;
      RECT 18026 1087.44 18054 1150.07 ;
      RECT 18026 1070.44 18054 1071.07 ;
      RECT 18033.475 1048.035 18054 1071.07 ;
      RECT 18026 1048.035 18054 1054.07 ;
      RECT 18010.48 1183.44 18023.48 1209.16 ;
      RECT 18012.145 1048.035 18023.48 1209.16 ;
      RECT 18010.48 1048.035 18023.48 1167.07 ;
      RECT 17993.5 1087.44 18006.5 1189.16 ;
      RECT 18000.13 1070.44 18006.5 1189.16 ;
      RECT 17993.5 1048.035 18003.455 1071.07 ;
      RECT 17993.5 1048.035 18006.5 1054.07 ;
      RECT 17976.52 1149.44 17989.52 1209.16 ;
      RECT 17984.63 1048.035 17989.52 1209.16 ;
      RECT 17982.865 1053.42 17989.52 1209.16 ;
      RECT 17976.52 1053.42 17989.52 1118.87 ;
      RECT 17976.52 1048.035 17981.85 1118.87 ;
      RECT 17976.52 1048.035 17989.52 1049.12 ;
      RECT 17946 1070.44 17974 1209.16 ;
      RECT 17956.865 1048.035 17974 1209.16 ;
      RECT 17946 1048.035 17951.955 1209.16 ;
      RECT 17946 1048.035 17974 1054.07 ;
      RECT 17930.48 1118.44 17943.48 1209.16 ;
      RECT 17938.375 1048.035 17943.48 1209.16 ;
      RECT 17930.48 1048.035 17943.48 1087.87 ;
      RECT 17913.5 1166.44 17926.5 1189.16 ;
      RECT 17924.43 1048.035 17926.5 1189.16 ;
      RECT 17920.475 1053.365 17926.5 1189.16 ;
      RECT 17913.5 1048.035 17915.565 1189.16 ;
      RECT 17913.5 1087.44 17926.5 1150.07 ;
      RECT 17913.5 1053.365 17926.5 1071.07 ;
      RECT 17913.5 1048.035 17918.81 1071.07 ;
      RECT 17913.5 1048.035 17926.5 1049.165 ;
      RECT 17896.52 1166.44 17909.52 1209.16 ;
      RECT 17898.145 1048.035 17909.52 1209.16 ;
      RECT 17896.52 1087.44 17909.52 1150.07 ;
      RECT 17896.52 1048.035 17909.52 1071.07 ;
      RECT 17866 1183.44 17894 1209.16 ;
      RECT 17872.145 1048.035 17888.565 1209.16 ;
      RECT 17866 1070.44 17867.235 1209.16 ;
      RECT 17866 1070.44 17893.235 1167.07 ;
      RECT 17866 1087.44 17894 1150.07 ;
      RECT 17868.365 1048.035 17888.565 1167.07 ;
      RECT 17866 1048.035 17894 1054.07 ;
      RECT 17850.48 1087.44 17863.48 1209.16 ;
      RECT 17850.48 1048.035 17856.835 1209.16 ;
      RECT 17850.48 1048.035 17863.48 1071.07 ;
      RECT 17833.5 1149.44 17846.5 1189.16 ;
      RECT 17844.63 1048.035 17846.5 1189.16 ;
      RECT 17842.865 1053.42 17846.5 1189.16 ;
      RECT 17833.5 1048.035 17835.115 1189.16 ;
      RECT 17833.5 1053.42 17846.5 1118.87 ;
      RECT 17833.5 1048.035 17841.85 1118.87 ;
      RECT 17833.5 1048.035 17846.5 1049.12 ;
      RECT 17816.52 1070.44 17829.52 1209.16 ;
      RECT 17816.865 1048.035 17829.52 1209.16 ;
      RECT 17816.52 1048.035 17829.52 1054.07 ;
      RECT 17786 1118.44 17814 1209.16 ;
      RECT 17798.375 1070.44 17814 1209.16 ;
      RECT 17786 1048.035 17790.625 1209.16 ;
      RECT 17786 1048.035 17811.955 1087.87 ;
      RECT 17786 1048.035 17814 1054.07 ;
      RECT 17770.48 1166.44 17783.48 1209.16 ;
      RECT 17780.475 1053.365 17783.48 1209.16 ;
      RECT 17770.48 1048.035 17775.565 1209.16 ;
      RECT 17770.48 1087.44 17783.48 1150.07 ;
      RECT 17770.48 1053.365 17783.48 1071.07 ;
      RECT 17770.48 1048.035 17778.81 1071.07 ;
      RECT 17770.48 1048.035 17783.48 1049.165 ;
      RECT 17753.5 1166.44 17766.5 1189.16 ;
      RECT 17758.145 1048.035 17766.5 1189.16 ;
      RECT 17757.98 1087.44 17766.5 1189.16 ;
      RECT 17753.5 1087.44 17766.5 1150.07 ;
      RECT 17753.5 1048.035 17766.5 1071.07 ;
      RECT 17736.52 1183.44 17749.52 1209.16 ;
      RECT 17736.52 1048.035 17748.565 1209.16 ;
      RECT 17736.52 1070.44 17749.52 1167.07 ;
      RECT 17736.52 1048.035 17749.52 1054.07 ;
      RECT 17706 1183.44 17734 1209.16 ;
      RECT 17732.145 1048.035 17734 1209.16 ;
      RECT 17706 1087.44 17727.235 1209.16 ;
      RECT 17729.555 1048.035 17734 1167.07 ;
      RECT 17712.55 1070.44 17734 1167.07 ;
      RECT 17706 1048.035 17724.645 1071.07 ;
      RECT 17706 1048.035 17734 1054.07 ;
      RECT 17690.48 1149.44 17703.48 1209.16 ;
      RECT 17702.865 1053.415 17703.48 1209.16 ;
      RECT 17690.48 1048.035 17695.115 1209.16 ;
      RECT 17690.48 1053.415 17703.48 1118.87 ;
      RECT 17690.48 1048.035 17701.85 1118.87 ;
      RECT 17690.48 1048.035 17703.48 1049.12 ;
      RECT 17673.5 1070.44 17686.5 1189.16 ;
      RECT 17676.865 1048.035 17686.5 1189.16 ;
      RECT 17673.5 1048.035 17686.5 1054.07 ;
      RECT 17656.52 1118.44 17669.52 1209.16 ;
      RECT 17658.375 1048.035 17669.52 1209.16 ;
      RECT 17656.52 1048.035 17669.52 1087.87 ;
      RECT 17626 1166.44 17654 1209.16 ;
      RECT 17640.475 1118.44 17654 1209.16 ;
      RECT 17626 1048.035 17635.565 1209.16 ;
      RECT 17626 1087.44 17650.625 1150.07 ;
      RECT 17644.53 1048.035 17654 1087.87 ;
      RECT 17640.475 1053.365 17654 1087.87 ;
      RECT 17626 1053.365 17654 1071.07 ;
      RECT 17626 1048.035 17638.81 1071.07 ;
      RECT 17626 1048.035 17654 1049.165 ;
      RECT 17610.48 1183.44 17623.48 1209.16 ;
      RECT 17618.145 1048.035 17623.48 1209.16 ;
      RECT 17613.475 1166.44 17623.48 1209.16 ;
      RECT 17610.48 1166.44 17623.48 1167.07 ;
      RECT 17610.48 1070.44 17613.235 1167.07 ;
      RECT 17610.48 1087.44 17623.48 1150.07 ;
      RECT 17610.48 1070.44 17623.48 1071.07 ;
      RECT 17613.475 1048.035 17623.48 1071.07 ;
      RECT 17610.48 1048.035 17623.48 1054.07 ;
      RECT 17576.52 1183.44 17589.52 1209.16 ;
      RECT 17576.52 1087.44 17587.235 1209.16 ;
      RECT 17581.75 1070.44 17589.52 1167.07 ;
      RECT 17576.52 1048.035 17584.565 1071.07 ;
      RECT 17576.52 1048.035 17589.52 1054.07 ;
      RECT 17546 1149.44 17574 1209.16 ;
      RECT 17564.63 1048.035 17574 1209.16 ;
      RECT 17562.865 1053.42 17574 1209.16 ;
      RECT 17546 1048.035 17555.115 1209.16 ;
      RECT 17546 1053.42 17574 1118.87 ;
      RECT 17546 1048.035 17561.85 1118.87 ;
      RECT 17546 1048.035 17574 1049.12 ;
      RECT 17530.48 1070.44 17543.48 1209.16 ;
      RECT 17536.865 1048.035 17543.48 1209.16 ;
      RECT 17530.48 1048.035 17531.955 1209.16 ;
      RECT 17530.48 1048.035 17543.48 1054.07 ;
      RECT 17513.5 1118.44 17526.5 1189.16 ;
      RECT 17518.375 1048.035 17526.5 1189.16 ;
      RECT 17513.5 1048.035 17526.5 1087.87 ;
      RECT 17496.52 1166.44 17509.52 1209.16 ;
      RECT 17504.53 1048.035 17509.52 1209.16 ;
      RECT 17500.475 1053.365 17509.52 1209.16 ;
      RECT 17496.52 1087.44 17509.52 1150.07 ;
      RECT 17496.52 1053.365 17509.52 1071.07 ;
      RECT 17496.52 1048.035 17498.81 1071.07 ;
      RECT 17496.52 1048.035 17509.52 1049.375 ;
      RECT 17466 1183.44 17494 1209.16 ;
      RECT 17478.145 1048.035 17494 1209.16 ;
      RECT 17473.475 1166.44 17494 1209.16 ;
      RECT 17466 1048.035 17468.565 1209.16 ;
      RECT 17466 1166.44 17494 1167.07 ;
      RECT 17466 1070.44 17473.235 1167.07 ;
      RECT 17466 1087.44 17494 1150.07 ;
      RECT 17466 1070.44 17494 1071.07 ;
      RECT 17473.475 1048.035 17494 1071.07 ;
      RECT 17466 1048.035 17494 1054.07 ;
      RECT 17450.48 1183.44 17463.48 1209.16 ;
      RECT 17452.145 1048.035 17463.48 1209.16 ;
      RECT 17450.48 1048.035 17463.48 1167.07 ;
      RECT 17433.5 1087.44 17446.5 1189.16 ;
      RECT 17440.13 1070.44 17446.5 1189.16 ;
      RECT 17433.5 1048.035 17443.455 1071.07 ;
      RECT 17433.5 1048.035 17446.5 1054.07 ;
      RECT 17416.52 1149.44 17429.52 1209.16 ;
      RECT 17424.63 1048.035 17429.52 1209.16 ;
      RECT 17422.865 1053.42 17429.52 1209.16 ;
      RECT 17416.52 1053.42 17429.52 1118.87 ;
      RECT 17416.52 1048.035 17421.85 1118.87 ;
      RECT 17416.52 1048.035 17429.52 1049.12 ;
      RECT 17386 1070.44 17414 1209.16 ;
      RECT 17396.865 1048.035 17414 1209.16 ;
      RECT 17386 1048.035 17391.955 1209.16 ;
      RECT 17386 1048.035 17414 1054.07 ;
      RECT 17370.48 1118.44 17383.48 1209.16 ;
      RECT 17378.375 1048.035 17383.48 1209.16 ;
      RECT 17370.48 1048.035 17383.48 1087.87 ;
      RECT 17353.5 1166.44 17366.5 1189.16 ;
      RECT 17364.43 1048.035 17366.5 1189.16 ;
      RECT 17360.475 1053.365 17366.5 1189.16 ;
      RECT 17353.5 1048.035 17355.565 1189.16 ;
      RECT 17353.5 1087.44 17366.5 1150.07 ;
      RECT 17353.5 1053.365 17366.5 1071.07 ;
      RECT 17353.5 1048.035 17358.81 1071.07 ;
      RECT 17353.5 1048.035 17366.5 1049.165 ;
      RECT 17336.52 1166.44 17349.52 1209.16 ;
      RECT 17338.145 1048.035 17349.52 1209.16 ;
      RECT 17336.52 1087.44 17349.52 1150.07 ;
      RECT 17336.52 1048.035 17349.52 1071.07 ;
      RECT 17306 1183.44 17334 1209.16 ;
      RECT 17312.145 1048.035 17328.565 1209.16 ;
      RECT 17306 1070.44 17307.235 1209.16 ;
      RECT 17306 1070.44 17333.235 1167.07 ;
      RECT 17306 1087.44 17334 1150.07 ;
      RECT 17308.365 1048.035 17328.565 1167.07 ;
      RECT 17306 1048.035 17334 1054.07 ;
      RECT 17290.48 1087.44 17303.48 1209.16 ;
      RECT 17290.48 1048.035 17296.835 1209.16 ;
      RECT 17290.48 1048.035 17303.48 1071.07 ;
      RECT 17273.5 1149.44 17286.5 1189.16 ;
      RECT 17284.63 1048.035 17286.5 1189.16 ;
      RECT 17282.865 1053.42 17286.5 1189.16 ;
      RECT 17273.5 1048.035 17275.115 1189.16 ;
      RECT 17273.5 1053.42 17286.5 1118.87 ;
      RECT 17273.5 1048.035 17281.85 1118.87 ;
      RECT 17273.5 1048.035 17286.5 1049.12 ;
      RECT 17256.52 1070.44 17269.52 1209.16 ;
      RECT 17256.865 1048.035 17269.52 1209.16 ;
      RECT 17256.52 1048.035 17269.52 1054.07 ;
      RECT 17226 1118.44 17254 1209.16 ;
      RECT 17238.375 1070.44 17254 1209.16 ;
      RECT 17226 1048.035 17230.625 1209.16 ;
      RECT 17226 1048.035 17251.955 1087.87 ;
      RECT 17226 1048.035 17254 1054.07 ;
      RECT 17210.48 1166.44 17223.48 1209.16 ;
      RECT 17220.475 1053.365 17223.48 1209.16 ;
      RECT 17210.48 1048.035 17215.565 1209.16 ;
      RECT 17210.48 1087.44 17223.48 1150.07 ;
      RECT 17210.48 1053.365 17223.48 1071.07 ;
      RECT 17210.48 1048.035 17218.81 1071.07 ;
      RECT 17210.48 1048.035 17223.48 1049.165 ;
      RECT 17193.5 1166.44 17206.5 1189.16 ;
      RECT 17198.145 1048.035 17206.5 1189.16 ;
      RECT 17197.98 1087.44 17206.5 1189.16 ;
      RECT 17193.5 1087.44 17206.5 1150.07 ;
      RECT 17193.5 1048.035 17206.5 1071.07 ;
      RECT 17176.52 1183.44 17189.52 1209.16 ;
      RECT 17176.52 1048.035 17188.565 1209.16 ;
      RECT 17176.52 1070.44 17189.52 1167.07 ;
      RECT 17176.52 1048.035 17189.52 1054.07 ;
      RECT 17146 1183.44 17174 1209.16 ;
      RECT 17172.145 1048.035 17174 1209.16 ;
      RECT 17146 1087.44 17167.235 1209.16 ;
      RECT 17169.555 1048.035 17174 1167.07 ;
      RECT 17152.55 1070.44 17174 1167.07 ;
      RECT 17146 1048.035 17164.645 1071.07 ;
      RECT 17146 1048.035 17174 1054.07 ;
      RECT 17130.48 1149.44 17143.48 1209.16 ;
      RECT 17142.865 1053.415 17143.48 1209.16 ;
      RECT 17130.48 1048.035 17135.115 1209.16 ;
      RECT 17130.48 1053.415 17143.48 1118.87 ;
      RECT 17130.48 1048.035 17141.85 1118.87 ;
      RECT 17130.48 1048.035 17143.48 1049.12 ;
      RECT 17113.5 1070.44 17126.5 1189.16 ;
      RECT 17116.865 1048.035 17126.5 1189.16 ;
      RECT 17113.5 1048.035 17126.5 1054.07 ;
      RECT 17096.52 1118.44 17109.52 1209.16 ;
      RECT 17098.375 1048.035 17109.52 1209.16 ;
      RECT 17096.52 1048.035 17109.52 1087.87 ;
      RECT 17066 1166.44 17094 1209.16 ;
      RECT 17080.475 1118.44 17094 1209.16 ;
      RECT 17066 1048.035 17075.565 1209.16 ;
      RECT 17066 1087.44 17090.625 1150.07 ;
      RECT 17084.53 1048.035 17094 1087.87 ;
      RECT 17080.475 1053.365 17094 1087.87 ;
      RECT 17066 1053.365 17094 1071.07 ;
      RECT 17066 1048.035 17078.81 1071.07 ;
      RECT 17066 1048.035 17094 1049.165 ;
      RECT 17050.48 1183.44 17063.48 1209.16 ;
      RECT 17058.145 1048.035 17063.48 1209.16 ;
      RECT 17053.475 1166.44 17063.48 1209.16 ;
      RECT 17050.48 1166.44 17063.48 1167.07 ;
      RECT 17050.48 1070.44 17053.235 1167.07 ;
      RECT 17050.48 1087.44 17063.48 1150.07 ;
      RECT 17050.48 1070.44 17063.48 1071.07 ;
      RECT 17053.475 1048.035 17063.48 1071.07 ;
      RECT 17050.48 1048.035 17063.48 1054.07 ;
      RECT 17016.52 1183.44 17029.52 1209.16 ;
      RECT 17016.52 1087.44 17027.235 1209.16 ;
      RECT 17021.75 1070.44 17029.52 1167.07 ;
      RECT 17016.52 1048.035 17024.565 1071.07 ;
      RECT 17016.52 1048.035 17029.52 1054.07 ;
      RECT 16986 1149.44 17014 1209.16 ;
      RECT 17004.63 1048.035 17014 1209.16 ;
      RECT 17002.865 1053.42 17014 1209.16 ;
      RECT 16986 1048.035 16995.115 1209.16 ;
      RECT 16986 1053.42 17014 1118.87 ;
      RECT 16986 1048.035 17001.85 1118.87 ;
      RECT 16986 1048.035 17014 1049.12 ;
      RECT 16970.48 1070.44 16983.48 1209.16 ;
      RECT 16976.865 1048.035 16983.48 1209.16 ;
      RECT 16970.48 1048.035 16971.955 1209.16 ;
      RECT 16970.48 1048.035 16983.48 1054.07 ;
      RECT 16953.5 1118.44 16966.5 1189.16 ;
      RECT 16958.375 1048.035 16966.5 1189.16 ;
      RECT 16953.5 1048.035 16966.5 1087.87 ;
      RECT 16936.52 1166.44 16949.52 1209.16 ;
      RECT 16944.53 1048.035 16949.52 1209.16 ;
      RECT 16940.475 1053.365 16949.52 1209.16 ;
      RECT 16936.52 1087.44 16949.52 1150.07 ;
      RECT 16936.52 1053.365 16949.52 1071.07 ;
      RECT 16936.52 1048.035 16938.81 1071.07 ;
      RECT 16936.52 1048.035 16949.52 1049.375 ;
      RECT 16906 1183.44 16934 1209.16 ;
      RECT 16918.145 1048.035 16934 1209.16 ;
      RECT 16913.475 1166.44 16934 1209.16 ;
      RECT 16906 1048.035 16908.565 1209.16 ;
      RECT 16906 1166.44 16934 1167.07 ;
      RECT 16906 1070.44 16913.235 1167.07 ;
      RECT 16906 1087.44 16934 1150.07 ;
      RECT 16906 1070.44 16934 1071.07 ;
      RECT 16913.475 1048.035 16934 1071.07 ;
      RECT 16906 1048.035 16934 1054.07 ;
      RECT 16890.48 1183.44 16903.48 1209.16 ;
      RECT 16892.145 1048.035 16903.48 1209.16 ;
      RECT 16890.48 1048.035 16903.48 1167.07 ;
      RECT 16873.5 1087.44 16886.5 1189.16 ;
      RECT 16880.13 1070.44 16886.5 1189.16 ;
      RECT 16873.5 1048.035 16883.455 1071.07 ;
      RECT 16873.5 1048.035 16886.5 1054.07 ;
      RECT 16856.52 1149.44 16869.52 1209.16 ;
      RECT 16864.63 1048.035 16869.52 1209.16 ;
      RECT 16862.865 1053.42 16869.52 1209.16 ;
      RECT 16856.52 1053.42 16869.52 1118.87 ;
      RECT 16856.52 1048.035 16861.85 1118.87 ;
      RECT 16856.52 1048.035 16869.52 1049.12 ;
      RECT 16826 1070.44 16854 1209.16 ;
      RECT 16836.865 1048.035 16854 1209.16 ;
      RECT 16826 1048.035 16831.955 1209.16 ;
      RECT 16826 1048.035 16854 1054.07 ;
      RECT 16810.48 1118.44 16823.48 1209.16 ;
      RECT 16818.375 1048.035 16823.48 1209.16 ;
      RECT 16810.48 1048.035 16823.48 1087.87 ;
      RECT 16793.5 1166.44 16806.5 1189.16 ;
      RECT 16804.43 1048.035 16806.5 1189.16 ;
      RECT 16800.475 1053.365 16806.5 1189.16 ;
      RECT 16793.5 1048.035 16795.565 1189.16 ;
      RECT 16793.5 1087.44 16806.5 1150.07 ;
      RECT 16793.5 1053.365 16806.5 1071.07 ;
      RECT 16793.5 1048.035 16798.81 1071.07 ;
      RECT 16793.5 1048.035 16806.5 1049.165 ;
      RECT 16776.52 1166.44 16789.52 1209.16 ;
      RECT 16778.145 1048.035 16789.52 1209.16 ;
      RECT 16776.52 1087.44 16789.52 1150.07 ;
      RECT 16776.52 1048.035 16789.52 1071.07 ;
      RECT 16746 1183.44 16774 1209.16 ;
      RECT 16752.145 1048.035 16768.565 1209.16 ;
      RECT 16746 1070.44 16747.235 1209.16 ;
      RECT 16746 1070.44 16773.235 1167.07 ;
      RECT 16746 1087.44 16774 1150.07 ;
      RECT 16748.365 1048.035 16768.565 1167.07 ;
      RECT 16746 1048.035 16774 1054.07 ;
      RECT 16730.48 1087.44 16743.48 1209.16 ;
      RECT 16730.48 1048.035 16736.835 1209.16 ;
      RECT 16730.48 1048.035 16743.48 1071.07 ;
      RECT 16713.5 1149.44 16726.5 1189.16 ;
      RECT 16724.63 1048.035 16726.5 1189.16 ;
      RECT 16722.865 1053.42 16726.5 1189.16 ;
      RECT 16713.5 1048.035 16715.115 1189.16 ;
      RECT 16713.5 1053.42 16726.5 1118.87 ;
      RECT 16713.5 1048.035 16721.85 1118.87 ;
      RECT 16713.5 1048.035 16726.5 1049.12 ;
      RECT 16696.52 1070.44 16709.52 1209.16 ;
      RECT 16696.865 1048.035 16709.52 1209.16 ;
      RECT 16696.52 1048.035 16709.52 1054.07 ;
      RECT 16666 1118.44 16694 1209.16 ;
      RECT 16678.375 1070.44 16694 1209.16 ;
      RECT 16666 1048.035 16670.625 1209.16 ;
      RECT 16666 1048.035 16691.955 1087.87 ;
      RECT 16666 1048.035 16694 1054.07 ;
      RECT 16650.48 1166.44 16663.48 1209.16 ;
      RECT 16660.475 1053.365 16663.48 1209.16 ;
      RECT 16650.48 1048.035 16655.565 1209.16 ;
      RECT 16650.48 1087.44 16663.48 1150.07 ;
      RECT 16650.48 1053.365 16663.48 1071.07 ;
      RECT 16650.48 1048.035 16658.81 1071.07 ;
      RECT 16650.48 1048.035 16663.48 1049.165 ;
      RECT 16633.5 1166.44 16646.5 1189.16 ;
      RECT 16638.145 1048.035 16646.5 1189.16 ;
      RECT 16637.98 1087.44 16646.5 1189.16 ;
      RECT 16633.5 1087.44 16646.5 1150.07 ;
      RECT 16633.5 1048.035 16646.5 1071.07 ;
      RECT 16616.52 1183.44 16629.52 1209.16 ;
      RECT 16616.52 1048.035 16628.565 1209.16 ;
      RECT 16616.52 1070.44 16629.52 1167.07 ;
      RECT 16616.52 1048.035 16629.52 1054.07 ;
      RECT 16586 1183.44 16614 1209.16 ;
      RECT 16612.145 1048.035 16614 1209.16 ;
      RECT 16586 1087.44 16607.235 1209.16 ;
      RECT 16609.555 1048.035 16614 1167.07 ;
      RECT 16592.55 1070.44 16614 1167.07 ;
      RECT 16586 1048.035 16604.645 1071.07 ;
      RECT 16586 1048.035 16614 1054.07 ;
      RECT 16570.48 1149.44 16583.48 1209.16 ;
      RECT 16582.865 1053.415 16583.48 1209.16 ;
      RECT 16570.48 1048.035 16575.115 1209.16 ;
      RECT 16570.48 1053.415 16583.48 1118.87 ;
      RECT 16570.48 1048.035 16581.85 1118.87 ;
      RECT 16570.48 1048.035 16583.48 1049.12 ;
      RECT 16553.5 1070.44 16566.5 1189.16 ;
      RECT 16556.865 1048.035 16566.5 1189.16 ;
      RECT 16553.5 1048.035 16566.5 1054.07 ;
      RECT 16536.52 1118.44 16549.52 1209.16 ;
      RECT 16538.375 1048.035 16549.52 1209.16 ;
      RECT 16536.52 1048.035 16549.52 1087.87 ;
      RECT 16506 1166.44 16534 1209.16 ;
      RECT 16520.475 1118.44 16534 1209.16 ;
      RECT 16506 1048.035 16515.565 1209.16 ;
      RECT 16506 1087.44 16530.625 1150.07 ;
      RECT 16524.53 1048.035 16534 1087.87 ;
      RECT 16520.475 1053.365 16534 1087.87 ;
      RECT 16506 1053.365 16534 1071.07 ;
      RECT 16506 1048.035 16518.81 1071.07 ;
      RECT 16506 1048.035 16534 1049.165 ;
      RECT 16490.48 1183.44 16503.48 1209.16 ;
      RECT 16498.145 1048.035 16503.48 1209.16 ;
      RECT 16493.475 1166.44 16503.48 1209.16 ;
      RECT 16490.48 1166.44 16503.48 1167.07 ;
      RECT 16490.48 1070.44 16493.235 1167.07 ;
      RECT 16490.48 1087.44 16503.48 1150.07 ;
      RECT 16490.48 1070.44 16503.48 1071.07 ;
      RECT 16493.475 1048.035 16503.48 1071.07 ;
      RECT 16490.48 1048.035 16503.48 1054.07 ;
      RECT 16456.52 1183.44 16469.52 1209.16 ;
      RECT 16456.52 1087.44 16467.235 1209.16 ;
      RECT 16461.75 1070.44 16469.52 1167.07 ;
      RECT 16456.52 1048.035 16464.565 1071.07 ;
      RECT 16456.52 1048.035 16469.52 1054.07 ;
      RECT 16426 1149.44 16454 1209.16 ;
      RECT 16444.63 1048.035 16454 1209.16 ;
      RECT 16442.865 1053.42 16454 1209.16 ;
      RECT 16426 1048.035 16435.115 1209.16 ;
      RECT 16426 1053.42 16454 1118.87 ;
      RECT 16426 1048.035 16441.85 1118.87 ;
      RECT 16426 1048.035 16454 1049.12 ;
      RECT 16410.48 1070.44 16423.48 1209.16 ;
      RECT 16416.865 1048.035 16423.48 1209.16 ;
      RECT 16410.48 1048.035 16411.955 1209.16 ;
      RECT 16410.48 1048.035 16423.48 1054.07 ;
      RECT 16393.5 1118.44 16406.5 1189.16 ;
      RECT 16398.375 1048.035 16406.5 1189.16 ;
      RECT 16393.5 1048.035 16406.5 1087.87 ;
      RECT 16376.52 1166.44 16389.52 1209.16 ;
      RECT 16384.53 1048.035 16389.52 1209.16 ;
      RECT 16380.475 1053.365 16389.52 1209.16 ;
      RECT 16376.52 1087.44 16389.52 1150.07 ;
      RECT 16376.52 1053.365 16389.52 1071.07 ;
      RECT 16376.52 1048.035 16378.81 1071.07 ;
      RECT 16376.52 1048.035 16389.52 1049.375 ;
      RECT 16346 1183.44 16374 1209.16 ;
      RECT 16358.145 1048.035 16374 1209.16 ;
      RECT 16353.475 1166.44 16374 1209.16 ;
      RECT 16346 1048.035 16348.565 1209.16 ;
      RECT 16346 1166.44 16374 1167.07 ;
      RECT 16346 1070.44 16353.235 1167.07 ;
      RECT 16346 1087.44 16374 1150.07 ;
      RECT 16346 1070.44 16374 1071.07 ;
      RECT 16353.475 1048.035 16374 1071.07 ;
      RECT 16346 1048.035 16374 1054.07 ;
      RECT 16330.48 1183.44 16343.48 1209.16 ;
      RECT 16332.145 1048.035 16343.48 1209.16 ;
      RECT 16330.48 1048.035 16343.48 1167.07 ;
      RECT 16313.5 1087.44 16326.5 1189.16 ;
      RECT 16320.13 1070.44 16326.5 1189.16 ;
      RECT 16313.5 1048.035 16323.455 1071.07 ;
      RECT 16313.5 1048.035 16326.5 1054.07 ;
      RECT 16296.52 1149.44 16309.52 1209.16 ;
      RECT 16304.63 1048.035 16309.52 1209.16 ;
      RECT 16302.865 1053.42 16309.52 1209.16 ;
      RECT 16296.52 1053.42 16309.52 1118.87 ;
      RECT 16296.52 1048.035 16301.85 1118.87 ;
      RECT 16296.52 1048.035 16309.52 1049.12 ;
      RECT 16266 1070.44 16294 1209.16 ;
      RECT 16276.865 1048.035 16294 1209.16 ;
      RECT 16266 1048.035 16271.955 1209.16 ;
      RECT 16266 1048.035 16294 1054.07 ;
      RECT 16250.48 1118.44 16263.48 1209.16 ;
      RECT 16258.375 1048.035 16263.48 1209.16 ;
      RECT 16250.48 1048.035 16263.48 1087.87 ;
      RECT 16233.5 1166.44 16246.5 1189.16 ;
      RECT 16244.43 1048.035 16246.5 1189.16 ;
      RECT 16240.475 1053.365 16246.5 1189.16 ;
      RECT 16233.5 1048.035 16235.565 1189.16 ;
      RECT 16233.5 1087.44 16246.5 1150.07 ;
      RECT 16233.5 1053.365 16246.5 1071.07 ;
      RECT 16233.5 1048.035 16238.81 1071.07 ;
      RECT 16233.5 1048.035 16246.5 1049.165 ;
      RECT 16216.52 1166.44 16229.52 1209.16 ;
      RECT 16218.145 1048.035 16229.52 1209.16 ;
      RECT 16216.52 1087.44 16229.52 1150.07 ;
      RECT 16216.52 1048.035 16229.52 1071.07 ;
      RECT 16186 1183.44 16214 1209.16 ;
      RECT 16192.145 1048.035 16208.565 1209.16 ;
      RECT 16186 1070.44 16187.235 1209.16 ;
      RECT 16186 1070.44 16213.235 1167.07 ;
      RECT 16186 1087.44 16214 1150.07 ;
      RECT 16188.365 1048.035 16208.565 1167.07 ;
      RECT 16186 1048.035 16214 1054.07 ;
      RECT 16170.48 1087.44 16183.48 1209.16 ;
      RECT 16170.48 1048.035 16176.835 1209.16 ;
      RECT 16170.48 1048.035 16183.48 1071.07 ;
      RECT 16153.5 1149.44 16166.5 1189.16 ;
      RECT 16164.63 1048.035 16166.5 1189.16 ;
      RECT 16162.865 1053.42 16166.5 1189.16 ;
      RECT 16153.5 1048.035 16155.115 1189.16 ;
      RECT 16153.5 1053.42 16166.5 1118.87 ;
      RECT 16153.5 1048.035 16161.85 1118.87 ;
      RECT 16153.5 1048.035 16166.5 1049.12 ;
      RECT 16136.52 1070.44 16149.52 1209.16 ;
      RECT 16136.865 1048.035 16149.52 1209.16 ;
      RECT 16136.52 1048.035 16149.52 1054.07 ;
      RECT 16106 1118.44 16134 1209.16 ;
      RECT 16118.375 1070.44 16134 1209.16 ;
      RECT 16106 1048.035 16110.625 1209.16 ;
      RECT 16106 1048.035 16131.955 1087.87 ;
      RECT 16106 1048.035 16134 1054.07 ;
      RECT 16090.48 1166.44 16103.48 1209.16 ;
      RECT 16100.475 1053.365 16103.48 1209.16 ;
      RECT 16090.48 1048.035 16095.565 1209.16 ;
      RECT 16090.48 1087.44 16103.48 1150.07 ;
      RECT 16090.48 1053.365 16103.48 1071.07 ;
      RECT 16090.48 1048.035 16098.81 1071.07 ;
      RECT 16090.48 1048.035 16103.48 1049.165 ;
      RECT 16073.5 1166.44 16086.5 1189.16 ;
      RECT 16078.145 1048.035 16086.5 1189.16 ;
      RECT 16077.98 1087.44 16086.5 1189.16 ;
      RECT 16073.5 1087.44 16086.5 1150.07 ;
      RECT 16073.5 1048.035 16086.5 1071.07 ;
      RECT 16056.52 1183.44 16069.52 1209.16 ;
      RECT 16056.52 1048.035 16068.565 1209.16 ;
      RECT 16056.52 1070.44 16069.52 1167.07 ;
      RECT 16056.52 1048.035 16069.52 1054.07 ;
      RECT 16026 1183.44 16054 1209.16 ;
      RECT 16052.145 1048.035 16054 1209.16 ;
      RECT 16026 1087.44 16047.235 1209.16 ;
      RECT 16049.555 1048.035 16054 1167.07 ;
      RECT 16032.55 1070.44 16054 1167.07 ;
      RECT 16026 1048.035 16044.645 1071.07 ;
      RECT 16026 1048.035 16054 1054.07 ;
      RECT 16010.48 1149.44 16023.48 1209.16 ;
      RECT 16022.865 1053.415 16023.48 1209.16 ;
      RECT 16010.48 1048.035 16015.115 1209.16 ;
      RECT 16010.48 1053.415 16023.48 1118.87 ;
      RECT 16010.48 1048.035 16021.85 1118.87 ;
      RECT 16010.48 1048.035 16023.48 1049.12 ;
      RECT 15993.5 1070.44 16006.5 1189.16 ;
      RECT 15996.865 1048.035 16006.5 1189.16 ;
      RECT 15993.5 1048.035 16006.5 1054.07 ;
      RECT 15976.52 1118.44 15989.52 1209.16 ;
      RECT 15978.375 1048.035 15989.52 1209.16 ;
      RECT 15976.52 1048.035 15989.52 1087.87 ;
      RECT 15946 1166.44 15974 1209.16 ;
      RECT 15960.475 1118.44 15974 1209.16 ;
      RECT 15946 1048.035 15955.565 1209.16 ;
      RECT 15946 1087.44 15970.625 1150.07 ;
      RECT 15964.53 1048.035 15974 1087.87 ;
      RECT 15960.475 1053.365 15974 1087.87 ;
      RECT 15946 1053.365 15974 1071.07 ;
      RECT 15946 1048.035 15958.81 1071.07 ;
      RECT 15946 1048.035 15974 1049.165 ;
      RECT 15930.48 1183.44 15943.48 1209.16 ;
      RECT 15938.145 1048.035 15943.48 1209.16 ;
      RECT 15933.475 1166.44 15943.48 1209.16 ;
      RECT 15930.48 1166.44 15943.48 1167.07 ;
      RECT 15930.48 1070.44 15933.235 1167.07 ;
      RECT 15930.48 1087.44 15943.48 1150.07 ;
      RECT 15930.48 1070.44 15943.48 1071.07 ;
      RECT 15933.475 1048.035 15943.48 1071.07 ;
      RECT 15930.48 1048.035 15943.48 1054.07 ;
      RECT 15896.52 1183.44 15909.52 1209.16 ;
      RECT 15896.52 1087.44 15907.235 1209.16 ;
      RECT 15901.75 1070.44 15909.52 1167.07 ;
      RECT 15896.52 1048.035 15904.565 1071.07 ;
      RECT 15896.52 1048.035 15909.52 1054.07 ;
      RECT 15866 1149.44 15894 1209.16 ;
      RECT 15884.63 1048.035 15894 1209.16 ;
      RECT 15882.865 1053.42 15894 1209.16 ;
      RECT 15866 1048.035 15875.115 1209.16 ;
      RECT 15866 1053.42 15894 1118.87 ;
      RECT 15866 1048.035 15881.85 1118.87 ;
      RECT 15866 1048.035 15894 1049.12 ;
      RECT 15850.48 1070.44 15863.48 1209.16 ;
      RECT 15856.865 1048.035 15863.48 1209.16 ;
      RECT 15850.48 1048.035 15851.955 1209.16 ;
      RECT 15850.48 1048.035 15863.48 1054.07 ;
      RECT 15833.5 1118.44 15846.5 1189.16 ;
      RECT 15838.375 1048.035 15846.5 1189.16 ;
      RECT 15833.5 1048.035 15846.5 1087.87 ;
      RECT 15816.52 1166.44 15829.52 1209.16 ;
      RECT 15824.53 1048.035 15829.52 1209.16 ;
      RECT 15820.475 1053.365 15829.52 1209.16 ;
      RECT 15816.52 1087.44 15829.52 1150.07 ;
      RECT 15816.52 1053.365 15829.52 1071.07 ;
      RECT 15816.52 1048.035 15818.81 1071.07 ;
      RECT 15816.52 1048.035 15829.52 1049.375 ;
      RECT 15786 1183.44 15814 1209.16 ;
      RECT 15798.145 1048.035 15814 1209.16 ;
      RECT 15793.475 1166.44 15814 1209.16 ;
      RECT 15786 1048.035 15788.565 1209.16 ;
      RECT 15786 1166.44 15814 1167.07 ;
      RECT 15786 1070.44 15793.235 1167.07 ;
      RECT 15786 1087.44 15814 1150.07 ;
      RECT 15786 1070.44 15814 1071.07 ;
      RECT 15793.475 1048.035 15814 1071.07 ;
      RECT 15786 1048.035 15814 1054.07 ;
      RECT 15770.48 1183.44 15783.48 1209.16 ;
      RECT 15772.145 1048.035 15783.48 1209.16 ;
      RECT 15770.48 1048.035 15783.48 1167.07 ;
      RECT 15753.5 1087.44 15766.5 1189.16 ;
      RECT 15760.13 1070.44 15766.5 1189.16 ;
      RECT 15753.5 1048.035 15763.455 1071.07 ;
      RECT 15753.5 1048.035 15766.5 1054.07 ;
      RECT 15736.52 1149.44 15749.52 1209.16 ;
      RECT 15744.63 1048.035 15749.52 1209.16 ;
      RECT 15742.865 1053.42 15749.52 1209.16 ;
      RECT 15736.52 1053.42 15749.52 1118.87 ;
      RECT 15736.52 1048.035 15741.85 1118.87 ;
      RECT 15736.52 1048.035 15749.52 1049.12 ;
      RECT 15706 1070.44 15734 1209.16 ;
      RECT 15716.865 1048.035 15734 1209.16 ;
      RECT 15706 1048.035 15711.955 1209.16 ;
      RECT 15706 1048.035 15734 1054.07 ;
      RECT 15690.48 1118.44 15703.48 1209.16 ;
      RECT 15698.375 1048.035 15703.48 1209.16 ;
      RECT 15690.48 1048.035 15703.48 1087.87 ;
      RECT 15673.5 1166.44 15686.5 1189.16 ;
      RECT 15684.43 1048.035 15686.5 1189.16 ;
      RECT 15680.475 1053.365 15686.5 1189.16 ;
      RECT 15673.5 1048.035 15675.565 1189.16 ;
      RECT 15673.5 1087.44 15686.5 1150.07 ;
      RECT 15673.5 1053.365 15686.5 1071.07 ;
      RECT 15673.5 1048.035 15678.81 1071.07 ;
      RECT 15673.5 1048.035 15686.5 1049.165 ;
      RECT 15656.52 1166.44 15669.52 1209.16 ;
      RECT 15658.145 1048.035 15669.52 1209.16 ;
      RECT 15656.52 1087.44 15669.52 1150.07 ;
      RECT 15656.52 1048.035 15669.52 1071.07 ;
      RECT 15626 1183.44 15654 1209.16 ;
      RECT 15632.145 1048.035 15648.565 1209.16 ;
      RECT 15626 1070.44 15627.235 1209.16 ;
      RECT 15626 1070.44 15653.235 1167.07 ;
      RECT 15626 1087.44 15654 1150.07 ;
      RECT 15628.365 1048.035 15648.565 1167.07 ;
      RECT 15626 1048.035 15654 1054.07 ;
      RECT 15610.48 1087.44 15623.48 1209.16 ;
      RECT 15610.48 1048.035 15616.835 1209.16 ;
      RECT 15610.48 1048.035 15623.48 1071.07 ;
      RECT 15593.5 1149.44 15606.5 1189.16 ;
      RECT 15604.63 1048.035 15606.5 1189.16 ;
      RECT 15602.865 1053.42 15606.5 1189.16 ;
      RECT 15593.5 1048.035 15595.115 1189.16 ;
      RECT 15593.5 1053.42 15606.5 1118.87 ;
      RECT 15593.5 1048.035 15601.85 1118.87 ;
      RECT 15593.5 1048.035 15606.5 1049.12 ;
      RECT 15576.52 1070.44 15589.52 1209.16 ;
      RECT 15576.865 1048.035 15589.52 1209.16 ;
      RECT 15576.52 1048.035 15589.52 1054.07 ;
      RECT 15546 1118.44 15574 1209.16 ;
      RECT 15558.375 1070.44 15574 1209.16 ;
      RECT 15546 1048.035 15550.625 1209.16 ;
      RECT 15546 1048.035 15571.955 1087.87 ;
      RECT 15546 1048.035 15574 1054.07 ;
      RECT 15530.48 1166.44 15543.48 1209.16 ;
      RECT 15540.475 1053.365 15543.48 1209.16 ;
      RECT 15530.48 1048.035 15535.565 1209.16 ;
      RECT 15530.48 1087.44 15543.48 1150.07 ;
      RECT 15530.48 1053.365 15543.48 1071.07 ;
      RECT 15530.48 1048.035 15538.81 1071.07 ;
      RECT 15530.48 1048.035 15543.48 1049.165 ;
      RECT 15513.5 1166.44 15526.5 1189.16 ;
      RECT 15518.145 1048.035 15526.5 1189.16 ;
      RECT 15517.98 1087.44 15526.5 1189.16 ;
      RECT 15513.5 1087.44 15526.5 1150.07 ;
      RECT 15513.5 1048.035 15526.5 1071.07 ;
      RECT 15496.52 1183.44 15509.52 1209.16 ;
      RECT 15496.52 1048.035 15508.565 1209.16 ;
      RECT 15496.52 1070.44 15509.52 1167.07 ;
      RECT 15496.52 1048.035 15509.52 1054.07 ;
      RECT 15466 1183.44 15494 1209.16 ;
      RECT 15492.145 1048.035 15494 1209.16 ;
      RECT 15466 1087.44 15487.235 1209.16 ;
      RECT 15489.555 1048.035 15494 1167.07 ;
      RECT 15472.55 1070.44 15494 1167.07 ;
      RECT 15466 1048.035 15484.645 1071.07 ;
      RECT 15466 1048.035 15494 1054.07 ;
      RECT 15450.48 1149.44 15463.48 1209.16 ;
      RECT 15462.865 1053.415 15463.48 1209.16 ;
      RECT 15450.48 1048.035 15455.115 1209.16 ;
      RECT 15450.48 1053.415 15463.48 1118.87 ;
      RECT 15450.48 1048.035 15461.85 1118.87 ;
      RECT 15450.48 1048.035 15463.48 1049.12 ;
      RECT 15433.5 1070.44 15446.5 1189.16 ;
      RECT 15436.865 1048.035 15446.5 1189.16 ;
      RECT 15433.5 1048.035 15446.5 1054.07 ;
      RECT 15416.52 1118.44 15429.52 1209.16 ;
      RECT 15418.375 1048.035 15429.52 1209.16 ;
      RECT 15416.52 1048.035 15429.52 1087.87 ;
      RECT 15386 1166.44 15414 1209.16 ;
      RECT 15400.475 1118.44 15414 1209.16 ;
      RECT 15386 1048.035 15395.565 1209.16 ;
      RECT 15386 1087.44 15410.625 1150.07 ;
      RECT 15404.53 1048.035 15414 1087.87 ;
      RECT 15400.475 1053.365 15414 1087.87 ;
      RECT 15386 1053.365 15414 1071.07 ;
      RECT 15386 1048.035 15398.81 1071.07 ;
      RECT 15386 1048.035 15414 1049.165 ;
      RECT 15370.48 1183.44 15383.48 1209.16 ;
      RECT 15378.145 1048.035 15383.48 1209.16 ;
      RECT 15373.475 1166.44 15383.48 1209.16 ;
      RECT 15370.48 1166.44 15383.48 1167.07 ;
      RECT 15370.48 1070.44 15373.235 1167.07 ;
      RECT 15370.48 1087.44 15383.48 1150.07 ;
      RECT 15370.48 1070.44 15383.48 1071.07 ;
      RECT 15373.475 1048.035 15383.48 1071.07 ;
      RECT 15370.48 1048.035 15383.48 1054.07 ;
      RECT 15336.52 1183.44 15349.52 1209.16 ;
      RECT 15336.52 1087.44 15347.235 1209.16 ;
      RECT 15341.75 1070.44 15349.52 1167.07 ;
      RECT 15336.52 1048.035 15344.565 1071.07 ;
      RECT 15336.52 1048.035 15349.52 1054.07 ;
      RECT 15306 1149.44 15334 1209.16 ;
      RECT 15324.63 1048.035 15334 1209.16 ;
      RECT 15322.865 1053.42 15334 1209.16 ;
      RECT 15306 1048.035 15315.115 1209.16 ;
      RECT 15306 1053.42 15334 1118.87 ;
      RECT 15306 1048.035 15321.85 1118.87 ;
      RECT 15306 1048.035 15334 1049.12 ;
      RECT 15290.48 1070.44 15303.48 1209.16 ;
      RECT 15296.865 1048.035 15303.48 1209.16 ;
      RECT 15290.48 1048.035 15291.955 1209.16 ;
      RECT 15290.48 1048.035 15303.48 1054.07 ;
      RECT 15273.5 1118.44 15286.5 1189.16 ;
      RECT 15278.375 1048.035 15286.5 1189.16 ;
      RECT 15273.5 1048.035 15286.5 1087.87 ;
      RECT 15256.52 1166.44 15269.52 1209.16 ;
      RECT 15264.53 1048.035 15269.52 1209.16 ;
      RECT 15260.475 1053.365 15269.52 1209.16 ;
      RECT 15256.52 1087.44 15269.52 1150.07 ;
      RECT 15256.52 1053.365 15269.52 1071.07 ;
      RECT 15256.52 1048.035 15258.81 1071.07 ;
      RECT 15256.52 1048.035 15269.52 1049.375 ;
      RECT 15226 1183.44 15254 1209.16 ;
      RECT 15238.145 1048.035 15254 1209.16 ;
      RECT 15233.475 1166.44 15254 1209.16 ;
      RECT 15226 1048.035 15228.565 1209.16 ;
      RECT 15226 1166.44 15254 1167.07 ;
      RECT 15226 1070.44 15233.235 1167.07 ;
      RECT 15226 1087.44 15254 1150.07 ;
      RECT 15226 1070.44 15254 1071.07 ;
      RECT 15233.475 1048.035 15254 1071.07 ;
      RECT 15226 1048.035 15254 1054.07 ;
      RECT 15210.48 1183.44 15223.48 1209.16 ;
      RECT 15212.145 1048.035 15223.48 1209.16 ;
      RECT 15210.48 1048.035 15223.48 1167.07 ;
      RECT 15193.5 1087.44 15206.5 1189.16 ;
      RECT 15200.13 1070.44 15206.5 1189.16 ;
      RECT 15193.5 1048.035 15203.455 1071.07 ;
      RECT 15193.5 1048.035 15206.5 1054.07 ;
      RECT 15176.52 1149.44 15189.52 1209.16 ;
      RECT 15184.63 1048.035 15189.52 1209.16 ;
      RECT 15182.865 1053.42 15189.52 1209.16 ;
      RECT 15176.52 1053.42 15189.52 1118.87 ;
      RECT 15176.52 1048.035 15181.85 1118.87 ;
      RECT 15176.52 1048.035 15189.52 1049.12 ;
      RECT 15146 1070.44 15174 1209.16 ;
      RECT 15156.865 1048.035 15174 1209.16 ;
      RECT 15146 1048.035 15151.955 1209.16 ;
      RECT 15146 1048.035 15174 1054.07 ;
      RECT 15130.48 1118.44 15143.48 1209.16 ;
      RECT 15138.375 1048.035 15143.48 1209.16 ;
      RECT 15130.48 1048.035 15143.48 1087.87 ;
      RECT 15113.5 1166.44 15126.5 1189.16 ;
      RECT 15124.43 1048.035 15126.5 1189.16 ;
      RECT 15120.475 1053.365 15126.5 1189.16 ;
      RECT 15113.5 1048.035 15115.565 1189.16 ;
      RECT 15113.5 1087.44 15126.5 1150.07 ;
      RECT 15113.5 1053.365 15126.5 1071.07 ;
      RECT 15113.5 1048.035 15118.81 1071.07 ;
      RECT 15113.5 1048.035 15126.5 1049.165 ;
      RECT 15096.52 1166.44 15109.52 1209.16 ;
      RECT 15098.145 1048.035 15109.52 1209.16 ;
      RECT 15096.52 1087.44 15109.52 1150.07 ;
      RECT 15096.52 1048.035 15109.52 1071.07 ;
      RECT 15066 1183.44 15094 1209.16 ;
      RECT 15072.145 1048.035 15088.565 1209.16 ;
      RECT 15066 1070.44 15067.235 1209.16 ;
      RECT 15066 1070.44 15093.235 1167.07 ;
      RECT 15066 1087.44 15094 1150.07 ;
      RECT 15068.365 1048.035 15088.565 1167.07 ;
      RECT 15066 1048.035 15094 1054.07 ;
      RECT 15050.48 1087.44 15063.48 1209.16 ;
      RECT 15050.48 1048.035 15056.835 1209.16 ;
      RECT 15050.48 1048.035 15063.48 1071.07 ;
      RECT 15033.5 1149.44 15046.5 1189.16 ;
      RECT 15044.63 1048.035 15046.5 1189.16 ;
      RECT 15042.865 1053.42 15046.5 1189.16 ;
      RECT 15033.5 1048.035 15035.115 1189.16 ;
      RECT 15033.5 1053.42 15046.5 1118.87 ;
      RECT 15033.5 1048.035 15041.85 1118.87 ;
      RECT 15033.5 1048.035 15046.5 1049.12 ;
      RECT 15016.52 1070.44 15029.52 1209.16 ;
      RECT 15016.865 1048.035 15029.52 1209.16 ;
      RECT 15016.52 1048.035 15029.52 1054.07 ;
      RECT 14986 1118.44 15014 1209.16 ;
      RECT 14998.375 1070.44 15014 1209.16 ;
      RECT 14986 1048.035 14990.625 1209.16 ;
      RECT 14986 1048.035 15011.955 1087.87 ;
      RECT 14986 1048.035 15014 1054.07 ;
      RECT 14970.48 1166.44 14983.48 1209.16 ;
      RECT 14980.475 1053.365 14983.48 1209.16 ;
      RECT 14970.48 1048.035 14975.565 1209.16 ;
      RECT 14970.48 1087.44 14983.48 1150.07 ;
      RECT 14970.48 1053.365 14983.48 1071.07 ;
      RECT 14970.48 1048.035 14978.81 1071.07 ;
      RECT 14970.48 1048.035 14983.48 1049.165 ;
      RECT 14953.5 1166.44 14966.5 1189.16 ;
      RECT 14958.145 1048.035 14966.5 1189.16 ;
      RECT 14957.98 1087.44 14966.5 1189.16 ;
      RECT 14953.5 1087.44 14966.5 1150.07 ;
      RECT 14953.5 1048.035 14966.5 1071.07 ;
      RECT 14936.52 1183.44 14949.52 1209.16 ;
      RECT 14936.52 1048.035 14948.565 1209.16 ;
      RECT 14936.52 1070.44 14949.52 1167.07 ;
      RECT 14936.52 1048.035 14949.52 1054.07 ;
      RECT 14906 1183.44 14934 1209.16 ;
      RECT 14932.145 1048.035 14934 1209.16 ;
      RECT 14906 1087.44 14927.235 1209.16 ;
      RECT 14929.555 1048.035 14934 1167.07 ;
      RECT 14912.55 1070.44 14934 1167.07 ;
      RECT 14906 1048.035 14924.645 1071.07 ;
      RECT 14906 1048.035 14934 1054.07 ;
      RECT 14890.48 1149.44 14903.48 1209.16 ;
      RECT 14902.865 1053.415 14903.48 1209.16 ;
      RECT 14890.48 1048.035 14895.115 1209.16 ;
      RECT 14890.48 1053.415 14903.48 1118.87 ;
      RECT 14890.48 1048.035 14901.85 1118.87 ;
      RECT 14890.48 1048.035 14903.48 1049.12 ;
      RECT 14873.5 1070.44 14886.5 1189.16 ;
      RECT 14876.865 1048.035 14886.5 1189.16 ;
      RECT 14873.5 1048.035 14886.5 1054.07 ;
      RECT 14856.52 1118.44 14869.52 1209.16 ;
      RECT 14858.375 1048.035 14869.52 1209.16 ;
      RECT 14856.52 1048.035 14869.52 1087.87 ;
      RECT 14826 1166.44 14854 1209.16 ;
      RECT 14840.475 1118.44 14854 1209.16 ;
      RECT 14826 1048.035 14835.565 1209.16 ;
      RECT 14826 1087.44 14850.625 1150.07 ;
      RECT 14844.53 1048.035 14854 1087.87 ;
      RECT 14840.475 1053.365 14854 1087.87 ;
      RECT 14826 1053.365 14854 1071.07 ;
      RECT 14826 1048.035 14838.81 1071.07 ;
      RECT 14826 1048.035 14854 1049.165 ;
      RECT 14810.48 1183.44 14823.48 1209.16 ;
      RECT 14818.145 1048.035 14823.48 1209.16 ;
      RECT 14813.475 1166.44 14823.48 1209.16 ;
      RECT 14810.48 1166.44 14823.48 1167.07 ;
      RECT 14810.48 1070.44 14813.235 1167.07 ;
      RECT 14810.48 1087.44 14823.48 1150.07 ;
      RECT 14810.48 1070.44 14823.48 1071.07 ;
      RECT 14813.475 1048.035 14823.48 1071.07 ;
      RECT 14810.48 1048.035 14823.48 1054.07 ;
      RECT 14776.52 1183.44 14789.52 1209.16 ;
      RECT 14776.52 1087.44 14787.235 1209.16 ;
      RECT 14781.75 1070.44 14789.52 1167.07 ;
      RECT 14776.52 1048.035 14784.565 1071.07 ;
      RECT 14776.52 1048.035 14789.52 1054.07 ;
      RECT 14746 1149.44 14774 1209.16 ;
      RECT 14764.63 1048.035 14774 1209.16 ;
      RECT 14762.865 1053.42 14774 1209.16 ;
      RECT 14746 1048.035 14755.115 1209.16 ;
      RECT 14746 1053.42 14774 1118.87 ;
      RECT 14746 1048.035 14761.85 1118.87 ;
      RECT 14746 1048.035 14774 1049.12 ;
      RECT 14730.48 1070.44 14743.48 1209.16 ;
      RECT 14736.865 1048.035 14743.48 1209.16 ;
      RECT 14730.48 1048.035 14731.955 1209.16 ;
      RECT 14730.48 1048.035 14743.48 1054.07 ;
      RECT 14713.5 1118.44 14726.5 1189.16 ;
      RECT 14718.375 1048.035 14726.5 1189.16 ;
      RECT 14713.5 1048.035 14726.5 1087.87 ;
      RECT 14696.52 1166.44 14709.52 1209.16 ;
      RECT 14704.53 1048.035 14709.52 1209.16 ;
      RECT 14700.475 1053.365 14709.52 1209.16 ;
      RECT 14696.52 1087.44 14709.52 1150.07 ;
      RECT 14696.52 1053.365 14709.52 1071.07 ;
      RECT 14696.52 1048.035 14698.81 1071.07 ;
      RECT 14696.52 1048.035 14709.52 1049.375 ;
      RECT 14666 1183.44 14694 1209.16 ;
      RECT 14678.145 1048.035 14694 1209.16 ;
      RECT 14673.475 1166.44 14694 1209.16 ;
      RECT 14666 1048.035 14668.565 1209.16 ;
      RECT 14666 1166.44 14694 1167.07 ;
      RECT 14666 1070.44 14673.235 1167.07 ;
      RECT 14666 1087.44 14694 1150.07 ;
      RECT 14666 1070.44 14694 1071.07 ;
      RECT 14673.475 1048.035 14694 1071.07 ;
      RECT 14666 1048.035 14694 1054.07 ;
      RECT 14650.48 1183.44 14663.48 1209.16 ;
      RECT 14652.145 1048.035 14663.48 1209.16 ;
      RECT 14650.48 1048.035 14663.48 1167.07 ;
      RECT 14633.5 1087.44 14646.5 1189.16 ;
      RECT 14640.13 1070.44 14646.5 1189.16 ;
      RECT 14633.5 1048.035 14643.455 1071.07 ;
      RECT 14633.5 1048.035 14646.5 1054.07 ;
      RECT 14616.52 1149.44 14629.52 1209.16 ;
      RECT 14624.63 1048.035 14629.52 1209.16 ;
      RECT 14622.865 1053.42 14629.52 1209.16 ;
      RECT 14616.52 1053.42 14629.52 1118.87 ;
      RECT 14616.52 1048.035 14621.85 1118.87 ;
      RECT 14616.52 1048.035 14629.52 1049.12 ;
      RECT 14586 1070.44 14614 1209.16 ;
      RECT 14596.865 1048.035 14614 1209.16 ;
      RECT 14586 1048.035 14591.955 1209.16 ;
      RECT 14586 1048.035 14614 1054.07 ;
      RECT 14570.48 1118.44 14583.48 1209.16 ;
      RECT 14578.375 1048.035 14583.48 1209.16 ;
      RECT 14570.48 1048.035 14583.48 1087.87 ;
      RECT 14553.5 1166.44 14566.5 1189.16 ;
      RECT 14564.43 1048.035 14566.5 1189.16 ;
      RECT 14560.475 1053.365 14566.5 1189.16 ;
      RECT 14553.5 1048.035 14555.565 1189.16 ;
      RECT 14553.5 1087.44 14566.5 1150.07 ;
      RECT 14553.5 1053.365 14566.5 1071.07 ;
      RECT 14553.5 1048.035 14558.81 1071.07 ;
      RECT 14553.5 1048.035 14566.5 1049.165 ;
      RECT 14536.52 1166.44 14549.52 1209.16 ;
      RECT 14538.145 1048.035 14549.52 1209.16 ;
      RECT 14536.52 1087.44 14549.52 1150.07 ;
      RECT 14536.52 1048.035 14549.52 1071.07 ;
      RECT 14506 1183.44 14534 1209.16 ;
      RECT 14512.145 1048.035 14528.565 1209.16 ;
      RECT 14506 1070.44 14507.235 1209.16 ;
      RECT 14506 1070.44 14533.235 1167.07 ;
      RECT 14506 1087.44 14534 1150.07 ;
      RECT 14508.365 1048.035 14528.565 1167.07 ;
      RECT 14506 1048.035 14534 1054.07 ;
      RECT 14490.48 1087.44 14503.48 1209.16 ;
      RECT 14490.48 1048.035 14496.835 1209.16 ;
      RECT 14490.48 1048.035 14503.48 1071.07 ;
      RECT 14473.5 1149.44 14486.5 1189.16 ;
      RECT 14484.63 1048.035 14486.5 1189.16 ;
      RECT 14482.865 1053.42 14486.5 1189.16 ;
      RECT 14473.5 1048.035 14475.115 1189.16 ;
      RECT 14473.5 1053.42 14486.5 1118.87 ;
      RECT 14473.5 1048.035 14481.85 1118.87 ;
      RECT 14473.5 1048.035 14486.5 1049.12 ;
      RECT 14456.52 1070.44 14469.52 1209.16 ;
      RECT 14456.865 1048.035 14469.52 1209.16 ;
      RECT 14456.52 1048.035 14469.52 1054.07 ;
      RECT 14426 1118.44 14454 1209.16 ;
      RECT 14438.375 1070.44 14454 1209.16 ;
      RECT 14426 1048.035 14430.625 1209.16 ;
      RECT 14426 1048.035 14451.955 1087.87 ;
      RECT 14426 1048.035 14454 1054.07 ;
      RECT 14410.48 1166.44 14423.48 1209.16 ;
      RECT 14420.475 1053.365 14423.48 1209.16 ;
      RECT 14410.48 1048.035 14415.565 1209.16 ;
      RECT 14410.48 1087.44 14423.48 1150.07 ;
      RECT 14410.48 1053.365 14423.48 1071.07 ;
      RECT 14410.48 1048.035 14418.81 1071.07 ;
      RECT 14410.48 1048.035 14423.48 1049.165 ;
      RECT 14393.5 1166.44 14406.5 1189.16 ;
      RECT 14398.145 1048.035 14406.5 1189.16 ;
      RECT 14397.98 1087.44 14406.5 1189.16 ;
      RECT 14393.5 1087.44 14406.5 1150.07 ;
      RECT 14393.5 1048.035 14406.5 1071.07 ;
      RECT 14376.52 1183.44 14389.52 1209.16 ;
      RECT 14376.52 1048.035 14388.565 1209.16 ;
      RECT 14376.52 1070.44 14389.52 1167.07 ;
      RECT 14376.52 1048.035 14389.52 1054.07 ;
      RECT 14346 1183.44 14374 1209.16 ;
      RECT 14372.145 1048.035 14374 1209.16 ;
      RECT 14346 1087.44 14367.235 1209.16 ;
      RECT 14369.555 1048.035 14374 1167.07 ;
      RECT 14352.55 1070.44 14374 1167.07 ;
      RECT 14346 1048.035 14364.645 1071.07 ;
      RECT 14346 1048.035 14374 1054.07 ;
      RECT 14330.48 1149.44 14343.48 1209.16 ;
      RECT 14342.865 1053.415 14343.48 1209.16 ;
      RECT 14330.48 1048.035 14335.115 1209.16 ;
      RECT 14330.48 1053.415 14343.48 1118.87 ;
      RECT 14330.48 1048.035 14341.85 1118.87 ;
      RECT 14330.48 1048.035 14343.48 1049.12 ;
      RECT 14313.5 1070.44 14326.5 1189.16 ;
      RECT 14316.865 1048.035 14326.5 1189.16 ;
      RECT 14313.5 1048.035 14326.5 1054.07 ;
      RECT 14296.52 1118.44 14309.52 1209.16 ;
      RECT 14298.375 1048.035 14309.52 1209.16 ;
      RECT 14296.52 1048.035 14309.52 1087.87 ;
      RECT 14266 1166.44 14294 1209.16 ;
      RECT 14280.475 1118.44 14294 1209.16 ;
      RECT 14266 1048.035 14275.565 1209.16 ;
      RECT 14266 1087.44 14290.625 1150.07 ;
      RECT 14284.53 1048.035 14294 1087.87 ;
      RECT 14280.475 1053.365 14294 1087.87 ;
      RECT 14266 1053.365 14294 1071.07 ;
      RECT 14266 1048.035 14278.81 1071.07 ;
      RECT 14266 1048.035 14294 1049.165 ;
      RECT 14250.48 1183.44 14263.48 1209.16 ;
      RECT 14258.145 1048.035 14263.48 1209.16 ;
      RECT 14253.475 1166.44 14263.48 1209.16 ;
      RECT 14250.48 1166.44 14263.48 1167.07 ;
      RECT 14250.48 1070.44 14253.235 1167.07 ;
      RECT 14250.48 1087.44 14263.48 1150.07 ;
      RECT 14250.48 1070.44 14263.48 1071.07 ;
      RECT 14253.475 1048.035 14263.48 1071.07 ;
      RECT 14250.48 1048.035 14263.48 1054.07 ;
      RECT 14216.52 1183.44 14229.52 1209.16 ;
      RECT 14216.52 1087.44 14227.235 1209.16 ;
      RECT 14221.75 1070.44 14229.52 1167.07 ;
      RECT 14216.52 1048.035 14224.565 1071.07 ;
      RECT 14216.52 1048.035 14229.52 1054.07 ;
      RECT 14186 1149.44 14214 1209.16 ;
      RECT 14204.63 1048.035 14214 1209.16 ;
      RECT 14202.865 1053.42 14214 1209.16 ;
      RECT 14186 1048.035 14195.115 1209.16 ;
      RECT 14186 1053.42 14214 1118.87 ;
      RECT 14186 1048.035 14201.85 1118.87 ;
      RECT 14186 1048.035 14214 1049.12 ;
      RECT 14170.48 1070.44 14183.48 1209.16 ;
      RECT 14176.865 1048.035 14183.48 1209.16 ;
      RECT 14170.48 1048.035 14171.955 1209.16 ;
      RECT 14170.48 1048.035 14183.48 1054.07 ;
      RECT 14153.5 1118.44 14166.5 1189.16 ;
      RECT 14158.375 1048.035 14166.5 1189.16 ;
      RECT 14153.5 1048.035 14166.5 1087.87 ;
      RECT 14136.52 1166.44 14149.52 1209.16 ;
      RECT 14144.53 1048.035 14149.52 1209.16 ;
      RECT 14140.475 1053.365 14149.52 1209.16 ;
      RECT 14136.52 1087.44 14149.52 1150.07 ;
      RECT 14136.52 1053.365 14149.52 1071.07 ;
      RECT 14136.52 1048.035 14138.81 1071.07 ;
      RECT 14136.52 1048.035 14149.52 1049.375 ;
      RECT 14106 1183.44 14134 1209.16 ;
      RECT 14118.145 1048.035 14134 1209.16 ;
      RECT 14113.475 1166.44 14134 1209.16 ;
      RECT 14106 1048.035 14108.565 1209.16 ;
      RECT 14106 1166.44 14134 1167.07 ;
      RECT 14106 1070.44 14113.235 1167.07 ;
      RECT 14106 1087.44 14134 1150.07 ;
      RECT 14106 1070.44 14134 1071.07 ;
      RECT 14113.475 1048.035 14134 1071.07 ;
      RECT 14106 1048.035 14134 1054.07 ;
      RECT 14090.48 1183.44 14103.48 1209.16 ;
      RECT 14092.145 1048.035 14103.48 1209.16 ;
      RECT 14090.48 1048.035 14103.48 1167.07 ;
      RECT 14073.5 1087.44 14086.5 1189.16 ;
      RECT 14080.13 1070.44 14086.5 1189.16 ;
      RECT 14073.5 1048.035 14083.455 1071.07 ;
      RECT 14073.5 1048.035 14086.5 1054.07 ;
      RECT 14056.52 1149.44 14069.52 1209.16 ;
      RECT 14064.63 1048.035 14069.52 1209.16 ;
      RECT 14062.865 1053.42 14069.52 1209.16 ;
      RECT 14056.52 1053.42 14069.52 1118.87 ;
      RECT 14056.52 1048.035 14061.85 1118.87 ;
      RECT 14056.52 1048.035 14069.52 1049.12 ;
      RECT 14026 1070.44 14054 1209.16 ;
      RECT 14036.865 1048.035 14054 1209.16 ;
      RECT 14026 1048.035 14031.955 1209.16 ;
      RECT 14026 1048.035 14054 1054.07 ;
      RECT 14010.48 1118.44 14023.48 1209.16 ;
      RECT 14018.375 1048.035 14023.48 1209.16 ;
      RECT 14010.48 1048.035 14023.48 1087.87 ;
      RECT 13993.5 1166.44 14006.5 1189.16 ;
      RECT 14004.43 1048.035 14006.5 1189.16 ;
      RECT 14000.475 1053.365 14006.5 1189.16 ;
      RECT 13993.5 1048.035 13995.565 1189.16 ;
      RECT 13993.5 1087.44 14006.5 1150.07 ;
      RECT 13993.5 1053.365 14006.5 1071.07 ;
      RECT 13993.5 1048.035 13998.81 1071.07 ;
      RECT 13993.5 1048.035 14006.5 1049.165 ;
      RECT 13976.52 1166.44 13989.52 1209.16 ;
      RECT 13978.145 1048.035 13989.52 1209.16 ;
      RECT 13976.52 1087.44 13989.52 1150.07 ;
      RECT 13976.52 1048.035 13989.52 1071.07 ;
      RECT 13946 1183.44 13974 1209.16 ;
      RECT 13952.145 1048.035 13968.565 1209.16 ;
      RECT 13946 1070.44 13947.235 1209.16 ;
      RECT 13946 1070.44 13973.235 1167.07 ;
      RECT 13946 1087.44 13974 1150.07 ;
      RECT 13948.365 1048.035 13968.565 1167.07 ;
      RECT 13946 1048.035 13974 1054.07 ;
      RECT 13930.48 1087.44 13943.48 1209.16 ;
      RECT 13930.48 1048.035 13936.835 1209.16 ;
      RECT 13930.48 1048.035 13943.48 1071.07 ;
      RECT 13913.5 1149.44 13926.5 1189.16 ;
      RECT 13924.63 1048.035 13926.5 1189.16 ;
      RECT 13922.865 1053.42 13926.5 1189.16 ;
      RECT 13913.5 1048.035 13915.115 1189.16 ;
      RECT 13913.5 1053.42 13926.5 1118.87 ;
      RECT 13913.5 1048.035 13921.85 1118.87 ;
      RECT 13913.5 1048.035 13926.5 1049.12 ;
      RECT 13896.52 1070.44 13909.52 1209.16 ;
      RECT 13896.865 1048.035 13909.52 1209.16 ;
      RECT 13896.52 1048.035 13909.52 1054.07 ;
      RECT 13866 1118.44 13894 1209.16 ;
      RECT 13878.375 1070.44 13894 1209.16 ;
      RECT 13866 1048.035 13870.625 1209.16 ;
      RECT 13866 1048.035 13891.955 1087.87 ;
      RECT 13866 1048.035 13894 1054.07 ;
      RECT 13850.48 1166.44 13863.48 1209.16 ;
      RECT 13860.475 1053.365 13863.48 1209.16 ;
      RECT 13850.48 1048.035 13855.565 1209.16 ;
      RECT 13850.48 1087.44 13863.48 1150.07 ;
      RECT 13850.48 1053.365 13863.48 1071.07 ;
      RECT 13850.48 1048.035 13858.81 1071.07 ;
      RECT 13850.48 1048.035 13863.48 1049.165 ;
      RECT 13833.5 1166.44 13846.5 1189.16 ;
      RECT 13838.145 1048.035 13846.5 1189.16 ;
      RECT 13837.98 1087.44 13846.5 1189.16 ;
      RECT 13833.5 1087.44 13846.5 1150.07 ;
      RECT 13833.5 1048.035 13846.5 1071.07 ;
      RECT 13816.52 1183.44 13829.52 1209.16 ;
      RECT 13816.52 1048.035 13828.565 1209.16 ;
      RECT 13816.52 1070.44 13829.52 1167.07 ;
      RECT 13816.52 1048.035 13829.52 1054.07 ;
      RECT 13786 1183.44 13814 1209.16 ;
      RECT 13812.145 1048.035 13814 1209.16 ;
      RECT 13786 1087.44 13807.235 1209.16 ;
      RECT 13809.555 1048.035 13814 1167.07 ;
      RECT 13792.55 1070.44 13814 1167.07 ;
      RECT 13786 1048.035 13804.645 1071.07 ;
      RECT 13786 1048.035 13814 1054.07 ;
      RECT 13770.48 1149.44 13783.48 1209.16 ;
      RECT 13782.865 1053.415 13783.48 1209.16 ;
      RECT 13770.48 1048.035 13775.115 1209.16 ;
      RECT 13770.48 1053.415 13783.48 1118.87 ;
      RECT 13770.48 1048.035 13781.85 1118.87 ;
      RECT 13770.48 1048.035 13783.48 1049.12 ;
      RECT 13753.5 1070.44 13766.5 1189.16 ;
      RECT 13756.865 1048.035 13766.5 1189.16 ;
      RECT 13753.5 1048.035 13766.5 1054.07 ;
      RECT 13736.52 1118.44 13749.52 1209.16 ;
      RECT 13738.375 1048.035 13749.52 1209.16 ;
      RECT 13736.52 1048.035 13749.52 1087.87 ;
      RECT 13706 1166.44 13734 1209.16 ;
      RECT 13720.475 1118.44 13734 1209.16 ;
      RECT 13706 1048.035 13715.565 1209.16 ;
      RECT 13706 1087.44 13730.625 1150.07 ;
      RECT 13724.53 1048.035 13734 1087.87 ;
      RECT 13720.475 1053.365 13734 1087.87 ;
      RECT 13706 1053.365 13734 1071.07 ;
      RECT 13706 1048.035 13718.81 1071.07 ;
      RECT 13706 1048.035 13734 1049.165 ;
      RECT 13690.48 1183.44 13703.48 1209.16 ;
      RECT 13698.145 1048.035 13703.48 1209.16 ;
      RECT 13693.475 1166.44 13703.48 1209.16 ;
      RECT 13690.48 1166.44 13703.48 1167.07 ;
      RECT 13690.48 1070.44 13693.235 1167.07 ;
      RECT 13690.48 1087.44 13703.48 1150.07 ;
      RECT 13690.48 1070.44 13703.48 1071.07 ;
      RECT 13693.475 1048.035 13703.48 1071.07 ;
      RECT 13690.48 1048.035 13703.48 1054.07 ;
      RECT 13656.52 1183.44 13669.52 1209.16 ;
      RECT 13656.52 1087.44 13667.235 1209.16 ;
      RECT 13661.75 1070.44 13669.52 1167.07 ;
      RECT 13656.52 1048.035 13664.565 1071.07 ;
      RECT 13656.52 1048.035 13669.52 1054.07 ;
      RECT 13626 1149.44 13654 1209.16 ;
      RECT 13644.63 1048.035 13654 1209.16 ;
      RECT 13642.865 1053.42 13654 1209.16 ;
      RECT 13626 1048.035 13635.115 1209.16 ;
      RECT 13626 1053.42 13654 1118.87 ;
      RECT 13626 1048.035 13641.85 1118.87 ;
      RECT 13626 1048.035 13654 1049.12 ;
      RECT 13610.48 1070.44 13623.48 1209.16 ;
      RECT 13616.865 1048.035 13623.48 1209.16 ;
      RECT 13610.48 1048.035 13611.955 1209.16 ;
      RECT 13610.48 1048.035 13623.48 1054.07 ;
      RECT 13593.5 1118.44 13606.5 1189.16 ;
      RECT 13598.375 1048.035 13606.5 1189.16 ;
      RECT 13593.5 1048.035 13606.5 1087.87 ;
      RECT 13576.52 1166.44 13589.52 1209.16 ;
      RECT 13584.53 1048.035 13589.52 1209.16 ;
      RECT 13580.475 1053.365 13589.52 1209.16 ;
      RECT 13576.52 1087.44 13589.52 1150.07 ;
      RECT 13576.52 1053.365 13589.52 1071.07 ;
      RECT 13576.52 1048.035 13578.81 1071.07 ;
      RECT 13576.52 1048.035 13589.52 1049.375 ;
      RECT 13546 1183.44 13574 1209.16 ;
      RECT 13558.145 1048.035 13574 1209.16 ;
      RECT 13553.475 1166.44 13574 1209.16 ;
      RECT 13546 1048.035 13548.565 1209.16 ;
      RECT 13546 1166.44 13574 1167.07 ;
      RECT 13546 1070.44 13553.235 1167.07 ;
      RECT 13546 1087.44 13574 1150.07 ;
      RECT 13546 1070.44 13574 1071.07 ;
      RECT 13553.475 1048.035 13574 1071.07 ;
      RECT 13546 1048.035 13574 1054.07 ;
      RECT 13530.48 1183.44 13543.48 1209.16 ;
      RECT 13532.145 1048.035 13543.48 1209.16 ;
      RECT 13530.48 1048.035 13543.48 1167.07 ;
      RECT 13513.5 1087.44 13526.5 1189.16 ;
      RECT 13520.13 1070.44 13526.5 1189.16 ;
      RECT 13513.5 1048.035 13523.455 1071.07 ;
      RECT 13513.5 1048.035 13526.5 1054.07 ;
      RECT 13496.52 1149.44 13509.52 1209.16 ;
      RECT 13504.63 1048.035 13509.52 1209.16 ;
      RECT 13502.865 1053.42 13509.52 1209.16 ;
      RECT 13496.52 1053.42 13509.52 1118.87 ;
      RECT 13496.52 1048.035 13501.85 1118.87 ;
      RECT 13496.52 1048.035 13509.52 1049.12 ;
      RECT 13466 1070.44 13494 1209.16 ;
      RECT 13476.865 1048.035 13494 1209.16 ;
      RECT 13466 1048.035 13471.955 1209.16 ;
      RECT 13466 1048.035 13494 1054.07 ;
      RECT 13450.48 1118.44 13463.48 1209.16 ;
      RECT 13458.375 1048.035 13463.48 1209.16 ;
      RECT 13450.48 1048.035 13463.48 1087.87 ;
      RECT 13433.5 1166.44 13446.5 1189.16 ;
      RECT 13444.43 1048.035 13446.5 1189.16 ;
      RECT 13440.475 1053.365 13446.5 1189.16 ;
      RECT 13433.5 1048.035 13435.565 1189.16 ;
      RECT 13433.5 1087.44 13446.5 1150.07 ;
      RECT 13433.5 1053.365 13446.5 1071.07 ;
      RECT 13433.5 1048.035 13438.81 1071.07 ;
      RECT 13433.5 1048.035 13446.5 1049.165 ;
      RECT 13416.52 1166.44 13429.52 1209.16 ;
      RECT 13418.145 1048.035 13429.52 1209.16 ;
      RECT 13416.52 1087.44 13429.52 1150.07 ;
      RECT 13416.52 1048.035 13429.52 1071.07 ;
      RECT 13386 1183.44 13414 1209.16 ;
      RECT 13392.145 1048.035 13408.565 1209.16 ;
      RECT 13386 1070.44 13387.235 1209.16 ;
      RECT 13386 1070.44 13413.235 1167.07 ;
      RECT 13386 1087.44 13414 1150.07 ;
      RECT 13388.365 1048.035 13408.565 1167.07 ;
      RECT 13386 1048.035 13414 1054.07 ;
      RECT 13370.48 1087.44 13383.48 1209.16 ;
      RECT 13370.48 1048.035 13376.835 1209.16 ;
      RECT 13370.48 1048.035 13383.48 1071.07 ;
      RECT 13353.5 1149.44 13366.5 1189.16 ;
      RECT 13364.63 1048.035 13366.5 1189.16 ;
      RECT 13362.865 1053.42 13366.5 1189.16 ;
      RECT 13353.5 1048.035 13355.115 1189.16 ;
      RECT 13353.5 1053.42 13366.5 1118.87 ;
      RECT 13353.5 1048.035 13361.85 1118.87 ;
      RECT 13353.5 1048.035 13366.5 1049.12 ;
      RECT 13336.52 1070.44 13349.52 1209.16 ;
      RECT 13336.865 1048.035 13349.52 1209.16 ;
      RECT 13336.52 1048.035 13349.52 1054.07 ;
      RECT 13306 1118.44 13334 1209.16 ;
      RECT 13318.375 1070.44 13334 1209.16 ;
      RECT 13306 1048.035 13310.625 1209.16 ;
      RECT 13306 1048.035 13331.955 1087.87 ;
      RECT 13306 1048.035 13334 1054.07 ;
      RECT 13290.48 1166.44 13303.48 1209.16 ;
      RECT 13300.475 1053.365 13303.48 1209.16 ;
      RECT 13290.48 1048.035 13295.565 1209.16 ;
      RECT 13290.48 1087.44 13303.48 1150.07 ;
      RECT 13290.48 1053.365 13303.48 1071.07 ;
      RECT 13290.48 1048.035 13298.81 1071.07 ;
      RECT 13290.48 1048.035 13303.48 1049.165 ;
      RECT 13273.5 1166.44 13286.5 1189.16 ;
      RECT 13278.145 1048.035 13286.5 1189.16 ;
      RECT 13277.98 1087.44 13286.5 1189.16 ;
      RECT 13273.5 1087.44 13286.5 1150.07 ;
      RECT 13273.5 1048.035 13286.5 1071.07 ;
      RECT 13256.52 1183.44 13269.52 1209.16 ;
      RECT 13256.52 1048.035 13268.565 1209.16 ;
      RECT 13256.52 1070.44 13269.52 1167.07 ;
      RECT 13256.52 1048.035 13269.52 1054.07 ;
      RECT 13226 1183.44 13254 1209.16 ;
      RECT 13252.145 1048.035 13254 1209.16 ;
      RECT 13226 1087.44 13247.235 1209.16 ;
      RECT 13249.555 1048.035 13254 1167.07 ;
      RECT 13232.55 1070.44 13254 1167.07 ;
      RECT 13226 1048.035 13244.645 1071.07 ;
      RECT 13226 1048.035 13254 1054.07 ;
      RECT 13210.48 1149.44 13223.48 1209.16 ;
      RECT 13222.865 1053.415 13223.48 1209.16 ;
      RECT 13210.48 1048.035 13215.115 1209.16 ;
      RECT 13210.48 1053.415 13223.48 1118.87 ;
      RECT 13210.48 1048.035 13221.85 1118.87 ;
      RECT 13210.48 1048.035 13223.48 1049.12 ;
      RECT 13193.5 1070.44 13206.5 1189.16 ;
      RECT 13196.865 1048.035 13206.5 1189.16 ;
      RECT 13193.5 1048.035 13206.5 1054.07 ;
      RECT 13176.52 1118.44 13189.52 1209.16 ;
      RECT 13178.375 1048.035 13189.52 1209.16 ;
      RECT 13176.52 1048.035 13189.52 1087.87 ;
      RECT 13146 1166.44 13174 1209.16 ;
      RECT 13160.475 1118.44 13174 1209.16 ;
      RECT 13146 1048.035 13155.565 1209.16 ;
      RECT 13146 1087.44 13170.625 1150.07 ;
      RECT 13164.53 1048.035 13174 1087.87 ;
      RECT 13160.475 1053.365 13174 1087.87 ;
      RECT 13146 1053.365 13174 1071.07 ;
      RECT 13146 1048.035 13158.81 1071.07 ;
      RECT 13146 1048.035 13174 1049.165 ;
      RECT 13130.48 1183.44 13143.48 1209.16 ;
      RECT 13138.145 1048.035 13143.48 1209.16 ;
      RECT 13133.475 1166.44 13143.48 1209.16 ;
      RECT 13130.48 1166.44 13143.48 1167.07 ;
      RECT 13130.48 1070.44 13133.235 1167.07 ;
      RECT 13130.48 1087.44 13143.48 1150.07 ;
      RECT 13130.48 1070.44 13143.48 1071.07 ;
      RECT 13133.475 1048.035 13143.48 1071.07 ;
      RECT 13130.48 1048.035 13143.48 1054.07 ;
      RECT 13096.52 1183.44 13109.52 1209.16 ;
      RECT 13096.52 1087.44 13107.235 1209.16 ;
      RECT 13101.75 1070.44 13109.52 1167.07 ;
      RECT 13096.52 1048.035 13104.565 1071.07 ;
      RECT 13096.52 1048.035 13109.52 1054.07 ;
      RECT 13066 1149.44 13094 1209.16 ;
      RECT 13084.63 1048.035 13094 1209.16 ;
      RECT 13082.865 1053.42 13094 1209.16 ;
      RECT 13066 1048.035 13075.115 1209.16 ;
      RECT 13066 1053.42 13094 1118.87 ;
      RECT 13066 1048.035 13081.85 1118.87 ;
      RECT 13066 1048.035 13094 1049.12 ;
      RECT 13050.48 1070.44 13063.48 1209.16 ;
      RECT 13056.865 1048.035 13063.48 1209.16 ;
      RECT 13050.48 1048.035 13051.955 1209.16 ;
      RECT 13050.48 1048.035 13063.48 1054.07 ;
      RECT 13033.5 1118.44 13046.5 1189.16 ;
      RECT 13038.375 1048.035 13046.5 1189.16 ;
      RECT 13033.5 1048.035 13046.5 1087.87 ;
      RECT 13016.52 1166.44 13029.52 1209.16 ;
      RECT 13024.53 1048.035 13029.52 1209.16 ;
      RECT 13020.475 1053.365 13029.52 1209.16 ;
      RECT 13016.52 1087.44 13029.52 1150.07 ;
      RECT 13016.52 1053.365 13029.52 1071.07 ;
      RECT 13016.52 1048.035 13018.81 1071.07 ;
      RECT 13016.52 1048.035 13029.52 1049.375 ;
      RECT 12986 1183.44 13014 1209.16 ;
      RECT 12998.145 1048.035 13014 1209.16 ;
      RECT 12993.475 1166.44 13014 1209.16 ;
      RECT 12986 1048.035 12988.565 1209.16 ;
      RECT 12986 1166.44 13014 1167.07 ;
      RECT 12986 1070.44 12993.235 1167.07 ;
      RECT 12986 1087.44 13014 1150.07 ;
      RECT 12986 1070.44 13014 1071.07 ;
      RECT 12993.475 1048.035 13014 1071.07 ;
      RECT 12986 1048.035 13014 1054.07 ;
      RECT 12970.48 1183.44 12983.48 1209.16 ;
      RECT 12972.145 1048.035 12983.48 1209.16 ;
      RECT 12970.48 1048.035 12983.48 1167.07 ;
      RECT 12953.5 1087.44 12966.5 1189.16 ;
      RECT 12960.13 1070.44 12966.5 1189.16 ;
      RECT 12953.5 1048.035 12963.455 1071.07 ;
      RECT 12953.5 1048.035 12966.5 1054.07 ;
      RECT 12936.52 1149.44 12949.52 1209.16 ;
      RECT 12944.63 1048.035 12949.52 1209.16 ;
      RECT 12942.865 1053.42 12949.52 1209.16 ;
      RECT 12936.52 1053.42 12949.52 1118.87 ;
      RECT 12936.52 1048.035 12941.85 1118.87 ;
      RECT 12936.52 1048.035 12949.52 1049.12 ;
      RECT 12906 1070.44 12934 1209.16 ;
      RECT 12916.865 1048.035 12934 1209.16 ;
      RECT 12906 1048.035 12911.955 1209.16 ;
      RECT 12906 1048.035 12934 1054.07 ;
      RECT 12890.48 1118.44 12903.48 1209.16 ;
      RECT 12898.375 1048.035 12903.48 1209.16 ;
      RECT 12890.48 1048.035 12903.48 1087.87 ;
      RECT 12873.5 1166.44 12886.5 1189.16 ;
      RECT 12884.43 1048.035 12886.5 1189.16 ;
      RECT 12880.475 1053.365 12886.5 1189.16 ;
      RECT 12873.5 1048.035 12875.565 1189.16 ;
      RECT 12873.5 1087.44 12886.5 1150.07 ;
      RECT 12873.5 1053.365 12886.5 1071.07 ;
      RECT 12873.5 1048.035 12878.81 1071.07 ;
      RECT 12873.5 1048.035 12886.5 1049.165 ;
      RECT 12856.52 1166.44 12869.52 1209.16 ;
      RECT 12858.145 1048.035 12869.52 1209.16 ;
      RECT 12856.52 1087.44 12869.52 1150.07 ;
      RECT 12856.52 1048.035 12869.52 1071.07 ;
      RECT 12826 1183.44 12854 1209.16 ;
      RECT 12832.145 1048.035 12848.565 1209.16 ;
      RECT 12826 1070.44 12827.235 1209.16 ;
      RECT 12826 1070.44 12853.235 1167.07 ;
      RECT 12826 1087.44 12854 1150.07 ;
      RECT 12828.365 1048.035 12848.565 1167.07 ;
      RECT 12826 1048.035 12854 1054.07 ;
      RECT 12810.48 1087.44 12823.48 1209.16 ;
      RECT 12810.48 1048.035 12816.835 1209.16 ;
      RECT 12810.48 1048.035 12823.48 1071.07 ;
      RECT 12793.5 1149.44 12806.5 1189.16 ;
      RECT 12804.63 1048.035 12806.5 1189.16 ;
      RECT 12802.865 1053.42 12806.5 1189.16 ;
      RECT 12793.5 1048.035 12795.115 1189.16 ;
      RECT 12793.5 1053.42 12806.5 1118.87 ;
      RECT 12793.5 1048.035 12801.85 1118.87 ;
      RECT 12793.5 1048.035 12806.5 1049.12 ;
      RECT 12776.52 1070.44 12789.52 1209.16 ;
      RECT 12776.865 1048.035 12789.52 1209.16 ;
      RECT 12776.52 1048.035 12789.52 1054.07 ;
      RECT 12746 1118.44 12774 1209.16 ;
      RECT 12758.375 1070.44 12774 1209.16 ;
      RECT 12746 1048.035 12750.625 1209.16 ;
      RECT 12746 1048.035 12771.955 1087.87 ;
      RECT 12746 1048.035 12774 1054.07 ;
      RECT 12730.48 1166.44 12743.48 1209.16 ;
      RECT 12740.475 1053.365 12743.48 1209.16 ;
      RECT 12730.48 1048.035 12735.565 1209.16 ;
      RECT 12730.48 1087.44 12743.48 1150.07 ;
      RECT 12730.48 1053.365 12743.48 1071.07 ;
      RECT 12730.48 1048.035 12738.81 1071.07 ;
      RECT 12730.48 1048.035 12743.48 1049.165 ;
      RECT 12713.5 1166.44 12726.5 1189.16 ;
      RECT 12718.145 1048.035 12726.5 1189.16 ;
      RECT 12717.98 1087.44 12726.5 1189.16 ;
      RECT 12713.5 1087.44 12726.5 1150.07 ;
      RECT 12713.5 1048.035 12726.5 1071.07 ;
      RECT 12696.52 1183.44 12709.52 1209.16 ;
      RECT 12696.52 1048.035 12708.565 1209.16 ;
      RECT 12696.52 1070.44 12709.52 1167.07 ;
      RECT 12696.52 1048.035 12709.52 1054.07 ;
      RECT 12666 1183.44 12694 1209.16 ;
      RECT 12692.145 1048.035 12694 1209.16 ;
      RECT 12666 1087.44 12687.235 1209.16 ;
      RECT 12689.555 1048.035 12694 1167.07 ;
      RECT 12672.55 1070.44 12694 1167.07 ;
      RECT 12666 1048.035 12684.645 1071.07 ;
      RECT 12666 1048.035 12694 1054.07 ;
      RECT 12650.48 1149.44 12663.48 1209.16 ;
      RECT 12662.865 1053.415 12663.48 1209.16 ;
      RECT 12650.48 1048.035 12655.115 1209.16 ;
      RECT 12650.48 1053.415 12663.48 1118.87 ;
      RECT 12650.48 1048.035 12661.85 1118.87 ;
      RECT 12650.48 1048.035 12663.48 1049.12 ;
      RECT 12633.5 1070.44 12646.5 1189.16 ;
      RECT 12636.865 1048.035 12646.5 1189.16 ;
      RECT 12633.5 1048.035 12646.5 1054.07 ;
      RECT 12616.52 1118.44 12629.52 1209.16 ;
      RECT 12618.375 1048.035 12629.52 1209.16 ;
      RECT 12616.52 1048.035 12629.52 1087.87 ;
      RECT 12586 1166.44 12614 1209.16 ;
      RECT 12600.475 1118.44 12614 1209.16 ;
      RECT 12586 1048.035 12595.565 1209.16 ;
      RECT 12586 1087.44 12610.625 1150.07 ;
      RECT 12604.53 1048.035 12614 1087.87 ;
      RECT 12600.475 1053.365 12614 1087.87 ;
      RECT 12586 1053.365 12614 1071.07 ;
      RECT 12586 1048.035 12598.81 1071.07 ;
      RECT 12586 1048.035 12614 1049.165 ;
      RECT 12570.48 1183.44 12583.48 1209.16 ;
      RECT 12578.145 1048.035 12583.48 1209.16 ;
      RECT 12573.475 1166.44 12583.48 1209.16 ;
      RECT 12570.48 1166.44 12583.48 1167.07 ;
      RECT 12570.48 1070.44 12573.235 1167.07 ;
      RECT 12570.48 1087.44 12583.48 1150.07 ;
      RECT 12570.48 1070.44 12583.48 1071.07 ;
      RECT 12573.475 1048.035 12583.48 1071.07 ;
      RECT 12570.48 1048.035 12583.48 1054.07 ;
      RECT 12536.52 1183.44 12549.52 1209.16 ;
      RECT 12536.52 1087.44 12547.235 1209.16 ;
      RECT 12541.75 1070.44 12549.52 1167.07 ;
      RECT 12536.52 1048.035 12544.565 1071.07 ;
      RECT 12536.52 1048.035 12549.52 1054.07 ;
      RECT 12506 1149.44 12534 1209.16 ;
      RECT 12524.63 1048.035 12534 1209.16 ;
      RECT 12522.865 1053.42 12534 1209.16 ;
      RECT 12506 1048.035 12515.115 1209.16 ;
      RECT 12506 1053.42 12534 1118.87 ;
      RECT 12506 1048.035 12521.85 1118.87 ;
      RECT 12506 1048.035 12534 1049.12 ;
      RECT 12490.48 1070.44 12503.48 1209.16 ;
      RECT 12496.865 1048.035 12503.48 1209.16 ;
      RECT 12490.48 1048.035 12491.955 1209.16 ;
      RECT 12490.48 1048.035 12503.48 1054.07 ;
      RECT 12473.5 1118.44 12486.5 1189.16 ;
      RECT 12478.375 1048.035 12486.5 1189.16 ;
      RECT 12473.5 1048.035 12486.5 1087.87 ;
      RECT 12456.52 1166.44 12469.52 1209.16 ;
      RECT 12464.53 1048.035 12469.52 1209.16 ;
      RECT 12460.475 1053.365 12469.52 1209.16 ;
      RECT 12456.52 1087.44 12469.52 1150.07 ;
      RECT 12456.52 1053.365 12469.52 1071.07 ;
      RECT 12456.52 1048.035 12458.81 1071.07 ;
      RECT 12456.52 1048.035 12469.52 1049.375 ;
      RECT 12426 1183.44 12454 1209.16 ;
      RECT 12438.145 1048.035 12454 1209.16 ;
      RECT 12433.475 1166.44 12454 1209.16 ;
      RECT 12426 1048.035 12428.565 1209.16 ;
      RECT 12426 1166.44 12454 1167.07 ;
      RECT 12426 1070.44 12433.235 1167.07 ;
      RECT 12426 1087.44 12454 1150.07 ;
      RECT 12426 1070.44 12454 1071.07 ;
      RECT 12433.475 1048.035 12454 1071.07 ;
      RECT 12426 1048.035 12454 1054.07 ;
      RECT 12410.48 1183.44 12423.48 1209.16 ;
      RECT 12412.145 1048.035 12423.48 1209.16 ;
      RECT 12410.48 1048.035 12423.48 1167.07 ;
      RECT 12393.5 1087.44 12406.5 1189.16 ;
      RECT 12400.13 1070.44 12406.5 1189.16 ;
      RECT 12393.5 1048.035 12403.455 1071.07 ;
      RECT 12393.5 1048.035 12406.5 1054.07 ;
      RECT 12376.52 1149.44 12389.52 1209.16 ;
      RECT 12384.63 1048.035 12389.52 1209.16 ;
      RECT 12382.865 1053.42 12389.52 1209.16 ;
      RECT 12376.52 1053.42 12389.52 1118.87 ;
      RECT 12376.52 1048.035 12381.85 1118.87 ;
      RECT 12376.52 1048.035 12389.52 1049.12 ;
      RECT 12346 1070.44 12374 1209.16 ;
      RECT 12356.865 1048.035 12374 1209.16 ;
      RECT 12346 1048.035 12351.955 1209.16 ;
      RECT 12346 1048.035 12374 1054.07 ;
      RECT 12330.48 1118.44 12343.48 1209.16 ;
      RECT 12338.375 1048.035 12343.48 1209.16 ;
      RECT 12330.48 1048.035 12343.48 1087.87 ;
      RECT 12313.5 1166.44 12326.5 1189.16 ;
      RECT 12324.43 1048.035 12326.5 1189.16 ;
      RECT 12320.475 1053.365 12326.5 1189.16 ;
      RECT 12313.5 1048.035 12315.565 1189.16 ;
      RECT 12313.5 1087.44 12326.5 1150.07 ;
      RECT 12313.5 1053.365 12326.5 1071.07 ;
      RECT 12313.5 1048.035 12318.81 1071.07 ;
      RECT 12313.5 1048.035 12326.5 1049.165 ;
      RECT 12296.52 1166.44 12309.52 1209.16 ;
      RECT 12298.145 1048.035 12309.52 1209.16 ;
      RECT 12296.52 1087.44 12309.52 1150.07 ;
      RECT 12296.52 1048.035 12309.52 1071.07 ;
      RECT 12266 1183.44 12294 1209.16 ;
      RECT 12272.145 1048.035 12288.565 1209.16 ;
      RECT 12266 1070.44 12267.235 1209.16 ;
      RECT 12266 1070.44 12293.235 1167.07 ;
      RECT 12266 1087.44 12294 1150.07 ;
      RECT 12268.365 1048.035 12288.565 1167.07 ;
      RECT 12266 1048.035 12294 1054.07 ;
      RECT 12250.48 1087.44 12263.48 1209.16 ;
      RECT 12250.48 1048.035 12256.835 1209.16 ;
      RECT 12250.48 1048.035 12263.48 1071.07 ;
      RECT 12233.5 1149.44 12246.5 1189.16 ;
      RECT 12244.63 1048.035 12246.5 1189.16 ;
      RECT 12242.865 1053.42 12246.5 1189.16 ;
      RECT 12233.5 1048.035 12235.115 1189.16 ;
      RECT 12233.5 1053.42 12246.5 1118.87 ;
      RECT 12233.5 1048.035 12241.85 1118.87 ;
      RECT 12233.5 1048.035 12246.5 1049.12 ;
      RECT 12216.52 1070.44 12229.52 1209.16 ;
      RECT 12216.865 1048.035 12229.52 1209.16 ;
      RECT 12216.52 1048.035 12229.52 1054.07 ;
      RECT 12186 1118.44 12214 1209.16 ;
      RECT 12198.375 1070.44 12214 1209.16 ;
      RECT 12186 1048.035 12190.625 1209.16 ;
      RECT 12186 1048.035 12211.955 1087.87 ;
      RECT 12186 1048.035 12214 1054.07 ;
      RECT 12170.48 1166.44 12183.48 1209.16 ;
      RECT 12180.475 1053.365 12183.48 1209.16 ;
      RECT 12170.48 1048.035 12175.565 1209.16 ;
      RECT 12170.48 1087.44 12183.48 1150.07 ;
      RECT 12170.48 1053.365 12183.48 1071.07 ;
      RECT 12170.48 1048.035 12178.81 1071.07 ;
      RECT 12170.48 1048.035 12183.48 1049.165 ;
      RECT 12153.5 1166.44 12166.5 1189.16 ;
      RECT 12158.145 1048.035 12166.5 1189.16 ;
      RECT 12157.98 1087.44 12166.5 1189.16 ;
      RECT 12153.5 1087.44 12166.5 1150.07 ;
      RECT 12153.5 1048.035 12166.5 1071.07 ;
      RECT 12136.52 1183.44 12149.52 1209.16 ;
      RECT 12136.52 1048.035 12148.565 1209.16 ;
      RECT 12136.52 1070.44 12149.52 1167.07 ;
      RECT 12136.52 1048.035 12149.52 1054.07 ;
      RECT 12106 1183.44 12134 1209.16 ;
      RECT 12132.145 1048.035 12134 1209.16 ;
      RECT 12106 1087.44 12127.235 1209.16 ;
      RECT 12129.555 1048.035 12134 1167.07 ;
      RECT 12112.55 1070.44 12134 1167.07 ;
      RECT 12106 1048.035 12124.645 1071.07 ;
      RECT 12106 1048.035 12134 1054.07 ;
      RECT 12090.48 1149.44 12103.48 1209.16 ;
      RECT 12102.865 1053.415 12103.48 1209.16 ;
      RECT 12090.48 1048.035 12095.115 1209.16 ;
      RECT 12090.48 1053.415 12103.48 1118.87 ;
      RECT 12090.48 1048.035 12101.85 1118.87 ;
      RECT 12090.48 1048.035 12103.48 1049.12 ;
      RECT 12073.5 1070.44 12086.5 1189.16 ;
      RECT 12076.865 1048.035 12086.5 1189.16 ;
      RECT 12073.5 1048.035 12086.5 1054.07 ;
      RECT 12056.52 1118.44 12069.52 1209.16 ;
      RECT 12058.375 1048.035 12069.52 1209.16 ;
      RECT 12056.52 1048.035 12069.52 1087.87 ;
      RECT 12026 1166.44 12054 1209.16 ;
      RECT 12040.475 1118.44 12054 1209.16 ;
      RECT 12026 1048.035 12035.565 1209.16 ;
      RECT 12026 1087.44 12050.625 1150.07 ;
      RECT 12044.53 1048.035 12054 1087.87 ;
      RECT 12040.475 1053.365 12054 1087.87 ;
      RECT 12026 1053.365 12054 1071.07 ;
      RECT 12026 1048.035 12038.81 1071.07 ;
      RECT 12026 1048.035 12054 1049.165 ;
      RECT 12010.48 1183.44 12023.48 1209.16 ;
      RECT 12018.145 1048.035 12023.48 1209.16 ;
      RECT 12013.475 1166.44 12023.48 1209.16 ;
      RECT 12010.48 1166.44 12023.48 1167.07 ;
      RECT 12010.48 1070.44 12013.235 1167.07 ;
      RECT 12010.48 1087.44 12023.48 1150.07 ;
      RECT 12010.48 1070.44 12023.48 1071.07 ;
      RECT 12013.475 1048.035 12023.48 1071.07 ;
      RECT 12010.48 1048.035 12023.48 1054.07 ;
      RECT 11976.52 1183.44 11989.52 1209.16 ;
      RECT 11976.52 1087.44 11987.235 1209.16 ;
      RECT 11981.75 1070.44 11989.52 1167.07 ;
      RECT 11976.52 1048.035 11984.565 1071.07 ;
      RECT 11976.52 1048.035 11989.52 1054.07 ;
      RECT 11946 1149.44 11974 1209.16 ;
      RECT 11964.63 1048.035 11974 1209.16 ;
      RECT 11962.865 1053.42 11974 1209.16 ;
      RECT 11946 1048.035 11955.115 1209.16 ;
      RECT 11946 1053.42 11974 1118.87 ;
      RECT 11946 1048.035 11961.85 1118.87 ;
      RECT 11946 1048.035 11974 1049.12 ;
      RECT 11930.48 1070.44 11943.48 1209.16 ;
      RECT 11936.865 1048.035 11943.48 1209.16 ;
      RECT 11930.48 1048.035 11931.955 1209.16 ;
      RECT 11930.48 1048.035 11943.48 1054.07 ;
      RECT 11913.5 1118.44 11926.5 1189.16 ;
      RECT 11918.375 1048.035 11926.5 1189.16 ;
      RECT 11913.5 1048.035 11926.5 1087.87 ;
      RECT 11896.52 1166.44 11909.52 1209.16 ;
      RECT 11904.53 1048.035 11909.52 1209.16 ;
      RECT 11900.475 1053.365 11909.52 1209.16 ;
      RECT 11896.52 1087.44 11909.52 1150.07 ;
      RECT 11896.52 1053.365 11909.52 1071.07 ;
      RECT 11896.52 1048.035 11898.81 1071.07 ;
      RECT 11896.52 1048.035 11909.52 1049.375 ;
      RECT 11866 1183.44 11894 1209.16 ;
      RECT 11878.145 1048.035 11894 1209.16 ;
      RECT 11873.475 1166.44 11894 1209.16 ;
      RECT 11866 1048.035 11868.565 1209.16 ;
      RECT 11866 1166.44 11894 1167.07 ;
      RECT 11866 1070.44 11873.235 1167.07 ;
      RECT 11866 1087.44 11894 1150.07 ;
      RECT 11866 1070.44 11894 1071.07 ;
      RECT 11873.475 1048.035 11894 1071.07 ;
      RECT 11866 1048.035 11894 1054.07 ;
      RECT 11850.48 1183.44 11863.48 1209.16 ;
      RECT 11852.145 1048.035 11863.48 1209.16 ;
      RECT 11850.48 1048.035 11863.48 1167.07 ;
      RECT 11833.5 1087.44 11846.5 1189.16 ;
      RECT 11840.13 1070.44 11846.5 1189.16 ;
      RECT 11833.5 1048.035 11843.455 1071.07 ;
      RECT 11833.5 1048.035 11846.5 1054.07 ;
      RECT 11816.52 1149.44 11829.52 1209.16 ;
      RECT 11824.63 1048.035 11829.52 1209.16 ;
      RECT 11822.865 1053.42 11829.52 1209.16 ;
      RECT 11816.52 1053.42 11829.52 1118.87 ;
      RECT 11816.52 1048.035 11821.85 1118.87 ;
      RECT 11816.52 1048.035 11829.52 1049.12 ;
      RECT 11786 1070.44 11814 1209.16 ;
      RECT 11796.865 1048.035 11814 1209.16 ;
      RECT 11786 1048.035 11791.955 1209.16 ;
      RECT 11786 1048.035 11814 1054.07 ;
      RECT 11770.48 1118.44 11783.48 1209.16 ;
      RECT 11778.375 1048.035 11783.48 1209.16 ;
      RECT 11770.48 1048.035 11783.48 1087.87 ;
      RECT 11753.5 1166.44 11766.5 1189.16 ;
      RECT 11764.43 1048.035 11766.5 1189.16 ;
      RECT 11760.475 1053.365 11766.5 1189.16 ;
      RECT 11753.5 1048.035 11755.565 1189.16 ;
      RECT 11753.5 1087.44 11766.5 1150.07 ;
      RECT 11753.5 1053.365 11766.5 1071.07 ;
      RECT 11753.5 1048.035 11758.81 1071.07 ;
      RECT 11753.5 1048.035 11766.5 1049.165 ;
      RECT 11736.52 1166.44 11749.52 1209.16 ;
      RECT 11738.145 1048.035 11749.52 1209.16 ;
      RECT 11736.52 1087.44 11749.52 1150.07 ;
      RECT 11736.52 1048.035 11749.52 1071.07 ;
      RECT 11706 1183.44 11734 1209.16 ;
      RECT 11712.145 1048.035 11728.565 1209.16 ;
      RECT 11706 1070.44 11707.235 1209.16 ;
      RECT 11706 1070.44 11733.235 1167.07 ;
      RECT 11706 1087.44 11734 1150.07 ;
      RECT 11708.365 1048.035 11728.565 1167.07 ;
      RECT 11706 1048.035 11734 1054.07 ;
      RECT 11690.48 1087.44 11703.48 1209.16 ;
      RECT 11690.48 1048.035 11696.835 1209.16 ;
      RECT 11690.48 1048.035 11703.48 1071.07 ;
      RECT 11673.5 1149.44 11686.5 1189.16 ;
      RECT 11684.63 1048.035 11686.5 1189.16 ;
      RECT 11682.865 1053.42 11686.5 1189.16 ;
      RECT 11673.5 1048.035 11675.115 1189.16 ;
      RECT 11673.5 1053.42 11686.5 1118.87 ;
      RECT 11673.5 1048.035 11681.85 1118.87 ;
      RECT 11673.5 1048.035 11686.5 1049.12 ;
      RECT 11656.52 1070.44 11669.52 1209.16 ;
      RECT 11656.865 1048.035 11669.52 1209.16 ;
      RECT 11656.52 1048.035 11669.52 1054.07 ;
      RECT 11626 1118.44 11654 1209.16 ;
      RECT 11638.375 1070.44 11654 1209.16 ;
      RECT 11626 1048.035 11630.625 1209.16 ;
      RECT 11626 1048.035 11651.955 1087.87 ;
      RECT 11626 1048.035 11654 1054.07 ;
      RECT 11610.48 1166.44 11623.48 1209.16 ;
      RECT 11620.475 1053.365 11623.48 1209.16 ;
      RECT 11610.48 1048.035 11615.565 1209.16 ;
      RECT 11610.48 1087.44 11623.48 1150.07 ;
      RECT 11610.48 1053.365 11623.48 1071.07 ;
      RECT 11610.48 1048.035 11618.81 1071.07 ;
      RECT 11610.48 1048.035 11623.48 1049.165 ;
      RECT 11593.5 1166.44 11606.5 1189.16 ;
      RECT 11598.145 1048.035 11606.5 1189.16 ;
      RECT 11597.98 1087.44 11606.5 1189.16 ;
      RECT 11593.5 1087.44 11606.5 1150.07 ;
      RECT 11593.5 1048.035 11606.5 1071.07 ;
      RECT 11576.52 1183.44 11589.52 1209.16 ;
      RECT 11576.52 1048.035 11588.565 1209.16 ;
      RECT 11576.52 1070.44 11589.52 1167.07 ;
      RECT 11576.52 1048.035 11589.52 1054.07 ;
      RECT 11546 1183.44 11574 1209.16 ;
      RECT 11572.145 1048.035 11574 1209.16 ;
      RECT 11546 1087.44 11567.235 1209.16 ;
      RECT 11569.555 1048.035 11574 1167.07 ;
      RECT 11552.55 1070.44 11574 1167.07 ;
      RECT 11546 1048.035 11564.645 1071.07 ;
      RECT 11546 1048.035 11574 1054.07 ;
      RECT 11530.48 1149.44 11543.48 1209.16 ;
      RECT 11542.865 1053.415 11543.48 1209.16 ;
      RECT 11530.48 1048.035 11535.115 1209.16 ;
      RECT 11530.48 1053.415 11543.48 1118.87 ;
      RECT 11530.48 1048.035 11541.85 1118.87 ;
      RECT 11530.48 1048.035 11543.48 1049.12 ;
      RECT 11513.5 1070.44 11526.5 1189.16 ;
      RECT 11516.865 1048.035 11526.5 1189.16 ;
      RECT 11513.5 1048.035 11526.5 1054.07 ;
      RECT 11496.52 1118.44 11509.52 1209.16 ;
      RECT 11498.375 1048.035 11509.52 1209.16 ;
      RECT 11496.52 1048.035 11509.52 1087.87 ;
      RECT 11466 1166.44 11494 1209.16 ;
      RECT 11480.475 1118.44 11494 1209.16 ;
      RECT 11466 1048.035 11475.565 1209.16 ;
      RECT 11466 1087.44 11490.625 1150.07 ;
      RECT 11484.53 1048.035 11494 1087.87 ;
      RECT 11480.475 1053.365 11494 1087.87 ;
      RECT 11466 1053.365 11494 1071.07 ;
      RECT 11466 1048.035 11478.81 1071.07 ;
      RECT 11466 1048.035 11494 1049.165 ;
      RECT 11450.48 1183.44 11463.48 1209.16 ;
      RECT 11458.145 1048.035 11463.48 1209.16 ;
      RECT 11453.475 1166.44 11463.48 1209.16 ;
      RECT 11450.48 1166.44 11463.48 1167.07 ;
      RECT 11450.48 1070.44 11453.235 1167.07 ;
      RECT 11450.48 1087.44 11463.48 1150.07 ;
      RECT 11450.48 1070.44 11463.48 1071.07 ;
      RECT 11453.475 1048.035 11463.48 1071.07 ;
      RECT 11450.48 1048.035 11463.48 1054.07 ;
      RECT 11416.52 1183.44 11429.52 1209.16 ;
      RECT 11416.52 1087.44 11427.235 1209.16 ;
      RECT 11421.75 1070.44 11429.52 1167.07 ;
      RECT 11416.52 1048.035 11424.565 1071.07 ;
      RECT 11416.52 1048.035 11429.52 1054.07 ;
      RECT 11386 1149.44 11414 1209.16 ;
      RECT 11404.63 1048.035 11414 1209.16 ;
      RECT 11402.865 1053.42 11414 1209.16 ;
      RECT 11386 1048.035 11395.115 1209.16 ;
      RECT 11386 1053.42 11414 1118.87 ;
      RECT 11386 1048.035 11401.85 1118.87 ;
      RECT 11386 1048.035 11414 1049.12 ;
      RECT 11370.48 1070.44 11383.48 1209.16 ;
      RECT 11376.865 1048.035 11383.48 1209.16 ;
      RECT 11370.48 1048.035 11371.955 1209.16 ;
      RECT 11370.48 1048.035 11383.48 1054.07 ;
      RECT 11353.5 1118.44 11366.5 1189.16 ;
      RECT 11358.375 1048.035 11366.5 1189.16 ;
      RECT 11353.5 1048.035 11366.5 1087.87 ;
      RECT 11336.52 1166.44 11349.52 1209.16 ;
      RECT 11344.53 1048.035 11349.52 1209.16 ;
      RECT 11340.475 1053.365 11349.52 1209.16 ;
      RECT 11336.52 1087.44 11349.52 1150.07 ;
      RECT 11336.52 1053.365 11349.52 1071.07 ;
      RECT 11336.52 1048.035 11338.81 1071.07 ;
      RECT 11336.52 1048.035 11349.52 1049.375 ;
      RECT 11306 1183.44 11334 1209.16 ;
      RECT 11318.145 1048.035 11334 1209.16 ;
      RECT 11313.475 1166.44 11334 1209.16 ;
      RECT 11306 1048.035 11308.565 1209.16 ;
      RECT 11306 1166.44 11334 1167.07 ;
      RECT 11306 1070.44 11313.235 1167.07 ;
      RECT 11306 1087.44 11334 1150.07 ;
      RECT 11306 1070.44 11334 1071.07 ;
      RECT 11313.475 1048.035 11334 1071.07 ;
      RECT 11306 1048.035 11334 1054.07 ;
      RECT 11290.48 1183.44 11303.48 1209.16 ;
      RECT 11292.145 1048.035 11303.48 1209.16 ;
      RECT 11290.48 1048.035 11303.48 1167.07 ;
      RECT 11273.5 1087.44 11286.5 1189.16 ;
      RECT 11280.13 1070.44 11286.5 1189.16 ;
      RECT 11273.5 1048.035 11283.455 1071.07 ;
      RECT 11273.5 1048.035 11286.5 1054.07 ;
      RECT 11256.52 1149.44 11269.52 1209.16 ;
      RECT 11264.63 1048.035 11269.52 1209.16 ;
      RECT 11262.865 1053.42 11269.52 1209.16 ;
      RECT 11256.52 1053.42 11269.52 1118.87 ;
      RECT 11256.52 1048.035 11261.85 1118.87 ;
      RECT 11256.52 1048.035 11269.52 1049.12 ;
      RECT 11226 1070.44 11254 1209.16 ;
      RECT 11236.865 1048.035 11254 1209.16 ;
      RECT 11226 1048.035 11231.955 1209.16 ;
      RECT 11226 1048.035 11254 1054.07 ;
      RECT 11210.48 1118.44 11223.48 1209.16 ;
      RECT 11218.375 1048.035 11223.48 1209.16 ;
      RECT 11210.48 1048.035 11223.48 1087.87 ;
      RECT 11193.5 1166.44 11206.5 1189.16 ;
      RECT 11204.43 1048.035 11206.5 1189.16 ;
      RECT 11200.475 1053.365 11206.5 1189.16 ;
      RECT 11193.5 1048.035 11195.565 1189.16 ;
      RECT 11193.5 1087.44 11206.5 1150.07 ;
      RECT 11193.5 1053.365 11206.5 1071.07 ;
      RECT 11193.5 1048.035 11198.81 1071.07 ;
      RECT 11193.5 1048.035 11206.5 1049.165 ;
      RECT 11176.52 1166.44 11189.52 1209.16 ;
      RECT 11178.145 1048.035 11189.52 1209.16 ;
      RECT 11176.52 1087.44 11189.52 1150.07 ;
      RECT 11176.52 1048.035 11189.52 1071.07 ;
      RECT 11146 1183.44 11174 1209.16 ;
      RECT 11152.145 1048.035 11168.565 1209.16 ;
      RECT 11146 1070.44 11147.235 1209.16 ;
      RECT 11146 1070.44 11173.235 1167.07 ;
      RECT 11146 1087.44 11174 1150.07 ;
      RECT 11148.365 1048.035 11168.565 1167.07 ;
      RECT 11146 1048.035 11174 1054.07 ;
      RECT 11130.48 1087.44 11143.48 1209.16 ;
      RECT 11130.48 1048.035 11136.835 1209.16 ;
      RECT 11130.48 1048.035 11143.48 1071.07 ;
      RECT 11113.5 1149.44 11126.5 1189.16 ;
      RECT 11124.63 1048.035 11126.5 1189.16 ;
      RECT 11122.865 1053.42 11126.5 1189.16 ;
      RECT 11113.5 1048.035 11115.115 1189.16 ;
      RECT 11113.5 1053.42 11126.5 1118.87 ;
      RECT 11113.5 1048.035 11121.85 1118.87 ;
      RECT 11113.5 1048.035 11126.5 1049.12 ;
      RECT 11096.52 1070.44 11109.52 1209.16 ;
      RECT 11096.865 1048.035 11109.52 1209.16 ;
      RECT 11096.52 1048.035 11109.52 1054.07 ;
      RECT 11066 1118.44 11094 1209.16 ;
      RECT 11078.375 1070.44 11094 1209.16 ;
      RECT 11066 1048.035 11070.625 1209.16 ;
      RECT 11066 1048.035 11091.955 1087.87 ;
      RECT 11066 1048.035 11094 1054.07 ;
      RECT 11050.48 1166.44 11063.48 1209.16 ;
      RECT 11060.475 1053.365 11063.48 1209.16 ;
      RECT 11050.48 1048.035 11055.565 1209.16 ;
      RECT 11050.48 1087.44 11063.48 1150.07 ;
      RECT 11050.48 1053.365 11063.48 1071.07 ;
      RECT 11050.48 1048.035 11058.81 1071.07 ;
      RECT 11050.48 1048.035 11063.48 1049.165 ;
      RECT 11033.5 1166.44 11046.5 1189.16 ;
      RECT 11038.145 1048.035 11046.5 1189.16 ;
      RECT 11037.98 1087.44 11046.5 1189.16 ;
      RECT 11033.5 1087.44 11046.5 1150.07 ;
      RECT 11033.5 1048.035 11046.5 1071.07 ;
      RECT 11016.52 1183.44 11029.52 1209.16 ;
      RECT 11016.52 1048.035 11028.565 1209.16 ;
      RECT 11016.52 1070.44 11029.52 1167.07 ;
      RECT 11016.52 1048.035 11029.52 1054.07 ;
      RECT 10986 1183.44 11014 1209.16 ;
      RECT 11012.145 1048.035 11014 1209.16 ;
      RECT 10986 1087.44 11007.235 1209.16 ;
      RECT 11009.555 1048.035 11014 1167.07 ;
      RECT 10992.55 1070.44 11014 1167.07 ;
      RECT 10986 1048.035 11004.645 1071.07 ;
      RECT 10986 1048.035 11014 1054.07 ;
      RECT 10970.48 1149.44 10983.48 1209.16 ;
      RECT 10982.865 1053.415 10983.48 1209.16 ;
      RECT 10970.48 1048.035 10975.115 1209.16 ;
      RECT 10970.48 1053.415 10983.48 1118.87 ;
      RECT 10970.48 1048.035 10981.85 1118.87 ;
      RECT 10970.48 1048.035 10983.48 1049.12 ;
      RECT 10953.5 1070.44 10966.5 1189.16 ;
      RECT 10956.865 1048.035 10966.5 1189.16 ;
      RECT 10953.5 1048.035 10966.5 1054.07 ;
      RECT 10936.52 1118.44 10949.52 1209.16 ;
      RECT 10938.375 1048.035 10949.52 1209.16 ;
      RECT 10936.52 1048.035 10949.52 1087.87 ;
      RECT 10906 1166.44 10934 1209.16 ;
      RECT 10920.475 1118.44 10934 1209.16 ;
      RECT 10906 1048.035 10915.565 1209.16 ;
      RECT 10906 1087.44 10930.625 1150.07 ;
      RECT 10924.53 1048.035 10934 1087.87 ;
      RECT 10920.475 1053.365 10934 1087.87 ;
      RECT 10906 1053.365 10934 1071.07 ;
      RECT 10906 1048.035 10918.81 1071.07 ;
      RECT 10906 1048.035 10934 1049.165 ;
      RECT 10890.48 1183.44 10903.48 1209.16 ;
      RECT 10898.145 1048.035 10903.48 1209.16 ;
      RECT 10893.475 1166.44 10903.48 1209.16 ;
      RECT 10890.48 1166.44 10903.48 1167.07 ;
      RECT 10890.48 1070.44 10893.235 1167.07 ;
      RECT 10890.48 1087.44 10903.48 1150.07 ;
      RECT 10890.48 1070.44 10903.48 1071.07 ;
      RECT 10893.475 1048.035 10903.48 1071.07 ;
      RECT 10890.48 1048.035 10903.48 1054.07 ;
      RECT 10856.52 1183.44 10869.52 1209.16 ;
      RECT 10856.52 1087.44 10867.235 1209.16 ;
      RECT 10861.75 1070.44 10869.52 1167.07 ;
      RECT 10856.52 1048.035 10864.565 1071.07 ;
      RECT 10856.52 1048.035 10869.52 1054.07 ;
      RECT 10826 1149.44 10854 1209.16 ;
      RECT 10844.63 1048.035 10854 1209.16 ;
      RECT 10842.865 1053.42 10854 1209.16 ;
      RECT 10826 1048.035 10835.115 1209.16 ;
      RECT 10826 1053.42 10854 1118.87 ;
      RECT 10826 1048.035 10841.85 1118.87 ;
      RECT 10826 1048.035 10854 1049.12 ;
      RECT 10810.48 1070.44 10823.48 1209.16 ;
      RECT 10816.865 1048.035 10823.48 1209.16 ;
      RECT 10810.48 1048.035 10811.955 1209.16 ;
      RECT 10810.48 1048.035 10823.48 1054.07 ;
      RECT 10793.5 1118.44 10806.5 1189.16 ;
      RECT 10798.375 1048.035 10806.5 1189.16 ;
      RECT 10793.5 1048.035 10806.5 1087.87 ;
      RECT 10776.52 1166.44 10789.52 1209.16 ;
      RECT 10784.53 1048.035 10789.52 1209.16 ;
      RECT 10780.475 1053.365 10789.52 1209.16 ;
      RECT 10776.52 1087.44 10789.52 1150.07 ;
      RECT 10776.52 1053.365 10789.52 1071.07 ;
      RECT 10776.52 1048.035 10778.81 1071.07 ;
      RECT 10776.52 1048.035 10789.52 1049.375 ;
      RECT 10746 1183.44 10774 1209.16 ;
      RECT 10758.145 1048.035 10774 1209.16 ;
      RECT 10753.475 1166.44 10774 1209.16 ;
      RECT 10746 1048.035 10748.565 1209.16 ;
      RECT 10746 1166.44 10774 1167.07 ;
      RECT 10746 1070.44 10753.235 1167.07 ;
      RECT 10746 1087.44 10774 1150.07 ;
      RECT 10746 1070.44 10774 1071.07 ;
      RECT 10753.475 1048.035 10774 1071.07 ;
      RECT 10746 1048.035 10774 1054.07 ;
      RECT 10730.48 1183.44 10743.48 1209.16 ;
      RECT 10732.145 1048.035 10743.48 1209.16 ;
      RECT 10730.48 1048.035 10743.48 1167.07 ;
      RECT 10713.5 1087.44 10726.5 1189.16 ;
      RECT 10720.13 1070.44 10726.5 1189.16 ;
      RECT 10713.5 1048.035 10723.455 1071.07 ;
      RECT 10713.5 1048.035 10726.5 1054.07 ;
      RECT 10696.52 1149.44 10709.52 1209.16 ;
      RECT 10704.63 1048.035 10709.52 1209.16 ;
      RECT 10702.865 1053.42 10709.52 1209.16 ;
      RECT 10696.52 1053.42 10709.52 1118.87 ;
      RECT 10696.52 1048.035 10701.85 1118.87 ;
      RECT 10696.52 1048.035 10709.52 1049.12 ;
      RECT 10666 1070.44 10694 1209.16 ;
      RECT 10676.865 1048.035 10694 1209.16 ;
      RECT 10666 1048.035 10671.955 1209.16 ;
      RECT 10666 1048.035 10694 1054.07 ;
      RECT 10650.48 1118.44 10663.48 1209.16 ;
      RECT 10658.375 1048.035 10663.48 1209.16 ;
      RECT 10650.48 1048.035 10663.48 1087.87 ;
      RECT 10633.5 1166.44 10646.5 1189.16 ;
      RECT 10644.43 1048.035 10646.5 1189.16 ;
      RECT 10640.475 1053.365 10646.5 1189.16 ;
      RECT 10633.5 1048.035 10635.565 1189.16 ;
      RECT 10633.5 1087.44 10646.5 1150.07 ;
      RECT 10633.5 1053.365 10646.5 1071.07 ;
      RECT 10633.5 1048.035 10638.81 1071.07 ;
      RECT 10633.5 1048.035 10646.5 1049.165 ;
      RECT 10616.52 1166.44 10629.52 1209.16 ;
      RECT 10618.145 1048.035 10629.52 1209.16 ;
      RECT 10616.52 1087.44 10629.52 1150.07 ;
      RECT 10616.52 1048.035 10629.52 1071.07 ;
      RECT 10586 1183.44 10614 1209.16 ;
      RECT 10592.145 1048.035 10608.565 1209.16 ;
      RECT 10586 1070.44 10587.235 1209.16 ;
      RECT 10586 1070.44 10613.235 1167.07 ;
      RECT 10586 1087.44 10614 1150.07 ;
      RECT 10588.365 1048.035 10608.565 1167.07 ;
      RECT 10586 1048.035 10614 1054.07 ;
      RECT 10570.48 1087.44 10583.48 1209.16 ;
      RECT 10570.48 1048.035 10576.835 1209.16 ;
      RECT 10570.48 1048.035 10583.48 1071.07 ;
      RECT 10553.5 1149.44 10566.5 1189.16 ;
      RECT 10564.63 1048.035 10566.5 1189.16 ;
      RECT 10562.865 1053.42 10566.5 1189.16 ;
      RECT 10553.5 1048.035 10555.115 1189.16 ;
      RECT 10553.5 1053.42 10566.5 1118.87 ;
      RECT 10553.5 1048.035 10561.85 1118.87 ;
      RECT 10553.5 1048.035 10566.5 1049.12 ;
      RECT 10536.52 1070.44 10549.52 1209.16 ;
      RECT 10536.865 1048.035 10549.52 1209.16 ;
      RECT 10536.52 1048.035 10549.52 1054.07 ;
      RECT 10506 1118.44 10534 1209.16 ;
      RECT 10518.375 1070.44 10534 1209.16 ;
      RECT 10506 1048.035 10510.625 1209.16 ;
      RECT 10506 1048.035 10531.955 1087.87 ;
      RECT 10506 1048.035 10534 1054.07 ;
      RECT 10490.48 1166.44 10503.48 1209.16 ;
      RECT 10500.475 1053.365 10503.48 1209.16 ;
      RECT 10490.48 1048.035 10495.565 1209.16 ;
      RECT 10490.48 1087.44 10503.48 1150.07 ;
      RECT 10490.48 1053.365 10503.48 1071.07 ;
      RECT 10490.48 1048.035 10498.81 1071.07 ;
      RECT 10490.48 1048.035 10503.48 1049.165 ;
      RECT 10473.5 1166.44 10486.5 1189.16 ;
      RECT 10478.145 1048.035 10486.5 1189.16 ;
      RECT 10477.98 1087.44 10486.5 1189.16 ;
      RECT 10473.5 1087.44 10486.5 1150.07 ;
      RECT 10473.5 1048.035 10486.5 1071.07 ;
      RECT 10456.52 1183.44 10469.52 1209.16 ;
      RECT 10456.52 1048.035 10468.565 1209.16 ;
      RECT 10456.52 1070.44 10469.52 1167.07 ;
      RECT 10456.52 1048.035 10469.52 1054.07 ;
      RECT 10426 1183.44 10454 1209.16 ;
      RECT 10452.145 1048.035 10454 1209.16 ;
      RECT 10426 1087.44 10447.235 1209.16 ;
      RECT 10449.555 1048.035 10454 1167.07 ;
      RECT 10432.55 1070.44 10454 1167.07 ;
      RECT 10426 1048.035 10444.645 1071.07 ;
      RECT 10426 1048.035 10454 1054.07 ;
      RECT 10410.48 1149.44 10423.48 1209.16 ;
      RECT 10422.865 1053.415 10423.48 1209.16 ;
      RECT 10410.48 1048.035 10415.115 1209.16 ;
      RECT 10410.48 1053.415 10423.48 1118.87 ;
      RECT 10410.48 1048.035 10421.85 1118.87 ;
      RECT 10410.48 1048.035 10423.48 1049.12 ;
      RECT 10393.5 1070.44 10406.5 1189.16 ;
      RECT 10396.865 1048.035 10406.5 1189.16 ;
      RECT 10393.5 1048.035 10406.5 1054.07 ;
      RECT 10376.52 1118.44 10389.52 1209.16 ;
      RECT 10378.375 1048.035 10389.52 1209.16 ;
      RECT 10376.52 1048.035 10389.52 1087.87 ;
      RECT 10346 1166.44 10374 1209.16 ;
      RECT 10360.475 1118.44 10374 1209.16 ;
      RECT 10346 1048.035 10355.565 1209.16 ;
      RECT 10346 1087.44 10370.625 1150.07 ;
      RECT 10364.53 1048.035 10374 1087.87 ;
      RECT 10360.475 1053.365 10374 1087.87 ;
      RECT 10346 1053.365 10374 1071.07 ;
      RECT 10346 1048.035 10358.81 1071.07 ;
      RECT 10346 1048.035 10374 1049.165 ;
      RECT 10330.48 1183.44 10343.48 1209.16 ;
      RECT 10338.145 1048.035 10343.48 1209.16 ;
      RECT 10333.475 1166.44 10343.48 1209.16 ;
      RECT 10330.48 1166.44 10343.48 1167.07 ;
      RECT 10330.48 1070.44 10333.235 1167.07 ;
      RECT 10330.48 1087.44 10343.48 1150.07 ;
      RECT 10330.48 1070.44 10343.48 1071.07 ;
      RECT 10333.475 1048.035 10343.48 1071.07 ;
      RECT 10330.48 1048.035 10343.48 1054.07 ;
      RECT 10296.52 1183.44 10309.52 1209.16 ;
      RECT 10296.52 1087.44 10307.235 1209.16 ;
      RECT 10301.75 1070.44 10309.52 1167.07 ;
      RECT 10296.52 1048.035 10304.565 1071.07 ;
      RECT 10296.52 1048.035 10309.52 1054.07 ;
      RECT 10266 1149.44 10294 1209.16 ;
      RECT 10284.63 1048.035 10294 1209.16 ;
      RECT 10282.865 1053.42 10294 1209.16 ;
      RECT 10266 1048.035 10275.115 1209.16 ;
      RECT 10266 1053.42 10294 1118.87 ;
      RECT 10266 1048.035 10281.85 1118.87 ;
      RECT 10266 1048.035 10294 1049.12 ;
      RECT 10250.48 1070.44 10263.48 1209.16 ;
      RECT 10256.865 1048.035 10263.48 1209.16 ;
      RECT 10250.48 1048.035 10251.955 1209.16 ;
      RECT 10250.48 1048.035 10263.48 1054.07 ;
      RECT 10233.5 1118.44 10246.5 1189.16 ;
      RECT 10238.375 1048.035 10246.5 1189.16 ;
      RECT 10233.5 1048.035 10246.5 1087.87 ;
      RECT 10216.52 1166.44 10229.52 1209.16 ;
      RECT 10224.53 1048.035 10229.52 1209.16 ;
      RECT 10220.475 1053.365 10229.52 1209.16 ;
      RECT 10216.52 1087.44 10229.52 1150.07 ;
      RECT 10216.52 1053.365 10229.52 1071.07 ;
      RECT 10216.52 1048.035 10218.81 1071.07 ;
      RECT 10216.52 1048.035 10229.52 1049.375 ;
      RECT 10186 1183.44 10214 1209.16 ;
      RECT 10198.145 1048.035 10214 1209.16 ;
      RECT 10193.475 1166.44 10214 1209.16 ;
      RECT 10186 1048.035 10188.565 1209.16 ;
      RECT 10186 1166.44 10214 1167.07 ;
      RECT 10186 1070.44 10193.235 1167.07 ;
      RECT 10186 1087.44 10214 1150.07 ;
      RECT 10186 1070.44 10214 1071.07 ;
      RECT 10193.475 1048.035 10214 1071.07 ;
      RECT 10186 1048.035 10214 1054.07 ;
      RECT 10170.48 1183.44 10183.48 1209.16 ;
      RECT 10172.145 1048.035 10183.48 1209.16 ;
      RECT 10170.48 1048.035 10183.48 1167.07 ;
      RECT 10153.5 1087.44 10166.5 1189.16 ;
      RECT 10160.13 1070.44 10166.5 1189.16 ;
      RECT 10153.5 1048.035 10163.455 1071.07 ;
      RECT 10153.5 1048.035 10166.5 1054.07 ;
      RECT 10136.52 1149.44 10149.52 1209.16 ;
      RECT 10144.63 1048.035 10149.52 1209.16 ;
      RECT 10142.865 1053.42 10149.52 1209.16 ;
      RECT 10136.52 1053.42 10149.52 1118.87 ;
      RECT 10136.52 1048.035 10141.85 1118.87 ;
      RECT 10136.52 1048.035 10149.52 1049.12 ;
      RECT 10106 1070.44 10134 1209.16 ;
      RECT 10116.865 1048.035 10134 1209.16 ;
      RECT 10106 1048.035 10111.955 1209.16 ;
      RECT 10106 1048.035 10134 1054.07 ;
      RECT 10090.48 1118.44 10103.48 1209.16 ;
      RECT 10098.375 1048.035 10103.48 1209.16 ;
      RECT 10090.48 1048.035 10103.48 1087.87 ;
      RECT 10073.5 1166.44 10086.5 1189.16 ;
      RECT 10084.43 1048.035 10086.5 1189.16 ;
      RECT 10080.475 1053.365 10086.5 1189.16 ;
      RECT 10073.5 1048.035 10075.565 1189.16 ;
      RECT 10073.5 1087.44 10086.5 1150.07 ;
      RECT 10073.5 1053.365 10086.5 1071.07 ;
      RECT 10073.5 1048.035 10078.81 1071.07 ;
      RECT 10073.5 1048.035 10086.5 1049.165 ;
      RECT 10056.52 1166.44 10069.52 1209.16 ;
      RECT 10058.145 1048.035 10069.52 1209.16 ;
      RECT 10056.52 1087.44 10069.52 1150.07 ;
      RECT 10056.52 1048.035 10069.52 1071.07 ;
      RECT 10026 1183.44 10054 1209.16 ;
      RECT 10032.145 1048.035 10048.565 1209.16 ;
      RECT 10026 1070.44 10027.235 1209.16 ;
      RECT 10026 1070.44 10053.235 1167.07 ;
      RECT 10026 1087.44 10054 1150.07 ;
      RECT 10028.365 1048.035 10048.565 1167.07 ;
      RECT 10026 1048.035 10054 1054.07 ;
      RECT 10010.48 1087.44 10023.48 1209.16 ;
      RECT 10010.48 1048.035 10016.835 1209.16 ;
      RECT 10010.48 1048.035 10023.48 1071.07 ;
      RECT 9993.5 1149.44 10006.5 1189.16 ;
      RECT 10004.63 1048.035 10006.5 1189.16 ;
      RECT 10002.865 1053.42 10006.5 1189.16 ;
      RECT 9993.5 1048.035 9995.115 1189.16 ;
      RECT 9993.5 1053.42 10006.5 1118.87 ;
      RECT 9993.5 1048.035 10001.85 1118.87 ;
      RECT 9993.5 1048.035 10006.5 1049.12 ;
      RECT 9976.52 1070.44 9989.52 1209.16 ;
      RECT 9976.865 1048.035 9989.52 1209.16 ;
      RECT 9976.52 1048.035 9989.52 1054.07 ;
      RECT 9946 1118.44 9974 1209.16 ;
      RECT 9958.375 1070.44 9974 1209.16 ;
      RECT 9946 1048.035 9950.625 1209.16 ;
      RECT 9946 1048.035 9971.955 1087.87 ;
      RECT 9946 1048.035 9974 1054.07 ;
      RECT 9930.48 1166.44 9943.48 1209.16 ;
      RECT 9940.475 1053.365 9943.48 1209.16 ;
      RECT 9930.48 1048.035 9935.565 1209.16 ;
      RECT 9930.48 1087.44 9943.48 1150.07 ;
      RECT 9930.48 1053.365 9943.48 1071.07 ;
      RECT 9930.48 1048.035 9938.81 1071.07 ;
      RECT 9930.48 1048.035 9943.48 1049.165 ;
      RECT 9913.5 1166.44 9926.5 1189.16 ;
      RECT 9918.145 1048.035 9926.5 1189.16 ;
      RECT 9917.98 1087.44 9926.5 1189.16 ;
      RECT 9913.5 1087.44 9926.5 1150.07 ;
      RECT 9913.5 1048.035 9926.5 1071.07 ;
      RECT 9896.52 1183.44 9909.52 1209.16 ;
      RECT 9896.52 1048.035 9908.565 1209.16 ;
      RECT 9896.52 1070.44 9909.52 1167.07 ;
      RECT 9896.52 1048.035 9909.52 1054.07 ;
      RECT 9866 1183.44 9894 1209.16 ;
      RECT 9892.145 1048.035 9894 1209.16 ;
      RECT 9866 1087.44 9887.235 1209.16 ;
      RECT 9889.555 1048.035 9894 1167.07 ;
      RECT 9872.55 1070.44 9894 1167.07 ;
      RECT 9866 1048.035 9884.645 1071.07 ;
      RECT 9866 1048.035 9894 1054.07 ;
      RECT 9850.48 1149.44 9863.48 1209.16 ;
      RECT 9862.865 1053.415 9863.48 1209.16 ;
      RECT 9850.48 1048.035 9855.115 1209.16 ;
      RECT 9850.48 1053.415 9863.48 1118.87 ;
      RECT 9850.48 1048.035 9861.85 1118.87 ;
      RECT 9850.48 1048.035 9863.48 1049.12 ;
      RECT 9833.5 1070.44 9846.5 1189.16 ;
      RECT 9836.865 1048.035 9846.5 1189.16 ;
      RECT 9833.5 1048.035 9846.5 1054.07 ;
      RECT 9816.52 1118.44 9829.52 1209.16 ;
      RECT 9818.375 1048.035 9829.52 1209.16 ;
      RECT 9816.52 1048.035 9829.52 1087.87 ;
      RECT 9786 1166.44 9814 1209.16 ;
      RECT 9800.475 1118.44 9814 1209.16 ;
      RECT 9786 1048.035 9795.565 1209.16 ;
      RECT 9786 1087.44 9810.625 1150.07 ;
      RECT 9804.53 1048.035 9814 1087.87 ;
      RECT 9800.475 1053.365 9814 1087.87 ;
      RECT 9786 1053.365 9814 1071.07 ;
      RECT 9786 1048.035 9798.81 1071.07 ;
      RECT 9786 1048.035 9814 1049.165 ;
      RECT 9770.48 1183.44 9783.48 1209.16 ;
      RECT 9778.145 1048.035 9783.48 1209.16 ;
      RECT 9773.475 1166.44 9783.48 1209.16 ;
      RECT 9770.48 1166.44 9783.48 1167.07 ;
      RECT 9770.48 1070.44 9773.235 1167.07 ;
      RECT 9770.48 1087.44 9783.48 1150.07 ;
      RECT 9770.48 1070.44 9783.48 1071.07 ;
      RECT 9773.475 1048.035 9783.48 1071.07 ;
      RECT 9770.48 1048.035 9783.48 1054.07 ;
      RECT 9736.52 1183.44 9749.52 1209.16 ;
      RECT 9736.52 1087.44 9747.235 1209.16 ;
      RECT 9741.75 1070.44 9749.52 1167.07 ;
      RECT 9736.52 1048.035 9744.565 1071.07 ;
      RECT 9736.52 1048.035 9749.52 1054.07 ;
      RECT 9706 1149.44 9734 1209.16 ;
      RECT 9724.63 1048.035 9734 1209.16 ;
      RECT 9722.865 1053.42 9734 1209.16 ;
      RECT 9706 1048.035 9715.115 1209.16 ;
      RECT 9706 1053.42 9734 1118.87 ;
      RECT 9706 1048.035 9721.85 1118.87 ;
      RECT 9706 1048.035 9734 1049.12 ;
      RECT 9690.48 1070.44 9703.48 1209.16 ;
      RECT 9696.865 1048.035 9703.48 1209.16 ;
      RECT 9690.48 1048.035 9691.955 1209.16 ;
      RECT 9690.48 1048.035 9703.48 1054.07 ;
      RECT 9673.5 1118.44 9686.5 1189.16 ;
      RECT 9678.375 1048.035 9686.5 1189.16 ;
      RECT 9673.5 1048.035 9686.5 1087.87 ;
      RECT 9656.52 1166.44 9669.52 1209.16 ;
      RECT 9664.53 1048.035 9669.52 1209.16 ;
      RECT 9660.475 1053.365 9669.52 1209.16 ;
      RECT 9656.52 1087.44 9669.52 1150.07 ;
      RECT 9656.52 1053.365 9669.52 1071.07 ;
      RECT 9656.52 1048.035 9658.81 1071.07 ;
      RECT 9656.52 1048.035 9669.52 1049.375 ;
      RECT 9626 1183.44 9654 1209.16 ;
      RECT 9638.145 1048.035 9654 1209.16 ;
      RECT 9633.475 1166.44 9654 1209.16 ;
      RECT 9626 1048.035 9628.565 1209.16 ;
      RECT 9626 1166.44 9654 1167.07 ;
      RECT 9626 1070.44 9633.235 1167.07 ;
      RECT 9626 1087.44 9654 1150.07 ;
      RECT 9626 1070.44 9654 1071.07 ;
      RECT 9633.475 1048.035 9654 1071.07 ;
      RECT 9626 1048.035 9654 1054.07 ;
      RECT 9610.48 1183.44 9623.48 1209.16 ;
      RECT 9612.145 1048.035 9623.48 1209.16 ;
      RECT 9610.48 1048.035 9623.48 1167.07 ;
      RECT 9593.5 1087.44 9606.5 1189.16 ;
      RECT 9600.13 1070.44 9606.5 1189.16 ;
      RECT 9593.5 1048.035 9603.455 1071.07 ;
      RECT 9593.5 1048.035 9606.5 1054.07 ;
      RECT 9576.52 1149.44 9589.52 1209.16 ;
      RECT 9584.63 1048.035 9589.52 1209.16 ;
      RECT 9582.865 1053.42 9589.52 1209.16 ;
      RECT 9576.52 1053.42 9589.52 1118.87 ;
      RECT 9576.52 1048.035 9581.85 1118.87 ;
      RECT 9576.52 1048.035 9589.52 1049.12 ;
      RECT 9546 1070.44 9574 1209.16 ;
      RECT 9556.865 1048.035 9574 1209.16 ;
      RECT 9546 1048.035 9551.955 1209.16 ;
      RECT 9546 1048.035 9574 1054.07 ;
      RECT 9530.48 1118.44 9543.48 1209.16 ;
      RECT 9538.375 1048.035 9543.48 1209.16 ;
      RECT 9530.48 1048.035 9543.48 1087.87 ;
      RECT 9513.5 1166.44 9526.5 1189.16 ;
      RECT 9524.43 1048.035 9526.5 1189.16 ;
      RECT 9520.475 1053.365 9526.5 1189.16 ;
      RECT 9513.5 1048.035 9515.565 1189.16 ;
      RECT 9513.5 1087.44 9526.5 1150.07 ;
      RECT 9513.5 1053.365 9526.5 1071.07 ;
      RECT 9513.5 1048.035 9518.81 1071.07 ;
      RECT 9513.5 1048.035 9526.5 1049.165 ;
      RECT 9496.52 1166.44 9509.52 1209.16 ;
      RECT 9498.145 1048.035 9509.52 1209.16 ;
      RECT 9496.52 1087.44 9509.52 1150.07 ;
      RECT 9496.52 1048.035 9509.52 1071.07 ;
      RECT 9466 1183.44 9494 1209.16 ;
      RECT 9472.145 1048.035 9488.565 1209.16 ;
      RECT 9466 1070.44 9467.235 1209.16 ;
      RECT 9466 1070.44 9493.235 1167.07 ;
      RECT 9466 1087.44 9494 1150.07 ;
      RECT 9468.365 1048.035 9488.565 1167.07 ;
      RECT 9466 1048.035 9494 1054.07 ;
      RECT 9450.48 1087.44 9463.48 1209.16 ;
      RECT 9450.48 1048.035 9456.835 1209.16 ;
      RECT 9450.48 1048.035 9463.48 1071.07 ;
      RECT 9433.5 1149.44 9446.5 1189.16 ;
      RECT 9444.63 1048.035 9446.5 1189.16 ;
      RECT 9442.865 1053.42 9446.5 1189.16 ;
      RECT 9433.5 1048.035 9435.115 1189.16 ;
      RECT 9433.5 1053.42 9446.5 1118.87 ;
      RECT 9433.5 1048.035 9441.85 1118.87 ;
      RECT 9433.5 1048.035 9446.5 1049.12 ;
      RECT 9416.52 1070.44 9429.52 1209.16 ;
      RECT 9416.865 1048.035 9429.52 1209.16 ;
      RECT 9416.52 1048.035 9429.52 1054.07 ;
      RECT 9386 1118.44 9414 1209.16 ;
      RECT 9398.375 1070.44 9414 1209.16 ;
      RECT 9386 1048.035 9390.625 1209.16 ;
      RECT 9386 1048.035 9411.955 1087.87 ;
      RECT 9386 1048.035 9414 1054.07 ;
      RECT 9370.48 1166.44 9383.48 1209.16 ;
      RECT 9380.475 1053.365 9383.48 1209.16 ;
      RECT 9370.48 1048.035 9375.565 1209.16 ;
      RECT 9370.48 1087.44 9383.48 1150.07 ;
      RECT 9370.48 1053.365 9383.48 1071.07 ;
      RECT 9370.48 1048.035 9378.81 1071.07 ;
      RECT 9370.48 1048.035 9383.48 1049.165 ;
      RECT 9353.5 1166.44 9366.5 1189.16 ;
      RECT 9358.145 1048.035 9366.5 1189.16 ;
      RECT 9357.98 1087.44 9366.5 1189.16 ;
      RECT 9353.5 1087.44 9366.5 1150.07 ;
      RECT 9353.5 1048.035 9366.5 1071.07 ;
      RECT 9336.52 1183.44 9349.52 1209.16 ;
      RECT 9336.52 1048.035 9348.565 1209.16 ;
      RECT 9336.52 1070.44 9349.52 1167.07 ;
      RECT 9336.52 1048.035 9349.52 1054.07 ;
      RECT 9306 1183.44 9334 1209.16 ;
      RECT 9332.145 1048.035 9334 1209.16 ;
      RECT 9306 1087.44 9327.235 1209.16 ;
      RECT 9329.555 1048.035 9334 1167.07 ;
      RECT 9312.55 1070.44 9334 1167.07 ;
      RECT 9306 1048.035 9324.645 1071.07 ;
      RECT 9306 1048.035 9334 1054.07 ;
      RECT 9290.48 1149.44 9303.48 1209.16 ;
      RECT 9302.865 1053.415 9303.48 1209.16 ;
      RECT 9290.48 1048.035 9295.115 1209.16 ;
      RECT 9290.48 1053.415 9303.48 1118.87 ;
      RECT 9290.48 1048.035 9301.85 1118.87 ;
      RECT 9290.48 1048.035 9303.48 1049.12 ;
      RECT 9273.5 1070.44 9286.5 1189.16 ;
      RECT 9276.865 1048.035 9286.5 1189.16 ;
      RECT 9273.5 1048.035 9286.5 1054.07 ;
      RECT 9256.52 1118.44 9269.52 1209.16 ;
      RECT 9258.375 1048.035 9269.52 1209.16 ;
      RECT 9256.52 1048.035 9269.52 1087.87 ;
      RECT 9226 1166.44 9254 1209.16 ;
      RECT 9240.475 1118.44 9254 1209.16 ;
      RECT 9226 1048.035 9235.565 1209.16 ;
      RECT 9226 1087.44 9250.625 1150.07 ;
      RECT 9244.53 1048.035 9254 1087.87 ;
      RECT 9240.475 1053.365 9254 1087.87 ;
      RECT 9226 1053.365 9254 1071.07 ;
      RECT 9226 1048.035 9238.81 1071.07 ;
      RECT 9226 1048.035 9254 1049.165 ;
      RECT 9210.48 1183.44 9223.48 1209.16 ;
      RECT 9218.145 1048.035 9223.48 1209.16 ;
      RECT 9213.475 1166.44 9223.48 1209.16 ;
      RECT 9210.48 1166.44 9223.48 1167.07 ;
      RECT 9210.48 1070.44 9213.235 1167.07 ;
      RECT 9210.48 1087.44 9223.48 1150.07 ;
      RECT 9210.48 1070.44 9223.48 1071.07 ;
      RECT 9213.475 1048.035 9223.48 1071.07 ;
      RECT 9210.48 1048.035 9223.48 1054.07 ;
      RECT 9176.52 1183.44 9189.52 1209.16 ;
      RECT 9176.52 1087.44 9187.235 1209.16 ;
      RECT 9181.75 1070.44 9189.52 1167.07 ;
      RECT 9176.52 1048.035 9184.565 1071.07 ;
      RECT 9176.52 1048.035 9189.52 1054.07 ;
      RECT 9146 1149.44 9174 1209.16 ;
      RECT 9164.63 1048.035 9174 1209.16 ;
      RECT 9162.865 1053.42 9174 1209.16 ;
      RECT 9146 1048.035 9155.115 1209.16 ;
      RECT 9146 1053.42 9174 1118.87 ;
      RECT 9146 1048.035 9161.85 1118.87 ;
      RECT 9146 1048.035 9174 1049.12 ;
      RECT 9130.48 1070.44 9143.48 1209.16 ;
      RECT 9136.865 1048.035 9143.48 1209.16 ;
      RECT 9130.48 1048.035 9131.955 1209.16 ;
      RECT 9130.48 1048.035 9143.48 1054.07 ;
      RECT 9113.5 1118.44 9126.5 1189.16 ;
      RECT 9118.375 1048.035 9126.5 1189.16 ;
      RECT 9113.5 1048.035 9126.5 1087.87 ;
      RECT 9096.52 1166.44 9109.52 1209.16 ;
      RECT 9104.53 1048.035 9109.52 1209.16 ;
      RECT 9100.475 1053.365 9109.52 1209.16 ;
      RECT 9096.52 1087.44 9109.52 1150.07 ;
      RECT 9096.52 1053.365 9109.52 1071.07 ;
      RECT 9096.52 1048.035 9098.81 1071.07 ;
      RECT 9096.52 1048.035 9109.52 1049.375 ;
      RECT 9066 1183.44 9094 1209.16 ;
      RECT 9078.145 1048.035 9094 1209.16 ;
      RECT 9073.475 1166.44 9094 1209.16 ;
      RECT 9066 1048.035 9068.565 1209.16 ;
      RECT 9066 1166.44 9094 1167.07 ;
      RECT 9066 1070.44 9073.235 1167.07 ;
      RECT 9066 1087.44 9094 1150.07 ;
      RECT 9066 1070.44 9094 1071.07 ;
      RECT 9073.475 1048.035 9094 1071.07 ;
      RECT 9066 1048.035 9094 1054.07 ;
      RECT 9050.48 1183.44 9063.48 1209.16 ;
      RECT 9052.145 1048.035 9063.48 1209.16 ;
      RECT 9050.48 1048.035 9063.48 1167.07 ;
      RECT 9033.5 1087.44 9046.5 1189.16 ;
      RECT 9040.13 1070.44 9046.5 1189.16 ;
      RECT 9033.5 1048.035 9043.455 1071.07 ;
      RECT 9033.5 1048.035 9046.5 1054.07 ;
      RECT 9016.52 1149.44 9029.52 1209.16 ;
      RECT 9024.63 1048.035 9029.52 1209.16 ;
      RECT 9022.865 1053.42 9029.52 1209.16 ;
      RECT 9016.52 1053.42 9029.52 1118.87 ;
      RECT 9016.52 1048.035 9021.85 1118.87 ;
      RECT 9016.52 1048.035 9029.52 1049.12 ;
      RECT 8986 1070.44 9014 1209.16 ;
      RECT 8996.865 1048.035 9014 1209.16 ;
      RECT 8986 1048.035 8991.955 1209.16 ;
      RECT 8986 1048.035 9014 1054.07 ;
      RECT 8970.48 1118.44 8983.48 1209.16 ;
      RECT 8978.375 1048.035 8983.48 1209.16 ;
      RECT 8970.48 1048.035 8983.48 1087.87 ;
      RECT 8953.5 1166.44 8966.5 1189.16 ;
      RECT 8964.43 1048.035 8966.5 1189.16 ;
      RECT 8960.475 1053.365 8966.5 1189.16 ;
      RECT 8953.5 1048.035 8955.565 1189.16 ;
      RECT 8953.5 1087.44 8966.5 1150.07 ;
      RECT 8953.5 1053.365 8966.5 1071.07 ;
      RECT 8953.5 1048.035 8958.81 1071.07 ;
      RECT 8953.5 1048.035 8966.5 1049.165 ;
      RECT 8936.52 1166.44 8949.52 1209.16 ;
      RECT 8938.145 1048.035 8949.52 1209.16 ;
      RECT 8936.52 1087.44 8949.52 1150.07 ;
      RECT 8936.52 1048.035 8949.52 1071.07 ;
      RECT 8906 1183.44 8934 1209.16 ;
      RECT 8912.145 1048.035 8928.565 1209.16 ;
      RECT 8906 1070.44 8907.235 1209.16 ;
      RECT 8906 1070.44 8933.235 1167.07 ;
      RECT 8906 1087.44 8934 1150.07 ;
      RECT 8908.365 1048.035 8928.565 1167.07 ;
      RECT 8906 1048.035 8934 1054.07 ;
      RECT 8890.48 1087.44 8903.48 1209.16 ;
      RECT 8890.48 1048.035 8896.835 1209.16 ;
      RECT 8890.48 1048.035 8903.48 1071.07 ;
      RECT 8873.5 1149.44 8886.5 1189.16 ;
      RECT 8884.63 1048.035 8886.5 1189.16 ;
      RECT 8882.865 1053.42 8886.5 1189.16 ;
      RECT 8873.5 1048.035 8875.115 1189.16 ;
      RECT 8873.5 1053.42 8886.5 1118.87 ;
      RECT 8873.5 1048.035 8881.85 1118.87 ;
      RECT 8873.5 1048.035 8886.5 1049.12 ;
      RECT 8856.52 1070.44 8869.52 1209.16 ;
      RECT 8856.865 1048.035 8869.52 1209.16 ;
      RECT 8856.52 1048.035 8869.52 1054.07 ;
      RECT 8826 1118.44 8854 1209.16 ;
      RECT 8838.375 1070.44 8854 1209.16 ;
      RECT 8826 1048.035 8830.625 1209.16 ;
      RECT 8826 1048.035 8851.955 1087.87 ;
      RECT 8826 1048.035 8854 1054.07 ;
      RECT 8810.48 1166.44 8823.48 1209.16 ;
      RECT 8820.475 1053.365 8823.48 1209.16 ;
      RECT 8810.48 1048.035 8815.565 1209.16 ;
      RECT 8810.48 1087.44 8823.48 1150.07 ;
      RECT 8810.48 1053.365 8823.48 1071.07 ;
      RECT 8810.48 1048.035 8818.81 1071.07 ;
      RECT 8810.48 1048.035 8823.48 1049.165 ;
      RECT 8793.5 1166.44 8806.5 1189.16 ;
      RECT 8798.145 1048.035 8806.5 1189.16 ;
      RECT 8797.98 1087.44 8806.5 1189.16 ;
      RECT 8793.5 1087.44 8806.5 1150.07 ;
      RECT 8793.5 1048.035 8806.5 1071.07 ;
      RECT 8776.52 1183.44 8789.52 1209.16 ;
      RECT 8776.52 1048.035 8788.565 1209.16 ;
      RECT 8776.52 1070.44 8789.52 1167.07 ;
      RECT 8776.52 1048.035 8789.52 1054.07 ;
      RECT 8746 1183.44 8774 1209.16 ;
      RECT 8772.145 1048.035 8774 1209.16 ;
      RECT 8746 1087.44 8767.235 1209.16 ;
      RECT 8769.555 1048.035 8774 1167.07 ;
      RECT 8752.55 1070.44 8774 1167.07 ;
      RECT 8746 1048.035 8764.645 1071.07 ;
      RECT 8746 1048.035 8774 1054.07 ;
      RECT 8730.48 1149.44 8743.48 1209.16 ;
      RECT 8742.865 1053.415 8743.48 1209.16 ;
      RECT 8730.48 1048.035 8735.115 1209.16 ;
      RECT 8730.48 1053.415 8743.48 1118.87 ;
      RECT 8730.48 1048.035 8741.85 1118.87 ;
      RECT 8730.48 1048.035 8743.48 1049.12 ;
      RECT 8713.5 1070.44 8726.5 1189.16 ;
      RECT 8716.865 1048.035 8726.5 1189.16 ;
      RECT 8713.5 1048.035 8726.5 1054.07 ;
      RECT 8696.52 1118.44 8709.52 1209.16 ;
      RECT 8698.375 1048.035 8709.52 1209.16 ;
      RECT 8696.52 1048.035 8709.52 1087.87 ;
      RECT 8666 1166.44 8694 1209.16 ;
      RECT 8680.475 1118.44 8694 1209.16 ;
      RECT 8666 1048.035 8675.565 1209.16 ;
      RECT 8666 1087.44 8690.625 1150.07 ;
      RECT 8684.53 1048.035 8694 1087.87 ;
      RECT 8680.475 1053.365 8694 1087.87 ;
      RECT 8666 1053.365 8694 1071.07 ;
      RECT 8666 1048.035 8678.81 1071.07 ;
      RECT 8666 1048.035 8694 1049.165 ;
      RECT 8650.48 1183.44 8663.48 1209.16 ;
      RECT 8658.145 1048.035 8663.48 1209.16 ;
      RECT 8653.475 1166.44 8663.48 1209.16 ;
      RECT 8650.48 1166.44 8663.48 1167.07 ;
      RECT 8650.48 1070.44 8653.235 1167.07 ;
      RECT 8650.48 1087.44 8663.48 1150.07 ;
      RECT 8650.48 1070.44 8663.48 1071.07 ;
      RECT 8653.475 1048.035 8663.48 1071.07 ;
      RECT 8650.48 1048.035 8663.48 1054.07 ;
      RECT 8616.52 1183.44 8629.52 1209.16 ;
      RECT 8616.52 1087.44 8627.235 1209.16 ;
      RECT 8621.75 1070.44 8629.52 1167.07 ;
      RECT 8616.52 1048.035 8624.565 1071.07 ;
      RECT 8616.52 1048.035 8629.52 1054.07 ;
      RECT 8586 1149.44 8614 1209.16 ;
      RECT 8604.63 1048.035 8614 1209.16 ;
      RECT 8602.865 1053.42 8614 1209.16 ;
      RECT 8586 1048.035 8595.115 1209.16 ;
      RECT 8586 1053.42 8614 1118.87 ;
      RECT 8586 1048.035 8601.85 1118.87 ;
      RECT 8586 1048.035 8614 1049.12 ;
      RECT 8570.48 1070.44 8583.48 1209.16 ;
      RECT 8576.865 1048.035 8583.48 1209.16 ;
      RECT 8570.48 1048.035 8571.955 1209.16 ;
      RECT 8570.48 1048.035 8583.48 1054.07 ;
      RECT 8553.5 1118.44 8566.5 1189.16 ;
      RECT 8558.375 1048.035 8566.5 1189.16 ;
      RECT 8553.5 1048.035 8566.5 1087.87 ;
      RECT 8536.52 1166.44 8549.52 1209.16 ;
      RECT 8544.53 1048.035 8549.52 1209.16 ;
      RECT 8540.475 1053.365 8549.52 1209.16 ;
      RECT 8536.52 1087.44 8549.52 1150.07 ;
      RECT 8536.52 1053.365 8549.52 1071.07 ;
      RECT 8536.52 1048.035 8538.81 1071.07 ;
      RECT 8536.52 1048.035 8549.52 1049.375 ;
      RECT 8506 1183.44 8534 1209.16 ;
      RECT 8518.145 1048.035 8534 1209.16 ;
      RECT 8513.475 1166.44 8534 1209.16 ;
      RECT 8506 1048.035 8508.565 1209.16 ;
      RECT 8506 1166.44 8534 1167.07 ;
      RECT 8506 1070.44 8513.235 1167.07 ;
      RECT 8506 1087.44 8534 1150.07 ;
      RECT 8506 1070.44 8534 1071.07 ;
      RECT 8513.475 1048.035 8534 1071.07 ;
      RECT 8506 1048.035 8534 1054.07 ;
      RECT 8490.48 1183.44 8503.48 1209.16 ;
      RECT 8492.145 1048.035 8503.48 1209.16 ;
      RECT 8490.48 1048.035 8503.48 1167.07 ;
      RECT 8473.5 1087.44 8486.5 1189.16 ;
      RECT 8480.13 1070.44 8486.5 1189.16 ;
      RECT 8473.5 1048.035 8483.455 1071.07 ;
      RECT 8473.5 1048.035 8486.5 1054.07 ;
      RECT 8456.52 1149.44 8469.52 1209.16 ;
      RECT 8464.63 1048.035 8469.52 1209.16 ;
      RECT 8462.865 1053.42 8469.52 1209.16 ;
      RECT 8456.52 1053.42 8469.52 1118.87 ;
      RECT 8456.52 1048.035 8461.85 1118.87 ;
      RECT 8456.52 1048.035 8469.52 1049.12 ;
      RECT 8426 1070.44 8454 1209.16 ;
      RECT 8436.865 1048.035 8454 1209.16 ;
      RECT 8426 1048.035 8431.955 1209.16 ;
      RECT 8426 1048.035 8454 1054.07 ;
      RECT 8410.48 1118.44 8423.48 1209.16 ;
      RECT 8418.375 1048.035 8423.48 1209.16 ;
      RECT 8410.48 1048.035 8423.48 1087.87 ;
      RECT 8393.5 1166.44 8406.5 1189.16 ;
      RECT 8404.43 1048.035 8406.5 1189.16 ;
      RECT 8400.475 1053.365 8406.5 1189.16 ;
      RECT 8393.5 1048.035 8395.565 1189.16 ;
      RECT 8393.5 1087.44 8406.5 1150.07 ;
      RECT 8393.5 1053.365 8406.5 1071.07 ;
      RECT 8393.5 1048.035 8398.81 1071.07 ;
      RECT 8393.5 1048.035 8406.5 1049.165 ;
      RECT 8376.52 1166.44 8389.52 1209.16 ;
      RECT 8378.145 1048.035 8389.52 1209.16 ;
      RECT 8376.52 1087.44 8389.52 1150.07 ;
      RECT 8376.52 1048.035 8389.52 1071.07 ;
      RECT 8346 1183.44 8374 1209.16 ;
      RECT 8352.145 1048.035 8368.565 1209.16 ;
      RECT 8346 1070.44 8347.235 1209.16 ;
      RECT 8346 1070.44 8373.235 1167.07 ;
      RECT 8346 1087.44 8374 1150.07 ;
      RECT 8348.365 1048.035 8368.565 1167.07 ;
      RECT 8346 1048.035 8374 1054.07 ;
      RECT 8330.48 1087.44 8343.48 1209.16 ;
      RECT 8330.48 1048.035 8336.835 1209.16 ;
      RECT 8330.48 1048.035 8343.48 1071.07 ;
      RECT 8313.5 1149.44 8326.5 1189.16 ;
      RECT 8324.63 1048.035 8326.5 1189.16 ;
      RECT 8322.865 1053.42 8326.5 1189.16 ;
      RECT 8313.5 1048.035 8315.115 1189.16 ;
      RECT 8313.5 1053.42 8326.5 1118.87 ;
      RECT 8313.5 1048.035 8321.85 1118.87 ;
      RECT 8313.5 1048.035 8326.5 1049.12 ;
      RECT 8296.52 1070.44 8309.52 1209.16 ;
      RECT 8296.865 1048.035 8309.52 1209.16 ;
      RECT 8296.52 1048.035 8309.52 1054.07 ;
      RECT 8266 1118.44 8294 1209.16 ;
      RECT 8278.375 1070.44 8294 1209.16 ;
      RECT 8266 1048.035 8270.625 1209.16 ;
      RECT 8266 1048.035 8291.955 1087.87 ;
      RECT 8266 1048.035 8294 1054.07 ;
      RECT 8250.48 1166.44 8263.48 1209.16 ;
      RECT 8260.475 1053.365 8263.48 1209.16 ;
      RECT 8250.48 1048.035 8255.565 1209.16 ;
      RECT 8250.48 1087.44 8263.48 1150.07 ;
      RECT 8250.48 1053.365 8263.48 1071.07 ;
      RECT 8250.48 1048.035 8258.81 1071.07 ;
      RECT 8250.48 1048.035 8263.48 1049.165 ;
      RECT 8233.5 1166.44 8246.5 1189.16 ;
      RECT 8238.145 1048.035 8246.5 1189.16 ;
      RECT 8237.98 1087.44 8246.5 1189.16 ;
      RECT 8233.5 1087.44 8246.5 1150.07 ;
      RECT 8233.5 1048.035 8246.5 1071.07 ;
      RECT 8216.52 1183.44 8229.52 1209.16 ;
      RECT 8216.52 1048.035 8228.565 1209.16 ;
      RECT 8216.52 1070.44 8229.52 1167.07 ;
      RECT 8216.52 1048.035 8229.52 1054.07 ;
      RECT 8186 1183.44 8214 1209.16 ;
      RECT 8212.145 1048.035 8214 1209.16 ;
      RECT 8186 1087.44 8207.235 1209.16 ;
      RECT 8209.555 1048.035 8214 1167.07 ;
      RECT 8192.55 1070.44 8214 1167.07 ;
      RECT 8186 1048.035 8204.645 1071.07 ;
      RECT 8186 1048.035 8214 1054.07 ;
      RECT 8170.48 1149.44 8183.48 1209.16 ;
      RECT 8182.865 1053.415 8183.48 1209.16 ;
      RECT 8170.48 1048.035 8175.115 1209.16 ;
      RECT 8170.48 1053.415 8183.48 1118.87 ;
      RECT 8170.48 1048.035 8181.85 1118.87 ;
      RECT 8170.48 1048.035 8183.48 1049.12 ;
      RECT 8153.5 1070.44 8166.5 1189.16 ;
      RECT 8156.865 1048.035 8166.5 1189.16 ;
      RECT 8153.5 1048.035 8166.5 1054.07 ;
      RECT 8136.52 1118.44 8149.52 1209.16 ;
      RECT 8138.375 1048.035 8149.52 1209.16 ;
      RECT 8136.52 1048.035 8149.52 1087.87 ;
      RECT 8106 1166.44 8134 1209.16 ;
      RECT 8120.475 1118.44 8134 1209.16 ;
      RECT 8106 1048.035 8115.565 1209.16 ;
      RECT 8106 1087.44 8130.625 1150.07 ;
      RECT 8124.53 1048.035 8134 1087.87 ;
      RECT 8120.475 1053.365 8134 1087.87 ;
      RECT 8106 1053.365 8134 1071.07 ;
      RECT 8106 1048.035 8118.81 1071.07 ;
      RECT 8106 1048.035 8134 1049.165 ;
      RECT 8090.48 1183.44 8103.48 1209.16 ;
      RECT 8098.145 1048.035 8103.48 1209.16 ;
      RECT 8093.475 1166.44 8103.48 1209.16 ;
      RECT 8090.48 1166.44 8103.48 1167.07 ;
      RECT 8090.48 1070.44 8093.235 1167.07 ;
      RECT 8090.48 1087.44 8103.48 1150.07 ;
      RECT 8090.48 1070.44 8103.48 1071.07 ;
      RECT 8093.475 1048.035 8103.48 1071.07 ;
      RECT 8090.48 1048.035 8103.48 1054.07 ;
      RECT 8056.52 1183.44 8069.52 1209.16 ;
      RECT 8056.52 1087.44 8067.235 1209.16 ;
      RECT 8061.75 1070.44 8069.52 1167.07 ;
      RECT 8056.52 1048.035 8064.565 1071.07 ;
      RECT 8056.52 1048.035 8069.52 1054.07 ;
      RECT 8026 1149.44 8054 1209.16 ;
      RECT 8044.63 1048.035 8054 1209.16 ;
      RECT 8042.865 1053.42 8054 1209.16 ;
      RECT 8026 1048.035 8035.115 1209.16 ;
      RECT 8026 1053.42 8054 1118.87 ;
      RECT 8026 1048.035 8041.85 1118.87 ;
      RECT 8026 1048.035 8054 1049.12 ;
      RECT 8010.48 1070.44 8023.48 1209.16 ;
      RECT 8016.865 1048.035 8023.48 1209.16 ;
      RECT 8010.48 1048.035 8011.955 1209.16 ;
      RECT 8010.48 1048.035 8023.48 1054.07 ;
      RECT 7993.5 1118.44 8006.5 1189.16 ;
      RECT 7998.375 1048.035 8006.5 1189.16 ;
      RECT 7993.5 1048.035 8006.5 1087.87 ;
      RECT 7976.52 1166.44 7989.52 1209.16 ;
      RECT 7984.53 1048.035 7989.52 1209.16 ;
      RECT 7980.475 1053.365 7989.52 1209.16 ;
      RECT 7976.52 1087.44 7989.52 1150.07 ;
      RECT 7976.52 1053.365 7989.52 1071.07 ;
      RECT 7976.52 1048.035 7978.81 1071.07 ;
      RECT 7976.52 1048.035 7989.52 1049.375 ;
      RECT 7946 1183.44 7974 1209.16 ;
      RECT 7958.145 1048.035 7974 1209.16 ;
      RECT 7953.475 1166.44 7974 1209.16 ;
      RECT 7946 1048.035 7948.565 1209.16 ;
      RECT 7946 1166.44 7974 1167.07 ;
      RECT 7946 1070.44 7953.235 1167.07 ;
      RECT 7946 1087.44 7974 1150.07 ;
      RECT 7946 1070.44 7974 1071.07 ;
      RECT 7953.475 1048.035 7974 1071.07 ;
      RECT 7946 1048.035 7974 1054.07 ;
      RECT 7930.48 1183.44 7943.48 1209.16 ;
      RECT 7932.145 1048.035 7943.48 1209.16 ;
      RECT 7930.48 1048.035 7943.48 1167.07 ;
      RECT 7913.5 1087.44 7926.5 1189.16 ;
      RECT 7920.13 1070.44 7926.5 1189.16 ;
      RECT 7913.5 1048.035 7923.455 1071.07 ;
      RECT 7913.5 1048.035 7926.5 1054.07 ;
      RECT 7896.52 1149.44 7909.52 1209.16 ;
      RECT 7904.63 1048.035 7909.52 1209.16 ;
      RECT 7902.865 1053.42 7909.52 1209.16 ;
      RECT 7896.52 1053.42 7909.52 1118.87 ;
      RECT 7896.52 1048.035 7901.85 1118.87 ;
      RECT 7896.52 1048.035 7909.52 1049.12 ;
      RECT 7866 1070.44 7894 1209.16 ;
      RECT 7876.865 1048.035 7894 1209.16 ;
      RECT 7866 1048.035 7871.955 1209.16 ;
      RECT 7866 1048.035 7894 1054.07 ;
      RECT 7850.48 1118.44 7863.48 1209.16 ;
      RECT 7858.375 1048.035 7863.48 1209.16 ;
      RECT 7850.48 1048.035 7863.48 1087.87 ;
      RECT 7833.5 1166.44 7846.5 1189.16 ;
      RECT 7844.43 1048.035 7846.5 1189.16 ;
      RECT 7840.475 1053.365 7846.5 1189.16 ;
      RECT 7833.5 1048.035 7835.565 1189.16 ;
      RECT 7833.5 1087.44 7846.5 1150.07 ;
      RECT 7833.5 1053.365 7846.5 1071.07 ;
      RECT 7833.5 1048.035 7838.81 1071.07 ;
      RECT 7833.5 1048.035 7846.5 1049.165 ;
      RECT 7816.52 1166.44 7829.52 1209.16 ;
      RECT 7818.145 1048.035 7829.52 1209.16 ;
      RECT 7816.52 1087.44 7829.52 1150.07 ;
      RECT 7816.52 1048.035 7829.52 1071.07 ;
      RECT 7786 1183.44 7814 1209.16 ;
      RECT 7792.145 1048.035 7808.565 1209.16 ;
      RECT 7786 1070.44 7787.235 1209.16 ;
      RECT 7786 1070.44 7813.235 1167.07 ;
      RECT 7786 1087.44 7814 1150.07 ;
      RECT 7788.365 1048.035 7808.565 1167.07 ;
      RECT 7786 1048.035 7814 1054.07 ;
      RECT 7770.48 1087.44 7783.48 1209.16 ;
      RECT 7770.48 1048.035 7776.835 1209.16 ;
      RECT 7770.48 1048.035 7783.48 1071.07 ;
      RECT 7753.5 1149.44 7766.5 1189.16 ;
      RECT 7764.63 1048.035 7766.5 1189.16 ;
      RECT 7762.865 1053.42 7766.5 1189.16 ;
      RECT 7753.5 1048.035 7755.115 1189.16 ;
      RECT 7753.5 1053.42 7766.5 1118.87 ;
      RECT 7753.5 1048.035 7761.85 1118.87 ;
      RECT 7753.5 1048.035 7766.5 1049.12 ;
      RECT 7736.52 1070.44 7749.52 1209.16 ;
      RECT 7736.865 1048.035 7749.52 1209.16 ;
      RECT 7736.52 1048.035 7749.52 1054.07 ;
      RECT 7706 1118.44 7734 1209.16 ;
      RECT 7718.375 1070.44 7734 1209.16 ;
      RECT 7706 1048.035 7710.625 1209.16 ;
      RECT 7706 1048.035 7731.955 1087.87 ;
      RECT 7706 1048.035 7734 1054.07 ;
      RECT 7690.48 1166.44 7703.48 1209.16 ;
      RECT 7700.475 1053.365 7703.48 1209.16 ;
      RECT 7690.48 1048.035 7695.565 1209.16 ;
      RECT 7690.48 1087.44 7703.48 1150.07 ;
      RECT 7690.48 1053.365 7703.48 1071.07 ;
      RECT 7690.48 1048.035 7698.81 1071.07 ;
      RECT 7690.48 1048.035 7703.48 1049.165 ;
      RECT 7673.5 1166.44 7686.5 1189.16 ;
      RECT 7678.145 1048.035 7686.5 1189.16 ;
      RECT 7677.98 1087.44 7686.5 1189.16 ;
      RECT 7673.5 1087.44 7686.5 1150.07 ;
      RECT 7673.5 1048.035 7686.5 1071.07 ;
      RECT 7656.52 1183.44 7669.52 1209.16 ;
      RECT 7656.52 1048.035 7668.565 1209.16 ;
      RECT 7656.52 1070.44 7669.52 1167.07 ;
      RECT 7656.52 1048.035 7669.52 1054.07 ;
      RECT 7626 1183.44 7654 1209.16 ;
      RECT 7652.145 1048.035 7654 1209.16 ;
      RECT 7626 1087.44 7647.235 1209.16 ;
      RECT 7649.555 1048.035 7654 1167.07 ;
      RECT 7632.55 1070.44 7654 1167.07 ;
      RECT 7626 1048.035 7644.645 1071.07 ;
      RECT 7626 1048.035 7654 1054.07 ;
      RECT 7610.48 1149.44 7623.48 1209.16 ;
      RECT 7622.865 1053.415 7623.48 1209.16 ;
      RECT 7610.48 1048.035 7615.115 1209.16 ;
      RECT 7610.48 1053.415 7623.48 1118.87 ;
      RECT 7610.48 1048.035 7621.85 1118.87 ;
      RECT 7610.48 1048.035 7623.48 1049.12 ;
      RECT 7593.5 1070.44 7606.5 1189.16 ;
      RECT 7596.865 1048.035 7606.5 1189.16 ;
      RECT 7593.5 1048.035 7606.5 1054.07 ;
      RECT 7576.52 1118.44 7589.52 1209.16 ;
      RECT 7578.375 1048.035 7589.52 1209.16 ;
      RECT 7576.52 1048.035 7589.52 1087.87 ;
      RECT 7546 1166.44 7574 1209.16 ;
      RECT 7560.475 1118.44 7574 1209.16 ;
      RECT 7546 1048.035 7555.565 1209.16 ;
      RECT 7546 1087.44 7570.625 1150.07 ;
      RECT 7564.53 1048.035 7574 1087.87 ;
      RECT 7560.475 1053.365 7574 1087.87 ;
      RECT 7546 1053.365 7574 1071.07 ;
      RECT 7546 1048.035 7558.81 1071.07 ;
      RECT 7546 1048.035 7574 1049.165 ;
      RECT 7530.48 1183.44 7543.48 1209.16 ;
      RECT 7538.145 1048.035 7543.48 1209.16 ;
      RECT 7533.475 1166.44 7543.48 1209.16 ;
      RECT 7530.48 1166.44 7543.48 1167.07 ;
      RECT 7530.48 1070.44 7533.235 1167.07 ;
      RECT 7530.48 1087.44 7543.48 1150.07 ;
      RECT 7530.48 1070.44 7543.48 1071.07 ;
      RECT 7533.475 1048.035 7543.48 1071.07 ;
      RECT 7530.48 1048.035 7543.48 1054.07 ;
      RECT 7496.52 1183.44 7509.52 1209.16 ;
      RECT 7496.52 1087.44 7507.235 1209.16 ;
      RECT 7501.75 1070.44 7509.52 1167.07 ;
      RECT 7496.52 1048.035 7504.565 1071.07 ;
      RECT 7496.52 1048.035 7509.52 1054.07 ;
      RECT 7466 1149.44 7494 1209.16 ;
      RECT 7484.63 1048.035 7494 1209.16 ;
      RECT 7482.865 1053.42 7494 1209.16 ;
      RECT 7466 1048.035 7475.115 1209.16 ;
      RECT 7466 1053.42 7494 1118.87 ;
      RECT 7466 1048.035 7481.85 1118.87 ;
      RECT 7466 1048.035 7494 1049.12 ;
      RECT 7450.48 1070.44 7463.48 1209.16 ;
      RECT 7456.865 1048.035 7463.48 1209.16 ;
      RECT 7450.48 1048.035 7451.955 1209.16 ;
      RECT 7450.48 1048.035 7463.48 1054.07 ;
      RECT 7433.5 1118.44 7446.5 1189.16 ;
      RECT 7438.375 1048.035 7446.5 1189.16 ;
      RECT 7433.5 1048.035 7446.5 1087.87 ;
      RECT 7416.52 1166.44 7429.52 1209.16 ;
      RECT 7424.53 1048.035 7429.52 1209.16 ;
      RECT 7420.475 1053.365 7429.52 1209.16 ;
      RECT 7416.52 1087.44 7429.52 1150.07 ;
      RECT 7416.52 1053.365 7429.52 1071.07 ;
      RECT 7416.52 1048.035 7418.81 1071.07 ;
      RECT 7416.52 1048.035 7429.52 1049.375 ;
      RECT 7386 1183.44 7414 1209.16 ;
      RECT 7398.145 1048.035 7414 1209.16 ;
      RECT 7393.475 1166.44 7414 1209.16 ;
      RECT 7386 1048.035 7388.565 1209.16 ;
      RECT 7386 1166.44 7414 1167.07 ;
      RECT 7386 1070.44 7393.235 1167.07 ;
      RECT 7386 1087.44 7414 1150.07 ;
      RECT 7386 1070.44 7414 1071.07 ;
      RECT 7393.475 1048.035 7414 1071.07 ;
      RECT 7386 1048.035 7414 1054.07 ;
      RECT 7370.48 1183.44 7383.48 1209.16 ;
      RECT 7372.145 1048.035 7383.48 1209.16 ;
      RECT 7370.48 1048.035 7383.48 1167.07 ;
      RECT 7353.5 1087.44 7366.5 1189.16 ;
      RECT 7360.13 1070.44 7366.5 1189.16 ;
      RECT 7353.5 1048.035 7363.455 1071.07 ;
      RECT 7353.5 1048.035 7366.5 1054.07 ;
      RECT 7336.52 1149.44 7349.52 1209.16 ;
      RECT 7344.63 1048.035 7349.52 1209.16 ;
      RECT 7342.865 1053.42 7349.52 1209.16 ;
      RECT 7336.52 1053.42 7349.52 1118.87 ;
      RECT 7336.52 1048.035 7341.85 1118.87 ;
      RECT 7336.52 1048.035 7349.52 1049.12 ;
      RECT 7306 1070.44 7334 1209.16 ;
      RECT 7316.865 1048.035 7334 1209.16 ;
      RECT 7306 1048.035 7311.955 1209.16 ;
      RECT 7306 1048.035 7334 1054.07 ;
      RECT 7290.48 1118.44 7303.48 1209.16 ;
      RECT 7298.375 1048.035 7303.48 1209.16 ;
      RECT 7290.48 1048.035 7303.48 1087.87 ;
      RECT 7273.5 1166.44 7286.5 1189.16 ;
      RECT 7284.43 1048.035 7286.5 1189.16 ;
      RECT 7280.475 1053.365 7286.5 1189.16 ;
      RECT 7273.5 1048.035 7275.565 1189.16 ;
      RECT 7273.5 1087.44 7286.5 1150.07 ;
      RECT 7273.5 1053.365 7286.5 1071.07 ;
      RECT 7273.5 1048.035 7278.81 1071.07 ;
      RECT 7273.5 1048.035 7286.5 1049.165 ;
      RECT 7256.52 1166.44 7269.52 1209.16 ;
      RECT 7258.145 1048.035 7269.52 1209.16 ;
      RECT 7256.52 1087.44 7269.52 1150.07 ;
      RECT 7256.52 1048.035 7269.52 1071.07 ;
      RECT 7226 1183.44 7254 1209.16 ;
      RECT 7232.145 1048.035 7248.565 1209.16 ;
      RECT 7226 1070.44 7227.235 1209.16 ;
      RECT 7226 1070.44 7253.235 1167.07 ;
      RECT 7226 1087.44 7254 1150.07 ;
      RECT 7228.365 1048.035 7248.565 1167.07 ;
      RECT 7226 1048.035 7254 1054.07 ;
      RECT 7210.48 1087.44 7223.48 1209.16 ;
      RECT 7210.48 1048.035 7216.835 1209.16 ;
      RECT 7210.48 1048.035 7223.48 1071.07 ;
      RECT 7193.5 1149.44 7206.5 1189.16 ;
      RECT 7204.63 1048.035 7206.5 1189.16 ;
      RECT 7202.865 1053.42 7206.5 1189.16 ;
      RECT 7193.5 1048.035 7195.115 1189.16 ;
      RECT 7193.5 1053.42 7206.5 1118.87 ;
      RECT 7193.5 1048.035 7201.85 1118.87 ;
      RECT 7193.5 1048.035 7206.5 1049.12 ;
      RECT 7176.52 1070.44 7189.52 1209.16 ;
      RECT 7176.865 1048.035 7189.52 1209.16 ;
      RECT 7176.52 1048.035 7189.52 1054.07 ;
      RECT 7146 1118.44 7174 1209.16 ;
      RECT 7158.375 1070.44 7174 1209.16 ;
      RECT 7146 1048.035 7150.625 1209.16 ;
      RECT 7146 1048.035 7171.955 1087.87 ;
      RECT 7146 1048.035 7174 1054.07 ;
      RECT 7130.48 1166.44 7143.48 1209.16 ;
      RECT 7140.475 1053.365 7143.48 1209.16 ;
      RECT 7130.48 1048.035 7135.565 1209.16 ;
      RECT 7130.48 1087.44 7143.48 1150.07 ;
      RECT 7130.48 1053.365 7143.48 1071.07 ;
      RECT 7130.48 1048.035 7138.81 1071.07 ;
      RECT 7130.48 1048.035 7143.48 1049.165 ;
      RECT 7113.5 1166.44 7126.5 1189.16 ;
      RECT 7118.145 1048.035 7126.5 1189.16 ;
      RECT 7117.98 1087.44 7126.5 1189.16 ;
      RECT 7113.5 1087.44 7126.5 1150.07 ;
      RECT 7113.5 1048.035 7126.5 1071.07 ;
      RECT 7096.52 1183.44 7109.52 1209.16 ;
      RECT 7096.52 1048.035 7108.565 1209.16 ;
      RECT 7096.52 1070.44 7109.52 1167.07 ;
      RECT 7096.52 1048.035 7109.52 1054.07 ;
      RECT 7066 1183.44 7094 1209.16 ;
      RECT 7092.145 1048.035 7094 1209.16 ;
      RECT 7066 1087.44 7087.235 1209.16 ;
      RECT 7089.555 1048.035 7094 1167.07 ;
      RECT 7072.55 1070.44 7094 1167.07 ;
      RECT 7066 1048.035 7084.645 1071.07 ;
      RECT 7066 1048.035 7094 1054.07 ;
      RECT 7050.48 1149.44 7063.48 1209.16 ;
      RECT 7062.865 1053.415 7063.48 1209.16 ;
      RECT 7050.48 1048.035 7055.115 1209.16 ;
      RECT 7050.48 1053.415 7063.48 1118.87 ;
      RECT 7050.48 1048.035 7061.85 1118.87 ;
      RECT 7050.48 1048.035 7063.48 1049.12 ;
      RECT 7033.5 1070.44 7046.5 1189.16 ;
      RECT 7036.865 1048.035 7046.5 1189.16 ;
      RECT 7033.5 1048.035 7046.5 1054.07 ;
      RECT 7016.52 1118.44 7029.52 1209.16 ;
      RECT 7018.375 1048.035 7029.52 1209.16 ;
      RECT 7016.52 1048.035 7029.52 1087.87 ;
      RECT 6986 1166.44 7014 1209.16 ;
      RECT 7000.475 1118.44 7014 1209.16 ;
      RECT 6986 1048.035 6995.565 1209.16 ;
      RECT 6986 1087.44 7010.625 1150.07 ;
      RECT 7004.53 1048.035 7014 1087.87 ;
      RECT 7000.475 1053.365 7014 1087.87 ;
      RECT 6986 1053.365 7014 1071.07 ;
      RECT 6986 1048.035 6998.81 1071.07 ;
      RECT 6986 1048.035 7014 1049.165 ;
      RECT 6970.48 1183.44 6983.48 1209.16 ;
      RECT 6978.145 1048.035 6983.48 1209.16 ;
      RECT 6973.475 1166.44 6983.48 1209.16 ;
      RECT 6970.48 1166.44 6983.48 1167.07 ;
      RECT 6970.48 1070.44 6973.235 1167.07 ;
      RECT 6970.48 1087.44 6983.48 1150.07 ;
      RECT 6970.48 1070.44 6983.48 1071.07 ;
      RECT 6973.475 1048.035 6983.48 1071.07 ;
      RECT 6970.48 1048.035 6983.48 1054.07 ;
      RECT 6936.52 1183.44 6949.52 1209.16 ;
      RECT 6936.52 1087.44 6947.235 1209.16 ;
      RECT 6941.75 1070.44 6949.52 1167.07 ;
      RECT 6936.52 1048.035 6944.565 1071.07 ;
      RECT 6936.52 1048.035 6949.52 1054.07 ;
      RECT 6906 1149.44 6934 1209.16 ;
      RECT 6924.63 1048.035 6934 1209.16 ;
      RECT 6922.865 1053.42 6934 1209.16 ;
      RECT 6906 1048.035 6915.115 1209.16 ;
      RECT 6906 1053.42 6934 1118.87 ;
      RECT 6906 1048.035 6921.85 1118.87 ;
      RECT 6906 1048.035 6934 1049.12 ;
      RECT 6890.48 1070.44 6903.48 1209.16 ;
      RECT 6896.865 1048.035 6903.48 1209.16 ;
      RECT 6890.48 1048.035 6891.955 1209.16 ;
      RECT 6890.48 1048.035 6903.48 1054.07 ;
      RECT 6873.5 1118.44 6886.5 1189.16 ;
      RECT 6878.375 1048.035 6886.5 1189.16 ;
      RECT 6873.5 1048.035 6886.5 1087.87 ;
      RECT 6856.52 1166.44 6869.52 1209.16 ;
      RECT 6864.53 1048.035 6869.52 1209.16 ;
      RECT 6860.475 1053.365 6869.52 1209.16 ;
      RECT 6856.52 1087.44 6869.52 1150.07 ;
      RECT 6856.52 1053.365 6869.52 1071.07 ;
      RECT 6856.52 1048.035 6858.81 1071.07 ;
      RECT 6856.52 1048.035 6869.52 1049.375 ;
      RECT 6826 1183.44 6854 1209.16 ;
      RECT 6838.145 1048.035 6854 1209.16 ;
      RECT 6833.475 1166.44 6854 1209.16 ;
      RECT 6826 1048.035 6828.565 1209.16 ;
      RECT 6826 1166.44 6854 1167.07 ;
      RECT 6826 1070.44 6833.235 1167.07 ;
      RECT 6826 1087.44 6854 1150.07 ;
      RECT 6826 1070.44 6854 1071.07 ;
      RECT 6833.475 1048.035 6854 1071.07 ;
      RECT 6826 1048.035 6854 1054.07 ;
      RECT 6810.48 1183.44 6823.48 1209.16 ;
      RECT 6812.145 1048.035 6823.48 1209.16 ;
      RECT 6810.48 1048.035 6823.48 1167.07 ;
      RECT 6793.5 1087.44 6806.5 1189.16 ;
      RECT 6800.13 1070.44 6806.5 1189.16 ;
      RECT 6793.5 1048.035 6803.455 1071.07 ;
      RECT 6793.5 1048.035 6806.5 1054.07 ;
      RECT 6776.52 1149.44 6789.52 1209.16 ;
      RECT 6784.63 1048.035 6789.52 1209.16 ;
      RECT 6782.865 1053.42 6789.52 1209.16 ;
      RECT 6776.52 1053.42 6789.52 1118.87 ;
      RECT 6776.52 1048.035 6781.85 1118.87 ;
      RECT 6776.52 1048.035 6789.52 1049.12 ;
      RECT 6746 1070.44 6774 1209.16 ;
      RECT 6756.865 1048.035 6774 1209.16 ;
      RECT 6746 1048.035 6751.955 1209.16 ;
      RECT 6746 1048.035 6774 1054.07 ;
      RECT 6730.48 1118.44 6743.48 1209.16 ;
      RECT 6738.375 1048.035 6743.48 1209.16 ;
      RECT 6730.48 1048.035 6743.48 1087.87 ;
      RECT 6713.5 1166.44 6726.5 1189.16 ;
      RECT 6724.43 1048.035 6726.5 1189.16 ;
      RECT 6720.475 1053.365 6726.5 1189.16 ;
      RECT 6713.5 1048.035 6715.565 1189.16 ;
      RECT 6713.5 1087.44 6726.5 1150.07 ;
      RECT 6713.5 1053.365 6726.5 1071.07 ;
      RECT 6713.5 1048.035 6718.81 1071.07 ;
      RECT 6713.5 1048.035 6726.5 1049.165 ;
      RECT 6696.52 1166.44 6709.52 1209.16 ;
      RECT 6698.145 1048.035 6709.52 1209.16 ;
      RECT 6696.52 1087.44 6709.52 1150.07 ;
      RECT 6696.52 1048.035 6709.52 1071.07 ;
      RECT 6666 1183.44 6694 1209.16 ;
      RECT 6672.145 1048.035 6688.565 1209.16 ;
      RECT 6666 1070.44 6667.235 1209.16 ;
      RECT 6666 1070.44 6693.235 1167.07 ;
      RECT 6666 1087.44 6694 1150.07 ;
      RECT 6668.365 1048.035 6688.565 1167.07 ;
      RECT 6666 1048.035 6694 1054.07 ;
      RECT 6650.48 1087.44 6663.48 1209.16 ;
      RECT 6650.48 1048.035 6656.835 1209.16 ;
      RECT 6650.48 1048.035 6663.48 1071.07 ;
      RECT 6633.5 1149.44 6646.5 1189.16 ;
      RECT 6644.63 1048.035 6646.5 1189.16 ;
      RECT 6642.865 1053.42 6646.5 1189.16 ;
      RECT 6633.5 1048.035 6635.115 1189.16 ;
      RECT 6633.5 1053.42 6646.5 1118.87 ;
      RECT 6633.5 1048.035 6641.85 1118.87 ;
      RECT 6633.5 1048.035 6646.5 1049.12 ;
      RECT 6616.52 1070.44 6629.52 1209.16 ;
      RECT 6616.865 1048.035 6629.52 1209.16 ;
      RECT 6616.52 1048.035 6629.52 1054.07 ;
      RECT 6586 1118.44 6614 1209.16 ;
      RECT 6598.375 1070.44 6614 1209.16 ;
      RECT 6586 1048.035 6590.625 1209.16 ;
      RECT 6586 1048.035 6611.955 1087.87 ;
      RECT 6586 1048.035 6614 1054.07 ;
      RECT 6570.48 1166.44 6583.48 1209.16 ;
      RECT 6580.475 1053.365 6583.48 1209.16 ;
      RECT 6570.48 1048.035 6575.565 1209.16 ;
      RECT 6570.48 1087.44 6583.48 1150.07 ;
      RECT 6570.48 1053.365 6583.48 1071.07 ;
      RECT 6570.48 1048.035 6578.81 1071.07 ;
      RECT 6570.48 1048.035 6583.48 1049.165 ;
      RECT 6553.5 1166.44 6566.5 1189.16 ;
      RECT 6558.145 1048.035 6566.5 1189.16 ;
      RECT 6557.98 1087.44 6566.5 1189.16 ;
      RECT 6553.5 1087.44 6566.5 1150.07 ;
      RECT 6553.5 1048.035 6566.5 1071.07 ;
      RECT 6536.52 1183.44 6549.52 1209.16 ;
      RECT 6536.52 1048.035 6548.565 1209.16 ;
      RECT 6536.52 1070.44 6549.52 1167.07 ;
      RECT 6536.52 1048.035 6549.52 1054.07 ;
      RECT 6506 1183.44 6534 1209.16 ;
      RECT 6532.145 1048.035 6534 1209.16 ;
      RECT 6506 1087.44 6527.235 1209.16 ;
      RECT 6529.555 1048.035 6534 1167.07 ;
      RECT 6512.55 1070.44 6534 1167.07 ;
      RECT 6506 1048.035 6524.645 1071.07 ;
      RECT 6506 1048.035 6534 1054.07 ;
      RECT 6490.48 1149.44 6503.48 1209.16 ;
      RECT 6502.865 1053.415 6503.48 1209.16 ;
      RECT 6490.48 1048.035 6495.115 1209.16 ;
      RECT 6490.48 1053.415 6503.48 1118.87 ;
      RECT 6490.48 1048.035 6501.85 1118.87 ;
      RECT 6490.48 1048.035 6503.48 1049.12 ;
      RECT 6473.5 1070.44 6486.5 1189.16 ;
      RECT 6476.865 1048.035 6486.5 1189.16 ;
      RECT 6473.5 1048.035 6486.5 1054.07 ;
      RECT 6456.52 1118.44 6469.52 1209.16 ;
      RECT 6458.375 1048.035 6469.52 1209.16 ;
      RECT 6456.52 1048.035 6469.52 1087.87 ;
      RECT 6426 1166.44 6454 1209.16 ;
      RECT 6440.475 1118.44 6454 1209.16 ;
      RECT 6426 1048.035 6435.565 1209.16 ;
      RECT 6426 1087.44 6450.625 1150.07 ;
      RECT 6444.53 1048.035 6454 1087.87 ;
      RECT 6440.475 1053.365 6454 1087.87 ;
      RECT 6426 1053.365 6454 1071.07 ;
      RECT 6426 1048.035 6438.81 1071.07 ;
      RECT 6426 1048.035 6454 1049.165 ;
      RECT 6410.48 1183.44 6423.48 1209.16 ;
      RECT 6418.145 1048.035 6423.48 1209.16 ;
      RECT 6413.475 1166.44 6423.48 1209.16 ;
      RECT 6410.48 1166.44 6423.48 1167.07 ;
      RECT 6410.48 1070.44 6413.235 1167.07 ;
      RECT 6410.48 1087.44 6423.48 1150.07 ;
      RECT 6410.48 1070.44 6423.48 1071.07 ;
      RECT 6413.475 1048.035 6423.48 1071.07 ;
      RECT 6410.48 1048.035 6423.48 1054.07 ;
      RECT 6376.52 1183.44 6389.52 1209.16 ;
      RECT 6376.52 1087.44 6387.235 1209.16 ;
      RECT 6381.75 1070.44 6389.52 1167.07 ;
      RECT 6376.52 1048.035 6384.565 1071.07 ;
      RECT 6376.52 1048.035 6389.52 1054.07 ;
      RECT 6346 1149.44 6374 1209.16 ;
      RECT 6364.63 1048.035 6374 1209.16 ;
      RECT 6362.865 1053.42 6374 1209.16 ;
      RECT 6346 1048.035 6355.115 1209.16 ;
      RECT 6346 1053.42 6374 1118.87 ;
      RECT 6346 1048.035 6361.85 1118.87 ;
      RECT 6346 1048.035 6374 1049.12 ;
      RECT 6330.48 1070.44 6343.48 1209.16 ;
      RECT 6336.865 1048.035 6343.48 1209.16 ;
      RECT 6330.48 1048.035 6331.955 1209.16 ;
      RECT 6330.48 1048.035 6343.48 1054.07 ;
      RECT 6313.5 1118.44 6326.5 1189.16 ;
      RECT 6318.375 1048.035 6326.5 1189.16 ;
      RECT 6313.5 1048.035 6326.5 1087.87 ;
      RECT 6296.52 1166.44 6309.52 1209.16 ;
      RECT 6304.53 1048.035 6309.52 1209.16 ;
      RECT 6300.475 1053.365 6309.52 1209.16 ;
      RECT 6296.52 1087.44 6309.52 1150.07 ;
      RECT 6296.52 1053.365 6309.52 1071.07 ;
      RECT 6296.52 1048.035 6298.81 1071.07 ;
      RECT 6296.52 1048.035 6309.52 1049.375 ;
      RECT 6266 1183.44 6294 1209.16 ;
      RECT 6278.145 1048.035 6294 1209.16 ;
      RECT 6273.475 1166.44 6294 1209.16 ;
      RECT 6266 1048.035 6268.565 1209.16 ;
      RECT 6266 1166.44 6294 1167.07 ;
      RECT 6266 1070.44 6273.235 1167.07 ;
      RECT 6266 1087.44 6294 1150.07 ;
      RECT 6266 1070.44 6294 1071.07 ;
      RECT 6273.475 1048.035 6294 1071.07 ;
      RECT 6266 1048.035 6294 1054.07 ;
      RECT 6250.48 1183.44 6263.48 1209.16 ;
      RECT 6252.145 1048.035 6263.48 1209.16 ;
      RECT 6250.48 1048.035 6263.48 1167.07 ;
      RECT 6233.5 1087.44 6246.5 1189.16 ;
      RECT 6240.13 1070.44 6246.5 1189.16 ;
      RECT 6233.5 1048.035 6243.455 1071.07 ;
      RECT 6233.5 1048.035 6246.5 1054.07 ;
      RECT 6216.52 1149.44 6229.52 1209.16 ;
      RECT 6224.63 1048.035 6229.52 1209.16 ;
      RECT 6222.865 1053.42 6229.52 1209.16 ;
      RECT 6216.52 1053.42 6229.52 1118.87 ;
      RECT 6216.52 1048.035 6221.85 1118.87 ;
      RECT 6216.52 1048.035 6229.52 1049.12 ;
      RECT 6186 1070.44 6214 1209.16 ;
      RECT 6196.865 1048.035 6214 1209.16 ;
      RECT 6186 1048.035 6191.955 1209.16 ;
      RECT 6186 1048.035 6214 1054.07 ;
      RECT 6170.48 1118.44 6183.48 1209.16 ;
      RECT 6178.375 1048.035 6183.48 1209.16 ;
      RECT 6170.48 1048.035 6183.48 1087.87 ;
      RECT 6153.5 1166.44 6166.5 1189.16 ;
      RECT 6164.43 1048.035 6166.5 1189.16 ;
      RECT 6160.475 1053.365 6166.5 1189.16 ;
      RECT 6153.5 1048.035 6155.565 1189.16 ;
      RECT 6153.5 1087.44 6166.5 1150.07 ;
      RECT 6153.5 1053.365 6166.5 1071.07 ;
      RECT 6153.5 1048.035 6158.81 1071.07 ;
      RECT 6153.5 1048.035 6166.5 1049.165 ;
      RECT 6136.52 1166.44 6149.52 1209.16 ;
      RECT 6138.145 1048.035 6149.52 1209.16 ;
      RECT 6136.52 1087.44 6149.52 1150.07 ;
      RECT 6136.52 1048.035 6149.52 1071.07 ;
      RECT 6106 1183.44 6134 1209.16 ;
      RECT 6112.145 1048.035 6128.565 1209.16 ;
      RECT 6106 1070.44 6107.235 1209.16 ;
      RECT 6106 1070.44 6133.235 1167.07 ;
      RECT 6106 1087.44 6134 1150.07 ;
      RECT 6108.365 1048.035 6128.565 1167.07 ;
      RECT 6106 1048.035 6134 1054.07 ;
      RECT 6090.48 1087.44 6103.48 1209.16 ;
      RECT 6090.48 1048.035 6096.835 1209.16 ;
      RECT 6090.48 1048.035 6103.48 1071.07 ;
      RECT 6073.5 1149.44 6086.5 1189.16 ;
      RECT 6084.63 1048.035 6086.5 1189.16 ;
      RECT 6082.865 1053.42 6086.5 1189.16 ;
      RECT 6073.5 1048.035 6075.115 1189.16 ;
      RECT 6073.5 1053.42 6086.5 1118.87 ;
      RECT 6073.5 1048.035 6081.85 1118.87 ;
      RECT 6073.5 1048.035 6086.5 1049.12 ;
      RECT 6056.52 1070.44 6069.52 1209.16 ;
      RECT 6056.865 1048.035 6069.52 1209.16 ;
      RECT 6056.52 1048.035 6069.52 1054.07 ;
      RECT 6026 1118.44 6054 1209.16 ;
      RECT 6038.375 1070.44 6054 1209.16 ;
      RECT 6026 1048.035 6030.625 1209.16 ;
      RECT 6026 1048.035 6051.955 1087.87 ;
      RECT 6026 1048.035 6054 1054.07 ;
      RECT 6010.48 1166.44 6023.48 1209.16 ;
      RECT 6020.475 1053.365 6023.48 1209.16 ;
      RECT 6010.48 1048.035 6015.565 1209.16 ;
      RECT 6010.48 1087.44 6023.48 1150.07 ;
      RECT 6010.48 1053.365 6023.48 1071.07 ;
      RECT 6010.48 1048.035 6018.81 1071.07 ;
      RECT 6010.48 1048.035 6023.48 1049.165 ;
      RECT 5993.5 1166.44 6006.5 1189.16 ;
      RECT 5998.145 1048.035 6006.5 1189.16 ;
      RECT 5997.98 1087.44 6006.5 1189.16 ;
      RECT 5993.5 1087.44 6006.5 1150.07 ;
      RECT 5993.5 1048.035 6006.5 1071.07 ;
      RECT 5976.52 1183.44 5989.52 1209.16 ;
      RECT 5976.52 1048.035 5988.565 1209.16 ;
      RECT 5976.52 1070.44 5989.52 1167.07 ;
      RECT 5976.52 1048.035 5989.52 1054.07 ;
      RECT 5946 1183.44 5974 1209.16 ;
      RECT 5972.145 1048.035 5974 1209.16 ;
      RECT 5946 1087.44 5967.235 1209.16 ;
      RECT 5969.555 1048.035 5974 1167.07 ;
      RECT 5952.55 1070.44 5974 1167.07 ;
      RECT 5946 1048.035 5964.645 1071.07 ;
      RECT 5946 1048.035 5974 1054.07 ;
      RECT 5930.48 1149.44 5943.48 1209.16 ;
      RECT 5942.865 1053.415 5943.48 1209.16 ;
      RECT 5930.48 1048.035 5935.115 1209.16 ;
      RECT 5930.48 1053.415 5943.48 1118.87 ;
      RECT 5930.48 1048.035 5941.85 1118.87 ;
      RECT 5930.48 1048.035 5943.48 1049.12 ;
      RECT 5913.5 1070.44 5926.5 1189.16 ;
      RECT 5916.865 1048.035 5926.5 1189.16 ;
      RECT 5913.5 1048.035 5926.5 1054.07 ;
      RECT 5896.52 1118.44 5909.52 1209.16 ;
      RECT 5898.375 1048.035 5909.52 1209.16 ;
      RECT 5896.52 1048.035 5909.52 1087.87 ;
      RECT 5866 1166.44 5894 1209.16 ;
      RECT 5880.475 1118.44 5894 1209.16 ;
      RECT 5866 1048.035 5875.565 1209.16 ;
      RECT 5866 1087.44 5890.625 1150.07 ;
      RECT 5884.53 1048.035 5894 1087.87 ;
      RECT 5880.475 1053.365 5894 1087.87 ;
      RECT 5866 1053.365 5894 1071.07 ;
      RECT 5866 1048.035 5878.81 1071.07 ;
      RECT 5866 1048.035 5894 1049.165 ;
      RECT 5850.48 1183.44 5863.48 1209.16 ;
      RECT 5858.145 1048.035 5863.48 1209.16 ;
      RECT 5853.475 1166.44 5863.48 1209.16 ;
      RECT 5850.48 1166.44 5863.48 1167.07 ;
      RECT 5850.48 1070.44 5853.235 1167.07 ;
      RECT 5850.48 1087.44 5863.48 1150.07 ;
      RECT 5850.48 1070.44 5863.48 1071.07 ;
      RECT 5853.475 1048.035 5863.48 1071.07 ;
      RECT 5850.48 1048.035 5863.48 1054.07 ;
      RECT 5816.52 1183.44 5829.52 1209.16 ;
      RECT 5816.52 1087.44 5827.235 1209.16 ;
      RECT 5821.75 1070.44 5829.52 1167.07 ;
      RECT 5816.52 1048.035 5824.565 1071.07 ;
      RECT 5816.52 1048.035 5829.52 1054.07 ;
      RECT 5786 1149.44 5814 1209.16 ;
      RECT 5804.63 1048.035 5814 1209.16 ;
      RECT 5802.865 1053.42 5814 1209.16 ;
      RECT 5786 1048.035 5795.115 1209.16 ;
      RECT 5786 1053.42 5814 1118.87 ;
      RECT 5786 1048.035 5801.85 1118.87 ;
      RECT 5786 1048.035 5814 1049.12 ;
      RECT 5770.48 1070.44 5783.48 1209.16 ;
      RECT 5776.865 1048.035 5783.48 1209.16 ;
      RECT 5770.48 1048.035 5771.955 1209.16 ;
      RECT 5770.48 1048.035 5783.48 1054.07 ;
      RECT 5753.5 1118.44 5766.5 1189.16 ;
      RECT 5758.375 1048.035 5766.5 1189.16 ;
      RECT 5753.5 1048.035 5766.5 1087.87 ;
      RECT 5736.52 1166.44 5749.52 1209.16 ;
      RECT 5744.53 1048.035 5749.52 1209.16 ;
      RECT 5740.475 1053.365 5749.52 1209.16 ;
      RECT 5736.52 1087.44 5749.52 1150.07 ;
      RECT 5736.52 1053.365 5749.52 1071.07 ;
      RECT 5736.52 1048.035 5738.81 1071.07 ;
      RECT 5736.52 1048.035 5749.52 1049.375 ;
      RECT 5706 1183.44 5734 1209.16 ;
      RECT 5718.145 1048.035 5734 1209.16 ;
      RECT 5713.475 1166.44 5734 1209.16 ;
      RECT 5706 1048.035 5708.565 1209.16 ;
      RECT 5706 1166.44 5734 1167.07 ;
      RECT 5706 1070.44 5713.235 1167.07 ;
      RECT 5706 1087.44 5734 1150.07 ;
      RECT 5706 1070.44 5734 1071.07 ;
      RECT 5713.475 1048.035 5734 1071.07 ;
      RECT 5706 1048.035 5734 1054.07 ;
      RECT 5690.48 1183.44 5703.48 1209.16 ;
      RECT 5692.145 1048.035 5703.48 1209.16 ;
      RECT 5690.48 1048.035 5703.48 1167.07 ;
      RECT 5673.5 1087.44 5686.5 1189.16 ;
      RECT 5680.13 1070.44 5686.5 1189.16 ;
      RECT 5673.5 1048.035 5683.455 1071.07 ;
      RECT 5673.5 1048.035 5686.5 1054.07 ;
      RECT 5656.52 1149.44 5669.52 1209.16 ;
      RECT 5664.63 1048.035 5669.52 1209.16 ;
      RECT 5662.865 1053.42 5669.52 1209.16 ;
      RECT 5656.52 1053.42 5669.52 1118.87 ;
      RECT 5656.52 1048.035 5661.85 1118.87 ;
      RECT 5656.52 1048.035 5669.52 1049.12 ;
      RECT 5626 1070.44 5654 1209.16 ;
      RECT 5636.865 1048.035 5654 1209.16 ;
      RECT 5626 1048.035 5631.955 1209.16 ;
      RECT 5626 1048.035 5654 1054.07 ;
      RECT 5610.48 1118.44 5623.48 1209.16 ;
      RECT 5618.375 1048.035 5623.48 1209.16 ;
      RECT 5610.48 1048.035 5623.48 1087.87 ;
      RECT 5593.5 1166.44 5606.5 1189.16 ;
      RECT 5604.43 1048.035 5606.5 1189.16 ;
      RECT 5600.475 1053.365 5606.5 1189.16 ;
      RECT 5593.5 1048.035 5595.565 1189.16 ;
      RECT 5593.5 1087.44 5606.5 1150.07 ;
      RECT 5593.5 1053.365 5606.5 1071.07 ;
      RECT 5593.5 1048.035 5598.81 1071.07 ;
      RECT 5593.5 1048.035 5606.5 1049.165 ;
      RECT 5576.52 1166.44 5589.52 1209.16 ;
      RECT 5578.145 1048.035 5589.52 1209.16 ;
      RECT 5576.52 1087.44 5589.52 1150.07 ;
      RECT 5576.52 1048.035 5589.52 1071.07 ;
      RECT 5546 1183.44 5574 1209.16 ;
      RECT 5552.145 1048.035 5568.565 1209.16 ;
      RECT 5546 1070.44 5547.235 1209.16 ;
      RECT 5546 1070.44 5573.235 1167.07 ;
      RECT 5546 1087.44 5574 1150.07 ;
      RECT 5548.365 1048.035 5568.565 1167.07 ;
      RECT 5546 1048.035 5574 1054.07 ;
      RECT 5530.48 1087.44 5543.48 1209.16 ;
      RECT 5530.48 1048.035 5536.835 1209.16 ;
      RECT 5530.48 1048.035 5543.48 1071.07 ;
      RECT 5513.5 1149.44 5526.5 1189.16 ;
      RECT 5524.63 1048.035 5526.5 1189.16 ;
      RECT 5522.865 1053.42 5526.5 1189.16 ;
      RECT 5513.5 1048.035 5515.115 1189.16 ;
      RECT 5513.5 1053.42 5526.5 1118.87 ;
      RECT 5513.5 1048.035 5521.85 1118.87 ;
      RECT 5513.5 1048.035 5526.5 1049.12 ;
      RECT 5496.52 1070.44 5509.52 1209.16 ;
      RECT 5496.865 1048.035 5509.52 1209.16 ;
      RECT 5496.52 1048.035 5509.52 1054.07 ;
      RECT 5466 1118.44 5494 1209.16 ;
      RECT 5478.375 1070.44 5494 1209.16 ;
      RECT 5466 1048.035 5470.625 1209.16 ;
      RECT 5466 1048.035 5491.955 1087.87 ;
      RECT 5466 1048.035 5494 1054.07 ;
      RECT 5450.48 1166.44 5463.48 1209.16 ;
      RECT 5460.475 1053.365 5463.48 1209.16 ;
      RECT 5450.48 1048.035 5455.565 1209.16 ;
      RECT 5450.48 1087.44 5463.48 1150.07 ;
      RECT 5450.48 1053.365 5463.48 1071.07 ;
      RECT 5450.48 1048.035 5458.81 1071.07 ;
      RECT 5450.48 1048.035 5463.48 1049.165 ;
      RECT 5433.5 1166.44 5446.5 1189.16 ;
      RECT 5438.145 1048.035 5446.5 1189.16 ;
      RECT 5437.98 1087.44 5446.5 1189.16 ;
      RECT 5433.5 1087.44 5446.5 1150.07 ;
      RECT 5433.5 1048.035 5446.5 1071.07 ;
      RECT 5416.52 1183.44 5429.52 1209.16 ;
      RECT 5416.52 1048.035 5428.565 1209.16 ;
      RECT 5416.52 1070.44 5429.52 1167.07 ;
      RECT 5416.52 1048.035 5429.52 1054.07 ;
      RECT 5386 1183.44 5414 1209.16 ;
      RECT 5412.145 1048.035 5414 1209.16 ;
      RECT 5386 1087.44 5407.235 1209.16 ;
      RECT 5409.555 1048.035 5414 1167.07 ;
      RECT 5392.55 1070.44 5414 1167.07 ;
      RECT 5386 1048.035 5404.645 1071.07 ;
      RECT 5386 1048.035 5414 1054.07 ;
      RECT 5370.48 1149.44 5383.48 1209.16 ;
      RECT 5382.865 1053.415 5383.48 1209.16 ;
      RECT 5370.48 1048.035 5375.115 1209.16 ;
      RECT 5370.48 1053.415 5383.48 1118.87 ;
      RECT 5370.48 1048.035 5381.85 1118.87 ;
      RECT 5370.48 1048.035 5383.48 1049.12 ;
      RECT 5353.5 1070.44 5366.5 1189.16 ;
      RECT 5356.865 1048.035 5366.5 1189.16 ;
      RECT 5353.5 1048.035 5366.5 1054.07 ;
      RECT 5336.52 1118.44 5349.52 1209.16 ;
      RECT 5338.375 1048.035 5349.52 1209.16 ;
      RECT 5336.52 1048.035 5349.52 1087.87 ;
      RECT 5306 1166.44 5334 1209.16 ;
      RECT 5320.475 1118.44 5334 1209.16 ;
      RECT 5306 1048.035 5315.565 1209.16 ;
      RECT 5306 1087.44 5330.625 1150.07 ;
      RECT 5324.53 1048.035 5334 1087.87 ;
      RECT 5320.475 1053.365 5334 1087.87 ;
      RECT 5306 1053.365 5334 1071.07 ;
      RECT 5306 1048.035 5318.81 1071.07 ;
      RECT 5306 1048.035 5334 1049.165 ;
      RECT 5290.48 1183.44 5303.48 1209.16 ;
      RECT 5298.145 1048.035 5303.48 1209.16 ;
      RECT 5293.475 1166.44 5303.48 1209.16 ;
      RECT 5290.48 1166.44 5303.48 1167.07 ;
      RECT 5290.48 1070.44 5293.235 1167.07 ;
      RECT 5290.48 1087.44 5303.48 1150.07 ;
      RECT 5290.48 1070.44 5303.48 1071.07 ;
      RECT 5293.475 1048.035 5303.48 1071.07 ;
      RECT 5290.48 1048.035 5303.48 1054.07 ;
      RECT 5256.52 1183.44 5269.52 1209.16 ;
      RECT 5256.52 1087.44 5267.235 1209.16 ;
      RECT 5261.75 1070.44 5269.52 1167.07 ;
      RECT 5256.52 1048.035 5264.565 1071.07 ;
      RECT 5256.52 1048.035 5269.52 1054.07 ;
      RECT 5226 1149.44 5254 1209.16 ;
      RECT 5244.63 1048.035 5254 1209.16 ;
      RECT 5242.865 1053.42 5254 1209.16 ;
      RECT 5226 1048.035 5235.115 1209.16 ;
      RECT 5226 1053.42 5254 1118.87 ;
      RECT 5226 1048.035 5241.85 1118.87 ;
      RECT 5226 1048.035 5254 1049.12 ;
      RECT 5210.48 1070.44 5223.48 1209.16 ;
      RECT 5216.865 1048.035 5223.48 1209.16 ;
      RECT 5210.48 1048.035 5211.955 1209.16 ;
      RECT 5210.48 1048.035 5223.48 1054.07 ;
      RECT 5193.5 1118.44 5206.5 1189.16 ;
      RECT 5198.375 1048.035 5206.5 1189.16 ;
      RECT 5193.5 1048.035 5206.5 1087.87 ;
      RECT 5176.52 1166.44 5189.52 1209.16 ;
      RECT 5184.53 1048.035 5189.52 1209.16 ;
      RECT 5180.475 1053.365 5189.52 1209.16 ;
      RECT 5176.52 1087.44 5189.52 1150.07 ;
      RECT 5176.52 1053.365 5189.52 1071.07 ;
      RECT 5176.52 1048.035 5178.81 1071.07 ;
      RECT 5176.52 1048.035 5189.52 1049.375 ;
      RECT 5146 1183.44 5174 1209.16 ;
      RECT 5158.145 1048.035 5174 1209.16 ;
      RECT 5153.475 1166.44 5174 1209.16 ;
      RECT 5146 1048.035 5148.565 1209.16 ;
      RECT 5146 1166.44 5174 1167.07 ;
      RECT 5146 1070.44 5153.235 1167.07 ;
      RECT 5146 1087.44 5174 1150.07 ;
      RECT 5146 1070.44 5174 1071.07 ;
      RECT 5153.475 1048.035 5174 1071.07 ;
      RECT 5146 1048.035 5174 1054.07 ;
      RECT 5130.48 1183.44 5143.48 1209.16 ;
      RECT 5132.145 1048.035 5143.48 1209.16 ;
      RECT 5130.48 1048.035 5143.48 1167.07 ;
      RECT 5113.5 1087.44 5126.5 1189.16 ;
      RECT 5120.13 1070.44 5126.5 1189.16 ;
      RECT 5113.5 1048.035 5123.455 1071.07 ;
      RECT 5113.5 1048.035 5126.5 1054.07 ;
      RECT 5096.52 1149.44 5109.52 1209.16 ;
      RECT 5104.63 1048.035 5109.52 1209.16 ;
      RECT 5102.865 1053.42 5109.52 1209.16 ;
      RECT 5096.52 1053.42 5109.52 1118.87 ;
      RECT 5096.52 1048.035 5101.85 1118.87 ;
      RECT 5096.52 1048.035 5109.52 1049.12 ;
      RECT 5066 1070.44 5094 1209.16 ;
      RECT 5076.865 1048.035 5094 1209.16 ;
      RECT 5066 1048.035 5071.955 1209.16 ;
      RECT 5066 1048.035 5094 1054.07 ;
      RECT 5050.48 1118.44 5063.48 1209.16 ;
      RECT 5058.375 1048.035 5063.48 1209.16 ;
      RECT 5050.48 1048.035 5063.48 1087.87 ;
      RECT 5033.5 1166.44 5046.5 1189.16 ;
      RECT 5044.43 1048.035 5046.5 1189.16 ;
      RECT 5040.475 1053.365 5046.5 1189.16 ;
      RECT 5033.5 1048.035 5035.565 1189.16 ;
      RECT 5033.5 1087.44 5046.5 1150.07 ;
      RECT 5033.5 1053.365 5046.5 1071.07 ;
      RECT 5033.5 1048.035 5038.81 1071.07 ;
      RECT 5033.5 1048.035 5046.5 1049.165 ;
      RECT 5016.52 1166.44 5029.52 1209.16 ;
      RECT 5018.145 1048.035 5029.52 1209.16 ;
      RECT 5016.52 1087.44 5029.52 1150.07 ;
      RECT 5016.52 1048.035 5029.52 1071.07 ;
      RECT 4986 1183.44 5014 1209.16 ;
      RECT 4992.145 1048.035 5008.565 1209.16 ;
      RECT 4986 1070.44 4987.235 1209.16 ;
      RECT 4986 1070.44 5013.235 1167.07 ;
      RECT 4986 1087.44 5014 1150.07 ;
      RECT 4988.365 1048.035 5008.565 1167.07 ;
      RECT 4986 1048.035 5014 1054.07 ;
      RECT 4970.48 1087.44 4983.48 1209.16 ;
      RECT 4970.48 1048.035 4976.835 1209.16 ;
      RECT 4970.48 1048.035 4983.48 1071.07 ;
      RECT 4953.5 1149.44 4966.5 1189.16 ;
      RECT 4964.63 1048.035 4966.5 1189.16 ;
      RECT 4962.865 1053.42 4966.5 1189.16 ;
      RECT 4953.5 1048.035 4955.115 1189.16 ;
      RECT 4953.5 1053.42 4966.5 1118.87 ;
      RECT 4953.5 1048.035 4961.85 1118.87 ;
      RECT 4953.5 1048.035 4966.5 1049.12 ;
      RECT 4936.52 1070.44 4949.52 1209.16 ;
      RECT 4936.865 1048.035 4949.52 1209.16 ;
      RECT 4936.52 1048.035 4949.52 1054.07 ;
      RECT 4906 1118.44 4934 1209.16 ;
      RECT 4918.375 1070.44 4934 1209.16 ;
      RECT 4906 1048.035 4910.625 1209.16 ;
      RECT 4906 1048.035 4931.955 1087.87 ;
      RECT 4906 1048.035 4934 1054.07 ;
      RECT 4890.48 1166.44 4903.48 1209.16 ;
      RECT 4900.475 1053.365 4903.48 1209.16 ;
      RECT 4890.48 1048.035 4895.565 1209.16 ;
      RECT 4890.48 1087.44 4903.48 1150.07 ;
      RECT 4890.48 1053.365 4903.48 1071.07 ;
      RECT 4890.48 1048.035 4898.81 1071.07 ;
      RECT 4890.48 1048.035 4903.48 1049.165 ;
      RECT 4873.5 1166.44 4886.5 1189.16 ;
      RECT 4878.145 1048.035 4886.5 1189.16 ;
      RECT 4877.98 1087.44 4886.5 1189.16 ;
      RECT 4873.5 1087.44 4886.5 1150.07 ;
      RECT 4873.5 1048.035 4886.5 1071.07 ;
      RECT 4856.52 1183.44 4869.52 1209.16 ;
      RECT 4856.52 1048.035 4868.565 1209.16 ;
      RECT 4856.52 1070.44 4869.52 1167.07 ;
      RECT 4856.52 1048.035 4869.52 1054.07 ;
      RECT 4826 1183.44 4854 1209.16 ;
      RECT 4852.145 1048.035 4854 1209.16 ;
      RECT 4826 1087.44 4847.235 1209.16 ;
      RECT 4849.555 1048.035 4854 1167.07 ;
      RECT 4832.55 1070.44 4854 1167.07 ;
      RECT 4826 1048.035 4844.645 1071.07 ;
      RECT 4826 1048.035 4854 1054.07 ;
      RECT 4810.48 1149.44 4823.48 1209.16 ;
      RECT 4822.865 1053.415 4823.48 1209.16 ;
      RECT 4810.48 1048.035 4815.115 1209.16 ;
      RECT 4810.48 1053.415 4823.48 1118.87 ;
      RECT 4810.48 1048.035 4821.85 1118.87 ;
      RECT 4810.48 1048.035 4823.48 1049.12 ;
      RECT 4793.5 1070.44 4806.5 1189.16 ;
      RECT 4796.865 1048.035 4806.5 1189.16 ;
      RECT 4793.5 1048.035 4806.5 1054.07 ;
      RECT 4776.52 1118.44 4789.52 1209.16 ;
      RECT 4778.375 1048.035 4789.52 1209.16 ;
      RECT 4776.52 1048.035 4789.52 1087.87 ;
      RECT 4746 1166.44 4774 1209.16 ;
      RECT 4760.475 1118.44 4774 1209.16 ;
      RECT 4746 1048.035 4755.565 1209.16 ;
      RECT 4746 1087.44 4770.625 1150.07 ;
      RECT 4764.53 1048.035 4774 1087.87 ;
      RECT 4760.475 1053.365 4774 1087.87 ;
      RECT 4746 1053.365 4774 1071.07 ;
      RECT 4746 1048.035 4758.81 1071.07 ;
      RECT 4746 1048.035 4774 1049.165 ;
      RECT 4730.48 1183.44 4743.48 1209.16 ;
      RECT 4738.145 1048.035 4743.48 1209.16 ;
      RECT 4733.475 1166.44 4743.48 1209.16 ;
      RECT 4730.48 1166.44 4743.48 1167.07 ;
      RECT 4730.48 1070.44 4733.235 1167.07 ;
      RECT 4730.48 1087.44 4743.48 1150.07 ;
      RECT 4730.48 1070.44 4743.48 1071.07 ;
      RECT 4733.475 1048.035 4743.48 1071.07 ;
      RECT 4730.48 1048.035 4743.48 1054.07 ;
      RECT 4696.52 1183.44 4709.52 1209.16 ;
      RECT 4696.52 1087.44 4707.235 1209.16 ;
      RECT 4701.75 1070.44 4709.52 1167.07 ;
      RECT 4696.52 1048.035 4704.565 1071.07 ;
      RECT 4696.52 1048.035 4709.52 1054.07 ;
      RECT 4666 1149.44 4694 1209.16 ;
      RECT 4684.63 1048.035 4694 1209.16 ;
      RECT 4682.865 1053.42 4694 1209.16 ;
      RECT 4666 1048.035 4675.115 1209.16 ;
      RECT 4666 1053.42 4694 1118.87 ;
      RECT 4666 1048.035 4681.85 1118.87 ;
      RECT 4666 1048.035 4694 1049.12 ;
      RECT 4650.48 1070.44 4663.48 1209.16 ;
      RECT 4656.865 1048.035 4663.48 1209.16 ;
      RECT 4650.48 1048.035 4651.955 1209.16 ;
      RECT 4650.48 1048.035 4663.48 1054.07 ;
      RECT 4633.5 1118.44 4646.5 1189.16 ;
      RECT 4638.375 1048.035 4646.5 1189.16 ;
      RECT 4633.5 1048.035 4646.5 1087.87 ;
      RECT 4616.52 1166.44 4629.52 1209.16 ;
      RECT 4624.53 1048.035 4629.52 1209.16 ;
      RECT 4620.475 1053.365 4629.52 1209.16 ;
      RECT 4616.52 1087.44 4629.52 1150.07 ;
      RECT 4616.52 1053.365 4629.52 1071.07 ;
      RECT 4616.52 1048.035 4618.81 1071.07 ;
      RECT 4616.52 1048.035 4629.52 1049.375 ;
      RECT 4586 1183.44 4614 1209.16 ;
      RECT 4598.145 1048.035 4614 1209.16 ;
      RECT 4593.475 1166.44 4614 1209.16 ;
      RECT 4586 1048.035 4588.565 1209.16 ;
      RECT 4586 1166.44 4614 1167.07 ;
      RECT 4586 1070.44 4593.235 1167.07 ;
      RECT 4586 1087.44 4614 1150.07 ;
      RECT 4586 1070.44 4614 1071.07 ;
      RECT 4593.475 1048.035 4614 1071.07 ;
      RECT 4586 1048.035 4614 1054.07 ;
      RECT 4570.48 1183.44 4583.48 1209.16 ;
      RECT 4572.145 1048.035 4583.48 1209.16 ;
      RECT 4570.48 1048.035 4583.48 1167.07 ;
      RECT 4553.5 1087.44 4566.5 1189.16 ;
      RECT 4560.13 1070.44 4566.5 1189.16 ;
      RECT 4553.5 1048.035 4563.455 1071.07 ;
      RECT 4553.5 1048.035 4566.5 1054.07 ;
      RECT 4536.52 1149.44 4549.52 1209.16 ;
      RECT 4544.63 1048.035 4549.52 1209.16 ;
      RECT 4542.865 1053.42 4549.52 1209.16 ;
      RECT 4536.52 1053.42 4549.52 1118.87 ;
      RECT 4536.52 1048.035 4541.85 1118.87 ;
      RECT 4536.52 1048.035 4549.52 1049.12 ;
      RECT 4506 1070.44 4534 1209.16 ;
      RECT 4516.865 1048.035 4534 1209.16 ;
      RECT 4506 1048.035 4511.955 1209.16 ;
      RECT 4506 1048.035 4534 1054.07 ;
      RECT 4490.48 1118.44 4503.48 1209.16 ;
      RECT 4498.375 1048.035 4503.48 1209.16 ;
      RECT 4490.48 1048.035 4503.48 1087.87 ;
      RECT 4473.5 1166.44 4486.5 1189.16 ;
      RECT 4484.43 1048.035 4486.5 1189.16 ;
      RECT 4480.475 1053.365 4486.5 1189.16 ;
      RECT 4473.5 1048.035 4475.565 1189.16 ;
      RECT 4473.5 1087.44 4486.5 1150.07 ;
      RECT 4473.5 1053.365 4486.5 1071.07 ;
      RECT 4473.5 1048.035 4478.81 1071.07 ;
      RECT 4473.5 1048.035 4486.5 1049.165 ;
      RECT 4456.52 1166.44 4469.52 1209.16 ;
      RECT 4458.145 1048.035 4469.52 1209.16 ;
      RECT 4456.52 1087.44 4469.52 1150.07 ;
      RECT 4456.52 1048.035 4469.52 1071.07 ;
      RECT 4426 1183.44 4454 1209.16 ;
      RECT 4432.145 1048.035 4448.565 1209.16 ;
      RECT 4426 1070.44 4427.235 1209.16 ;
      RECT 4426 1070.44 4453.235 1167.07 ;
      RECT 4426 1087.44 4454 1150.07 ;
      RECT 4428.365 1048.035 4448.565 1167.07 ;
      RECT 4426 1048.035 4454 1054.07 ;
      RECT 4410.48 1087.44 4423.48 1209.16 ;
      RECT 4410.48 1048.035 4416.835 1209.16 ;
      RECT 4410.48 1048.035 4423.48 1071.07 ;
      RECT 4393.5 1149.44 4406.5 1189.16 ;
      RECT 4404.63 1048.035 4406.5 1189.16 ;
      RECT 4402.865 1053.42 4406.5 1189.16 ;
      RECT 4393.5 1048.035 4395.115 1189.16 ;
      RECT 4393.5 1053.42 4406.5 1118.87 ;
      RECT 4393.5 1048.035 4401.85 1118.87 ;
      RECT 4393.5 1048.035 4406.5 1049.12 ;
      RECT 4376.52 1070.44 4389.52 1209.16 ;
      RECT 4376.865 1048.035 4389.52 1209.16 ;
      RECT 4376.52 1048.035 4389.52 1054.07 ;
      RECT 4346 1118.44 4374 1209.16 ;
      RECT 4358.375 1070.44 4374 1209.16 ;
      RECT 4346 1048.035 4350.625 1209.16 ;
      RECT 4346 1048.035 4371.955 1087.87 ;
      RECT 4346 1048.035 4374 1054.07 ;
      RECT 4330.48 1166.44 4343.48 1209.16 ;
      RECT 4340.475 1053.365 4343.48 1209.16 ;
      RECT 4330.48 1048.035 4335.565 1209.16 ;
      RECT 4330.48 1087.44 4343.48 1150.07 ;
      RECT 4330.48 1053.365 4343.48 1071.07 ;
      RECT 4330.48 1048.035 4338.81 1071.07 ;
      RECT 4330.48 1048.035 4343.48 1049.165 ;
      RECT 4313.5 1166.44 4326.5 1189.16 ;
      RECT 4318.145 1048.035 4326.5 1189.16 ;
      RECT 4317.98 1087.44 4326.5 1189.16 ;
      RECT 4313.5 1087.44 4326.5 1150.07 ;
      RECT 4313.5 1048.035 4326.5 1071.07 ;
      RECT 4296.52 1183.44 4309.52 1209.16 ;
      RECT 4296.52 1048.035 4308.565 1209.16 ;
      RECT 4296.52 1070.44 4309.52 1167.07 ;
      RECT 4296.52 1048.035 4309.52 1054.07 ;
      RECT 4266 1183.44 4294 1209.16 ;
      RECT 4292.145 1048.035 4294 1209.16 ;
      RECT 4266 1087.44 4287.235 1209.16 ;
      RECT 4289.555 1048.035 4294 1167.07 ;
      RECT 4272.55 1070.44 4294 1167.07 ;
      RECT 4266 1048.035 4284.645 1071.07 ;
      RECT 4266 1048.035 4294 1054.07 ;
      RECT 4250.48 1149.44 4263.48 1209.16 ;
      RECT 4262.865 1053.415 4263.48 1209.16 ;
      RECT 4250.48 1048.035 4255.115 1209.16 ;
      RECT 4250.48 1053.415 4263.48 1118.87 ;
      RECT 4250.48 1048.035 4261.85 1118.87 ;
      RECT 4250.48 1048.035 4263.48 1049.12 ;
      RECT 4233.5 1070.44 4246.5 1189.16 ;
      RECT 4236.865 1048.035 4246.5 1189.16 ;
      RECT 4233.5 1048.035 4246.5 1054.07 ;
      RECT 4216.52 1118.44 4229.52 1209.16 ;
      RECT 4218.375 1048.035 4229.52 1209.16 ;
      RECT 4216.52 1048.035 4229.52 1087.87 ;
      RECT 4186 1166.44 4214 1209.16 ;
      RECT 4200.475 1118.44 4214 1209.16 ;
      RECT 4186 1048.035 4195.565 1209.16 ;
      RECT 4186 1087.44 4210.625 1150.07 ;
      RECT 4204.53 1048.035 4214 1087.87 ;
      RECT 4200.475 1053.365 4214 1087.87 ;
      RECT 4186 1053.365 4214 1071.07 ;
      RECT 4186 1048.035 4198.81 1071.07 ;
      RECT 4186 1048.035 4214 1049.165 ;
      RECT 4170.48 1183.44 4183.48 1209.16 ;
      RECT 4178.145 1048.035 4183.48 1209.16 ;
      RECT 4173.475 1166.44 4183.48 1209.16 ;
      RECT 4170.48 1166.44 4183.48 1167.07 ;
      RECT 4170.48 1070.44 4173.235 1167.07 ;
      RECT 4170.48 1087.44 4183.48 1150.07 ;
      RECT 4170.48 1070.44 4183.48 1071.07 ;
      RECT 4173.475 1048.035 4183.48 1071.07 ;
      RECT 4170.48 1048.035 4183.48 1054.07 ;
      RECT 4136.52 1183.44 4149.52 1209.16 ;
      RECT 4136.52 1087.44 4147.235 1209.16 ;
      RECT 4141.75 1070.44 4149.52 1167.07 ;
      RECT 4136.52 1048.035 4144.565 1071.07 ;
      RECT 4136.52 1048.035 4149.52 1054.07 ;
      RECT 4106 1149.44 4134 1209.16 ;
      RECT 4124.63 1048.035 4134 1209.16 ;
      RECT 4122.865 1053.42 4134 1209.16 ;
      RECT 4106 1048.035 4115.115 1209.16 ;
      RECT 4106 1053.42 4134 1118.87 ;
      RECT 4106 1048.035 4121.85 1118.87 ;
      RECT 4106 1048.035 4134 1049.12 ;
      RECT 4090.48 1070.44 4103.48 1209.16 ;
      RECT 4096.865 1048.035 4103.48 1209.16 ;
      RECT 4090.48 1048.035 4091.955 1209.16 ;
      RECT 4090.48 1048.035 4103.48 1054.07 ;
      RECT 4073.5 1118.44 4086.5 1189.16 ;
      RECT 4078.375 1048.035 4086.5 1189.16 ;
      RECT 4073.5 1048.035 4086.5 1087.87 ;
      RECT 4056.52 1166.44 4069.52 1209.16 ;
      RECT 4064.53 1048.035 4069.52 1209.16 ;
      RECT 4060.475 1053.365 4069.52 1209.16 ;
      RECT 4056.52 1087.44 4069.52 1150.07 ;
      RECT 4056.52 1053.365 4069.52 1071.07 ;
      RECT 4056.52 1048.035 4058.81 1071.07 ;
      RECT 4056.52 1048.035 4069.52 1049.375 ;
      RECT 4026 1183.44 4054 1209.16 ;
      RECT 4038.145 1048.035 4054 1209.16 ;
      RECT 4033.475 1166.44 4054 1209.16 ;
      RECT 4026 1048.035 4028.565 1209.16 ;
      RECT 4026 1166.44 4054 1167.07 ;
      RECT 4026 1070.44 4033.235 1167.07 ;
      RECT 4026 1087.44 4054 1150.07 ;
      RECT 4026 1070.44 4054 1071.07 ;
      RECT 4033.475 1048.035 4054 1071.07 ;
      RECT 4026 1048.035 4054 1054.07 ;
      RECT 4010.48 1183.44 4023.48 1209.16 ;
      RECT 4012.145 1048.035 4023.48 1209.16 ;
      RECT 4010.48 1048.035 4023.48 1167.07 ;
      RECT 3993.5 1087.44 4006.5 1189.16 ;
      RECT 4000.13 1070.44 4006.5 1189.16 ;
      RECT 3993.5 1048.035 4003.455 1071.07 ;
      RECT 3993.5 1048.035 4006.5 1054.07 ;
      RECT 3976.52 1149.44 3989.52 1209.16 ;
      RECT 3984.63 1048.035 3989.52 1209.16 ;
      RECT 3982.865 1053.42 3989.52 1209.16 ;
      RECT 3976.52 1053.42 3989.52 1118.87 ;
      RECT 3976.52 1048.035 3981.85 1118.87 ;
      RECT 3976.52 1048.035 3989.52 1049.12 ;
      RECT 3946 1070.44 3974 1209.16 ;
      RECT 3956.865 1048.035 3974 1209.16 ;
      RECT 3946 1048.035 3951.955 1209.16 ;
      RECT 3946 1048.035 3974 1054.07 ;
      RECT 3930.48 1118.44 3943.48 1209.16 ;
      RECT 3938.375 1048.035 3943.48 1209.16 ;
      RECT 3930.48 1048.035 3943.48 1087.87 ;
      RECT 3913.5 1166.44 3926.5 1189.16 ;
      RECT 3924.43 1048.035 3926.5 1189.16 ;
      RECT 3920.475 1053.365 3926.5 1189.16 ;
      RECT 3913.5 1048.035 3915.565 1189.16 ;
      RECT 3913.5 1087.44 3926.5 1150.07 ;
      RECT 3913.5 1053.365 3926.5 1071.07 ;
      RECT 3913.5 1048.035 3918.81 1071.07 ;
      RECT 3913.5 1048.035 3926.5 1049.165 ;
      RECT 3896.52 1166.44 3909.52 1209.16 ;
      RECT 3898.145 1048.035 3909.52 1209.16 ;
      RECT 3896.52 1087.44 3909.52 1150.07 ;
      RECT 3896.52 1048.035 3909.52 1071.07 ;
      RECT 3866 1183.44 3894 1209.16 ;
      RECT 3872.145 1048.035 3888.565 1209.16 ;
      RECT 3866 1070.44 3867.235 1209.16 ;
      RECT 3866 1070.44 3893.235 1167.07 ;
      RECT 3866 1087.44 3894 1150.07 ;
      RECT 3868.365 1048.035 3888.565 1167.07 ;
      RECT 3866 1048.035 3894 1054.07 ;
      RECT 3850.48 1087.44 3863.48 1209.16 ;
      RECT 3850.48 1048.035 3856.835 1209.16 ;
      RECT 3850.48 1048.035 3863.48 1071.07 ;
      RECT 3833.5 1149.44 3846.5 1189.16 ;
      RECT 3844.63 1048.035 3846.5 1189.16 ;
      RECT 3842.865 1053.42 3846.5 1189.16 ;
      RECT 3833.5 1048.035 3835.115 1189.16 ;
      RECT 3833.5 1053.42 3846.5 1118.87 ;
      RECT 3833.5 1048.035 3841.85 1118.87 ;
      RECT 3833.5 1048.035 3846.5 1049.12 ;
      RECT 3816.52 1070.44 3829.52 1209.16 ;
      RECT 3816.865 1048.035 3829.52 1209.16 ;
      RECT 3816.52 1048.035 3829.52 1054.07 ;
      RECT 3786 1118.44 3814 1209.16 ;
      RECT 3798.375 1070.44 3814 1209.16 ;
      RECT 3786 1048.035 3790.625 1209.16 ;
      RECT 3786 1048.035 3811.955 1087.87 ;
      RECT 3786 1048.035 3814 1054.07 ;
      RECT 3770.48 1166.44 3783.48 1209.16 ;
      RECT 3780.475 1053.365 3783.48 1209.16 ;
      RECT 3770.48 1048.035 3775.565 1209.16 ;
      RECT 3770.48 1087.44 3783.48 1150.07 ;
      RECT 3770.48 1053.365 3783.48 1071.07 ;
      RECT 3770.48 1048.035 3778.81 1071.07 ;
      RECT 3770.48 1048.035 3783.48 1049.165 ;
      RECT 3753.5 1166.44 3766.5 1189.16 ;
      RECT 3758.145 1048.035 3766.5 1189.16 ;
      RECT 3757.98 1087.44 3766.5 1189.16 ;
      RECT 3753.5 1087.44 3766.5 1150.07 ;
      RECT 3753.5 1048.035 3766.5 1071.07 ;
      RECT 3736.52 1183.44 3749.52 1209.16 ;
      RECT 3736.52 1048.035 3748.565 1209.16 ;
      RECT 3736.52 1070.44 3749.52 1167.07 ;
      RECT 3736.52 1048.035 3749.52 1054.07 ;
      RECT 3706 1183.44 3734 1209.16 ;
      RECT 3732.145 1048.035 3734 1209.16 ;
      RECT 3706 1087.44 3727.235 1209.16 ;
      RECT 3729.555 1048.035 3734 1167.07 ;
      RECT 3712.55 1070.44 3734 1167.07 ;
      RECT 3706 1048.035 3724.645 1071.07 ;
      RECT 3706 1048.035 3734 1054.07 ;
      RECT 3690.48 1149.44 3703.48 1209.16 ;
      RECT 3702.865 1053.415 3703.48 1209.16 ;
      RECT 3690.48 1048.035 3695.115 1209.16 ;
      RECT 3690.48 1053.415 3703.48 1118.87 ;
      RECT 3690.48 1048.035 3701.85 1118.87 ;
      RECT 3690.48 1048.035 3703.48 1049.12 ;
      RECT 3673.5 1070.44 3686.5 1189.16 ;
      RECT 3676.865 1048.035 3686.5 1189.16 ;
      RECT 3673.5 1048.035 3686.5 1054.07 ;
      RECT 3656.52 1118.44 3669.52 1209.16 ;
      RECT 3658.375 1048.035 3669.52 1209.16 ;
      RECT 3656.52 1048.035 3669.52 1087.87 ;
      RECT 3626 1166.44 3654 1209.16 ;
      RECT 3640.475 1118.44 3654 1209.16 ;
      RECT 3626 1048.035 3635.565 1209.16 ;
      RECT 3626 1087.44 3650.625 1150.07 ;
      RECT 3644.53 1048.035 3654 1087.87 ;
      RECT 3640.475 1053.365 3654 1087.87 ;
      RECT 3626 1053.365 3654 1071.07 ;
      RECT 3626 1048.035 3638.81 1071.07 ;
      RECT 3626 1048.035 3654 1049.165 ;
      RECT 3610.48 1183.44 3623.48 1209.16 ;
      RECT 3618.145 1048.035 3623.48 1209.16 ;
      RECT 3613.475 1166.44 3623.48 1209.16 ;
      RECT 3610.48 1166.44 3623.48 1167.07 ;
      RECT 3610.48 1070.44 3613.235 1167.07 ;
      RECT 3610.48 1087.44 3623.48 1150.07 ;
      RECT 3610.48 1070.44 3623.48 1071.07 ;
      RECT 3613.475 1048.035 3623.48 1071.07 ;
      RECT 3610.48 1048.035 3623.48 1054.07 ;
      RECT 3576.52 1183.44 3589.52 1209.16 ;
      RECT 3576.52 1087.44 3587.235 1209.16 ;
      RECT 3581.75 1070.44 3589.52 1167.07 ;
      RECT 3576.52 1048.035 3584.565 1071.07 ;
      RECT 3576.52 1048.035 3589.52 1054.07 ;
      RECT 3546 1149.44 3574 1209.16 ;
      RECT 3564.63 1048.035 3574 1209.16 ;
      RECT 3562.865 1053.42 3574 1209.16 ;
      RECT 3546 1048.035 3555.115 1209.16 ;
      RECT 3546 1053.42 3574 1118.87 ;
      RECT 3546 1048.035 3561.85 1118.87 ;
      RECT 3546 1048.035 3574 1049.12 ;
      RECT 3530.48 1070.44 3543.48 1209.16 ;
      RECT 3536.865 1048.035 3543.48 1209.16 ;
      RECT 3530.48 1048.035 3531.955 1209.16 ;
      RECT 3530.48 1048.035 3543.48 1054.07 ;
      RECT 3513.5 1118.44 3526.5 1189.16 ;
      RECT 3518.375 1048.035 3526.5 1189.16 ;
      RECT 3513.5 1048.035 3526.5 1087.87 ;
      RECT 3496.52 1166.44 3509.52 1209.16 ;
      RECT 3504.53 1048.035 3509.52 1209.16 ;
      RECT 3500.475 1053.365 3509.52 1209.16 ;
      RECT 3496.52 1087.44 3509.52 1150.07 ;
      RECT 3496.52 1053.365 3509.52 1071.07 ;
      RECT 3496.52 1048.035 3498.81 1071.07 ;
      RECT 3496.52 1048.035 3509.52 1049.375 ;
      RECT 3466 1183.44 3494 1209.16 ;
      RECT 3478.145 1048.035 3494 1209.16 ;
      RECT 3473.475 1166.44 3494 1209.16 ;
      RECT 3466 1048.035 3468.565 1209.16 ;
      RECT 3466 1166.44 3494 1167.07 ;
      RECT 3466 1070.44 3473.235 1167.07 ;
      RECT 3466 1087.44 3494 1150.07 ;
      RECT 3466 1070.44 3494 1071.07 ;
      RECT 3473.475 1048.035 3494 1071.07 ;
      RECT 3466 1048.035 3494 1054.07 ;
      RECT 3450.48 1183.44 3463.48 1209.16 ;
      RECT 3452.145 1048.035 3463.48 1209.16 ;
      RECT 3450.48 1048.035 3463.48 1167.07 ;
      RECT 3433.5 1087.44 3446.5 1189.16 ;
      RECT 3440.13 1070.44 3446.5 1189.16 ;
      RECT 3433.5 1048.035 3443.455 1071.07 ;
      RECT 3433.5 1048.035 3446.5 1054.07 ;
      RECT 3416.52 1149.44 3429.52 1209.16 ;
      RECT 3424.63 1048.035 3429.52 1209.16 ;
      RECT 3422.865 1053.42 3429.52 1209.16 ;
      RECT 3416.52 1053.42 3429.52 1118.87 ;
      RECT 3416.52 1048.035 3421.85 1118.87 ;
      RECT 3416.52 1048.035 3429.52 1049.12 ;
      RECT 3386 1070.44 3414 1209.16 ;
      RECT 3396.865 1048.035 3414 1209.16 ;
      RECT 3386 1048.035 3391.955 1209.16 ;
      RECT 3386 1048.035 3414 1054.07 ;
      RECT 3370.48 1118.44 3383.48 1209.16 ;
      RECT 3378.375 1048.035 3383.48 1209.16 ;
      RECT 3370.48 1048.035 3383.48 1087.87 ;
      RECT 3353.5 1166.44 3366.5 1189.16 ;
      RECT 3364.43 1048.035 3366.5 1189.16 ;
      RECT 3360.475 1053.365 3366.5 1189.16 ;
      RECT 3353.5 1048.035 3355.565 1189.16 ;
      RECT 3353.5 1087.44 3366.5 1150.07 ;
      RECT 3353.5 1053.365 3366.5 1071.07 ;
      RECT 3353.5 1048.035 3358.81 1071.07 ;
      RECT 3353.5 1048.035 3366.5 1049.165 ;
      RECT 3336.52 1166.44 3349.52 1209.16 ;
      RECT 3338.145 1048.035 3349.52 1209.16 ;
      RECT 3336.52 1087.44 3349.52 1150.07 ;
      RECT 3336.52 1048.035 3349.52 1071.07 ;
      RECT 3306 1183.44 3334 1209.16 ;
      RECT 3312.145 1048.035 3328.565 1209.16 ;
      RECT 3306 1070.44 3307.235 1209.16 ;
      RECT 3306 1070.44 3333.235 1167.07 ;
      RECT 3306 1087.44 3334 1150.07 ;
      RECT 3308.365 1048.035 3328.565 1167.07 ;
      RECT 3306 1048.035 3334 1054.07 ;
      RECT 3290.48 1087.44 3303.48 1209.16 ;
      RECT 3290.48 1048.035 3296.835 1209.16 ;
      RECT 3290.48 1048.035 3303.48 1071.07 ;
      RECT 3273.5 1149.44 3286.5 1189.16 ;
      RECT 3284.63 1048.035 3286.5 1189.16 ;
      RECT 3282.865 1053.42 3286.5 1189.16 ;
      RECT 3273.5 1048.035 3275.115 1189.16 ;
      RECT 3273.5 1053.42 3286.5 1118.87 ;
      RECT 3273.5 1048.035 3281.85 1118.87 ;
      RECT 3273.5 1048.035 3286.5 1049.12 ;
      RECT 3256.52 1070.44 3269.52 1209.16 ;
      RECT 3256.865 1048.035 3269.52 1209.16 ;
      RECT 3256.52 1048.035 3269.52 1054.07 ;
      RECT 3226 1118.44 3254 1209.16 ;
      RECT 3238.375 1070.44 3254 1209.16 ;
      RECT 3226 1048.035 3230.625 1209.16 ;
      RECT 3226 1048.035 3251.955 1087.87 ;
      RECT 3226 1048.035 3254 1054.07 ;
      RECT 3210.48 1166.44 3223.48 1209.16 ;
      RECT 3220.475 1053.365 3223.48 1209.16 ;
      RECT 3210.48 1048.035 3215.565 1209.16 ;
      RECT 3210.48 1087.44 3223.48 1150.07 ;
      RECT 3210.48 1053.365 3223.48 1071.07 ;
      RECT 3210.48 1048.035 3218.81 1071.07 ;
      RECT 3210.48 1048.035 3223.48 1049.165 ;
      RECT 3193.5 1166.44 3206.5 1189.16 ;
      RECT 3198.145 1048.035 3206.5 1189.16 ;
      RECT 3197.98 1087.44 3206.5 1189.16 ;
      RECT 3193.5 1087.44 3206.5 1150.07 ;
      RECT 3193.5 1048.035 3206.5 1071.07 ;
      RECT 3176.52 1183.44 3189.52 1209.16 ;
      RECT 3176.52 1048.035 3188.565 1209.16 ;
      RECT 3176.52 1070.44 3189.52 1167.07 ;
      RECT 3176.52 1048.035 3189.52 1054.07 ;
      RECT 3146 1183.44 3174 1209.16 ;
      RECT 3172.145 1048.035 3174 1209.16 ;
      RECT 3146 1087.44 3167.235 1209.16 ;
      RECT 3169.555 1048.035 3174 1167.07 ;
      RECT 3152.55 1070.44 3174 1167.07 ;
      RECT 3146 1048.035 3164.645 1071.07 ;
      RECT 3146 1048.035 3174 1054.07 ;
      RECT 3130.48 1149.44 3143.48 1209.16 ;
      RECT 3142.865 1053.415 3143.48 1209.16 ;
      RECT 3130.48 1048.035 3135.115 1209.16 ;
      RECT 3130.48 1053.415 3143.48 1118.87 ;
      RECT 3130.48 1048.035 3141.85 1118.87 ;
      RECT 3130.48 1048.035 3143.48 1049.12 ;
      RECT 3113.5 1070.44 3126.5 1189.16 ;
      RECT 3116.865 1048.035 3126.5 1189.16 ;
      RECT 3113.5 1048.035 3126.5 1054.07 ;
      RECT 3096.52 1118.44 3109.52 1209.16 ;
      RECT 3098.375 1048.035 3109.52 1209.16 ;
      RECT 3096.52 1048.035 3109.52 1087.87 ;
      RECT 3066 1166.44 3094 1209.16 ;
      RECT 3080.475 1118.44 3094 1209.16 ;
      RECT 3066 1048.035 3075.565 1209.16 ;
      RECT 3066 1087.44 3090.625 1150.07 ;
      RECT 3084.53 1048.035 3094 1087.87 ;
      RECT 3080.475 1053.365 3094 1087.87 ;
      RECT 3066 1053.365 3094 1071.07 ;
      RECT 3066 1048.035 3078.81 1071.07 ;
      RECT 3066 1048.035 3094 1049.165 ;
      RECT 3050.48 1183.44 3063.48 1209.16 ;
      RECT 3058.145 1048.035 3063.48 1209.16 ;
      RECT 3053.475 1166.44 3063.48 1209.16 ;
      RECT 3050.48 1166.44 3063.48 1167.07 ;
      RECT 3050.48 1070.44 3053.235 1167.07 ;
      RECT 3050.48 1087.44 3063.48 1150.07 ;
      RECT 3050.48 1070.44 3063.48 1071.07 ;
      RECT 3053.475 1048.035 3063.48 1071.07 ;
      RECT 3050.48 1048.035 3063.48 1054.07 ;
      RECT 3016.52 1183.44 3029.52 1209.16 ;
      RECT 3016.52 1087.44 3027.235 1209.16 ;
      RECT 3021.75 1070.44 3029.52 1167.07 ;
      RECT 3016.52 1048.035 3024.565 1071.07 ;
      RECT 3016.52 1048.035 3029.52 1054.07 ;
      RECT 2986 1149.44 3014 1209.16 ;
      RECT 3004.63 1048.035 3014 1209.16 ;
      RECT 3002.865 1053.42 3014 1209.16 ;
      RECT 2986 1048.035 2995.115 1209.16 ;
      RECT 2986 1053.42 3014 1118.87 ;
      RECT 2986 1048.035 3001.85 1118.87 ;
      RECT 2986 1048.035 3014 1049.12 ;
      RECT 2970.48 1070.44 2983.48 1209.16 ;
      RECT 2976.865 1048.035 2983.48 1209.16 ;
      RECT 2970.48 1048.035 2971.955 1209.16 ;
      RECT 2970.48 1048.035 2983.48 1054.07 ;
      RECT 2953.5 1118.44 2966.5 1189.16 ;
      RECT 2958.375 1048.035 2966.5 1189.16 ;
      RECT 2953.5 1048.035 2966.5 1087.87 ;
      RECT 2936.52 1166.44 2949.52 1209.16 ;
      RECT 2944.53 1048.035 2949.52 1209.16 ;
      RECT 2940.475 1053.365 2949.52 1209.16 ;
      RECT 2936.52 1087.44 2949.52 1150.07 ;
      RECT 2936.52 1053.365 2949.52 1071.07 ;
      RECT 2936.52 1048.035 2938.81 1071.07 ;
      RECT 2936.52 1048.035 2949.52 1049.375 ;
      RECT 2906 1183.44 2934 1209.16 ;
      RECT 2918.145 1048.035 2934 1209.16 ;
      RECT 2913.475 1166.44 2934 1209.16 ;
      RECT 2906 1048.035 2908.565 1209.16 ;
      RECT 2906 1166.44 2934 1167.07 ;
      RECT 2906 1070.44 2913.235 1167.07 ;
      RECT 2906 1087.44 2934 1150.07 ;
      RECT 2906 1070.44 2934 1071.07 ;
      RECT 2913.475 1048.035 2934 1071.07 ;
      RECT 2906 1048.035 2934 1054.07 ;
      RECT 2890.48 1183.44 2903.48 1209.16 ;
      RECT 2892.145 1048.035 2903.48 1209.16 ;
      RECT 2890.48 1048.035 2903.48 1167.07 ;
      RECT 2873.5 1087.44 2886.5 1189.16 ;
      RECT 2880.13 1070.44 2886.5 1189.16 ;
      RECT 2873.5 1048.035 2883.455 1071.07 ;
      RECT 2873.5 1048.035 2886.5 1054.07 ;
      RECT 2856.52 1149.44 2869.52 1209.16 ;
      RECT 2864.63 1048.035 2869.52 1209.16 ;
      RECT 2862.865 1053.42 2869.52 1209.16 ;
      RECT 2856.52 1053.42 2869.52 1118.87 ;
      RECT 2856.52 1048.035 2861.85 1118.87 ;
      RECT 2856.52 1048.035 2869.52 1049.12 ;
      RECT 2826 1070.44 2854 1209.16 ;
      RECT 2836.865 1048.035 2854 1209.16 ;
      RECT 2826 1048.035 2831.955 1209.16 ;
      RECT 2826 1048.035 2854 1054.07 ;
      RECT 2810.48 1118.44 2823.48 1209.16 ;
      RECT 2818.375 1048.035 2823.48 1209.16 ;
      RECT 2810.48 1048.035 2823.48 1087.87 ;
      RECT 2793.5 1166.44 2806.5 1189.16 ;
      RECT 2804.43 1048.035 2806.5 1189.16 ;
      RECT 2800.475 1053.365 2806.5 1189.16 ;
      RECT 2793.5 1048.035 2795.565 1189.16 ;
      RECT 2793.5 1087.44 2806.5 1150.07 ;
      RECT 2793.5 1053.365 2806.5 1071.07 ;
      RECT 2793.5 1048.035 2798.81 1071.07 ;
      RECT 2793.5 1048.035 2806.5 1049.165 ;
      RECT 2776.52 1166.44 2789.52 1209.16 ;
      RECT 2778.145 1048.035 2789.52 1209.16 ;
      RECT 2776.52 1087.44 2789.52 1150.07 ;
      RECT 2776.52 1048.035 2789.52 1071.07 ;
      RECT 2746 1183.44 2774 1209.16 ;
      RECT 2752.145 1048.035 2768.565 1209.16 ;
      RECT 2746 1070.44 2747.235 1209.16 ;
      RECT 2746 1070.44 2773.235 1167.07 ;
      RECT 2746 1087.44 2774 1150.07 ;
      RECT 2748.365 1048.035 2768.565 1167.07 ;
      RECT 2746 1048.035 2774 1054.07 ;
      RECT 2730.48 1087.44 2743.48 1209.16 ;
      RECT 2730.48 1048.035 2736.835 1209.16 ;
      RECT 2730.48 1048.035 2743.48 1071.07 ;
      RECT 2713.5 1149.44 2726.5 1189.16 ;
      RECT 2724.63 1048.035 2726.5 1189.16 ;
      RECT 2722.865 1053.42 2726.5 1189.16 ;
      RECT 2713.5 1048.035 2715.115 1189.16 ;
      RECT 2713.5 1053.42 2726.5 1118.87 ;
      RECT 2713.5 1048.035 2721.85 1118.87 ;
      RECT 2713.5 1048.035 2726.5 1049.12 ;
      RECT 2696.52 1070.44 2709.52 1209.16 ;
      RECT 2696.865 1048.035 2709.52 1209.16 ;
      RECT 2696.52 1048.035 2709.52 1054.07 ;
      RECT 2666 1118.44 2694 1209.16 ;
      RECT 2678.375 1070.44 2694 1209.16 ;
      RECT 2666 1048.035 2670.625 1209.16 ;
      RECT 2666 1048.035 2691.955 1087.87 ;
      RECT 2666 1048.035 2694 1054.07 ;
      RECT 2650.48 1166.44 2663.48 1209.16 ;
      RECT 2660.475 1053.365 2663.48 1209.16 ;
      RECT 2650.48 1048.035 2655.565 1209.16 ;
      RECT 2650.48 1087.44 2663.48 1150.07 ;
      RECT 2650.48 1053.365 2663.48 1071.07 ;
      RECT 2650.48 1048.035 2658.81 1071.07 ;
      RECT 2650.48 1048.035 2663.48 1049.165 ;
      RECT 2633.5 1166.44 2646.5 1189.16 ;
      RECT 2638.145 1048.035 2646.5 1189.16 ;
      RECT 2637.98 1087.44 2646.5 1189.16 ;
      RECT 2633.5 1087.44 2646.5 1150.07 ;
      RECT 2633.5 1048.035 2646.5 1071.07 ;
      RECT 2616.52 1183.44 2629.52 1209.16 ;
      RECT 2616.52 1048.035 2628.565 1209.16 ;
      RECT 2616.52 1070.44 2629.52 1167.07 ;
      RECT 2616.52 1048.035 2629.52 1054.07 ;
      RECT 2586 1183.44 2614 1209.16 ;
      RECT 2612.145 1048.035 2614 1209.16 ;
      RECT 2586 1087.44 2607.235 1209.16 ;
      RECT 2609.555 1048.035 2614 1167.07 ;
      RECT 2592.55 1070.44 2614 1167.07 ;
      RECT 2586 1048.035 2604.645 1071.07 ;
      RECT 2586 1048.035 2614 1054.07 ;
      RECT 2570.48 1149.44 2583.48 1209.16 ;
      RECT 2582.865 1053.415 2583.48 1209.16 ;
      RECT 2570.48 1048.035 2575.115 1209.16 ;
      RECT 2570.48 1053.415 2583.48 1118.87 ;
      RECT 2570.48 1048.035 2581.85 1118.87 ;
      RECT 2570.48 1048.035 2583.48 1049.12 ;
      RECT 2553.5 1070.44 2566.5 1189.16 ;
      RECT 2556.865 1048.035 2566.5 1189.16 ;
      RECT 2553.5 1048.035 2566.5 1054.07 ;
      RECT 2536.52 1118.44 2549.52 1209.16 ;
      RECT 2538.375 1048.035 2549.52 1209.16 ;
      RECT 2536.52 1048.035 2549.52 1087.87 ;
      RECT 2506 1166.44 2534 1209.16 ;
      RECT 2520.475 1118.44 2534 1209.16 ;
      RECT 2506 1048.035 2515.565 1209.16 ;
      RECT 2506 1087.44 2530.625 1150.07 ;
      RECT 2524.53 1048.035 2534 1087.87 ;
      RECT 2520.475 1053.365 2534 1087.87 ;
      RECT 2506 1053.365 2534 1071.07 ;
      RECT 2506 1048.035 2518.81 1071.07 ;
      RECT 2506 1048.035 2534 1049.165 ;
      RECT 2490.48 1183.44 2503.48 1209.16 ;
      RECT 2498.145 1048.035 2503.48 1209.16 ;
      RECT 2493.475 1166.44 2503.48 1209.16 ;
      RECT 2490.48 1166.44 2503.48 1167.07 ;
      RECT 2490.48 1070.44 2493.235 1167.07 ;
      RECT 2490.48 1087.44 2503.48 1150.07 ;
      RECT 2490.48 1070.44 2503.48 1071.07 ;
      RECT 2493.475 1048.035 2503.48 1071.07 ;
      RECT 2490.48 1048.035 2503.48 1054.07 ;
      RECT 2456.52 1183.44 2469.52 1209.16 ;
      RECT 2456.52 1087.44 2467.235 1209.16 ;
      RECT 2461.75 1070.44 2469.52 1167.07 ;
      RECT 2456.52 1048.035 2464.565 1071.07 ;
      RECT 2456.52 1048.035 2469.52 1054.07 ;
      RECT 2426 1149.44 2454 1209.16 ;
      RECT 2444.63 1048.035 2454 1209.16 ;
      RECT 2442.865 1053.42 2454 1209.16 ;
      RECT 2426 1048.035 2435.115 1209.16 ;
      RECT 2426 1053.42 2454 1118.87 ;
      RECT 2426 1048.035 2441.85 1118.87 ;
      RECT 2426 1048.035 2454 1049.12 ;
      RECT 2410.48 1070.44 2423.48 1209.16 ;
      RECT 2416.865 1048.035 2423.48 1209.16 ;
      RECT 2410.48 1048.035 2411.955 1209.16 ;
      RECT 2410.48 1048.035 2423.48 1054.07 ;
      RECT 2393.5 1118.44 2406.5 1189.16 ;
      RECT 2398.375 1048.035 2406.5 1189.16 ;
      RECT 2393.5 1048.035 2406.5 1087.87 ;
      RECT 2376.52 1166.44 2389.52 1209.16 ;
      RECT 2384.53 1048.035 2389.52 1209.16 ;
      RECT 2380.475 1053.365 2389.52 1209.16 ;
      RECT 2376.52 1087.44 2389.52 1150.07 ;
      RECT 2376.52 1053.365 2389.52 1071.07 ;
      RECT 2376.52 1048.035 2378.81 1071.07 ;
      RECT 2376.52 1048.035 2389.52 1049.375 ;
      RECT 2346 1183.44 2374 1209.16 ;
      RECT 2358.145 1048.035 2374 1209.16 ;
      RECT 2353.475 1166.44 2374 1209.16 ;
      RECT 2346 1048.035 2348.565 1209.16 ;
      RECT 2346 1166.44 2374 1167.07 ;
      RECT 2346 1070.44 2353.235 1167.07 ;
      RECT 2346 1087.44 2374 1150.07 ;
      RECT 2346 1070.44 2374 1071.07 ;
      RECT 2353.475 1048.035 2374 1071.07 ;
      RECT 2346 1048.035 2374 1054.07 ;
      RECT 2330.48 1183.44 2343.48 1209.16 ;
      RECT 2332.145 1048.035 2343.48 1209.16 ;
      RECT 2330.48 1048.035 2343.48 1167.07 ;
      RECT 2313.5 1087.44 2326.5 1189.16 ;
      RECT 2320.13 1070.44 2326.5 1189.16 ;
      RECT 2313.5 1048.035 2323.455 1071.07 ;
      RECT 2313.5 1048.035 2326.5 1054.07 ;
      RECT 2296.52 1149.44 2309.52 1209.16 ;
      RECT 2304.63 1048.035 2309.52 1209.16 ;
      RECT 2302.865 1053.42 2309.52 1209.16 ;
      RECT 2296.52 1053.42 2309.52 1118.87 ;
      RECT 2296.52 1048.035 2301.85 1118.87 ;
      RECT 2296.52 1048.035 2309.52 1049.12 ;
      RECT 2266 1070.44 2294 1209.16 ;
      RECT 2276.865 1048.035 2294 1209.16 ;
      RECT 2266 1048.035 2271.955 1209.16 ;
      RECT 2266 1048.035 2294 1054.07 ;
      RECT 2250.48 1118.44 2263.48 1209.16 ;
      RECT 2258.375 1048.035 2263.48 1209.16 ;
      RECT 2250.48 1048.035 2263.48 1087.87 ;
      RECT 2233.5 1166.44 2246.5 1189.16 ;
      RECT 2244.43 1048.035 2246.5 1189.16 ;
      RECT 2240.475 1053.365 2246.5 1189.16 ;
      RECT 2233.5 1048.035 2235.565 1189.16 ;
      RECT 2233.5 1087.44 2246.5 1150.07 ;
      RECT 2233.5 1053.365 2246.5 1071.07 ;
      RECT 2233.5 1048.035 2238.81 1071.07 ;
      RECT 2233.5 1048.035 2246.5 1049.165 ;
      RECT 2216.52 1166.44 2229.52 1209.16 ;
      RECT 2218.145 1048.035 2229.52 1209.16 ;
      RECT 2216.52 1087.44 2229.52 1150.07 ;
      RECT 2216.52 1048.035 2229.52 1071.07 ;
      RECT 2186 1183.44 2214 1209.16 ;
      RECT 2192.145 1048.035 2208.565 1209.16 ;
      RECT 2186 1070.44 2187.235 1209.16 ;
      RECT 2186 1070.44 2213.235 1167.07 ;
      RECT 2186 1087.44 2214 1150.07 ;
      RECT 2188.365 1048.035 2208.565 1167.07 ;
      RECT 2186 1048.035 2214 1054.07 ;
      RECT 2170.48 1087.44 2183.48 1209.16 ;
      RECT 2170.48 1048.035 2176.835 1209.16 ;
      RECT 2170.48 1048.035 2183.48 1071.07 ;
      RECT 2153.5 1149.44 2166.5 1189.16 ;
      RECT 2164.63 1048.035 2166.5 1189.16 ;
      RECT 2162.865 1053.42 2166.5 1189.16 ;
      RECT 2153.5 1048.035 2155.115 1189.16 ;
      RECT 2153.5 1053.42 2166.5 1118.87 ;
      RECT 2153.5 1048.035 2161.85 1118.87 ;
      RECT 2153.5 1048.035 2166.5 1049.12 ;
      RECT 2136.52 1070.44 2149.52 1209.16 ;
      RECT 2136.865 1048.035 2149.52 1209.16 ;
      RECT 2136.52 1048.035 2149.52 1054.07 ;
      RECT 2106 1118.44 2134 1209.16 ;
      RECT 2118.375 1070.44 2134 1209.16 ;
      RECT 2106 1048.035 2110.625 1209.16 ;
      RECT 2106 1048.035 2131.955 1087.87 ;
      RECT 2106 1048.035 2134 1054.07 ;
      RECT 2090.48 1166.44 2103.48 1209.16 ;
      RECT 2100.475 1053.365 2103.48 1209.16 ;
      RECT 2090.48 1048.035 2095.565 1209.16 ;
      RECT 2090.48 1087.44 2103.48 1150.07 ;
      RECT 2090.48 1053.365 2103.48 1071.07 ;
      RECT 2090.48 1048.035 2098.81 1071.07 ;
      RECT 2090.48 1048.035 2103.48 1049.165 ;
      RECT 2073.5 1166.44 2086.5 1189.16 ;
      RECT 2078.145 1048.035 2086.5 1189.16 ;
      RECT 2077.98 1087.44 2086.5 1189.16 ;
      RECT 2073.5 1087.44 2086.5 1150.07 ;
      RECT 2073.5 1048.035 2086.5 1071.07 ;
      RECT 2056.52 1183.44 2069.52 1209.16 ;
      RECT 2056.52 1048.035 2068.565 1209.16 ;
      RECT 2056.52 1070.44 2069.52 1167.07 ;
      RECT 2056.52 1048.035 2069.52 1054.07 ;
      RECT 2026 1183.44 2054 1209.16 ;
      RECT 2052.145 1048.035 2054 1209.16 ;
      RECT 2026 1087.44 2047.235 1209.16 ;
      RECT 2049.555 1048.035 2054 1167.07 ;
      RECT 2032.55 1070.44 2054 1167.07 ;
      RECT 2026 1048.035 2044.645 1071.07 ;
      RECT 2026 1048.035 2054 1054.07 ;
      RECT 2010.48 1149.44 2023.48 1209.16 ;
      RECT 2022.865 1053.415 2023.48 1209.16 ;
      RECT 2010.48 1048.035 2015.115 1209.16 ;
      RECT 2010.48 1053.415 2023.48 1118.87 ;
      RECT 2010.48 1048.035 2021.85 1118.87 ;
      RECT 2010.48 1048.035 2023.48 1049.12 ;
      RECT 1993.5 1070.44 2006.5 1189.16 ;
      RECT 1996.865 1048.035 2006.5 1189.16 ;
      RECT 1993.5 1048.035 2006.5 1054.07 ;
      RECT 1976.52 1118.44 1989.52 1209.16 ;
      RECT 1978.375 1048.035 1989.52 1209.16 ;
      RECT 1976.52 1048.035 1989.52 1087.87 ;
      RECT 1946 1166.44 1974 1209.16 ;
      RECT 1960.475 1118.44 1974 1209.16 ;
      RECT 1946 1048.035 1955.565 1209.16 ;
      RECT 1946 1087.44 1970.625 1150.07 ;
      RECT 1964.53 1048.035 1974 1087.87 ;
      RECT 1960.475 1053.365 1974 1087.87 ;
      RECT 1946 1053.365 1974 1071.07 ;
      RECT 1946 1048.035 1958.81 1071.07 ;
      RECT 1946 1048.035 1974 1049.165 ;
      RECT 1930.48 1183.44 1943.48 1209.16 ;
      RECT 1938.145 1048.035 1943.48 1209.16 ;
      RECT 1933.475 1166.44 1943.48 1209.16 ;
      RECT 1930.48 1166.44 1943.48 1167.07 ;
      RECT 1930.48 1070.44 1933.235 1167.07 ;
      RECT 1930.48 1087.44 1943.48 1150.07 ;
      RECT 1930.48 1070.44 1943.48 1071.07 ;
      RECT 1933.475 1048.035 1943.48 1071.07 ;
      RECT 1930.48 1048.035 1943.48 1054.07 ;
      RECT 1896.52 1183.44 1909.52 1209.16 ;
      RECT 1896.52 1087.44 1907.235 1209.16 ;
      RECT 1901.75 1070.44 1909.52 1167.07 ;
      RECT 1896.52 1048.035 1904.565 1071.07 ;
      RECT 1896.52 1048.035 1909.52 1054.07 ;
      RECT 1866 1149.44 1894 1209.16 ;
      RECT 1884.63 1048.035 1894 1209.16 ;
      RECT 1882.865 1053.42 1894 1209.16 ;
      RECT 1866 1048.035 1875.115 1209.16 ;
      RECT 1866 1053.42 1894 1118.87 ;
      RECT 1866 1048.035 1881.85 1118.87 ;
      RECT 1866 1048.035 1894 1049.12 ;
      RECT 1850.48 1070.44 1863.48 1209.16 ;
      RECT 1856.865 1048.035 1863.48 1209.16 ;
      RECT 1850.48 1048.035 1851.955 1209.16 ;
      RECT 1850.48 1048.035 1863.48 1054.07 ;
      RECT 1833.5 1118.44 1846.5 1189.16 ;
      RECT 1838.375 1048.035 1846.5 1189.16 ;
      RECT 1833.5 1048.035 1846.5 1087.87 ;
      RECT 1816.52 1166.44 1829.52 1209.16 ;
      RECT 1824.53 1048.035 1829.52 1209.16 ;
      RECT 1820.475 1053.365 1829.52 1209.16 ;
      RECT 1816.52 1087.44 1829.52 1150.07 ;
      RECT 1816.52 1053.365 1829.52 1071.07 ;
      RECT 1816.52 1048.035 1818.81 1071.07 ;
      RECT 1816.52 1048.035 1829.52 1049.375 ;
      RECT 1786 1183.44 1814 1209.16 ;
      RECT 1798.145 1048.035 1814 1209.16 ;
      RECT 1793.475 1166.44 1814 1209.16 ;
      RECT 1786 1048.035 1788.565 1209.16 ;
      RECT 1786 1166.44 1814 1167.07 ;
      RECT 1786 1070.44 1793.235 1167.07 ;
      RECT 1786 1087.44 1814 1150.07 ;
      RECT 1786 1070.44 1814 1071.07 ;
      RECT 1793.475 1048.035 1814 1071.07 ;
      RECT 1786 1048.035 1814 1054.07 ;
      RECT 1770.48 1183.44 1783.48 1209.16 ;
      RECT 1772.145 1048.035 1783.48 1209.16 ;
      RECT 1770.48 1048.035 1783.48 1167.07 ;
      RECT 1753.5 1087.44 1766.5 1189.16 ;
      RECT 1760.13 1070.44 1766.5 1189.16 ;
      RECT 1753.5 1048.035 1763.455 1071.07 ;
      RECT 1753.5 1048.035 1766.5 1054.07 ;
      RECT 1736.52 1149.44 1749.52 1209.16 ;
      RECT 1744.63 1048.035 1749.52 1209.16 ;
      RECT 1742.865 1053.42 1749.52 1209.16 ;
      RECT 1736.52 1053.42 1749.52 1118.87 ;
      RECT 1736.52 1048.035 1741.85 1118.87 ;
      RECT 1736.52 1048.035 1749.52 1049.12 ;
      RECT 1706 1070.44 1734 1209.16 ;
      RECT 1716.865 1048.035 1734 1209.16 ;
      RECT 1706 1048.035 1711.955 1209.16 ;
      RECT 1706 1048.035 1734 1054.07 ;
      RECT 1690.48 1118.44 1703.48 1209.16 ;
      RECT 1698.375 1048.035 1703.48 1209.16 ;
      RECT 1690.48 1048.035 1703.48 1087.87 ;
      RECT 1673.5 1166.44 1686.5 1189.16 ;
      RECT 1684.43 1048.035 1686.5 1189.16 ;
      RECT 1680.475 1053.365 1686.5 1189.16 ;
      RECT 1673.5 1048.035 1675.565 1189.16 ;
      RECT 1673.5 1087.44 1686.5 1150.07 ;
      RECT 1673.5 1053.365 1686.5 1071.07 ;
      RECT 1673.5 1048.035 1678.81 1071.07 ;
      RECT 1673.5 1048.035 1686.5 1049.165 ;
      RECT 1656.52 1166.44 1669.52 1209.16 ;
      RECT 1658.145 1048.035 1669.52 1209.16 ;
      RECT 1656.52 1087.44 1669.52 1150.07 ;
      RECT 1656.52 1048.035 1669.52 1071.07 ;
      RECT 1626 1183.44 1654 1209.16 ;
      RECT 1632.145 1048.035 1648.565 1209.16 ;
      RECT 1626 1070.44 1627.235 1209.16 ;
      RECT 1626 1070.44 1653.235 1167.07 ;
      RECT 1626 1087.44 1654 1150.07 ;
      RECT 1628.365 1048.035 1648.565 1167.07 ;
      RECT 1626 1048.035 1654 1054.07 ;
      RECT 1610.48 1087.44 1623.48 1209.16 ;
      RECT 1610.48 1048.035 1616.835 1209.16 ;
      RECT 1610.48 1048.035 1623.48 1071.07 ;
      RECT 1593.5 1149.44 1606.5 1189.16 ;
      RECT 1604.63 1048.035 1606.5 1189.16 ;
      RECT 1602.865 1053.42 1606.5 1189.16 ;
      RECT 1593.5 1048.035 1595.115 1189.16 ;
      RECT 1593.5 1053.42 1606.5 1118.87 ;
      RECT 1593.5 1048.035 1601.85 1118.87 ;
      RECT 1593.5 1048.035 1606.5 1049.12 ;
      RECT 1576.52 1070.44 1589.52 1209.16 ;
      RECT 1576.865 1048.035 1589.52 1209.16 ;
      RECT 1576.52 1048.035 1589.52 1054.07 ;
      RECT 1546 1118.44 1574 1209.16 ;
      RECT 1558.375 1070.44 1574 1209.16 ;
      RECT 1546 1048.035 1550.625 1209.16 ;
      RECT 1546 1048.035 1571.955 1087.87 ;
      RECT 1546 1048.035 1574 1054.07 ;
      RECT 1530.48 1166.44 1543.48 1209.16 ;
      RECT 1540.475 1053.365 1543.48 1209.16 ;
      RECT 1530.48 1048.035 1535.565 1209.16 ;
      RECT 1530.48 1087.44 1543.48 1150.07 ;
      RECT 1530.48 1053.365 1543.48 1071.07 ;
      RECT 1530.48 1048.035 1538.81 1071.07 ;
      RECT 1530.48 1048.035 1543.48 1049.165 ;
      RECT 1513.5 1166.44 1526.5 1189.16 ;
      RECT 1518.145 1048.035 1526.5 1189.16 ;
      RECT 1517.98 1087.44 1526.5 1189.16 ;
      RECT 1513.5 1087.44 1526.5 1150.07 ;
      RECT 1513.5 1048.035 1526.5 1071.07 ;
      RECT 1496.52 1183.44 1509.52 1209.16 ;
      RECT 1496.52 1048.035 1508.565 1209.16 ;
      RECT 1496.52 1070.44 1509.52 1167.07 ;
      RECT 1496.52 1048.035 1509.52 1054.07 ;
      RECT 1466 1183.44 1494 1209.16 ;
      RECT 1492.145 1048.035 1494 1209.16 ;
      RECT 1466 1087.44 1487.235 1209.16 ;
      RECT 1489.555 1048.035 1494 1167.07 ;
      RECT 1472.55 1070.44 1494 1167.07 ;
      RECT 1466 1048.035 1484.645 1071.07 ;
      RECT 1466 1048.035 1494 1054.07 ;
      RECT 1450.48 1149.44 1463.48 1209.16 ;
      RECT 1462.865 1053.415 1463.48 1209.16 ;
      RECT 1450.48 1048.035 1455.115 1209.16 ;
      RECT 1450.48 1053.415 1463.48 1118.87 ;
      RECT 1450.48 1048.035 1461.85 1118.87 ;
      RECT 1450.48 1048.035 1463.48 1049.12 ;
      RECT 1433.5 1070.44 1446.5 1189.16 ;
      RECT 1436.865 1048.035 1446.5 1189.16 ;
      RECT 1433.5 1048.035 1446.5 1054.07 ;
      RECT 1416.52 1118.44 1429.52 1209.16 ;
      RECT 1418.375 1048.035 1429.52 1209.16 ;
      RECT 1416.52 1048.035 1429.52 1087.87 ;
      RECT 1386 1166.44 1414 1209.16 ;
      RECT 1400.475 1118.44 1414 1209.16 ;
      RECT 1386 1048.035 1395.565 1209.16 ;
      RECT 1386 1087.44 1410.625 1150.07 ;
      RECT 1404.53 1048.035 1414 1087.87 ;
      RECT 1400.475 1053.365 1414 1087.87 ;
      RECT 1386 1053.365 1414 1071.07 ;
      RECT 1386 1048.035 1398.81 1071.07 ;
      RECT 1386 1048.035 1414 1049.165 ;
      RECT 1370.48 1183.44 1383.48 1209.16 ;
      RECT 1378.145 1048.035 1383.48 1209.16 ;
      RECT 1373.475 1166.44 1383.48 1209.16 ;
      RECT 1370.48 1166.44 1383.48 1167.07 ;
      RECT 1370.48 1070.44 1373.235 1167.07 ;
      RECT 1370.48 1087.44 1383.48 1150.07 ;
      RECT 1370.48 1070.44 1383.48 1071.07 ;
      RECT 1373.475 1048.035 1383.48 1071.07 ;
      RECT 1370.48 1048.035 1383.48 1054.07 ;
      RECT 1336.52 1183.44 1349.52 1209.16 ;
      RECT 1336.52 1087.44 1347.235 1209.16 ;
      RECT 1341.75 1070.44 1349.52 1167.07 ;
      RECT 1336.52 1048.035 1344.565 1071.07 ;
      RECT 1336.52 1048.035 1349.52 1054.07 ;
      RECT 1306 1149.44 1334 1209.16 ;
      RECT 1324.63 1048.035 1334 1209.16 ;
      RECT 1322.865 1053.42 1334 1209.16 ;
      RECT 1306 1048.035 1315.115 1209.16 ;
      RECT 1306 1053.42 1334 1118.87 ;
      RECT 1306 1048.035 1321.85 1118.87 ;
      RECT 1306 1048.035 1334 1049.12 ;
      RECT 1290.48 1070.44 1303.48 1209.16 ;
      RECT 1296.865 1048.035 1303.48 1209.16 ;
      RECT 1290.48 1048.035 1291.955 1209.16 ;
      RECT 1290.48 1048.035 1303.48 1054.07 ;
      RECT 1273.5 1118.44 1286.5 1189.16 ;
      RECT 1278.375 1048.035 1286.5 1189.16 ;
      RECT 1273.5 1048.035 1286.5 1087.87 ;
      RECT 1256.52 1166.44 1269.52 1209.16 ;
      RECT 1264.53 1048.035 1269.52 1209.16 ;
      RECT 1260.475 1053.365 1269.52 1209.16 ;
      RECT 1256.52 1087.44 1269.52 1150.07 ;
      RECT 1256.52 1053.365 1269.52 1071.07 ;
      RECT 1256.52 1048.035 1258.81 1071.07 ;
      RECT 1256.52 1048.035 1269.52 1049.375 ;
      RECT 1226 1183.44 1254 1209.16 ;
      RECT 1238.145 1048.035 1254 1209.16 ;
      RECT 1233.475 1166.44 1254 1209.16 ;
      RECT 1226 1048.035 1228.565 1209.16 ;
      RECT 1226 1166.44 1254 1167.07 ;
      RECT 1226 1070.44 1233.235 1167.07 ;
      RECT 1226 1087.44 1254 1150.07 ;
      RECT 1226 1070.44 1254 1071.07 ;
      RECT 1233.475 1048.035 1254 1071.07 ;
      RECT 1226 1048.035 1254 1054.07 ;
      RECT 1210.48 1183.44 1223.48 1209.16 ;
      RECT 1212.145 1048.035 1223.48 1209.16 ;
      RECT 1210.48 1048.035 1223.48 1167.07 ;
      RECT 1193.5 1087.44 1206.5 1189.16 ;
      RECT 1200.13 1070.44 1206.5 1189.16 ;
      RECT 1193.5 1048.035 1203.455 1071.07 ;
      RECT 1193.5 1048.035 1206.5 1054.07 ;
      RECT 1176.52 1149.44 1189.52 1209.16 ;
      RECT 1184.63 1048.035 1189.52 1209.16 ;
      RECT 1182.865 1053.42 1189.52 1209.16 ;
      RECT 1176.52 1053.42 1189.52 1118.87 ;
      RECT 1176.52 1048.035 1181.85 1118.87 ;
      RECT 1176.52 1048.035 1189.52 1049.12 ;
      RECT 1146 1070.44 1174 1209.16 ;
      RECT 1156.865 1048.035 1174 1209.16 ;
      RECT 1146 1048.035 1151.955 1209.16 ;
      RECT 1146 1048.035 1174 1054.07 ;
      RECT 1130.48 1118.44 1143.48 1209.16 ;
      RECT 1138.375 1048.035 1143.48 1209.16 ;
      RECT 1130.48 1048.035 1143.48 1087.87 ;
      RECT 992.1 1116.585 999.1 1117.785 ;
      RECT 992.1 1116.79 1001.84 1117.59 ;
      RECT 992.1 1118.985 999.1 1120.185 ;
      RECT 992.1 1119.19 1001.84 1119.99 ;
      RECT 992.1 1121.385 999.1 1122.585 ;
      RECT 992.1 1121.59 1001.84 1122.39 ;
      RECT 992.1 1123.785 999.1 1124.985 ;
      RECT 992.1 1123.99 1001.84 1124.79 ;
      RECT 992.1 1126.185 999.1 1127.385 ;
      RECT 992.1 1126.39 1001.84 1127.19 ;
      RECT 19049.325 1053.685 19168.28 1054.485 ;
      RECT 19049.325 1055.685 19167.9 1056.485 ;
      RECT 19083.24 1088.01 19167.9 1088.81 ;
      RECT 19158.1 1364.41 19167.81 1365.5 ;
      RECT 19158.1 1367.39 19167.81 1368.48 ;
      RECT 19049.325 1051.685 19165.7 1052.485 ;
      RECT 18713.5 1048.035 18726.5 1189.16 ;
      RECT 18153.5 1048.035 18166.5 1189.16 ;
      RECT 17593.5 1048.035 17606.5 1189.16 ;
      RECT 17033.5 1048.035 17046.5 1189.16 ;
      RECT 16473.5 1048.035 16486.5 1189.16 ;
      RECT 15913.5 1048.035 15926.5 1189.16 ;
      RECT 15353.5 1048.035 15366.5 1189.16 ;
      RECT 14793.5 1048.035 14806.5 1189.16 ;
      RECT 14233.5 1048.035 14246.5 1189.16 ;
      RECT 13673.5 1048.035 13686.5 1189.16 ;
      RECT 13113.5 1048.035 13126.5 1189.16 ;
      RECT 12553.5 1048.035 12566.5 1189.16 ;
      RECT 11993.5 1048.035 12006.5 1189.16 ;
      RECT 11433.5 1048.035 11446.5 1189.16 ;
      RECT 10873.5 1048.035 10886.5 1189.16 ;
      RECT 10313.5 1048.035 10326.5 1189.16 ;
      RECT 9753.5 1048.035 9766.5 1189.16 ;
      RECT 9193.5 1048.035 9206.5 1189.16 ;
      RECT 8633.5 1048.035 8646.5 1189.16 ;
      RECT 8073.5 1048.035 8086.5 1189.16 ;
      RECT 7513.5 1048.035 7526.5 1189.16 ;
      RECT 6953.5 1048.035 6966.5 1189.16 ;
      RECT 6393.5 1048.035 6406.5 1189.16 ;
      RECT 5833.5 1048.035 5846.5 1189.16 ;
      RECT 5273.5 1048.035 5286.5 1189.16 ;
      RECT 4713.5 1048.035 4726.5 1189.16 ;
      RECT 4153.5 1048.035 4166.5 1189.16 ;
      RECT 3593.5 1048.035 3606.5 1189.16 ;
      RECT 3033.5 1048.035 3046.5 1189.16 ;
      RECT 2473.5 1048.035 2486.5 1189.16 ;
      RECT 1913.5 1048.035 1926.5 1189.16 ;
      RECT 1353.5 1048.035 1366.5 1189.16 ;
      RECT 994.79 1053.81 1118.225 1054.61 ;
      RECT 991.74 1055.81 1118.225 1056.61 ;
      RECT 992.1 1057.81 1118.225 1058.61 ;
      RECT 992.1 1090.38 1013.415 1091.18 ;
      RECT 992.1 1087.58 1011.415 1088.38 ;
    LAYER M5 SPACING 0.28 ;
      RECT 998.1 1047.905 19161.9 10000 ;
      RECT 19046.97 1046.435 19161.9 10000 ;
      RECT 19029.99 1047.855 19033.03 10000 ;
      RECT 19014.47 1046.435 19016.05 10000 ;
      RECT 18983.95 1046.435 18985.53 10000 ;
      RECT 18966.97 1046.435 18970.01 10000 ;
      RECT 18949.99 1047.855 18953.03 10000 ;
      RECT 18934.47 1046.435 18936.05 10000 ;
      RECT 18903.95 1046.435 18905.53 10000 ;
      RECT 18886.97 1047.855 18890.01 10000 ;
      RECT 18869.99 1046.435 18873.03 10000 ;
      RECT 18854.47 1047.855 18856.05 10000 ;
      RECT 18823.95 1046.435 18825.53 10000 ;
      RECT 18806.97 1047.855 18810.01 10000 ;
      RECT 18789.99 1047.855 18793.03 10000 ;
      RECT 18792.405 1046.435 18793.03 10000 ;
      RECT 18774.47 1046.435 18776.05 10000 ;
      RECT 18743.95 1047.855 18745.53 10000 ;
      RECT 18726.97 1046.435 18730.01 10000 ;
      RECT 18709.99 1046.435 18713.03 10000 ;
      RECT 18694.47 1046.435 18696.05 10000 ;
      RECT 18663.95 1047.855 18665.53 10000 ;
      RECT 18646.97 1047.855 18650.01 10000 ;
      RECT 18629.99 1046.435 18633.03 10000 ;
      RECT 18614.47 1046.435 18616.05 10000 ;
      RECT 18583.95 1047.855 18585.53 10000 ;
      RECT 18566.97 1046.435 18570.01 10000 ;
      RECT 18549.99 1046.435 18553.03 10000 ;
      RECT 18534.47 1046.435 18536.05 10000 ;
      RECT 18503.95 1047.855 18505.53 10000 ;
      RECT 18486.97 1046.435 18490.01 10000 ;
      RECT 18469.99 1047.855 18473.03 10000 ;
      RECT 18472.645 1046.435 18473.03 10000 ;
      RECT 18454.47 1046.435 18456.05 10000 ;
      RECT 18423.95 1046.435 18425.53 10000 ;
      RECT 18406.97 1046.435 18410.01 10000 ;
      RECT 18389.99 1047.855 18393.03 10000 ;
      RECT 18374.47 1046.435 18376.05 10000 ;
      RECT 18343.95 1046.435 18345.53 10000 ;
      RECT 18326.97 1047.855 18330.01 10000 ;
      RECT 18309.99 1046.435 18313.03 10000 ;
      RECT 18294.47 1047.855 18296.05 10000 ;
      RECT 18263.95 1046.435 18265.53 10000 ;
      RECT 18246.97 1047.855 18250.01 10000 ;
      RECT 18229.99 1047.855 18233.03 10000 ;
      RECT 18232.405 1046.435 18233.03 10000 ;
      RECT 18214.47 1046.435 18216.05 10000 ;
      RECT 18183.95 1047.855 18185.53 10000 ;
      RECT 18166.97 1046.435 18170.01 10000 ;
      RECT 18149.99 1046.435 18153.03 10000 ;
      RECT 18134.47 1046.435 18136.05 10000 ;
      RECT 18103.95 1047.855 18105.53 10000 ;
      RECT 18086.97 1047.855 18090.01 10000 ;
      RECT 18069.99 1046.435 18073.03 10000 ;
      RECT 18054.47 1046.435 18056.05 10000 ;
      RECT 18023.95 1047.855 18025.53 10000 ;
      RECT 18006.97 1046.435 18010.01 10000 ;
      RECT 17989.99 1046.435 17993.03 10000 ;
      RECT 17974.47 1046.435 17976.05 10000 ;
      RECT 17943.95 1047.855 17945.53 10000 ;
      RECT 17926.97 1046.435 17930.01 10000 ;
      RECT 17909.99 1047.855 17913.03 10000 ;
      RECT 17912.645 1046.435 17913.03 10000 ;
      RECT 17894.47 1046.435 17896.05 10000 ;
      RECT 17863.95 1046.435 17865.53 10000 ;
      RECT 17846.97 1046.435 17850.01 10000 ;
      RECT 17829.99 1047.855 17833.03 10000 ;
      RECT 17814.47 1046.435 17816.05 10000 ;
      RECT 17783.95 1046.435 17785.53 10000 ;
      RECT 17766.97 1047.855 17770.01 10000 ;
      RECT 17749.99 1046.435 17753.03 10000 ;
      RECT 17734.47 1047.855 17736.05 10000 ;
      RECT 17703.95 1046.435 17705.53 10000 ;
      RECT 17686.97 1047.855 17690.01 10000 ;
      RECT 17669.99 1047.855 17673.03 10000 ;
      RECT 17672.405 1046.435 17673.03 10000 ;
      RECT 17654.47 1046.435 17656.05 10000 ;
      RECT 17623.95 1047.855 17625.53 10000 ;
      RECT 17606.97 1046.435 17610.01 10000 ;
      RECT 17589.99 1046.435 17593.03 10000 ;
      RECT 17574.47 1046.435 17576.05 10000 ;
      RECT 17543.95 1047.855 17545.53 10000 ;
      RECT 17526.97 1047.855 17530.01 10000 ;
      RECT 17509.99 1046.435 17513.03 10000 ;
      RECT 17494.47 1046.435 17496.05 10000 ;
      RECT 17463.95 1047.855 17465.53 10000 ;
      RECT 17446.97 1046.435 17450.01 10000 ;
      RECT 17429.99 1046.435 17433.03 10000 ;
      RECT 17414.47 1046.435 17416.05 10000 ;
      RECT 17383.95 1047.855 17385.53 10000 ;
      RECT 17366.97 1046.435 17370.01 10000 ;
      RECT 17349.99 1047.855 17353.03 10000 ;
      RECT 17352.645 1046.435 17353.03 10000 ;
      RECT 17334.47 1046.435 17336.05 10000 ;
      RECT 17303.95 1046.435 17305.53 10000 ;
      RECT 17286.97 1046.435 17290.01 10000 ;
      RECT 17269.99 1047.855 17273.03 10000 ;
      RECT 17254.47 1046.435 17256.05 10000 ;
      RECT 17223.95 1046.435 17225.53 10000 ;
      RECT 17206.97 1047.855 17210.01 10000 ;
      RECT 17189.99 1046.435 17193.03 10000 ;
      RECT 17174.47 1047.855 17176.05 10000 ;
      RECT 17143.95 1046.435 17145.53 10000 ;
      RECT 17126.97 1047.855 17130.01 10000 ;
      RECT 17109.99 1047.855 17113.03 10000 ;
      RECT 17112.405 1046.435 17113.03 10000 ;
      RECT 17094.47 1046.435 17096.05 10000 ;
      RECT 17063.95 1047.855 17065.53 10000 ;
      RECT 17046.97 1046.435 17050.01 10000 ;
      RECT 17029.99 1046.435 17033.03 10000 ;
      RECT 17014.47 1046.435 17016.05 10000 ;
      RECT 16983.95 1047.855 16985.53 10000 ;
      RECT 16966.97 1047.855 16970.01 10000 ;
      RECT 16949.99 1046.435 16953.03 10000 ;
      RECT 16934.47 1046.435 16936.05 10000 ;
      RECT 16903.95 1047.855 16905.53 10000 ;
      RECT 16886.97 1046.435 16890.01 10000 ;
      RECT 16869.99 1046.435 16873.03 10000 ;
      RECT 16854.47 1046.435 16856.05 10000 ;
      RECT 16823.95 1047.855 16825.53 10000 ;
      RECT 16806.97 1046.435 16810.01 10000 ;
      RECT 16789.99 1047.855 16793.03 10000 ;
      RECT 16792.645 1046.435 16793.03 10000 ;
      RECT 16774.47 1046.435 16776.05 10000 ;
      RECT 16743.95 1046.435 16745.53 10000 ;
      RECT 16726.97 1046.435 16730.01 10000 ;
      RECT 16709.99 1047.855 16713.03 10000 ;
      RECT 16694.47 1046.435 16696.05 10000 ;
      RECT 16663.95 1046.435 16665.53 10000 ;
      RECT 16646.97 1047.855 16650.01 10000 ;
      RECT 16629.99 1046.435 16633.03 10000 ;
      RECT 16614.47 1047.855 16616.05 10000 ;
      RECT 16583.95 1046.435 16585.53 10000 ;
      RECT 16566.97 1047.855 16570.01 10000 ;
      RECT 16549.99 1047.855 16553.03 10000 ;
      RECT 16552.405 1046.435 16553.03 10000 ;
      RECT 16534.47 1046.435 16536.05 10000 ;
      RECT 16503.95 1047.855 16505.53 10000 ;
      RECT 16486.97 1046.435 16490.01 10000 ;
      RECT 16469.99 1046.435 16473.03 10000 ;
      RECT 16454.47 1046.435 16456.05 10000 ;
      RECT 16423.95 1047.855 16425.53 10000 ;
      RECT 16406.97 1047.855 16410.01 10000 ;
      RECT 16389.99 1046.435 16393.03 10000 ;
      RECT 16374.47 1046.435 16376.05 10000 ;
      RECT 16343.95 1047.855 16345.53 10000 ;
      RECT 16326.97 1046.435 16330.01 10000 ;
      RECT 16309.99 1046.435 16313.03 10000 ;
      RECT 16294.47 1046.435 16296.05 10000 ;
      RECT 16263.95 1047.855 16265.53 10000 ;
      RECT 16246.97 1046.435 16250.01 10000 ;
      RECT 16229.99 1047.855 16233.03 10000 ;
      RECT 16232.645 1046.435 16233.03 10000 ;
      RECT 16214.47 1046.435 16216.05 10000 ;
      RECT 16183.95 1046.435 16185.53 10000 ;
      RECT 16166.97 1046.435 16170.01 10000 ;
      RECT 16149.99 1047.855 16153.03 10000 ;
      RECT 16134.47 1046.435 16136.05 10000 ;
      RECT 16103.95 1046.435 16105.53 10000 ;
      RECT 16086.97 1047.855 16090.01 10000 ;
      RECT 16069.99 1046.435 16073.03 10000 ;
      RECT 16054.47 1047.855 16056.05 10000 ;
      RECT 16023.95 1046.435 16025.53 10000 ;
      RECT 16006.97 1047.855 16010.01 10000 ;
      RECT 15989.99 1047.855 15993.03 10000 ;
      RECT 15992.405 1046.435 15993.03 10000 ;
      RECT 15974.47 1046.435 15976.05 10000 ;
      RECT 15943.95 1047.855 15945.53 10000 ;
      RECT 15926.97 1046.435 15930.01 10000 ;
      RECT 15909.99 1046.435 15913.03 10000 ;
      RECT 15894.47 1046.435 15896.05 10000 ;
      RECT 15863.95 1047.855 15865.53 10000 ;
      RECT 15846.97 1047.855 15850.01 10000 ;
      RECT 15829.99 1046.435 15833.03 10000 ;
      RECT 15814.47 1046.435 15816.05 10000 ;
      RECT 15783.95 1047.855 15785.53 10000 ;
      RECT 15766.97 1046.435 15770.01 10000 ;
      RECT 15749.99 1046.435 15753.03 10000 ;
      RECT 15734.47 1046.435 15736.05 10000 ;
      RECT 15703.95 1047.855 15705.53 10000 ;
      RECT 15686.97 1046.435 15690.01 10000 ;
      RECT 15669.99 1047.855 15673.03 10000 ;
      RECT 15672.645 1046.435 15673.03 10000 ;
      RECT 15654.47 1046.435 15656.05 10000 ;
      RECT 15623.95 1046.435 15625.53 10000 ;
      RECT 15606.97 1046.435 15610.01 10000 ;
      RECT 15589.99 1047.855 15593.03 10000 ;
      RECT 15574.47 1046.435 15576.05 10000 ;
      RECT 15543.95 1046.435 15545.53 10000 ;
      RECT 15526.97 1047.855 15530.01 10000 ;
      RECT 15509.99 1046.435 15513.03 10000 ;
      RECT 15494.47 1047.855 15496.05 10000 ;
      RECT 15463.95 1046.435 15465.53 10000 ;
      RECT 15446.97 1047.855 15450.01 10000 ;
      RECT 15429.99 1047.855 15433.03 10000 ;
      RECT 15432.405 1046.435 15433.03 10000 ;
      RECT 15414.47 1046.435 15416.05 10000 ;
      RECT 15383.95 1047.855 15385.53 10000 ;
      RECT 15366.97 1046.435 15370.01 10000 ;
      RECT 15349.99 1046.435 15353.03 10000 ;
      RECT 15334.47 1046.435 15336.05 10000 ;
      RECT 15303.95 1047.855 15305.53 10000 ;
      RECT 15286.97 1047.855 15290.01 10000 ;
      RECT 15269.99 1046.435 15273.03 10000 ;
      RECT 15254.47 1046.435 15256.05 10000 ;
      RECT 15223.95 1047.855 15225.53 10000 ;
      RECT 15206.97 1046.435 15210.01 10000 ;
      RECT 15189.99 1046.435 15193.03 10000 ;
      RECT 15174.47 1046.435 15176.05 10000 ;
      RECT 15143.95 1047.855 15145.53 10000 ;
      RECT 15126.97 1046.435 15130.01 10000 ;
      RECT 15109.99 1047.855 15113.03 10000 ;
      RECT 15112.645 1046.435 15113.03 10000 ;
      RECT 15094.47 1046.435 15096.05 10000 ;
      RECT 15063.95 1046.435 15065.53 10000 ;
      RECT 15046.97 1046.435 15050.01 10000 ;
      RECT 15029.99 1047.855 15033.03 10000 ;
      RECT 15014.47 1046.435 15016.05 10000 ;
      RECT 14983.95 1046.435 14985.53 10000 ;
      RECT 14966.97 1047.855 14970.01 10000 ;
      RECT 14949.99 1046.435 14953.03 10000 ;
      RECT 14934.47 1047.855 14936.05 10000 ;
      RECT 14903.95 1046.435 14905.53 10000 ;
      RECT 14886.97 1047.855 14890.01 10000 ;
      RECT 14869.99 1047.855 14873.03 10000 ;
      RECT 14872.405 1046.435 14873.03 10000 ;
      RECT 14854.47 1046.435 14856.05 10000 ;
      RECT 14823.95 1047.855 14825.53 10000 ;
      RECT 14806.97 1046.435 14810.01 10000 ;
      RECT 14789.99 1046.435 14793.03 10000 ;
      RECT 14774.47 1046.435 14776.05 10000 ;
      RECT 14743.95 1047.855 14745.53 10000 ;
      RECT 14726.97 1047.855 14730.01 10000 ;
      RECT 14709.99 1046.435 14713.03 10000 ;
      RECT 14694.47 1046.435 14696.05 10000 ;
      RECT 14663.95 1047.855 14665.53 10000 ;
      RECT 14646.97 1046.435 14650.01 10000 ;
      RECT 14629.99 1046.435 14633.03 10000 ;
      RECT 14614.47 1046.435 14616.05 10000 ;
      RECT 14583.95 1047.855 14585.53 10000 ;
      RECT 14566.97 1046.435 14570.01 10000 ;
      RECT 14549.99 1047.855 14553.03 10000 ;
      RECT 14552.645 1046.435 14553.03 10000 ;
      RECT 14534.47 1046.435 14536.05 10000 ;
      RECT 14503.95 1046.435 14505.53 10000 ;
      RECT 14486.97 1046.435 14490.01 10000 ;
      RECT 14469.99 1047.855 14473.03 10000 ;
      RECT 14454.47 1046.435 14456.05 10000 ;
      RECT 14423.95 1046.435 14425.53 10000 ;
      RECT 14406.97 1047.855 14410.01 10000 ;
      RECT 14389.99 1046.435 14393.03 10000 ;
      RECT 14374.47 1047.855 14376.05 10000 ;
      RECT 14343.95 1046.435 14345.53 10000 ;
      RECT 14326.97 1047.855 14330.01 10000 ;
      RECT 14309.99 1047.855 14313.03 10000 ;
      RECT 14312.405 1046.435 14313.03 10000 ;
      RECT 14294.47 1046.435 14296.05 10000 ;
      RECT 14263.95 1047.855 14265.53 10000 ;
      RECT 14246.97 1046.435 14250.01 10000 ;
      RECT 14229.99 1046.435 14233.03 10000 ;
      RECT 14214.47 1046.435 14216.05 10000 ;
      RECT 14183.95 1047.855 14185.53 10000 ;
      RECT 14166.97 1047.855 14170.01 10000 ;
      RECT 14149.99 1046.435 14153.03 10000 ;
      RECT 14134.47 1046.435 14136.05 10000 ;
      RECT 14103.95 1047.855 14105.53 10000 ;
      RECT 14086.97 1046.435 14090.01 10000 ;
      RECT 14069.99 1046.435 14073.03 10000 ;
      RECT 14054.47 1046.435 14056.05 10000 ;
      RECT 14023.95 1047.855 14025.53 10000 ;
      RECT 14006.97 1046.435 14010.01 10000 ;
      RECT 13989.99 1047.855 13993.03 10000 ;
      RECT 13992.645 1046.435 13993.03 10000 ;
      RECT 13974.47 1046.435 13976.05 10000 ;
      RECT 13943.95 1046.435 13945.53 10000 ;
      RECT 13926.97 1046.435 13930.01 10000 ;
      RECT 13909.99 1047.855 13913.03 10000 ;
      RECT 13894.47 1046.435 13896.05 10000 ;
      RECT 13863.95 1046.435 13865.53 10000 ;
      RECT 13846.97 1047.855 13850.01 10000 ;
      RECT 13829.99 1046.435 13833.03 10000 ;
      RECT 13814.47 1047.855 13816.05 10000 ;
      RECT 13783.95 1046.435 13785.53 10000 ;
      RECT 13766.97 1047.855 13770.01 10000 ;
      RECT 13749.99 1047.855 13753.03 10000 ;
      RECT 13752.405 1046.435 13753.03 10000 ;
      RECT 13734.47 1046.435 13736.05 10000 ;
      RECT 13703.95 1047.855 13705.53 10000 ;
      RECT 13686.97 1046.435 13690.01 10000 ;
      RECT 13669.99 1046.435 13673.03 10000 ;
      RECT 13654.47 1046.435 13656.05 10000 ;
      RECT 13623.95 1047.855 13625.53 10000 ;
      RECT 13606.97 1047.855 13610.01 10000 ;
      RECT 13589.99 1046.435 13593.03 10000 ;
      RECT 13574.47 1046.435 13576.05 10000 ;
      RECT 13543.95 1047.855 13545.53 10000 ;
      RECT 13526.97 1046.435 13530.01 10000 ;
      RECT 13509.99 1046.435 13513.03 10000 ;
      RECT 13494.47 1046.435 13496.05 10000 ;
      RECT 13463.95 1047.855 13465.53 10000 ;
      RECT 13446.97 1046.435 13450.01 10000 ;
      RECT 13429.99 1047.855 13433.03 10000 ;
      RECT 13432.645 1046.435 13433.03 10000 ;
      RECT 13414.47 1046.435 13416.05 10000 ;
      RECT 13383.95 1046.435 13385.53 10000 ;
      RECT 13366.97 1046.435 13370.01 10000 ;
      RECT 13349.99 1047.855 13353.03 10000 ;
      RECT 13334.47 1046.435 13336.05 10000 ;
      RECT 13303.95 1046.435 13305.53 10000 ;
      RECT 13286.97 1047.855 13290.01 10000 ;
      RECT 13269.99 1046.435 13273.03 10000 ;
      RECT 13254.47 1047.855 13256.05 10000 ;
      RECT 13223.95 1046.435 13225.53 10000 ;
      RECT 13206.97 1047.855 13210.01 10000 ;
      RECT 13189.99 1047.855 13193.03 10000 ;
      RECT 13192.405 1046.435 13193.03 10000 ;
      RECT 13174.47 1046.435 13176.05 10000 ;
      RECT 13143.95 1047.855 13145.53 10000 ;
      RECT 13126.97 1046.435 13130.01 10000 ;
      RECT 13109.99 1046.435 13113.03 10000 ;
      RECT 13094.47 1046.435 13096.05 10000 ;
      RECT 13063.95 1047.855 13065.53 10000 ;
      RECT 13046.97 1047.855 13050.01 10000 ;
      RECT 13029.99 1046.435 13033.03 10000 ;
      RECT 13014.47 1046.435 13016.05 10000 ;
      RECT 12983.95 1047.855 12985.53 10000 ;
      RECT 12966.97 1046.435 12970.01 10000 ;
      RECT 12949.99 1046.435 12953.03 10000 ;
      RECT 12934.47 1046.435 12936.05 10000 ;
      RECT 12903.95 1047.855 12905.53 10000 ;
      RECT 12886.97 1046.435 12890.01 10000 ;
      RECT 12869.99 1047.855 12873.03 10000 ;
      RECT 12872.645 1046.435 12873.03 10000 ;
      RECT 12854.47 1046.435 12856.05 10000 ;
      RECT 12823.95 1046.435 12825.53 10000 ;
      RECT 12806.97 1046.435 12810.01 10000 ;
      RECT 12789.99 1047.855 12793.03 10000 ;
      RECT 12774.47 1046.435 12776.05 10000 ;
      RECT 12743.95 1046.435 12745.53 10000 ;
      RECT 12726.97 1047.855 12730.01 10000 ;
      RECT 12709.99 1046.435 12713.03 10000 ;
      RECT 12694.47 1047.855 12696.05 10000 ;
      RECT 12663.95 1046.435 12665.53 10000 ;
      RECT 12646.97 1047.855 12650.01 10000 ;
      RECT 12629.99 1047.855 12633.03 10000 ;
      RECT 12632.405 1046.435 12633.03 10000 ;
      RECT 12614.47 1046.435 12616.05 10000 ;
      RECT 12583.95 1047.855 12585.53 10000 ;
      RECT 12566.97 1046.435 12570.01 10000 ;
      RECT 12549.99 1046.435 12553.03 10000 ;
      RECT 12534.47 1046.435 12536.05 10000 ;
      RECT 12503.95 1047.855 12505.53 10000 ;
      RECT 12486.97 1047.855 12490.01 10000 ;
      RECT 12469.99 1046.435 12473.03 10000 ;
      RECT 12454.47 1046.435 12456.05 10000 ;
      RECT 12423.95 1047.855 12425.53 10000 ;
      RECT 12406.97 1046.435 12410.01 10000 ;
      RECT 12389.99 1046.435 12393.03 10000 ;
      RECT 12374.47 1046.435 12376.05 10000 ;
      RECT 12343.95 1047.855 12345.53 10000 ;
      RECT 12326.97 1046.435 12330.01 10000 ;
      RECT 12309.99 1047.855 12313.03 10000 ;
      RECT 12312.645 1046.435 12313.03 10000 ;
      RECT 12294.47 1046.435 12296.05 10000 ;
      RECT 12263.95 1046.435 12265.53 10000 ;
      RECT 12246.97 1046.435 12250.01 10000 ;
      RECT 12229.99 1047.855 12233.03 10000 ;
      RECT 12214.47 1046.435 12216.05 10000 ;
      RECT 12183.95 1046.435 12185.53 10000 ;
      RECT 12166.97 1047.855 12170.01 10000 ;
      RECT 12149.99 1046.435 12153.03 10000 ;
      RECT 12134.47 1047.855 12136.05 10000 ;
      RECT 12103.95 1046.435 12105.53 10000 ;
      RECT 12086.97 1047.855 12090.01 10000 ;
      RECT 12069.99 1047.855 12073.03 10000 ;
      RECT 12072.405 1046.435 12073.03 10000 ;
      RECT 12054.47 1046.435 12056.05 10000 ;
      RECT 12023.95 1047.855 12025.53 10000 ;
      RECT 12006.97 1046.435 12010.01 10000 ;
      RECT 11989.99 1046.435 11993.03 10000 ;
      RECT 11974.47 1046.435 11976.05 10000 ;
      RECT 11943.95 1047.855 11945.53 10000 ;
      RECT 11926.97 1047.855 11930.01 10000 ;
      RECT 11909.99 1046.435 11913.03 10000 ;
      RECT 11894.47 1046.435 11896.05 10000 ;
      RECT 11863.95 1047.855 11865.53 10000 ;
      RECT 11846.97 1046.435 11850.01 10000 ;
      RECT 11829.99 1046.435 11833.03 10000 ;
      RECT 11814.47 1046.435 11816.05 10000 ;
      RECT 11783.95 1047.855 11785.53 10000 ;
      RECT 11766.97 1046.435 11770.01 10000 ;
      RECT 11749.99 1047.855 11753.03 10000 ;
      RECT 11752.645 1046.435 11753.03 10000 ;
      RECT 11734.47 1046.435 11736.05 10000 ;
      RECT 11703.95 1046.435 11705.53 10000 ;
      RECT 11686.97 1046.435 11690.01 10000 ;
      RECT 11669.99 1047.855 11673.03 10000 ;
      RECT 11654.47 1046.435 11656.05 10000 ;
      RECT 11623.95 1046.435 11625.53 10000 ;
      RECT 11606.97 1047.855 11610.01 10000 ;
      RECT 11589.99 1046.435 11593.03 10000 ;
      RECT 11574.47 1047.855 11576.05 10000 ;
      RECT 11543.95 1046.435 11545.53 10000 ;
      RECT 11526.97 1047.855 11530.01 10000 ;
      RECT 11509.99 1047.855 11513.03 10000 ;
      RECT 11512.405 1046.435 11513.03 10000 ;
      RECT 11494.47 1046.435 11496.05 10000 ;
      RECT 11463.95 1047.855 11465.53 10000 ;
      RECT 11446.97 1046.435 11450.01 10000 ;
      RECT 11429.99 1046.435 11433.03 10000 ;
      RECT 11414.47 1046.435 11416.05 10000 ;
      RECT 11383.95 1047.855 11385.53 10000 ;
      RECT 11366.97 1047.855 11370.01 10000 ;
      RECT 11349.99 1046.435 11353.03 10000 ;
      RECT 11334.47 1046.435 11336.05 10000 ;
      RECT 11303.95 1047.855 11305.53 10000 ;
      RECT 11286.97 1046.435 11290.01 10000 ;
      RECT 11269.99 1046.435 11273.03 10000 ;
      RECT 11254.47 1046.435 11256.05 10000 ;
      RECT 11223.95 1047.855 11225.53 10000 ;
      RECT 11206.97 1046.435 11210.01 10000 ;
      RECT 11189.99 1047.855 11193.03 10000 ;
      RECT 11192.645 1046.435 11193.03 10000 ;
      RECT 11174.47 1046.435 11176.05 10000 ;
      RECT 11143.95 1046.435 11145.53 10000 ;
      RECT 11126.97 1046.435 11130.01 10000 ;
      RECT 11109.99 1047.855 11113.03 10000 ;
      RECT 11094.47 1046.435 11096.05 10000 ;
      RECT 11063.95 1046.435 11065.53 10000 ;
      RECT 11046.97 1047.855 11050.01 10000 ;
      RECT 11029.99 1046.435 11033.03 10000 ;
      RECT 11014.47 1047.855 11016.05 10000 ;
      RECT 10983.95 1046.435 10985.53 10000 ;
      RECT 10966.97 1047.855 10970.01 10000 ;
      RECT 10949.99 1047.855 10953.03 10000 ;
      RECT 10952.405 1046.435 10953.03 10000 ;
      RECT 10934.47 1046.435 10936.05 10000 ;
      RECT 10903.95 1047.855 10905.53 10000 ;
      RECT 10886.97 1046.435 10890.01 10000 ;
      RECT 10869.99 1046.435 10873.03 10000 ;
      RECT 10854.47 1046.435 10856.05 10000 ;
      RECT 10823.95 1047.855 10825.53 10000 ;
      RECT 10806.97 1047.855 10810.01 10000 ;
      RECT 10789.99 1046.435 10793.03 10000 ;
      RECT 10774.47 1046.435 10776.05 10000 ;
      RECT 10743.95 1047.855 10745.53 10000 ;
      RECT 10726.97 1046.435 10730.01 10000 ;
      RECT 10709.99 1046.435 10713.03 10000 ;
      RECT 10694.47 1046.435 10696.05 10000 ;
      RECT 10663.95 1047.855 10665.53 10000 ;
      RECT 10646.97 1046.435 10650.01 10000 ;
      RECT 10629.99 1047.855 10633.03 10000 ;
      RECT 10632.645 1046.435 10633.03 10000 ;
      RECT 10614.47 1046.435 10616.05 10000 ;
      RECT 10583.95 1046.435 10585.53 10000 ;
      RECT 10566.97 1046.435 10570.01 10000 ;
      RECT 10549.99 1047.855 10553.03 10000 ;
      RECT 10534.47 1046.435 10536.05 10000 ;
      RECT 10503.95 1046.435 10505.53 10000 ;
      RECT 10486.97 1047.855 10490.01 10000 ;
      RECT 10469.99 1046.435 10473.03 10000 ;
      RECT 10454.47 1047.855 10456.05 10000 ;
      RECT 10423.95 1046.435 10425.53 10000 ;
      RECT 10406.97 1047.855 10410.01 10000 ;
      RECT 10389.99 1047.855 10393.03 10000 ;
      RECT 10392.405 1046.435 10393.03 10000 ;
      RECT 10374.47 1046.435 10376.05 10000 ;
      RECT 10343.95 1047.855 10345.53 10000 ;
      RECT 10326.97 1046.435 10330.01 10000 ;
      RECT 10309.99 1046.435 10313.03 10000 ;
      RECT 10294.47 1046.435 10296.05 10000 ;
      RECT 10263.95 1047.855 10265.53 10000 ;
      RECT 10246.97 1047.855 10250.01 10000 ;
      RECT 10229.99 1046.435 10233.03 10000 ;
      RECT 10214.47 1046.435 10216.05 10000 ;
      RECT 10183.95 1047.855 10185.53 10000 ;
      RECT 10166.97 1046.435 10170.01 10000 ;
      RECT 10149.99 1046.435 10153.03 10000 ;
      RECT 10134.47 1046.435 10136.05 10000 ;
      RECT 10103.95 1047.855 10105.53 10000 ;
      RECT 10086.97 1046.435 10090.01 10000 ;
      RECT 10069.99 1047.855 10073.03 10000 ;
      RECT 10072.645 1046.435 10073.03 10000 ;
      RECT 10054.47 1046.435 10056.05 10000 ;
      RECT 10023.95 1046.435 10025.53 10000 ;
      RECT 10006.97 1046.435 10010.01 10000 ;
      RECT 9989.99 1047.855 9993.03 10000 ;
      RECT 9974.47 1046.435 9976.05 10000 ;
      RECT 9943.95 1046.435 9945.53 10000 ;
      RECT 9926.97 1047.855 9930.01 10000 ;
      RECT 9909.99 1046.435 9913.03 10000 ;
      RECT 9894.47 1047.855 9896.05 10000 ;
      RECT 9863.95 1046.435 9865.53 10000 ;
      RECT 9846.97 1047.855 9850.01 10000 ;
      RECT 9829.99 1047.855 9833.03 10000 ;
      RECT 9832.405 1046.435 9833.03 10000 ;
      RECT 9814.47 1046.435 9816.05 10000 ;
      RECT 9783.95 1047.855 9785.53 10000 ;
      RECT 9766.97 1046.435 9770.01 10000 ;
      RECT 9749.99 1046.435 9753.03 10000 ;
      RECT 9734.47 1046.435 9736.05 10000 ;
      RECT 9703.95 1047.855 9705.53 10000 ;
      RECT 9686.97 1047.855 9690.01 10000 ;
      RECT 9669.99 1046.435 9673.03 10000 ;
      RECT 9654.47 1046.435 9656.05 10000 ;
      RECT 9623.95 1047.855 9625.53 10000 ;
      RECT 9606.97 1046.435 9610.01 10000 ;
      RECT 9589.99 1046.435 9593.03 10000 ;
      RECT 9574.47 1046.435 9576.05 10000 ;
      RECT 9543.95 1047.855 9545.53 10000 ;
      RECT 9526.97 1046.435 9530.01 10000 ;
      RECT 9509.99 1047.855 9513.03 10000 ;
      RECT 9512.645 1046.435 9513.03 10000 ;
      RECT 9494.47 1046.435 9496.05 10000 ;
      RECT 9463.95 1046.435 9465.53 10000 ;
      RECT 9446.97 1046.435 9450.01 10000 ;
      RECT 9429.99 1047.855 9433.03 10000 ;
      RECT 9414.47 1046.435 9416.05 10000 ;
      RECT 9383.95 1046.435 9385.53 10000 ;
      RECT 9366.97 1047.855 9370.01 10000 ;
      RECT 9349.99 1046.435 9353.03 10000 ;
      RECT 9334.47 1047.855 9336.05 10000 ;
      RECT 9303.95 1046.435 9305.53 10000 ;
      RECT 9286.97 1047.855 9290.01 10000 ;
      RECT 9269.99 1047.855 9273.03 10000 ;
      RECT 9272.405 1046.435 9273.03 10000 ;
      RECT 9254.47 1046.435 9256.05 10000 ;
      RECT 9223.95 1047.855 9225.53 10000 ;
      RECT 9206.97 1046.435 9210.01 10000 ;
      RECT 9189.99 1046.435 9193.03 10000 ;
      RECT 9174.47 1046.435 9176.05 10000 ;
      RECT 9143.95 1047.855 9145.53 10000 ;
      RECT 9126.97 1047.855 9130.01 10000 ;
      RECT 9109.99 1046.435 9113.03 10000 ;
      RECT 9094.47 1046.435 9096.05 10000 ;
      RECT 9063.95 1047.855 9065.53 10000 ;
      RECT 9046.97 1046.435 9050.01 10000 ;
      RECT 9029.99 1046.435 9033.03 10000 ;
      RECT 9014.47 1046.435 9016.05 10000 ;
      RECT 8983.95 1047.855 8985.53 10000 ;
      RECT 8966.97 1046.435 8970.01 10000 ;
      RECT 8949.99 1047.855 8953.03 10000 ;
      RECT 8952.645 1046.435 8953.03 10000 ;
      RECT 8934.47 1046.435 8936.05 10000 ;
      RECT 8903.95 1046.435 8905.53 10000 ;
      RECT 8886.97 1046.435 8890.01 10000 ;
      RECT 8869.99 1047.855 8873.03 10000 ;
      RECT 8854.47 1046.435 8856.05 10000 ;
      RECT 8823.95 1046.435 8825.53 10000 ;
      RECT 8806.97 1047.855 8810.01 10000 ;
      RECT 8789.99 1046.435 8793.03 10000 ;
      RECT 8774.47 1047.855 8776.05 10000 ;
      RECT 8743.95 1046.435 8745.53 10000 ;
      RECT 8726.97 1047.855 8730.01 10000 ;
      RECT 8709.99 1047.855 8713.03 10000 ;
      RECT 8712.405 1046.435 8713.03 10000 ;
      RECT 8694.47 1046.435 8696.05 10000 ;
      RECT 8663.95 1047.855 8665.53 10000 ;
      RECT 8646.97 1046.435 8650.01 10000 ;
      RECT 8629.99 1046.435 8633.03 10000 ;
      RECT 8614.47 1046.435 8616.05 10000 ;
      RECT 8583.95 1047.855 8585.53 10000 ;
      RECT 8566.97 1047.855 8570.01 10000 ;
      RECT 8549.99 1046.435 8553.03 10000 ;
      RECT 8534.47 1046.435 8536.05 10000 ;
      RECT 8503.95 1047.855 8505.53 10000 ;
      RECT 8486.97 1046.435 8490.01 10000 ;
      RECT 8469.99 1046.435 8473.03 10000 ;
      RECT 8454.47 1046.435 8456.05 10000 ;
      RECT 8423.95 1047.855 8425.53 10000 ;
      RECT 8406.97 1046.435 8410.01 10000 ;
      RECT 8389.99 1047.855 8393.03 10000 ;
      RECT 8392.645 1046.435 8393.03 10000 ;
      RECT 8374.47 1046.435 8376.05 10000 ;
      RECT 8343.95 1046.435 8345.53 10000 ;
      RECT 8326.97 1046.435 8330.01 10000 ;
      RECT 8309.99 1047.855 8313.03 10000 ;
      RECT 8294.47 1046.435 8296.05 10000 ;
      RECT 8263.95 1046.435 8265.53 10000 ;
      RECT 8246.97 1047.855 8250.01 10000 ;
      RECT 8229.99 1046.435 8233.03 10000 ;
      RECT 8214.47 1047.855 8216.05 10000 ;
      RECT 8183.95 1046.435 8185.53 10000 ;
      RECT 8166.97 1047.855 8170.01 10000 ;
      RECT 8149.99 1047.855 8153.03 10000 ;
      RECT 8152.405 1046.435 8153.03 10000 ;
      RECT 8134.47 1046.435 8136.05 10000 ;
      RECT 8103.95 1047.855 8105.53 10000 ;
      RECT 8086.97 1046.435 8090.01 10000 ;
      RECT 8069.99 1046.435 8073.03 10000 ;
      RECT 8054.47 1046.435 8056.05 10000 ;
      RECT 8023.95 1047.855 8025.53 10000 ;
      RECT 8006.97 1047.855 8010.01 10000 ;
      RECT 7989.99 1046.435 7993.03 10000 ;
      RECT 7974.47 1046.435 7976.05 10000 ;
      RECT 7943.95 1047.855 7945.53 10000 ;
      RECT 7926.97 1046.435 7930.01 10000 ;
      RECT 7909.99 1046.435 7913.03 10000 ;
      RECT 7894.47 1046.435 7896.05 10000 ;
      RECT 7863.95 1047.855 7865.53 10000 ;
      RECT 7846.97 1046.435 7850.01 10000 ;
      RECT 7829.99 1047.855 7833.03 10000 ;
      RECT 7832.645 1046.435 7833.03 10000 ;
      RECT 7814.47 1046.435 7816.05 10000 ;
      RECT 7783.95 1046.435 7785.53 10000 ;
      RECT 7766.97 1046.435 7770.01 10000 ;
      RECT 7749.99 1047.855 7753.03 10000 ;
      RECT 7734.47 1046.435 7736.05 10000 ;
      RECT 7703.95 1046.435 7705.53 10000 ;
      RECT 7686.97 1047.855 7690.01 10000 ;
      RECT 7669.99 1046.435 7673.03 10000 ;
      RECT 7654.47 1047.855 7656.05 10000 ;
      RECT 7623.95 1046.435 7625.53 10000 ;
      RECT 7606.97 1047.855 7610.01 10000 ;
      RECT 7589.99 1047.855 7593.03 10000 ;
      RECT 7592.405 1046.435 7593.03 10000 ;
      RECT 7574.47 1046.435 7576.05 10000 ;
      RECT 7543.95 1047.855 7545.53 10000 ;
      RECT 7526.97 1046.435 7530.01 10000 ;
      RECT 7509.99 1046.435 7513.03 10000 ;
      RECT 7494.47 1046.435 7496.05 10000 ;
      RECT 7463.95 1047.855 7465.53 10000 ;
      RECT 7446.97 1047.855 7450.01 10000 ;
      RECT 7429.99 1046.435 7433.03 10000 ;
      RECT 7414.47 1046.435 7416.05 10000 ;
      RECT 7383.95 1047.855 7385.53 10000 ;
      RECT 7366.97 1046.435 7370.01 10000 ;
      RECT 7349.99 1046.435 7353.03 10000 ;
      RECT 7334.47 1046.435 7336.05 10000 ;
      RECT 7303.95 1047.855 7305.53 10000 ;
      RECT 7286.97 1046.435 7290.01 10000 ;
      RECT 7269.99 1047.855 7273.03 10000 ;
      RECT 7272.645 1046.435 7273.03 10000 ;
      RECT 7254.47 1046.435 7256.05 10000 ;
      RECT 7223.95 1046.435 7225.53 10000 ;
      RECT 7206.97 1046.435 7210.01 10000 ;
      RECT 7189.99 1047.855 7193.03 10000 ;
      RECT 7174.47 1046.435 7176.05 10000 ;
      RECT 7143.95 1046.435 7145.53 10000 ;
      RECT 7126.97 1047.855 7130.01 10000 ;
      RECT 7109.99 1046.435 7113.03 10000 ;
      RECT 7094.47 1047.855 7096.05 10000 ;
      RECT 7063.95 1046.435 7065.53 10000 ;
      RECT 7046.97 1047.855 7050.01 10000 ;
      RECT 7029.99 1047.855 7033.03 10000 ;
      RECT 7032.405 1046.435 7033.03 10000 ;
      RECT 7014.47 1046.435 7016.05 10000 ;
      RECT 6983.95 1047.855 6985.53 10000 ;
      RECT 6966.97 1046.435 6970.01 10000 ;
      RECT 6949.99 1046.435 6953.03 10000 ;
      RECT 6934.47 1046.435 6936.05 10000 ;
      RECT 6903.95 1047.855 6905.53 10000 ;
      RECT 6886.97 1047.855 6890.01 10000 ;
      RECT 6869.99 1046.435 6873.03 10000 ;
      RECT 6854.47 1046.435 6856.05 10000 ;
      RECT 6823.95 1047.855 6825.53 10000 ;
      RECT 6806.97 1046.435 6810.01 10000 ;
      RECT 6789.99 1046.435 6793.03 10000 ;
      RECT 6774.47 1046.435 6776.05 10000 ;
      RECT 6743.95 1047.855 6745.53 10000 ;
      RECT 6726.97 1046.435 6730.01 10000 ;
      RECT 6709.99 1047.855 6713.03 10000 ;
      RECT 6712.645 1046.435 6713.03 10000 ;
      RECT 6694.47 1046.435 6696.05 10000 ;
      RECT 6663.95 1046.435 6665.53 10000 ;
      RECT 6646.97 1046.435 6650.01 10000 ;
      RECT 6629.99 1047.855 6633.03 10000 ;
      RECT 6614.47 1046.435 6616.05 10000 ;
      RECT 6583.95 1046.435 6585.53 10000 ;
      RECT 6566.97 1047.855 6570.01 10000 ;
      RECT 6549.99 1046.435 6553.03 10000 ;
      RECT 6534.47 1047.855 6536.05 10000 ;
      RECT 6503.95 1046.435 6505.53 10000 ;
      RECT 6486.97 1047.855 6490.01 10000 ;
      RECT 6469.99 1047.855 6473.03 10000 ;
      RECT 6472.405 1046.435 6473.03 10000 ;
      RECT 6454.47 1046.435 6456.05 10000 ;
      RECT 6423.95 1047.855 6425.53 10000 ;
      RECT 6406.97 1046.435 6410.01 10000 ;
      RECT 6389.99 1046.435 6393.03 10000 ;
      RECT 6374.47 1046.435 6376.05 10000 ;
      RECT 6343.95 1047.855 6345.53 10000 ;
      RECT 6326.97 1047.855 6330.01 10000 ;
      RECT 6309.99 1046.435 6313.03 10000 ;
      RECT 6294.47 1046.435 6296.05 10000 ;
      RECT 6263.95 1047.855 6265.53 10000 ;
      RECT 6246.97 1046.435 6250.01 10000 ;
      RECT 6229.99 1046.435 6233.03 10000 ;
      RECT 6214.47 1046.435 6216.05 10000 ;
      RECT 6183.95 1047.855 6185.53 10000 ;
      RECT 6166.97 1046.435 6170.01 10000 ;
      RECT 6149.99 1047.855 6153.03 10000 ;
      RECT 6152.645 1046.435 6153.03 10000 ;
      RECT 6134.47 1046.435 6136.05 10000 ;
      RECT 6103.95 1046.435 6105.53 10000 ;
      RECT 6086.97 1046.435 6090.01 10000 ;
      RECT 6069.99 1047.855 6073.03 10000 ;
      RECT 6054.47 1046.435 6056.05 10000 ;
      RECT 6023.95 1046.435 6025.53 10000 ;
      RECT 6006.97 1047.855 6010.01 10000 ;
      RECT 5989.99 1046.435 5993.03 10000 ;
      RECT 5974.47 1047.855 5976.05 10000 ;
      RECT 5943.95 1046.435 5945.53 10000 ;
      RECT 5926.97 1047.855 5930.01 10000 ;
      RECT 5909.99 1047.855 5913.03 10000 ;
      RECT 5912.405 1046.435 5913.03 10000 ;
      RECT 5894.47 1046.435 5896.05 10000 ;
      RECT 5863.95 1047.855 5865.53 10000 ;
      RECT 5846.97 1046.435 5850.01 10000 ;
      RECT 5829.99 1046.435 5833.03 10000 ;
      RECT 5814.47 1046.435 5816.05 10000 ;
      RECT 5783.95 1047.855 5785.53 10000 ;
      RECT 5766.97 1047.855 5770.01 10000 ;
      RECT 5749.99 1046.435 5753.03 10000 ;
      RECT 5734.47 1046.435 5736.05 10000 ;
      RECT 5703.95 1047.855 5705.53 10000 ;
      RECT 5686.97 1046.435 5690.01 10000 ;
      RECT 5669.99 1046.435 5673.03 10000 ;
      RECT 5654.47 1046.435 5656.05 10000 ;
      RECT 5623.95 1047.855 5625.53 10000 ;
      RECT 5606.97 1046.435 5610.01 10000 ;
      RECT 5589.99 1047.855 5593.03 10000 ;
      RECT 5592.645 1046.435 5593.03 10000 ;
      RECT 5574.47 1046.435 5576.05 10000 ;
      RECT 5543.95 1046.435 5545.53 10000 ;
      RECT 5526.97 1046.435 5530.01 10000 ;
      RECT 5509.99 1047.855 5513.03 10000 ;
      RECT 5494.47 1046.435 5496.05 10000 ;
      RECT 5463.95 1046.435 5465.53 10000 ;
      RECT 5446.97 1047.855 5450.01 10000 ;
      RECT 5429.99 1046.435 5433.03 10000 ;
      RECT 5414.47 1047.855 5416.05 10000 ;
      RECT 5383.95 1046.435 5385.53 10000 ;
      RECT 5366.97 1047.855 5370.01 10000 ;
      RECT 5349.99 1047.855 5353.03 10000 ;
      RECT 5352.405 1046.435 5353.03 10000 ;
      RECT 5334.47 1046.435 5336.05 10000 ;
      RECT 5303.95 1047.855 5305.53 10000 ;
      RECT 5286.97 1046.435 5290.01 10000 ;
      RECT 5269.99 1046.435 5273.03 10000 ;
      RECT 5254.47 1046.435 5256.05 10000 ;
      RECT 5223.95 1047.855 5225.53 10000 ;
      RECT 5206.97 1047.855 5210.01 10000 ;
      RECT 5189.99 1046.435 5193.03 10000 ;
      RECT 5174.47 1046.435 5176.05 10000 ;
      RECT 5143.95 1047.855 5145.53 10000 ;
      RECT 5126.97 1046.435 5130.01 10000 ;
      RECT 5109.99 1046.435 5113.03 10000 ;
      RECT 5094.47 1046.435 5096.05 10000 ;
      RECT 5063.95 1047.855 5065.53 10000 ;
      RECT 5046.97 1046.435 5050.01 10000 ;
      RECT 5029.99 1047.855 5033.03 10000 ;
      RECT 5032.645 1046.435 5033.03 10000 ;
      RECT 5014.47 1046.435 5016.05 10000 ;
      RECT 4983.95 1046.435 4985.53 10000 ;
      RECT 4966.97 1046.435 4970.01 10000 ;
      RECT 4949.99 1047.855 4953.03 10000 ;
      RECT 4934.47 1046.435 4936.05 10000 ;
      RECT 4903.95 1046.435 4905.53 10000 ;
      RECT 4886.97 1047.855 4890.01 10000 ;
      RECT 4869.99 1046.435 4873.03 10000 ;
      RECT 4854.47 1047.855 4856.05 10000 ;
      RECT 4823.95 1046.435 4825.53 10000 ;
      RECT 4806.97 1047.855 4810.01 10000 ;
      RECT 4789.99 1047.855 4793.03 10000 ;
      RECT 4792.405 1046.435 4793.03 10000 ;
      RECT 4774.47 1046.435 4776.05 10000 ;
      RECT 4743.95 1047.855 4745.53 10000 ;
      RECT 4726.97 1046.435 4730.01 10000 ;
      RECT 4709.99 1046.435 4713.03 10000 ;
      RECT 4694.47 1046.435 4696.05 10000 ;
      RECT 4663.95 1047.855 4665.53 10000 ;
      RECT 4646.97 1047.855 4650.01 10000 ;
      RECT 4629.99 1046.435 4633.03 10000 ;
      RECT 4614.47 1046.435 4616.05 10000 ;
      RECT 4583.95 1047.855 4585.53 10000 ;
      RECT 4566.97 1046.435 4570.01 10000 ;
      RECT 4549.99 1046.435 4553.03 10000 ;
      RECT 4534.47 1046.435 4536.05 10000 ;
      RECT 4503.95 1047.855 4505.53 10000 ;
      RECT 4486.97 1046.435 4490.01 10000 ;
      RECT 4469.99 1047.855 4473.03 10000 ;
      RECT 4472.645 1046.435 4473.03 10000 ;
      RECT 4454.47 1046.435 4456.05 10000 ;
      RECT 4423.95 1046.435 4425.53 10000 ;
      RECT 4406.97 1046.435 4410.01 10000 ;
      RECT 4389.99 1047.855 4393.03 10000 ;
      RECT 4374.47 1046.435 4376.05 10000 ;
      RECT 4343.95 1046.435 4345.53 10000 ;
      RECT 4326.97 1047.855 4330.01 10000 ;
      RECT 4309.99 1046.435 4313.03 10000 ;
      RECT 4294.47 1047.855 4296.05 10000 ;
      RECT 4263.95 1046.435 4265.53 10000 ;
      RECT 4246.97 1047.855 4250.01 10000 ;
      RECT 4229.99 1047.855 4233.03 10000 ;
      RECT 4232.405 1046.435 4233.03 10000 ;
      RECT 4214.47 1046.435 4216.05 10000 ;
      RECT 4183.95 1047.855 4185.53 10000 ;
      RECT 4166.97 1046.435 4170.01 10000 ;
      RECT 4149.99 1046.435 4153.03 10000 ;
      RECT 4134.47 1046.435 4136.05 10000 ;
      RECT 4103.95 1047.855 4105.53 10000 ;
      RECT 4086.97 1047.855 4090.01 10000 ;
      RECT 4069.99 1046.435 4073.03 10000 ;
      RECT 4054.47 1046.435 4056.05 10000 ;
      RECT 4023.95 1047.855 4025.53 10000 ;
      RECT 4006.97 1046.435 4010.01 10000 ;
      RECT 3989.99 1046.435 3993.03 10000 ;
      RECT 3974.47 1046.435 3976.05 10000 ;
      RECT 3943.95 1047.855 3945.53 10000 ;
      RECT 3926.97 1046.435 3930.01 10000 ;
      RECT 3909.99 1047.855 3913.03 10000 ;
      RECT 3912.645 1046.435 3913.03 10000 ;
      RECT 3894.47 1046.435 3896.05 10000 ;
      RECT 3863.95 1046.435 3865.53 10000 ;
      RECT 3846.97 1046.435 3850.01 10000 ;
      RECT 3829.99 1047.855 3833.03 10000 ;
      RECT 3814.47 1046.435 3816.05 10000 ;
      RECT 3783.95 1046.435 3785.53 10000 ;
      RECT 3766.97 1047.855 3770.01 10000 ;
      RECT 3749.99 1046.435 3753.03 10000 ;
      RECT 3734.47 1047.855 3736.05 10000 ;
      RECT 3703.95 1046.435 3705.53 10000 ;
      RECT 3686.97 1047.855 3690.01 10000 ;
      RECT 3669.99 1047.855 3673.03 10000 ;
      RECT 3672.405 1046.435 3673.03 10000 ;
      RECT 3654.47 1046.435 3656.05 10000 ;
      RECT 3623.95 1047.855 3625.53 10000 ;
      RECT 3606.97 1046.435 3610.01 10000 ;
      RECT 3589.99 1046.435 3593.03 10000 ;
      RECT 3574.47 1046.435 3576.05 10000 ;
      RECT 3543.95 1047.855 3545.53 10000 ;
      RECT 3526.97 1047.855 3530.01 10000 ;
      RECT 3509.99 1046.435 3513.03 10000 ;
      RECT 3494.47 1046.435 3496.05 10000 ;
      RECT 3463.95 1047.855 3465.53 10000 ;
      RECT 3446.97 1046.435 3450.01 10000 ;
      RECT 3429.99 1046.435 3433.03 10000 ;
      RECT 3414.47 1046.435 3416.05 10000 ;
      RECT 3383.95 1047.855 3385.53 10000 ;
      RECT 3366.97 1046.435 3370.01 10000 ;
      RECT 3349.99 1047.855 3353.03 10000 ;
      RECT 3352.645 1046.435 3353.03 10000 ;
      RECT 3334.47 1046.435 3336.05 10000 ;
      RECT 3303.95 1046.435 3305.53 10000 ;
      RECT 3286.97 1046.435 3290.01 10000 ;
      RECT 3269.99 1047.855 3273.03 10000 ;
      RECT 3254.47 1046.435 3256.05 10000 ;
      RECT 3223.95 1046.435 3225.53 10000 ;
      RECT 3206.97 1047.855 3210.01 10000 ;
      RECT 3189.99 1046.435 3193.03 10000 ;
      RECT 3174.47 1047.855 3176.05 10000 ;
      RECT 3143.95 1046.435 3145.53 10000 ;
      RECT 3126.97 1047.855 3130.01 10000 ;
      RECT 3109.99 1047.855 3113.03 10000 ;
      RECT 3112.405 1046.435 3113.03 10000 ;
      RECT 3094.47 1046.435 3096.05 10000 ;
      RECT 3063.95 1047.855 3065.53 10000 ;
      RECT 3046.97 1046.435 3050.01 10000 ;
      RECT 3029.99 1046.435 3033.03 10000 ;
      RECT 3014.47 1046.435 3016.05 10000 ;
      RECT 2983.95 1047.855 2985.53 10000 ;
      RECT 2966.97 1047.855 2970.01 10000 ;
      RECT 2949.99 1046.435 2953.03 10000 ;
      RECT 2934.47 1046.435 2936.05 10000 ;
      RECT 2903.95 1047.855 2905.53 10000 ;
      RECT 2886.97 1046.435 2890.01 10000 ;
      RECT 2869.99 1046.435 2873.03 10000 ;
      RECT 2854.47 1046.435 2856.05 10000 ;
      RECT 2823.95 1047.855 2825.53 10000 ;
      RECT 2806.97 1046.435 2810.01 10000 ;
      RECT 2789.99 1047.855 2793.03 10000 ;
      RECT 2792.645 1046.435 2793.03 10000 ;
      RECT 2774.47 1046.435 2776.05 10000 ;
      RECT 2743.95 1046.435 2745.53 10000 ;
      RECT 2726.97 1046.435 2730.01 10000 ;
      RECT 2709.99 1047.855 2713.03 10000 ;
      RECT 2694.47 1046.435 2696.05 10000 ;
      RECT 2663.95 1046.435 2665.53 10000 ;
      RECT 2646.97 1047.855 2650.01 10000 ;
      RECT 2629.99 1046.435 2633.03 10000 ;
      RECT 2614.47 1047.855 2616.05 10000 ;
      RECT 2583.95 1046.435 2585.53 10000 ;
      RECT 2566.97 1047.855 2570.01 10000 ;
      RECT 2549.99 1047.855 2553.03 10000 ;
      RECT 2552.405 1046.435 2553.03 10000 ;
      RECT 2534.47 1046.435 2536.05 10000 ;
      RECT 2503.95 1047.855 2505.53 10000 ;
      RECT 2486.97 1046.435 2490.01 10000 ;
      RECT 2469.99 1046.435 2473.03 10000 ;
      RECT 2454.47 1046.435 2456.05 10000 ;
      RECT 2423.95 1047.855 2425.53 10000 ;
      RECT 2406.97 1047.855 2410.01 10000 ;
      RECT 2389.99 1046.435 2393.03 10000 ;
      RECT 2374.47 1046.435 2376.05 10000 ;
      RECT 2343.95 1047.855 2345.53 10000 ;
      RECT 2326.97 1046.435 2330.01 10000 ;
      RECT 2309.99 1046.435 2313.03 10000 ;
      RECT 2294.47 1046.435 2296.05 10000 ;
      RECT 2263.95 1047.855 2265.53 10000 ;
      RECT 2246.97 1046.435 2250.01 10000 ;
      RECT 2229.99 1047.855 2233.03 10000 ;
      RECT 2232.645 1046.435 2233.03 10000 ;
      RECT 2214.47 1046.435 2216.05 10000 ;
      RECT 2183.95 1046.435 2185.53 10000 ;
      RECT 2166.97 1046.435 2170.01 10000 ;
      RECT 2149.99 1047.855 2153.03 10000 ;
      RECT 2134.47 1046.435 2136.05 10000 ;
      RECT 2103.95 1046.435 2105.53 10000 ;
      RECT 2086.97 1047.855 2090.01 10000 ;
      RECT 2069.99 1046.435 2073.03 10000 ;
      RECT 2054.47 1047.855 2056.05 10000 ;
      RECT 2023.95 1046.435 2025.53 10000 ;
      RECT 2006.97 1047.855 2010.01 10000 ;
      RECT 1989.99 1047.855 1993.03 10000 ;
      RECT 1992.405 1046.435 1993.03 10000 ;
      RECT 1974.47 1046.435 1976.05 10000 ;
      RECT 1943.95 1047.855 1945.53 10000 ;
      RECT 1926.97 1046.435 1930.01 10000 ;
      RECT 1909.99 1046.435 1913.03 10000 ;
      RECT 1894.47 1046.435 1896.05 10000 ;
      RECT 1863.95 1047.855 1865.53 10000 ;
      RECT 1846.97 1047.855 1850.01 10000 ;
      RECT 1829.99 1046.435 1833.03 10000 ;
      RECT 1814.47 1046.435 1816.05 10000 ;
      RECT 1783.95 1047.855 1785.53 10000 ;
      RECT 1766.97 1046.435 1770.01 10000 ;
      RECT 1749.99 1046.435 1753.03 10000 ;
      RECT 1734.47 1046.435 1736.05 10000 ;
      RECT 1703.95 1047.855 1705.53 10000 ;
      RECT 1686.97 1046.435 1690.01 10000 ;
      RECT 1669.99 1047.855 1673.03 10000 ;
      RECT 1672.645 1046.435 1673.03 10000 ;
      RECT 1654.47 1046.435 1656.05 10000 ;
      RECT 1623.95 1046.435 1625.53 10000 ;
      RECT 1606.97 1046.435 1610.01 10000 ;
      RECT 1589.99 1047.855 1593.03 10000 ;
      RECT 1574.47 1046.435 1576.05 10000 ;
      RECT 1543.95 1046.435 1545.53 10000 ;
      RECT 1526.97 1047.855 1530.01 10000 ;
      RECT 1509.99 1046.435 1513.03 10000 ;
      RECT 1494.47 1047.855 1496.05 10000 ;
      RECT 1463.95 1046.435 1465.53 10000 ;
      RECT 1446.97 1047.855 1450.01 10000 ;
      RECT 1429.99 1047.855 1433.03 10000 ;
      RECT 1432.405 1046.435 1433.03 10000 ;
      RECT 1414.47 1046.435 1416.05 10000 ;
      RECT 1383.95 1047.855 1385.53 10000 ;
      RECT 1366.97 1046.435 1370.01 10000 ;
      RECT 1349.99 1046.435 1353.03 10000 ;
      RECT 1334.47 1046.435 1336.05 10000 ;
      RECT 1303.95 1047.855 1305.53 10000 ;
      RECT 1286.97 1047.855 1290.01 10000 ;
      RECT 1269.99 1046.435 1273.03 10000 ;
      RECT 1254.47 1046.435 1256.05 10000 ;
      RECT 1223.95 1047.855 1225.53 10000 ;
      RECT 1206.97 1046.435 1210.01 10000 ;
      RECT 1189.99 1046.435 1193.03 10000 ;
      RECT 1174.47 1046.435 1176.05 10000 ;
      RECT 1143.95 1047.855 1145.53 10000 ;
      RECT 998.1 1046.435 1130.01 10000 ;
      RECT 18503.95 1046.435 18504.565 10000 ;
      RECT 17943.95 1046.435 17944.565 10000 ;
      RECT 17383.95 1046.435 17384.565 10000 ;
      RECT 16823.95 1046.435 16824.565 10000 ;
      RECT 16263.95 1046.435 16264.565 10000 ;
      RECT 15703.95 1046.435 15704.565 10000 ;
      RECT 15143.95 1046.435 15144.565 10000 ;
      RECT 14583.95 1046.435 14584.565 10000 ;
      RECT 14023.95 1046.435 14024.565 10000 ;
      RECT 13463.95 1046.435 13464.565 10000 ;
      RECT 12903.95 1046.435 12904.565 10000 ;
      RECT 12343.95 1046.435 12344.565 10000 ;
      RECT 11783.95 1046.435 11784.565 10000 ;
      RECT 11223.95 1046.435 11224.565 10000 ;
      RECT 10663.95 1046.435 10664.565 10000 ;
      RECT 10103.95 1046.435 10104.565 10000 ;
      RECT 9543.95 1046.435 9544.565 10000 ;
      RECT 8983.95 1046.435 8984.565 10000 ;
      RECT 8423.95 1046.435 8424.565 10000 ;
      RECT 7863.95 1046.435 7864.565 10000 ;
      RECT 7303.95 1046.435 7304.565 10000 ;
      RECT 6743.95 1046.435 6744.565 10000 ;
      RECT 6183.95 1046.435 6184.565 10000 ;
      RECT 5623.95 1046.435 5624.565 10000 ;
      RECT 5063.95 1046.435 5064.565 10000 ;
      RECT 4503.95 1046.435 4504.565 10000 ;
      RECT 3943.95 1046.435 3944.565 10000 ;
      RECT 3383.95 1046.435 3384.565 10000 ;
      RECT 2823.95 1046.435 2824.565 10000 ;
      RECT 2263.95 1046.435 2264.565 10000 ;
      RECT 1703.95 1046.435 1704.565 10000 ;
      RECT 1143.95 1046.435 1144.565 10000 ;
    LAYER TOP_M ;
      RECT 0.5 9996.5 20199.5 9999.5 ;
      RECT 20196.5 0.5 20199.5 9999.5 ;
      RECT 0.5 0.5 3.5 9999.5 ;
      RECT 0.5 0.5 20199.5 3.5 ;
      RECT 4.1 9989 20195.9 9995.9 ;
      RECT 20189 4.1 20195.9 9995.9 ;
      RECT 4.1 4.1 11 9995.9 ;
      RECT 4.1 4.1 20195.9 11 ;
      RECT 19475.9 617.18 19567.9 709.18 ;
      RECT 19454.5 638.18 19567.9 688.18 ;
      RECT 19454.5 657.18 19697.905 669.18 ;
      RECT 19475.9 9377.18 19567.9 9469.18 ;
      RECT 19454.5 9398.18 19567.9 9448.18 ;
      RECT 19454.5 9417.18 19697.905 9429.18 ;
      RECT 19605.9 677.18 19697.9 769.18 ;
      RECT 19584.5 680.155 19697.9 715.155 ;
      RECT 19605.9 797.18 19697.9 889.18 ;
      RECT 19584.5 800.155 19697.9 835.155 ;
      RECT 19605.9 917.18 19697.9 1009.18 ;
      RECT 19584.5 920.155 19697.9 955.155 ;
      RECT 19605.9 1037.18 19697.9 1129.18 ;
      RECT 19584.5 1040.155 19697.9 1075.155 ;
      RECT 19605.9 1277.18 19697.9 1369.18 ;
      RECT 19584.5 1280.155 19697.9 1315.155 ;
      RECT 19605.9 1397.18 19697.9 1489.18 ;
      RECT 19584.5 1400.155 19697.9 1435.155 ;
      RECT 19605.9 8717.18 19697.9 8809.18 ;
      RECT 19584.5 8720.155 19697.9 8755.155 ;
      RECT 19605.9 8837.18 19697.9 8929.18 ;
      RECT 19584.5 8840.155 19697.9 8875.155 ;
      RECT 19605.9 8957.18 19697.9 9049.18 ;
      RECT 19584.5 8960.155 19697.9 8995.155 ;
      RECT 19605.9 9077.18 19697.9 9169.18 ;
      RECT 19584.5 9080.155 19697.9 9115.155 ;
      RECT 19605.9 9197.18 19697.9 9289.18 ;
      RECT 19584.5 9200.155 19697.9 9235.155 ;
      RECT 19605.9 9317.18 19697.9 9409.18 ;
      RECT 19584.5 9320.155 19697.9 9355.155 ;
      RECT 19475.9 857.18 19567.9 949.18 ;
      RECT 19454.5 878.18 19567.9 928.18 ;
      RECT 19454.5 897.18 19691.9 909.18 ;
      RECT 19475.9 1097.18 19567.9 1189.18 ;
      RECT 19454.5 1118.18 19567.9 1168.18 ;
      RECT 19454.5 1137.18 19691.9 1149.18 ;
      RECT 19475.9 1337.18 19567.9 1429.18 ;
      RECT 19454.5 1358.18 19567.9 1408.18 ;
      RECT 19454.5 1377.18 19691.9 1389.18 ;
      RECT 19475.9 1937.18 19567.9 2029.18 ;
      RECT 19454.5 1958.18 19567.9 2008.18 ;
      RECT 19454.5 1977.18 19691.9 1989.18 ;
      RECT 19475.9 2417.18 19567.9 2509.18 ;
      RECT 19454.5 2438.18 19567.9 2488.18 ;
      RECT 19454.5 2457.18 19691.9 2469.18 ;
      RECT 19475.9 2897.18 19567.9 2989.18 ;
      RECT 19454.5 2918.18 19567.9 2968.18 ;
      RECT 19454.5 2937.18 19691.9 2949.18 ;
      RECT 19475.9 3377.18 19567.9 3469.18 ;
      RECT 19454.5 3398.18 19567.9 3448.18 ;
      RECT 19454.5 3417.18 19691.9 3429.18 ;
      RECT 19475.9 3857.18 19567.9 3949.18 ;
      RECT 19454.5 3878.18 19567.9 3928.18 ;
      RECT 19454.5 3897.18 19691.9 3909.18 ;
      RECT 19475.9 4337.18 19567.9 4429.18 ;
      RECT 19454.5 4358.18 19567.9 4408.18 ;
      RECT 19454.5 4377.18 19691.9 4389.18 ;
      RECT 19475.9 4817.18 19567.9 4909.18 ;
      RECT 19454.5 4838.18 19567.9 4888.18 ;
      RECT 19454.5 4857.18 19691.9 4869.18 ;
      RECT 19475.9 5297.18 19567.9 5389.18 ;
      RECT 19454.5 5318.18 19567.9 5368.18 ;
      RECT 19454.5 5337.18 19691.9 5349.18 ;
      RECT 19475.9 5777.18 19567.9 5869.18 ;
      RECT 19454.5 5798.18 19567.9 5848.18 ;
      RECT 19454.5 5817.18 19691.9 5829.18 ;
      RECT 19475.9 6257.18 19567.9 6349.18 ;
      RECT 19454.5 6278.18 19567.9 6328.18 ;
      RECT 19454.5 6297.18 19691.9 6309.18 ;
      RECT 19475.9 6737.18 19567.9 6829.18 ;
      RECT 19454.5 6758.18 19567.9 6808.18 ;
      RECT 19454.5 6777.18 19691.9 6789.18 ;
      RECT 19475.9 7217.18 19567.9 7309.18 ;
      RECT 19454.5 7238.18 19567.9 7288.18 ;
      RECT 19454.5 7257.18 19691.9 7269.18 ;
      RECT 19475.9 7697.18 19567.9 7789.18 ;
      RECT 19454.5 7718.18 19567.9 7768.18 ;
      RECT 19454.5 7737.18 19691.9 7749.18 ;
      RECT 19475.9 8177.18 19567.9 8269.18 ;
      RECT 19454.5 8198.18 19567.9 8248.18 ;
      RECT 19454.5 8217.18 19691.9 8229.18 ;
      RECT 19475.9 8657.18 19567.9 8749.18 ;
      RECT 19454.5 8678.18 19567.9 8728.18 ;
      RECT 19454.5 8697.18 19691.9 8709.18 ;
      RECT 19475.9 9137.18 19567.9 9229.18 ;
      RECT 19454.5 9158.18 19567.9 9208.18 ;
      RECT 19454.5 9177.18 19691.9 9189.18 ;
      RECT 19475.9 737.18 19567.9 829.18 ;
      RECT 19454.5 758.18 19567.9 808.18 ;
      RECT 19454.5 777.18 19679.9 789.18 ;
      RECT 19475.9 977.18 19567.9 1069.18 ;
      RECT 19454.5 998.18 19567.9 1048.18 ;
      RECT 19454.5 1017.18 19679.9 1029.18 ;
      RECT 19040 1292.55 19475.9 1317.55 ;
      RECT 19475.9 1217.18 19567.9 1309.18 ;
      RECT 19040 1284.55 19196.9 1317.55 ;
      RECT 19161.9 1238.18 19196.9 1317.55 ;
      RECT 19040 1288.78 19567.9 1290.55 ;
      RECT 19454.5 1238.18 19567.9 1290.55 ;
      RECT 19161.9 1265.55 19451.3 1290.55 ;
      RECT 19454.5 1257.18 19679.9 1269.18 ;
      RECT 19161.9 1238.18 19451.3 1263.55 ;
      RECT 19475.9 1817.18 19567.9 1909.18 ;
      RECT 19454.5 1838.18 19567.9 1888.18 ;
      RECT 19454.5 1857.18 19679.9 1869.18 ;
      RECT 19475.9 2297.18 19567.9 2389.18 ;
      RECT 19454.5 2318.18 19567.9 2368.18 ;
      RECT 19454.5 2337.18 19679.9 2349.18 ;
      RECT 19475.9 2777.18 19567.9 2869.18 ;
      RECT 19454.5 2798.18 19567.9 2848.18 ;
      RECT 19454.5 2817.18 19679.9 2829.18 ;
      RECT 19475.9 3257.18 19567.9 3349.18 ;
      RECT 19454.5 3278.18 19567.9 3328.18 ;
      RECT 19454.5 3297.18 19679.9 3309.18 ;
      RECT 19475.9 3737.18 19567.9 3829.18 ;
      RECT 19454.5 3758.18 19567.9 3808.18 ;
      RECT 19454.5 3777.18 19679.9 3789.18 ;
      RECT 19475.9 4217.18 19567.9 4309.18 ;
      RECT 19454.5 4238.18 19567.9 4288.18 ;
      RECT 19454.5 4257.18 19679.9 4269.18 ;
      RECT 19475.9 4697.18 19567.9 4789.18 ;
      RECT 19454.5 4718.18 19567.9 4768.18 ;
      RECT 19454.5 4737.18 19679.9 4749.18 ;
      RECT 19475.9 5177.18 19567.9 5269.18 ;
      RECT 19454.5 5198.18 19567.9 5248.18 ;
      RECT 19454.5 5217.18 19679.9 5229.18 ;
      RECT 19475.9 5657.18 19567.9 5749.18 ;
      RECT 19454.5 5678.18 19567.9 5728.18 ;
      RECT 19454.5 5697.18 19679.9 5709.18 ;
      RECT 19475.9 6137.18 19567.9 6229.18 ;
      RECT 19454.5 6158.18 19567.9 6208.18 ;
      RECT 19454.5 6177.18 19679.9 6189.18 ;
      RECT 19475.9 6617.18 19567.9 6709.18 ;
      RECT 19454.5 6638.18 19567.9 6688.18 ;
      RECT 19454.5 6657.18 19679.9 6669.18 ;
      RECT 19475.9 7097.18 19567.9 7189.18 ;
      RECT 19454.5 7118.18 19567.9 7168.18 ;
      RECT 19454.5 7137.18 19679.9 7149.18 ;
      RECT 19475.9 7577.18 19567.9 7669.18 ;
      RECT 19454.5 7598.18 19567.9 7648.18 ;
      RECT 19454.5 7617.18 19679.9 7629.18 ;
      RECT 19475.9 8057.18 19567.9 8149.18 ;
      RECT 19454.5 8078.18 19567.9 8128.18 ;
      RECT 19454.5 8097.18 19679.9 8109.18 ;
      RECT 19475.9 8537.18 19567.9 8629.18 ;
      RECT 19454.5 8558.18 19567.9 8608.18 ;
      RECT 19454.5 8577.18 19679.9 8589.18 ;
      RECT 19475.9 9017.18 19567.9 9109.18 ;
      RECT 19454.5 9038.18 19567.9 9088.18 ;
      RECT 19454.5 9057.18 19679.9 9069.18 ;
      RECT 19475.9 1697.18 19567.9 1789.18 ;
      RECT 19454.5 1718.18 19567.9 1768.18 ;
      RECT 19454.5 1737.18 19667.905 1749.18 ;
      RECT 19475.9 2177.18 19567.9 2269.18 ;
      RECT 19454.5 2198.18 19567.9 2248.18 ;
      RECT 19454.5 2217.18 19667.905 2229.18 ;
      RECT 19475.9 2657.18 19567.9 2749.18 ;
      RECT 19454.5 2678.18 19567.9 2728.18 ;
      RECT 19454.5 2697.18 19667.905 2709.18 ;
      RECT 19475.9 3137.18 19567.9 3229.18 ;
      RECT 19454.5 3158.18 19567.9 3208.18 ;
      RECT 19454.5 3177.18 19667.905 3189.18 ;
      RECT 19475.9 3617.18 19567.9 3709.18 ;
      RECT 19454.5 3638.18 19567.9 3688.18 ;
      RECT 19454.5 3657.18 19667.905 3669.18 ;
      RECT 19475.9 4097.18 19567.9 4189.18 ;
      RECT 19454.5 4118.18 19567.9 4168.18 ;
      RECT 19454.5 4137.18 19667.905 4149.18 ;
      RECT 19475.9 4577.18 19567.9 4669.18 ;
      RECT 19454.5 4598.18 19567.9 4648.18 ;
      RECT 19454.5 4617.18 19667.905 4629.18 ;
      RECT 19475.9 5057.18 19567.9 5149.18 ;
      RECT 19454.5 5078.18 19567.9 5128.18 ;
      RECT 19454.5 5097.18 19667.905 5109.18 ;
      RECT 19475.9 6017.18 19567.9 6109.18 ;
      RECT 19454.5 6038.18 19567.9 6088.18 ;
      RECT 19454.5 6057.18 19667.905 6069.18 ;
      RECT 19475.9 6497.18 19567.9 6589.18 ;
      RECT 19454.5 6518.18 19567.9 6568.18 ;
      RECT 19454.5 6537.18 19667.905 6549.18 ;
      RECT 19475.9 6977.18 19567.9 7069.18 ;
      RECT 19454.5 6998.18 19567.9 7048.18 ;
      RECT 19454.5 7017.18 19667.905 7029.18 ;
      RECT 19475.9 7457.18 19567.9 7549.18 ;
      RECT 19454.5 7478.18 19567.9 7528.18 ;
      RECT 19454.5 7497.18 19667.905 7509.18 ;
      RECT 19475.9 7937.18 19567.9 8029.18 ;
      RECT 19454.5 7958.18 19567.9 8008.18 ;
      RECT 19454.5 7977.18 19667.905 7989.18 ;
      RECT 19475.9 8417.18 19567.9 8509.18 ;
      RECT 19454.5 8438.18 19567.9 8488.18 ;
      RECT 19454.5 8457.18 19667.905 8469.18 ;
      RECT 19475.9 8897.18 19567.9 8989.18 ;
      RECT 19454.5 8918.18 19567.9 8968.18 ;
      RECT 19454.5 8937.18 19667.905 8949.18 ;
      RECT 19475.9 1577.18 19567.9 1669.18 ;
      RECT 19454.5 1598.18 19567.9 1648.18 ;
      RECT 19454.5 1617.18 19635.9 1629.18 ;
      RECT 19475.9 2057.18 19567.9 2149.18 ;
      RECT 19454.5 2078.18 19567.9 2128.18 ;
      RECT 19454.5 2097.18 19635.9 2109.18 ;
      RECT 19475.9 2537.18 19567.9 2629.18 ;
      RECT 19454.5 2558.18 19567.9 2608.18 ;
      RECT 19454.5 2577.18 19635.9 2589.18 ;
      RECT 19475.9 3017.18 19567.9 3109.18 ;
      RECT 19454.5 3038.18 19567.9 3088.18 ;
      RECT 19454.5 3057.18 19635.9 3069.18 ;
      RECT 19475.9 3497.18 19567.9 3589.18 ;
      RECT 19454.5 3518.18 19567.9 3568.18 ;
      RECT 19454.5 3537.18 19635.9 3549.18 ;
      RECT 19475.9 3977.18 19567.9 4069.18 ;
      RECT 19454.5 3998.18 19567.9 4048.18 ;
      RECT 19454.5 4017.18 19635.9 4029.18 ;
      RECT 19475.9 4457.18 19567.9 4549.18 ;
      RECT 19454.5 4478.18 19567.9 4528.18 ;
      RECT 19454.5 4497.18 19635.9 4509.18 ;
      RECT 19475.9 4937.18 19567.9 5029.18 ;
      RECT 19454.5 4958.18 19567.9 5008.18 ;
      RECT 19454.5 4977.18 19635.9 4989.18 ;
      RECT 19475.9 5897.18 19567.9 5989.18 ;
      RECT 19454.5 5918.18 19567.9 5968.18 ;
      RECT 19454.5 5937.18 19635.9 5949.18 ;
      RECT 19475.9 6377.18 19567.9 6469.18 ;
      RECT 19454.5 6398.18 19567.9 6448.18 ;
      RECT 19454.5 6417.18 19635.9 6429.18 ;
      RECT 19475.9 6857.18 19567.9 6949.18 ;
      RECT 19454.5 6878.18 19567.9 6928.18 ;
      RECT 19454.5 6897.18 19635.9 6909.18 ;
      RECT 19475.9 7337.18 19567.9 7429.18 ;
      RECT 19454.5 7358.18 19567.9 7408.18 ;
      RECT 19454.5 7377.18 19635.9 7389.18 ;
      RECT 19475.9 7817.18 19567.9 7909.18 ;
      RECT 19454.5 7838.18 19567.9 7888.18 ;
      RECT 19454.5 7857.18 19635.9 7869.18 ;
      RECT 19475.9 8297.18 19567.9 8389.18 ;
      RECT 19454.5 8318.18 19567.9 8368.18 ;
      RECT 19454.5 8337.18 19635.9 8349.18 ;
      RECT 19475.9 8777.18 19567.9 8869.18 ;
      RECT 19454.5 8798.18 19567.9 8848.18 ;
      RECT 19454.5 8817.18 19635.9 8829.18 ;
      RECT 19475.9 1457.18 19567.9 1549.18 ;
      RECT 19454.5 1478.18 19567.9 1528.18 ;
      RECT 19475.9 5417.18 19567.9 5509.18 ;
      RECT 19454.5 5438.18 19567.9 5488.18 ;
      RECT 19475.9 5537.18 19567.9 5629.18 ;
      RECT 19454.5 5558.18 19567.9 5608.18 ;
      RECT 19475.9 9257.18 19567.9 9349.18 ;
      RECT 19454.5 9278.18 19567.9 9328.18 ;
      RECT 19161.9 1380.63 19406.9 1381.75 ;
      RECT 19160.9 1380.555 19161.9 1381.675 ;
      RECT 19040 1327.55 19161.9 1360.55 ;
      RECT 19040 1327.55 19246.9 1355.26 ;
      RECT 19158.07 1364.33 19167.84 1365.58 ;
      RECT 19158.07 1364.44 19167.9 1365.44 ;
      RECT 19158.07 1367.31 19167.84 1368.56 ;
      RECT 19158.07 1367.44 19167.9 1368.44 ;
      RECT 724.1 1292.55 1120 1317.55 ;
      RECT 963.1 1284.55 1120 1317.55 ;
      RECT 632.1 1217.18 724.1 1309.18 ;
      RECT 632.1 1288.78 1120 1290.55 ;
      RECT 748.7 1265.55 998.1 1290.55 ;
      RECT 632.1 1238.18 745.5 1290.55 ;
      RECT 520.1 1257.18 745.5 1269.18 ;
      RECT 963.1 1238.18 998.1 1317.55 ;
      RECT 748.7 1238.18 998.1 1263.55 ;
      RECT 793.1 1380.63 998.1 1381.75 ;
      RECT 998.1 1380.555 999.1 1381.675 ;
      RECT 632.1 617.18 724.1 709.18 ;
      RECT 632.1 638.18 745.5 688.18 ;
      RECT 502.095 657.18 745.5 669.18 ;
      RECT 632.1 737.18 724.1 829.18 ;
      RECT 632.1 758.18 745.5 808.18 ;
      RECT 520.1 777.18 745.5 789.18 ;
      RECT 632.1 857.18 724.1 949.18 ;
      RECT 632.1 878.18 745.5 928.18 ;
      RECT 508.1 897.18 745.5 909.18 ;
      RECT 632.1 977.18 724.1 1069.18 ;
      RECT 632.1 998.18 745.5 1048.18 ;
      RECT 520.1 1017.18 745.5 1029.18 ;
      RECT 632.1 1097.18 724.1 1189.18 ;
      RECT 632.1 1118.18 745.5 1168.18 ;
      RECT 508.1 1137.18 745.5 1149.18 ;
      RECT 632.1 1337.18 724.1 1429.18 ;
      RECT 632.1 1358.18 745.5 1408.18 ;
      RECT 508.1 1377.18 745.5 1389.18 ;
      RECT 632.1 1457.18 724.1 1549.18 ;
      RECT 632.1 1478.18 745.5 1528.18 ;
      RECT 632.1 1577.18 724.1 1669.18 ;
      RECT 632.1 1598.18 745.5 1648.18 ;
      RECT 564.1 1617.18 745.5 1629.18 ;
      RECT 632.1 1697.18 724.1 1789.18 ;
      RECT 632.1 1718.18 745.5 1768.18 ;
      RECT 532.095 1737.18 745.5 1749.18 ;
      RECT 632.1 1817.18 724.1 1909.18 ;
      RECT 632.1 1838.18 745.5 1888.18 ;
      RECT 520.1 1857.18 745.5 1869.18 ;
      RECT 632.1 1937.18 724.1 2029.18 ;
      RECT 632.1 1958.18 745.5 2008.18 ;
      RECT 508.1 1977.18 745.5 1989.18 ;
      RECT 632.1 2057.18 724.1 2149.18 ;
      RECT 632.1 2078.18 745.5 2128.18 ;
      RECT 564.1 2097.18 745.5 2109.18 ;
      RECT 632.1 2177.18 724.1 2269.18 ;
      RECT 632.1 2198.18 745.5 2248.18 ;
      RECT 532.095 2217.18 745.5 2229.18 ;
      RECT 632.1 2297.18 724.1 2389.18 ;
      RECT 632.1 2318.18 745.5 2368.18 ;
      RECT 520.1 2337.18 745.5 2349.18 ;
      RECT 632.1 2417.18 724.1 2509.18 ;
      RECT 632.1 2438.18 745.5 2488.18 ;
      RECT 508.1 2457.18 745.5 2469.18 ;
      RECT 632.1 2537.18 724.1 2629.18 ;
      RECT 632.1 2558.18 745.5 2608.18 ;
      RECT 564.1 2577.18 745.5 2589.18 ;
      RECT 632.1 2657.18 724.1 2749.18 ;
      RECT 632.1 2678.18 745.5 2728.18 ;
      RECT 532.095 2697.18 745.5 2709.18 ;
      RECT 632.1 2777.18 724.1 2869.18 ;
      RECT 632.1 2798.18 745.5 2848.18 ;
      RECT 520.1 2817.18 745.5 2829.18 ;
      RECT 632.1 2897.18 724.1 2989.18 ;
      RECT 632.1 2918.18 745.5 2968.18 ;
      RECT 508.1 2937.18 745.5 2949.18 ;
      RECT 632.1 3017.18 724.1 3109.18 ;
      RECT 632.1 3038.18 745.5 3088.18 ;
      RECT 564.1 3057.18 745.5 3069.18 ;
      RECT 632.1 3137.18 724.1 3229.18 ;
      RECT 632.1 3158.18 745.5 3208.18 ;
      RECT 532.095 3177.18 745.5 3189.18 ;
      RECT 632.1 3257.18 724.1 3349.18 ;
      RECT 632.1 3278.18 745.5 3328.18 ;
      RECT 520.1 3297.18 745.5 3309.18 ;
      RECT 632.1 3377.18 724.1 3469.18 ;
      RECT 632.1 3398.18 745.5 3448.18 ;
      RECT 508.1 3417.18 745.5 3429.18 ;
      RECT 632.1 3497.18 724.1 3589.18 ;
      RECT 632.1 3518.18 745.5 3568.18 ;
      RECT 564.1 3537.18 745.5 3549.18 ;
      RECT 632.1 3617.18 724.1 3709.18 ;
      RECT 632.1 3638.18 745.5 3688.18 ;
      RECT 532.095 3657.18 745.5 3669.18 ;
      RECT 632.1 3737.18 724.1 3829.18 ;
      RECT 632.1 3758.18 745.5 3808.18 ;
      RECT 520.1 3777.18 745.5 3789.18 ;
      RECT 632.1 3857.18 724.1 3949.18 ;
      RECT 632.1 3878.18 745.5 3928.18 ;
      RECT 508.1 3897.18 745.5 3909.18 ;
      RECT 632.1 3977.18 724.1 4069.18 ;
      RECT 632.1 3998.18 745.5 4048.18 ;
      RECT 564.1 4017.18 745.5 4029.18 ;
      RECT 632.1 4097.18 724.1 4189.18 ;
      RECT 632.1 4118.18 745.5 4168.18 ;
      RECT 532.095 4137.18 745.5 4149.18 ;
      RECT 632.1 4217.18 724.1 4309.18 ;
      RECT 632.1 4238.18 745.5 4288.18 ;
      RECT 520.1 4257.18 745.5 4269.18 ;
      RECT 632.1 4337.18 724.1 4429.18 ;
      RECT 632.1 4358.18 745.5 4408.18 ;
      RECT 508.1 4377.18 745.5 4389.18 ;
      RECT 632.1 4457.18 724.1 4549.18 ;
      RECT 632.1 4478.18 745.5 4528.18 ;
      RECT 564.1 4497.18 745.5 4509.18 ;
      RECT 632.1 4577.18 724.1 4669.18 ;
      RECT 632.1 4598.18 745.5 4648.18 ;
      RECT 532.095 4617.18 745.5 4629.18 ;
      RECT 632.1 4697.18 724.1 4789.18 ;
      RECT 632.1 4718.18 745.5 4768.18 ;
      RECT 520.1 4737.18 745.5 4749.18 ;
      RECT 632.1 4817.18 724.1 4909.18 ;
      RECT 632.1 4838.18 745.5 4888.18 ;
      RECT 508.1 4857.18 745.5 4869.18 ;
      RECT 632.1 4937.18 724.1 5029.18 ;
      RECT 632.1 4958.18 745.5 5008.18 ;
      RECT 564.1 4977.18 745.5 4989.18 ;
      RECT 632.1 5057.18 724.1 5149.18 ;
      RECT 632.1 5078.18 745.5 5128.18 ;
      RECT 532.095 5097.18 745.5 5109.18 ;
      RECT 632.1 5177.18 724.1 5269.18 ;
      RECT 632.1 5198.18 745.5 5248.18 ;
      RECT 520.1 5217.18 745.5 5229.18 ;
      RECT 632.1 5297.18 724.1 5389.18 ;
      RECT 632.1 5318.18 745.5 5368.18 ;
      RECT 508.1 5337.18 745.5 5349.18 ;
      RECT 632.1 5417.18 724.1 5509.18 ;
      RECT 632.1 5438.18 745.5 5488.18 ;
      RECT 632.1 5537.18 724.1 5629.18 ;
      RECT 632.1 5558.18 745.5 5608.18 ;
      RECT 532.095 5577.18 745.5 5589.18 ;
      RECT 632.1 5657.18 724.1 5749.18 ;
      RECT 632.1 5678.18 745.5 5728.18 ;
      RECT 520.1 5697.18 745.5 5709.18 ;
      RECT 632.1 5777.18 724.1 5869.18 ;
      RECT 632.1 5798.18 745.5 5848.18 ;
      RECT 508.1 5817.18 745.5 5829.18 ;
      RECT 632.1 5897.18 724.1 5989.18 ;
      RECT 632.1 5918.18 745.5 5968.18 ;
      RECT 564.1 5937.18 745.5 5949.18 ;
      RECT 632.1 6017.18 724.1 6109.18 ;
      RECT 632.1 6038.18 745.5 6088.18 ;
      RECT 532.095 6057.18 745.5 6069.18 ;
      RECT 632.1 6137.18 724.1 6229.18 ;
      RECT 632.1 6158.18 745.5 6208.18 ;
      RECT 520.1 6177.18 745.5 6189.18 ;
      RECT 632.1 6257.18 724.1 6349.18 ;
      RECT 632.1 6278.18 745.5 6328.18 ;
      RECT 508.1 6297.18 745.5 6309.18 ;
      RECT 632.1 6377.18 724.1 6469.18 ;
      RECT 632.1 6398.18 745.5 6448.18 ;
      RECT 564.1 6417.18 745.5 6429.18 ;
      RECT 632.1 6497.18 724.1 6589.18 ;
      RECT 632.1 6518.18 745.5 6568.18 ;
      RECT 532.095 6537.18 745.5 6549.18 ;
      RECT 632.1 6617.18 724.1 6709.18 ;
      RECT 632.1 6638.18 745.5 6688.18 ;
      RECT 520.1 6657.18 745.5 6669.18 ;
      RECT 632.1 6737.18 724.1 6829.18 ;
      RECT 632.1 6758.18 745.5 6808.18 ;
      RECT 508.1 6777.18 745.5 6789.18 ;
      RECT 632.1 6857.18 724.1 6949.18 ;
      RECT 632.1 6878.18 745.5 6928.18 ;
      RECT 564.1 6897.18 745.5 6909.18 ;
      RECT 632.1 6977.18 724.1 7069.18 ;
      RECT 632.1 6998.18 745.5 7048.18 ;
      RECT 532.095 7017.18 745.5 7029.18 ;
      RECT 632.1 7097.18 724.1 7189.18 ;
      RECT 632.1 7118.18 745.5 7168.18 ;
      RECT 520.1 7137.18 745.5 7149.18 ;
      RECT 632.1 7217.18 724.1 7309.18 ;
      RECT 632.1 7238.18 745.5 7288.18 ;
      RECT 508.1 7257.18 745.5 7269.18 ;
      RECT 632.1 7337.18 724.1 7429.18 ;
      RECT 632.1 7358.18 745.5 7408.18 ;
      RECT 564.1 7377.18 745.5 7389.18 ;
      RECT 632.1 7457.18 724.1 7549.18 ;
      RECT 632.1 7478.18 745.5 7528.18 ;
      RECT 532.095 7497.18 745.5 7509.18 ;
      RECT 632.1 7577.18 724.1 7669.18 ;
      RECT 632.1 7598.18 745.5 7648.18 ;
      RECT 520.1 7617.18 745.5 7629.18 ;
      RECT 632.1 7697.18 724.1 7789.18 ;
      RECT 632.1 7718.18 745.5 7768.18 ;
      RECT 508.1 7737.18 745.5 7749.18 ;
      RECT 632.1 7817.18 724.1 7909.18 ;
      RECT 632.1 7838.18 745.5 7888.18 ;
      RECT 564.1 7857.18 745.5 7869.18 ;
      RECT 632.1 7937.18 724.1 8029.18 ;
      RECT 632.1 7958.18 745.5 8008.18 ;
      RECT 532.095 7977.18 745.5 7989.18 ;
      RECT 632.1 8057.18 724.1 8149.18 ;
      RECT 632.1 8078.18 745.5 8128.18 ;
      RECT 520.1 8097.18 745.5 8109.18 ;
      RECT 632.1 8177.18 724.1 8269.18 ;
      RECT 632.1 8198.18 745.5 8248.18 ;
      RECT 508.1 8217.18 745.5 8229.18 ;
      RECT 632.1 8297.18 724.1 8389.18 ;
      RECT 632.1 8318.18 745.5 8368.18 ;
      RECT 564.1 8337.18 745.5 8349.18 ;
      RECT 632.1 8417.18 724.1 8509.18 ;
      RECT 632.1 8438.18 745.5 8488.18 ;
      RECT 532.095 8457.18 745.5 8469.18 ;
      RECT 632.1 8537.18 724.1 8629.18 ;
      RECT 632.1 8558.18 745.5 8608.18 ;
      RECT 520.1 8577.18 745.5 8589.18 ;
      RECT 632.1 8657.18 724.1 8749.18 ;
      RECT 632.1 8678.18 745.5 8728.18 ;
      RECT 508.1 8697.18 745.5 8709.18 ;
      RECT 632.1 8777.18 724.1 8869.18 ;
      RECT 632.1 8798.18 745.5 8848.18 ;
      RECT 564.1 8817.18 745.5 8829.18 ;
      RECT 632.1 8897.18 724.1 8989.18 ;
      RECT 632.1 8918.18 745.5 8968.18 ;
      RECT 532.095 8937.18 745.5 8949.18 ;
      RECT 632.1 9017.18 724.1 9109.18 ;
      RECT 632.1 9038.18 745.5 9088.18 ;
      RECT 520.1 9057.18 745.5 9069.18 ;
      RECT 632.1 9137.18 724.1 9229.18 ;
      RECT 632.1 9158.18 745.5 9208.18 ;
      RECT 508.1 9177.18 745.5 9189.18 ;
      RECT 632.1 9257.18 724.1 9349.18 ;
      RECT 632.1 9278.18 745.5 9328.18 ;
      RECT 632.1 9377.18 724.1 9469.18 ;
      RECT 632.1 9398.18 745.5 9448.18 ;
      RECT 502.095 9417.18 745.5 9429.18 ;
      RECT 502.1 677.18 594.1 769.18 ;
      RECT 502.1 680.155 615.5 715.155 ;
      RECT 502.1 797.18 594.1 889.18 ;
      RECT 502.1 800.155 615.5 835.155 ;
      RECT 502.1 917.18 594.1 1009.18 ;
      RECT 502.1 920.155 615.5 955.155 ;
      RECT 502.1 1037.18 594.1 1129.18 ;
      RECT 502.1 1040.155 615.5 1075.155 ;
      RECT 502.1 1157.18 594.1 1249.18 ;
      RECT 502.1 1160.155 615.5 1195.155 ;
      RECT 502.1 1277.18 594.1 1369.18 ;
      RECT 502.1 1298.18 615.5 1348.18 ;
      RECT 502.1 8717.18 594.1 8809.18 ;
      RECT 502.1 8720.155 615.5 8755.155 ;
      RECT 502.1 8837.18 594.1 8929.18 ;
      RECT 502.1 8840.155 615.5 8875.155 ;
      RECT 502.1 8957.18 594.1 9049.18 ;
      RECT 502.1 8960.155 615.5 8995.155 ;
      RECT 502.1 9077.18 594.1 9169.18 ;
      RECT 502.1 9080.155 615.5 9115.155 ;
      RECT 502.1 9197.18 594.1 9289.18 ;
      RECT 502.1 9200.155 615.5 9235.155 ;
      RECT 502.1 9317.18 594.1 9409.18 ;
      RECT 502.1 9320.155 615.5 9355.155 ;
      RECT 19160.9 1050.27 19446.9 1052.27 ;
      RECT 19160.9 1371.26 19446.9 1373.26 ;
      RECT 753.1 9470.56 19446.9 9472.56 ;
      RECT 19160.9 1408.19 19406.9 1409.31 ;
      RECT 19160.9 1452.63 19406.9 1453.75 ;
      RECT 19160.9 1480.19 19406.9 1481.31 ;
      RECT 19160.9 1524.63 19406.9 1525.75 ;
      RECT 19160.9 1552.19 19406.9 1553.31 ;
      RECT 19160.9 1596.63 19406.9 1597.75 ;
      RECT 19160.9 1624.19 19406.9 1625.31 ;
      RECT 19160.9 1668.63 19406.9 1669.75 ;
      RECT 19160.9 1696.19 19406.9 1697.31 ;
      RECT 19160.9 1740.63 19406.9 1741.75 ;
      RECT 19160.9 1768.19 19406.9 1769.31 ;
      RECT 19160.9 1812.63 19406.9 1813.75 ;
      RECT 19160.9 1840.19 19406.9 1841.31 ;
      RECT 19160.9 1884.63 19406.9 1885.75 ;
      RECT 19160.9 1912.19 19406.9 1913.31 ;
      RECT 19160.9 1956.63 19406.9 1957.75 ;
      RECT 19160.9 1984.19 19406.9 1985.31 ;
      RECT 19160.9 2028.63 19406.9 2029.75 ;
      RECT 19160.9 2056.19 19406.9 2057.31 ;
      RECT 19160.9 2100.63 19406.9 2101.75 ;
      RECT 19160.9 2128.19 19406.9 2129.31 ;
      RECT 19160.9 2172.63 19406.9 2173.75 ;
      RECT 19160.9 2200.19 19406.9 2201.31 ;
      RECT 19160.9 2244.63 19406.9 2245.75 ;
      RECT 19160.9 2272.19 19406.9 2273.31 ;
      RECT 19160.9 2316.63 19406.9 2317.75 ;
      RECT 19160.9 2344.19 19406.9 2345.31 ;
      RECT 19160.9 2388.63 19406.9 2389.75 ;
      RECT 19160.9 2416.19 19406.9 2417.31 ;
      RECT 19160.9 2460.63 19406.9 2461.75 ;
      RECT 19160.9 2488.19 19406.9 2489.31 ;
      RECT 19160.9 2532.63 19406.9 2533.75 ;
      RECT 19160.9 2560.19 19406.9 2561.31 ;
      RECT 19160.9 2604.63 19406.9 2605.75 ;
      RECT 19160.9 2632.19 19406.9 2633.31 ;
      RECT 19160.9 2676.63 19406.9 2677.75 ;
      RECT 19160.9 2704.19 19406.9 2705.31 ;
      RECT 19160.9 2748.63 19406.9 2749.75 ;
      RECT 19160.9 2776.19 19406.9 2777.31 ;
      RECT 19160.9 2820.63 19406.9 2821.75 ;
      RECT 19160.9 2848.19 19406.9 2849.31 ;
      RECT 19160.9 2892.63 19406.9 2893.75 ;
      RECT 19160.9 2920.19 19406.9 2921.31 ;
      RECT 19160.9 2964.63 19406.9 2965.75 ;
      RECT 19160.9 2992.19 19406.9 2993.31 ;
      RECT 19160.9 3036.63 19406.9 3037.75 ;
      RECT 19160.9 3064.19 19406.9 3065.31 ;
      RECT 19160.9 3108.63 19406.9 3109.75 ;
      RECT 19160.9 3136.19 19406.9 3137.31 ;
      RECT 19160.9 3180.63 19406.9 3181.75 ;
      RECT 19160.9 3208.19 19406.9 3209.31 ;
      RECT 19160.9 3252.63 19406.9 3253.75 ;
      RECT 19160.9 3280.19 19406.9 3281.31 ;
      RECT 19160.9 3324.63 19406.9 3325.75 ;
      RECT 19160.9 3352.19 19406.9 3353.31 ;
      RECT 19160.9 3396.63 19406.9 3397.75 ;
      RECT 19160.9 3424.19 19406.9 3425.31 ;
      RECT 19160.9 3468.63 19406.9 3469.75 ;
      RECT 19160.9 3496.19 19406.9 3497.31 ;
      RECT 19160.9 3540.63 19406.9 3541.75 ;
      RECT 19160.9 3568.19 19406.9 3569.31 ;
      RECT 19160.9 3612.63 19406.9 3613.75 ;
      RECT 19160.9 3640.19 19406.9 3641.31 ;
      RECT 19160.9 3684.63 19406.9 3685.75 ;
      RECT 19160.9 3712.19 19406.9 3713.31 ;
      RECT 19160.9 3756.63 19406.9 3757.75 ;
      RECT 19160.9 3784.19 19406.9 3785.31 ;
      RECT 19160.9 3828.63 19406.9 3829.75 ;
      RECT 19160.9 3856.19 19406.9 3857.31 ;
      RECT 19160.9 3900.63 19406.9 3901.75 ;
      RECT 19160.9 3928.19 19406.9 3929.31 ;
      RECT 19160.9 3972.63 19406.9 3973.75 ;
      RECT 19160.9 4000.19 19406.9 4001.31 ;
      RECT 19160.9 4044.63 19406.9 4045.75 ;
      RECT 19160.9 4072.19 19406.9 4073.31 ;
      RECT 19160.9 4116.63 19406.9 4117.75 ;
      RECT 19160.9 4144.19 19406.9 4145.31 ;
      RECT 19160.9 4188.63 19406.9 4189.75 ;
      RECT 19160.9 4216.19 19406.9 4217.31 ;
      RECT 19160.9 4260.63 19406.9 4261.75 ;
      RECT 19160.9 4288.19 19406.9 4289.31 ;
      RECT 19160.9 4332.63 19406.9 4333.75 ;
      RECT 19160.9 4360.19 19406.9 4361.31 ;
      RECT 19160.9 4404.63 19406.9 4405.75 ;
      RECT 19160.9 4432.19 19406.9 4433.31 ;
      RECT 19160.9 4476.63 19406.9 4477.75 ;
      RECT 19160.9 4504.19 19406.9 4505.31 ;
      RECT 19160.9 4548.63 19406.9 4549.75 ;
      RECT 19160.9 4576.19 19406.9 4577.31 ;
      RECT 19160.9 4620.63 19406.9 4621.75 ;
      RECT 19160.9 4648.19 19406.9 4649.31 ;
      RECT 19160.9 4692.63 19406.9 4693.75 ;
      RECT 19160.9 4720.19 19406.9 4721.31 ;
      RECT 19160.9 4764.63 19406.9 4765.75 ;
      RECT 19160.9 4792.19 19406.9 4793.31 ;
      RECT 19160.9 4836.63 19406.9 4837.75 ;
      RECT 19160.9 4864.19 19406.9 4865.31 ;
      RECT 19160.9 4908.63 19406.9 4909.75 ;
      RECT 19160.9 4936.19 19406.9 4937.31 ;
      RECT 19160.9 4980.63 19406.9 4981.75 ;
      RECT 19160.9 5008.19 19406.9 5009.31 ;
      RECT 19160.9 5052.63 19406.9 5053.75 ;
      RECT 19160.9 5080.19 19406.9 5081.31 ;
      RECT 19160.9 5124.63 19406.9 5125.75 ;
      RECT 19160.9 5152.19 19406.9 5153.31 ;
      RECT 19160.9 5196.63 19406.9 5197.75 ;
      RECT 19160.9 5224.19 19406.9 5225.31 ;
      RECT 19160.9 5268.63 19406.9 5269.75 ;
      RECT 19160.9 5296.19 19406.9 5297.31 ;
      RECT 19160.9 5340.63 19406.9 5341.75 ;
      RECT 19160.9 5368.19 19406.9 5369.31 ;
      RECT 19160.9 5412.63 19406.9 5413.75 ;
      RECT 19160.9 5440.19 19406.9 5441.31 ;
      RECT 19160.9 5484.63 19406.9 5485.75 ;
      RECT 19160.9 5512.19 19406.9 5513.31 ;
      RECT 19160.9 5556.63 19406.9 5557.75 ;
      RECT 19160.9 5584.19 19406.9 5585.31 ;
      RECT 19160.9 5628.63 19406.9 5629.75 ;
      RECT 19160.9 5656.19 19406.9 5657.31 ;
      RECT 19160.9 5700.63 19406.9 5701.75 ;
      RECT 19160.9 5728.19 19406.9 5729.31 ;
      RECT 19160.9 5772.63 19406.9 5773.75 ;
      RECT 19160.9 5800.19 19406.9 5801.31 ;
      RECT 19160.9 5844.63 19406.9 5845.75 ;
      RECT 19160.9 5872.19 19406.9 5873.31 ;
      RECT 19160.9 5916.63 19406.9 5917.75 ;
      RECT 19160.9 5944.19 19406.9 5945.31 ;
      RECT 19160.9 5988.63 19406.9 5989.75 ;
      RECT 19160.9 6016.19 19406.9 6017.31 ;
      RECT 19160.9 6060.63 19406.9 6061.75 ;
      RECT 19160.9 6088.19 19406.9 6089.31 ;
      RECT 19160.9 6132.63 19406.9 6133.75 ;
      RECT 19160.9 6160.19 19406.9 6161.31 ;
      RECT 19160.9 6204.63 19406.9 6205.75 ;
      RECT 19160.9 6232.19 19406.9 6233.31 ;
      RECT 19160.9 6276.63 19406.9 6277.75 ;
      RECT 19160.9 6304.19 19406.9 6305.31 ;
      RECT 19160.9 6348.63 19406.9 6349.75 ;
      RECT 19160.9 6376.19 19406.9 6377.31 ;
      RECT 19160.9 6420.63 19406.9 6421.75 ;
      RECT 19160.9 6448.19 19406.9 6449.31 ;
      RECT 19160.9 6492.63 19406.9 6493.75 ;
      RECT 19160.9 6520.19 19406.9 6521.31 ;
      RECT 19160.9 6564.63 19406.9 6565.75 ;
      RECT 19160.9 6592.19 19406.9 6593.31 ;
      RECT 19160.9 6636.63 19406.9 6637.75 ;
      RECT 19160.9 6664.19 19406.9 6665.31 ;
      RECT 19160.9 6708.63 19406.9 6709.75 ;
      RECT 19160.9 6736.19 19406.9 6737.31 ;
      RECT 19160.9 6780.63 19406.9 6781.75 ;
      RECT 19160.9 6808.19 19406.9 6809.31 ;
      RECT 19160.9 6852.63 19406.9 6853.75 ;
      RECT 19160.9 6880.19 19406.9 6881.31 ;
      RECT 19160.9 6924.63 19406.9 6925.75 ;
      RECT 19160.9 6952.19 19406.9 6953.31 ;
      RECT 19160.9 6996.63 19406.9 6997.75 ;
      RECT 19160.9 7024.19 19406.9 7025.31 ;
      RECT 19160.9 7068.63 19406.9 7069.75 ;
      RECT 19160.9 7096.19 19406.9 7097.31 ;
      RECT 19160.9 7140.63 19406.9 7141.75 ;
      RECT 19160.9 7168.19 19406.9 7169.31 ;
      RECT 19160.9 7212.63 19406.9 7213.75 ;
      RECT 19160.9 7240.19 19406.9 7241.31 ;
      RECT 19160.9 7284.63 19406.9 7285.75 ;
      RECT 19160.9 7312.19 19406.9 7313.31 ;
      RECT 19160.9 7356.63 19406.9 7357.75 ;
      RECT 19160.9 7384.19 19406.9 7385.31 ;
      RECT 19160.9 7428.63 19406.9 7429.75 ;
      RECT 19160.9 7456.19 19406.9 7457.31 ;
      RECT 19160.9 7500.63 19406.9 7501.75 ;
      RECT 19160.9 7528.19 19406.9 7529.31 ;
      RECT 19160.9 7572.63 19406.9 7573.75 ;
      RECT 19160.9 7600.19 19406.9 7601.31 ;
      RECT 19160.9 7644.63 19406.9 7645.75 ;
      RECT 19160.9 7672.19 19406.9 7673.31 ;
      RECT 19160.9 7716.63 19406.9 7717.75 ;
      RECT 19160.9 7744.19 19406.9 7745.31 ;
      RECT 19160.9 7788.63 19406.9 7789.75 ;
      RECT 19160.9 7816.19 19406.9 7817.31 ;
      RECT 19160.9 7860.63 19406.9 7861.75 ;
      RECT 19160.9 7888.19 19406.9 7889.31 ;
      RECT 19160.9 7932.63 19406.9 7933.75 ;
      RECT 19160.9 7960.19 19406.9 7961.31 ;
      RECT 19160.9 8004.63 19406.9 8005.75 ;
      RECT 19160.9 8032.19 19406.9 8033.31 ;
      RECT 19160.9 8076.63 19406.9 8077.75 ;
      RECT 19160.9 8104.19 19406.9 8105.31 ;
      RECT 19160.9 8148.63 19406.9 8149.75 ;
      RECT 19160.9 8176.19 19406.9 8177.31 ;
      RECT 19160.9 8220.63 19406.9 8221.75 ;
      RECT 19160.9 8248.19 19406.9 8249.31 ;
      RECT 19160.9 8292.63 19406.9 8293.75 ;
      RECT 19160.9 8320.19 19406.9 8321.31 ;
      RECT 19160.9 8364.63 19406.9 8365.75 ;
      RECT 19160.9 8392.19 19406.9 8393.31 ;
      RECT 19160.9 8436.63 19406.9 8437.75 ;
      RECT 19160.9 8464.19 19406.9 8465.31 ;
      RECT 19160.9 8508.63 19406.9 8509.75 ;
      RECT 19160.9 8536.19 19406.9 8537.31 ;
      RECT 19160.9 8580.63 19406.9 8581.75 ;
      RECT 19160.9 8608.19 19406.9 8609.31 ;
      RECT 19160.9 8652.63 19406.9 8653.75 ;
      RECT 19160.9 8680.19 19406.9 8681.31 ;
      RECT 19160.9 8724.63 19406.9 8725.75 ;
      RECT 19160.9 8752.19 19406.9 8753.31 ;
      RECT 19160.9 8796.63 19406.9 8797.75 ;
      RECT 19160.9 8824.19 19406.9 8825.31 ;
      RECT 19160.9 8868.63 19406.9 8869.75 ;
      RECT 19160.9 8896.19 19406.9 8897.31 ;
      RECT 19160.9 8940.63 19406.9 8941.75 ;
      RECT 19160.9 8968.19 19406.9 8969.31 ;
      RECT 19160.9 9012.63 19406.9 9013.75 ;
      RECT 19160.9 9040.19 19406.9 9041.31 ;
      RECT 19160.9 9084.63 19406.9 9085.75 ;
      RECT 19160.9 9112.19 19406.9 9113.31 ;
      RECT 19160.9 9156.63 19406.9 9157.75 ;
      RECT 19160.9 9184.19 19406.9 9185.31 ;
      RECT 19160.9 9228.63 19406.9 9229.75 ;
      RECT 19160.9 9256.19 19406.9 9257.31 ;
      RECT 19160.9 9300.63 19406.9 9301.75 ;
      RECT 19160.9 9328.19 19406.9 9329.31 ;
      RECT 19160.9 9372.63 19406.9 9373.75 ;
      RECT 19160.9 9400.19 19406.9 9401.31 ;
      RECT 19160.9 9444.63 19406.9 9445.75 ;
      RECT 19160.4 1411.31 19366.9 1411.87 ;
      RECT 19160.4 1450.07 19366.9 1450.63 ;
      RECT 19160.4 1483.31 19366.9 1483.87 ;
      RECT 19160.4 1522.07 19366.9 1522.63 ;
      RECT 19160.4 1555.31 19366.9 1555.87 ;
      RECT 19160.4 1594.07 19366.9 1594.63 ;
      RECT 19160.4 1627.31 19366.9 1627.87 ;
      RECT 19160.4 1666.07 19366.9 1666.63 ;
      RECT 19160.4 1699.31 19366.9 1699.87 ;
      RECT 19160.4 1738.07 19366.9 1738.63 ;
      RECT 19160.4 1771.31 19366.9 1771.87 ;
      RECT 19160.4 1810.07 19366.9 1810.63 ;
      RECT 19160.4 1843.31 19366.9 1843.87 ;
      RECT 19160.4 1882.07 19366.9 1882.63 ;
      RECT 19160.4 1915.31 19366.9 1915.87 ;
      RECT 19160.4 1954.07 19366.9 1954.63 ;
      RECT 19160.4 1987.31 19366.9 1987.87 ;
      RECT 19160.4 2026.07 19366.9 2026.63 ;
      RECT 19160.4 2059.31 19366.9 2059.87 ;
      RECT 19160.4 2098.07 19366.9 2098.63 ;
      RECT 19160.4 2131.31 19366.9 2131.87 ;
      RECT 19160.4 2170.07 19366.9 2170.63 ;
      RECT 19160.4 2203.31 19366.9 2203.87 ;
      RECT 19160.4 2242.07 19366.9 2242.63 ;
      RECT 19160.4 2275.31 19366.9 2275.87 ;
      RECT 19160.4 2314.07 19366.9 2314.63 ;
      RECT 19160.4 2347.31 19366.9 2347.87 ;
      RECT 19160.4 2386.07 19366.9 2386.63 ;
      RECT 19160.4 2419.31 19366.9 2419.87 ;
      RECT 19160.4 2458.07 19366.9 2458.63 ;
      RECT 19160.4 2491.31 19366.9 2491.87 ;
      RECT 19160.4 2530.07 19366.9 2530.63 ;
      RECT 19160.4 2563.31 19366.9 2563.87 ;
      RECT 19160.4 2602.07 19366.9 2602.63 ;
      RECT 19160.4 2635.31 19366.9 2635.87 ;
      RECT 19160.4 2674.07 19366.9 2674.63 ;
      RECT 19160.4 2707.31 19366.9 2707.87 ;
      RECT 19160.4 2746.07 19366.9 2746.63 ;
      RECT 19160.4 2779.31 19366.9 2779.87 ;
      RECT 19160.4 2818.07 19366.9 2818.63 ;
      RECT 19160.4 2851.31 19366.9 2851.87 ;
      RECT 19160.4 2890.07 19366.9 2890.63 ;
      RECT 19160.4 2923.31 19366.9 2923.87 ;
      RECT 19160.4 2962.07 19366.9 2962.63 ;
      RECT 19160.4 2995.31 19366.9 2995.87 ;
      RECT 19160.4 3034.07 19366.9 3034.63 ;
      RECT 19160.4 3067.31 19366.9 3067.87 ;
      RECT 19160.4 3106.07 19366.9 3106.63 ;
      RECT 19160.4 3139.31 19366.9 3139.87 ;
      RECT 19160.4 3178.07 19366.9 3178.63 ;
      RECT 19160.4 3211.31 19366.9 3211.87 ;
      RECT 19160.4 3250.07 19366.9 3250.63 ;
      RECT 19160.4 3283.31 19366.9 3283.87 ;
      RECT 19160.4 3322.07 19366.9 3322.63 ;
      RECT 19160.4 3355.31 19366.9 3355.87 ;
      RECT 19160.4 3394.07 19366.9 3394.63 ;
      RECT 19160.4 3427.31 19366.9 3427.87 ;
      RECT 19160.4 3466.07 19366.9 3466.63 ;
      RECT 19160.4 3499.31 19366.9 3499.87 ;
      RECT 19160.4 3538.07 19366.9 3538.63 ;
      RECT 19160.4 3571.31 19366.9 3571.87 ;
      RECT 19160.4 3610.07 19366.9 3610.63 ;
      RECT 19160.4 3643.31 19366.9 3643.87 ;
      RECT 19160.4 3682.07 19366.9 3682.63 ;
      RECT 19160.4 3715.31 19366.9 3715.87 ;
      RECT 19160.4 3754.07 19366.9 3754.63 ;
      RECT 19160.4 3787.31 19366.9 3787.87 ;
      RECT 19160.4 3826.07 19366.9 3826.63 ;
      RECT 19160.4 3859.31 19366.9 3859.87 ;
      RECT 19160.4 3898.07 19366.9 3898.63 ;
      RECT 19160.4 3931.31 19366.9 3931.87 ;
      RECT 19160.4 3970.07 19366.9 3970.63 ;
      RECT 19160.4 4003.31 19366.9 4003.87 ;
      RECT 19160.4 4042.07 19366.9 4042.63 ;
      RECT 19160.4 4075.31 19366.9 4075.87 ;
      RECT 19160.4 4114.07 19366.9 4114.63 ;
      RECT 19160.4 4147.31 19366.9 4147.87 ;
      RECT 19160.4 4186.07 19366.9 4186.63 ;
      RECT 19160.4 4219.31 19366.9 4219.87 ;
      RECT 19160.4 4258.07 19366.9 4258.63 ;
      RECT 19160.4 4291.31 19366.9 4291.87 ;
      RECT 19160.4 4330.07 19366.9 4330.63 ;
      RECT 19160.4 4363.31 19366.9 4363.87 ;
      RECT 19160.4 4402.07 19366.9 4402.63 ;
      RECT 19160.4 4435.31 19366.9 4435.87 ;
      RECT 19160.4 4474.07 19366.9 4474.63 ;
      RECT 19160.4 4507.31 19366.9 4507.87 ;
      RECT 19160.4 4546.07 19366.9 4546.63 ;
      RECT 19160.4 4579.31 19366.9 4579.87 ;
      RECT 19160.4 4618.07 19366.9 4618.63 ;
      RECT 19160.4 4651.31 19366.9 4651.87 ;
      RECT 19160.4 4690.07 19366.9 4690.63 ;
      RECT 19160.4 4723.31 19366.9 4723.87 ;
      RECT 19160.4 4762.07 19366.9 4762.63 ;
      RECT 19160.4 4795.31 19366.9 4795.87 ;
      RECT 19160.4 4834.07 19366.9 4834.63 ;
      RECT 19160.4 4867.31 19366.9 4867.87 ;
      RECT 19160.4 4906.07 19366.9 4906.63 ;
      RECT 19160.4 4939.31 19366.9 4939.87 ;
      RECT 19160.4 4978.07 19366.9 4978.63 ;
      RECT 19160.4 5011.31 19366.9 5011.87 ;
      RECT 19160.4 5050.07 19366.9 5050.63 ;
      RECT 19160.4 5083.31 19366.9 5083.87 ;
      RECT 19160.4 5122.07 19366.9 5122.63 ;
      RECT 19160.4 5155.31 19366.9 5155.87 ;
      RECT 19160.4 5194.07 19366.9 5194.63 ;
      RECT 19160.4 5227.31 19366.9 5227.87 ;
      RECT 19160.4 5266.07 19366.9 5266.63 ;
      RECT 19160.4 5299.31 19366.9 5299.87 ;
      RECT 19160.4 5338.07 19366.9 5338.63 ;
      RECT 19160.4 5371.31 19366.9 5371.87 ;
      RECT 19160.4 5410.07 19366.9 5410.63 ;
      RECT 19160.4 5443.31 19366.9 5443.87 ;
      RECT 19160.4 5482.07 19366.9 5482.63 ;
      RECT 19160.4 5515.31 19366.9 5515.87 ;
      RECT 19160.4 5554.07 19366.9 5554.63 ;
      RECT 19160.4 5587.31 19366.9 5587.87 ;
      RECT 19160.4 5626.07 19366.9 5626.63 ;
      RECT 19160.4 5659.31 19366.9 5659.87 ;
      RECT 19160.4 5698.07 19366.9 5698.63 ;
      RECT 19160.4 5731.31 19366.9 5731.87 ;
      RECT 19160.4 5770.07 19366.9 5770.63 ;
      RECT 19160.4 5803.31 19366.9 5803.87 ;
      RECT 19160.4 5842.07 19366.9 5842.63 ;
      RECT 19160.4 5875.31 19366.9 5875.87 ;
      RECT 19160.4 5914.07 19366.9 5914.63 ;
      RECT 19160.4 5947.31 19366.9 5947.87 ;
      RECT 19160.4 5986.07 19366.9 5986.63 ;
      RECT 19160.4 6019.31 19366.9 6019.87 ;
      RECT 19160.4 6058.07 19366.9 6058.63 ;
      RECT 19160.4 6091.31 19366.9 6091.87 ;
      RECT 19160.4 6130.07 19366.9 6130.63 ;
      RECT 19160.4 6163.31 19366.9 6163.87 ;
      RECT 19160.4 6202.07 19366.9 6202.63 ;
      RECT 19160.4 6235.31 19366.9 6235.87 ;
      RECT 19160.4 6274.07 19366.9 6274.63 ;
      RECT 19160.4 6307.31 19366.9 6307.87 ;
      RECT 19160.4 6346.07 19366.9 6346.63 ;
      RECT 19160.4 6379.31 19366.9 6379.87 ;
      RECT 19160.4 6418.07 19366.9 6418.63 ;
      RECT 19160.4 6451.31 19366.9 6451.87 ;
      RECT 19160.4 6490.07 19366.9 6490.63 ;
      RECT 19160.4 6523.31 19366.9 6523.87 ;
      RECT 19160.4 6562.07 19366.9 6562.63 ;
      RECT 19160.4 6595.31 19366.9 6595.87 ;
      RECT 19160.4 6634.07 19366.9 6634.63 ;
      RECT 19160.4 6667.31 19366.9 6667.87 ;
      RECT 19160.4 6706.07 19366.9 6706.63 ;
      RECT 19160.4 6739.31 19366.9 6739.87 ;
      RECT 19160.4 6778.07 19366.9 6778.63 ;
      RECT 19160.4 6811.31 19366.9 6811.87 ;
      RECT 19160.4 6850.07 19366.9 6850.63 ;
      RECT 19160.4 6883.31 19366.9 6883.87 ;
      RECT 19160.4 6922.07 19366.9 6922.63 ;
      RECT 19160.4 6955.31 19366.9 6955.87 ;
      RECT 19160.4 6994.07 19366.9 6994.63 ;
      RECT 19160.4 7027.31 19366.9 7027.87 ;
      RECT 19160.4 7066.07 19366.9 7066.63 ;
      RECT 19160.4 7099.31 19366.9 7099.87 ;
      RECT 19160.4 7138.07 19366.9 7138.63 ;
      RECT 19160.4 7171.31 19366.9 7171.87 ;
      RECT 19160.4 7210.07 19366.9 7210.63 ;
      RECT 19160.4 7243.31 19366.9 7243.87 ;
      RECT 19160.4 7282.07 19366.9 7282.63 ;
      RECT 19160.4 7315.31 19366.9 7315.87 ;
      RECT 19160.4 7354.07 19366.9 7354.63 ;
      RECT 19160.4 7387.31 19366.9 7387.87 ;
      RECT 19160.4 7426.07 19366.9 7426.63 ;
      RECT 19160.4 7459.31 19366.9 7459.87 ;
      RECT 19160.4 7498.07 19366.9 7498.63 ;
      RECT 19160.4 7531.31 19366.9 7531.87 ;
      RECT 19160.4 7570.07 19366.9 7570.63 ;
      RECT 19160.4 7603.31 19366.9 7603.87 ;
      RECT 19160.4 7642.07 19366.9 7642.63 ;
      RECT 19160.4 7675.31 19366.9 7675.87 ;
      RECT 19160.4 7714.07 19366.9 7714.63 ;
      RECT 19160.4 7747.31 19366.9 7747.87 ;
      RECT 19160.4 7786.07 19366.9 7786.63 ;
      RECT 19160.4 7819.31 19366.9 7819.87 ;
      RECT 19160.4 7858.07 19366.9 7858.63 ;
      RECT 19160.4 7891.31 19366.9 7891.87 ;
      RECT 19160.4 7930.07 19366.9 7930.63 ;
      RECT 19160.4 7963.31 19366.9 7963.87 ;
      RECT 19160.4 8002.07 19366.9 8002.63 ;
      RECT 19160.4 8035.31 19366.9 8035.87 ;
      RECT 19160.4 8074.07 19366.9 8074.63 ;
      RECT 19160.4 8107.31 19366.9 8107.87 ;
      RECT 19160.4 8146.07 19366.9 8146.63 ;
      RECT 19160.4 8179.31 19366.9 8179.87 ;
      RECT 19160.4 8218.07 19366.9 8218.63 ;
      RECT 19160.4 8251.31 19366.9 8251.87 ;
      RECT 19160.4 8290.07 19366.9 8290.63 ;
      RECT 19160.4 8323.31 19366.9 8323.87 ;
      RECT 19160.4 8362.07 19366.9 8362.63 ;
      RECT 19160.4 8395.31 19366.9 8395.87 ;
      RECT 19160.4 8434.07 19366.9 8434.63 ;
      RECT 19160.4 8467.31 19366.9 8467.87 ;
      RECT 19160.4 8506.07 19366.9 8506.63 ;
      RECT 19160.4 8539.31 19366.9 8539.87 ;
      RECT 19160.4 8578.07 19366.9 8578.63 ;
      RECT 19160.4 8611.31 19366.9 8611.87 ;
      RECT 19160.4 8650.07 19366.9 8650.63 ;
      RECT 19160.4 8683.31 19366.9 8683.87 ;
      RECT 19160.4 8722.07 19366.9 8722.63 ;
      RECT 19160.4 8755.31 19366.9 8755.87 ;
      RECT 19160.4 8794.07 19366.9 8794.63 ;
      RECT 19160.4 8827.31 19366.9 8827.87 ;
      RECT 19160.4 8866.07 19366.9 8866.63 ;
      RECT 19160.4 8899.31 19366.9 8899.87 ;
      RECT 19160.4 8938.07 19366.9 8938.63 ;
      RECT 19160.4 8971.31 19366.9 8971.87 ;
      RECT 19160.4 9010.07 19366.9 9010.63 ;
      RECT 19160.4 9043.31 19366.9 9043.87 ;
      RECT 19160.4 9082.07 19366.9 9082.63 ;
      RECT 19160.4 9115.31 19366.9 9115.87 ;
      RECT 19160.4 9154.07 19366.9 9154.63 ;
      RECT 19160.4 9187.31 19366.9 9187.87 ;
      RECT 19160.4 9226.07 19366.9 9226.63 ;
      RECT 19160.4 9259.31 19366.9 9259.87 ;
      RECT 19160.4 9298.07 19366.9 9298.63 ;
      RECT 19160.4 9331.31 19366.9 9331.87 ;
      RECT 19160.4 9370.07 19366.9 9370.63 ;
      RECT 19160.4 9403.31 19366.9 9403.87 ;
      RECT 19160.4 9442.07 19366.9 9442.63 ;
      RECT 19160.9 1055.24 19326.9 1069.27 ;
      RECT 19160.9 1120.24 19326.9 1148.27 ;
      RECT 19160.9 1168.24 19326.9 1182.27 ;
      RECT 19160.9 1394.97 19326.9 1399.58 ;
      RECT 19160.9 1462.36 19326.9 1471.58 ;
      RECT 19160.9 1534.36 19326.9 1543.58 ;
      RECT 19160.9 1606.36 19326.9 1615.58 ;
      RECT 19160.9 1678.36 19326.9 1687.58 ;
      RECT 19160.9 1750.36 19326.9 1759.58 ;
      RECT 19160.9 1822.36 19326.9 1831.58 ;
      RECT 19160.9 1894.36 19326.9 1903.58 ;
      RECT 19160.9 1966.36 19326.9 1975.58 ;
      RECT 19160.9 2038.36 19326.9 2047.58 ;
      RECT 19160.9 2110.36 19326.9 2119.58 ;
      RECT 19160.9 2182.36 19326.9 2191.58 ;
      RECT 19160.9 2254.36 19326.9 2263.58 ;
      RECT 19160.9 2326.36 19326.9 2335.58 ;
      RECT 19160.9 2398.36 19326.9 2407.58 ;
      RECT 19160.9 2470.36 19326.9 2479.58 ;
      RECT 19160.9 2542.36 19326.9 2551.58 ;
      RECT 19160.9 2614.36 19326.9 2623.58 ;
      RECT 19160.9 2686.36 19326.9 2695.58 ;
      RECT 19160.9 2758.36 19326.9 2767.58 ;
      RECT 19160.9 2830.36 19326.9 2839.58 ;
      RECT 19160.9 2902.36 19326.9 2911.58 ;
      RECT 19160.9 2974.36 19326.9 2983.58 ;
      RECT 19160.9 3046.36 19326.9 3055.58 ;
      RECT 19160.9 3118.36 19326.9 3127.58 ;
      RECT 19160.9 3190.36 19326.9 3199.58 ;
      RECT 19160.9 3262.36 19326.9 3271.58 ;
      RECT 19160.9 3334.36 19326.9 3343.58 ;
      RECT 19160.9 3406.36 19326.9 3415.58 ;
      RECT 19160.9 3478.36 19326.9 3487.58 ;
      RECT 19160.9 3550.36 19326.9 3559.58 ;
      RECT 19160.9 3622.36 19326.9 3631.58 ;
      RECT 19160.9 3694.36 19326.9 3703.58 ;
      RECT 19160.9 3766.36 19326.9 3775.58 ;
      RECT 19160.9 3838.36 19326.9 3847.58 ;
      RECT 19160.9 3910.36 19326.9 3919.58 ;
      RECT 19160.9 3982.36 19326.9 3991.58 ;
      RECT 19160.9 4054.36 19326.9 4063.58 ;
      RECT 19160.9 4126.36 19326.9 4135.58 ;
      RECT 19160.9 4198.36 19326.9 4207.58 ;
      RECT 19160.9 4270.36 19326.9 4279.58 ;
      RECT 19160.9 4342.36 19326.9 4351.58 ;
      RECT 19160.9 4414.36 19326.9 4423.58 ;
      RECT 19160.9 4486.36 19326.9 4495.58 ;
      RECT 19160.9 4558.36 19326.9 4567.58 ;
      RECT 19160.9 4630.36 19326.9 4639.58 ;
      RECT 19160.9 4702.36 19326.9 4711.58 ;
      RECT 19160.9 4774.36 19326.9 4783.58 ;
      RECT 19160.9 4846.36 19326.9 4855.58 ;
      RECT 19160.9 4918.36 19326.9 4927.58 ;
      RECT 19160.9 4990.36 19326.9 4999.58 ;
      RECT 19160.9 5062.36 19326.9 5071.58 ;
      RECT 19160.9 5134.36 19326.9 5143.58 ;
      RECT 19160.9 5206.36 19326.9 5215.58 ;
      RECT 19160.9 5278.36 19326.9 5287.58 ;
      RECT 19160.9 5350.36 19326.9 5359.58 ;
      RECT 19160.9 5422.36 19326.9 5431.58 ;
      RECT 19160.9 5494.36 19326.9 5503.58 ;
      RECT 19160.9 5566.36 19326.9 5575.58 ;
      RECT 19160.9 5638.36 19326.9 5647.58 ;
      RECT 19160.9 5710.36 19326.9 5719.58 ;
      RECT 19160.9 5782.36 19326.9 5791.58 ;
      RECT 19160.9 5854.36 19326.9 5863.58 ;
      RECT 19160.9 5926.36 19326.9 5935.58 ;
      RECT 19160.9 5998.36 19326.9 6007.58 ;
      RECT 19160.9 6070.36 19326.9 6079.58 ;
      RECT 19160.9 6142.36 19326.9 6151.58 ;
      RECT 19160.9 6214.36 19326.9 6223.58 ;
      RECT 19160.9 6286.36 19326.9 6295.58 ;
      RECT 19160.9 6358.36 19326.9 6367.58 ;
      RECT 19160.9 6430.36 19326.9 6439.58 ;
      RECT 19160.9 6502.36 19326.9 6511.58 ;
      RECT 19160.9 6574.36 19326.9 6583.58 ;
      RECT 19160.9 6646.36 19326.9 6655.58 ;
      RECT 19160.9 6718.36 19326.9 6727.58 ;
      RECT 19160.9 6790.36 19326.9 6799.58 ;
      RECT 19160.9 6862.36 19326.9 6871.58 ;
      RECT 19160.9 6934.36 19326.9 6943.58 ;
      RECT 19160.9 7006.36 19326.9 7015.58 ;
      RECT 19160.9 7078.36 19326.9 7087.58 ;
      RECT 19160.9 7150.36 19326.9 7159.58 ;
      RECT 19160.9 7222.36 19326.9 7231.58 ;
      RECT 19160.9 7294.36 19326.9 7303.58 ;
      RECT 19160.9 7366.36 19326.9 7375.58 ;
      RECT 19160.9 7438.36 19326.9 7447.58 ;
      RECT 19160.9 7510.36 19326.9 7519.58 ;
      RECT 19160.9 7582.36 19326.9 7591.58 ;
      RECT 19160.9 7654.36 19326.9 7663.58 ;
      RECT 19160.9 7726.36 19326.9 7735.58 ;
      RECT 19160.9 7798.36 19326.9 7807.58 ;
      RECT 19160.9 7870.36 19326.9 7879.58 ;
      RECT 19160.9 7942.36 19326.9 7951.58 ;
      RECT 19160.9 8014.36 19326.9 8023.58 ;
      RECT 19160.9 8086.36 19326.9 8095.58 ;
      RECT 19160.9 8158.36 19326.9 8167.58 ;
      RECT 19160.9 8230.36 19326.9 8239.58 ;
      RECT 19160.9 8302.36 19326.9 8311.58 ;
      RECT 19160.9 8374.36 19326.9 8383.58 ;
      RECT 19160.9 8446.36 19326.9 8455.58 ;
      RECT 19160.9 8518.36 19326.9 8527.58 ;
      RECT 19160.9 8590.36 19326.9 8599.58 ;
      RECT 19160.9 8662.36 19326.9 8671.58 ;
      RECT 19160.9 8734.36 19326.9 8743.58 ;
      RECT 19160.9 8806.36 19326.9 8815.58 ;
      RECT 19160.9 8878.36 19326.9 8887.58 ;
      RECT 19160.9 8950.36 19326.9 8959.58 ;
      RECT 19160.9 9022.36 19326.9 9031.58 ;
      RECT 19160.9 9094.36 19326.9 9103.58 ;
      RECT 19160.9 9166.36 19326.9 9175.58 ;
      RECT 19160.9 9238.36 19326.9 9247.58 ;
      RECT 19160.9 9310.36 19326.9 9319.58 ;
      RECT 19160.9 9382.36 19326.9 9391.58 ;
      RECT 19160.9 9454.36 19326.9 9458.97 ;
      RECT 19160.9 1401.58 19286.9 1406.19 ;
      RECT 19160.9 1455.75 19286.9 1460.36 ;
      RECT 19160.9 1473.58 19286.9 1478.19 ;
      RECT 19160.9 1527.75 19286.9 1532.36 ;
      RECT 19160.9 1545.58 19286.9 1550.19 ;
      RECT 19160.9 1599.75 19286.9 1604.36 ;
      RECT 19160.9 1617.58 19286.9 1622.19 ;
      RECT 19160.9 1671.75 19286.9 1676.36 ;
      RECT 19160.9 1689.58 19286.9 1694.19 ;
      RECT 19160.9 1743.75 19286.9 1748.36 ;
      RECT 19160.9 1761.58 19286.9 1766.19 ;
      RECT 19160.9 1815.75 19286.9 1820.36 ;
      RECT 19160.9 1833.58 19286.9 1838.19 ;
      RECT 19160.9 1887.75 19286.9 1892.36 ;
      RECT 19160.9 1905.58 19286.9 1910.19 ;
      RECT 19160.9 1959.75 19286.9 1964.36 ;
      RECT 19160.9 1977.58 19286.9 1982.19 ;
      RECT 19160.9 2031.75 19286.9 2036.36 ;
      RECT 19160.9 2049.58 19286.9 2054.19 ;
      RECT 19160.9 2103.75 19286.9 2108.36 ;
      RECT 19160.9 2121.58 19286.9 2126.19 ;
      RECT 19160.9 2175.75 19286.9 2180.36 ;
      RECT 19160.9 2193.58 19286.9 2198.19 ;
      RECT 19160.9 2247.75 19286.9 2252.36 ;
      RECT 19160.9 2265.58 19286.9 2270.19 ;
      RECT 19160.9 2319.75 19286.9 2324.36 ;
      RECT 19160.9 2337.58 19286.9 2342.19 ;
      RECT 19160.9 2391.75 19286.9 2396.36 ;
      RECT 19160.9 2409.58 19286.9 2414.19 ;
      RECT 19160.9 2463.75 19286.9 2468.36 ;
      RECT 19160.9 2481.58 19286.9 2486.19 ;
      RECT 19160.9 2535.75 19286.9 2540.36 ;
      RECT 19160.9 2553.58 19286.9 2558.19 ;
      RECT 19160.9 2607.75 19286.9 2612.36 ;
      RECT 19160.9 2625.58 19286.9 2630.19 ;
      RECT 19160.9 2679.75 19286.9 2684.36 ;
      RECT 19160.9 2697.58 19286.9 2702.19 ;
      RECT 19160.9 2751.75 19286.9 2756.36 ;
      RECT 19160.9 2769.58 19286.9 2774.19 ;
      RECT 19160.9 2823.75 19286.9 2828.36 ;
      RECT 19160.9 2841.58 19286.9 2846.19 ;
      RECT 19160.9 2895.75 19286.9 2900.36 ;
      RECT 19160.9 2913.58 19286.9 2918.19 ;
      RECT 19160.9 2967.75 19286.9 2972.36 ;
      RECT 19160.9 2985.58 19286.9 2990.19 ;
      RECT 19160.9 3039.75 19286.9 3044.36 ;
      RECT 19160.9 3057.58 19286.9 3062.19 ;
      RECT 19160.9 3111.75 19286.9 3116.36 ;
      RECT 19160.9 3129.58 19286.9 3134.19 ;
      RECT 19160.9 3183.75 19286.9 3188.36 ;
      RECT 19160.9 3201.58 19286.9 3206.19 ;
      RECT 19160.9 3255.75 19286.9 3260.36 ;
      RECT 19160.9 3273.58 19286.9 3278.19 ;
      RECT 19160.9 3327.75 19286.9 3332.36 ;
      RECT 19160.9 3345.58 19286.9 3350.19 ;
      RECT 19160.9 3399.75 19286.9 3404.36 ;
      RECT 19160.9 3417.58 19286.9 3422.19 ;
      RECT 19160.9 3471.75 19286.9 3476.36 ;
      RECT 19160.9 3489.58 19286.9 3494.19 ;
      RECT 19160.9 3543.75 19286.9 3548.36 ;
      RECT 19160.9 3561.58 19286.9 3566.19 ;
      RECT 19160.9 3615.75 19286.9 3620.36 ;
      RECT 19160.9 3633.58 19286.9 3638.19 ;
      RECT 19160.9 3687.75 19286.9 3692.36 ;
      RECT 19160.9 3705.58 19286.9 3710.19 ;
      RECT 19160.9 3759.75 19286.9 3764.36 ;
      RECT 19160.9 3777.58 19286.9 3782.19 ;
      RECT 19160.9 3831.75 19286.9 3836.36 ;
      RECT 19160.9 3849.58 19286.9 3854.19 ;
      RECT 19160.9 3903.75 19286.9 3908.36 ;
      RECT 19160.9 3921.58 19286.9 3926.19 ;
      RECT 19160.9 3975.75 19286.9 3980.36 ;
      RECT 19160.9 3993.58 19286.9 3998.19 ;
      RECT 19160.9 4047.75 19286.9 4052.36 ;
      RECT 19160.9 4065.58 19286.9 4070.19 ;
      RECT 19160.9 4119.75 19286.9 4124.36 ;
      RECT 19160.9 4137.58 19286.9 4142.19 ;
      RECT 19160.9 4191.75 19286.9 4196.36 ;
      RECT 19160.9 4209.58 19286.9 4214.19 ;
      RECT 19160.9 4263.75 19286.9 4268.36 ;
      RECT 19160.9 4281.58 19286.9 4286.19 ;
      RECT 19160.9 4335.75 19286.9 4340.36 ;
      RECT 19160.9 4353.58 19286.9 4358.19 ;
      RECT 19160.9 4407.75 19286.9 4412.36 ;
      RECT 19160.9 4425.58 19286.9 4430.19 ;
      RECT 19160.9 4479.75 19286.9 4484.36 ;
      RECT 19160.9 4497.58 19286.9 4502.19 ;
      RECT 19160.9 4551.75 19286.9 4556.36 ;
      RECT 19160.9 4569.58 19286.9 4574.19 ;
      RECT 19160.9 4623.75 19286.9 4628.36 ;
      RECT 19160.9 4641.58 19286.9 4646.19 ;
      RECT 19160.9 4695.75 19286.9 4700.36 ;
      RECT 19160.9 4713.58 19286.9 4718.19 ;
      RECT 19160.9 4767.75 19286.9 4772.36 ;
      RECT 19160.9 4785.58 19286.9 4790.19 ;
      RECT 19160.9 4839.75 19286.9 4844.36 ;
      RECT 19160.9 4857.58 19286.9 4862.19 ;
      RECT 19160.9 4911.75 19286.9 4916.36 ;
      RECT 19160.9 4929.58 19286.9 4934.19 ;
      RECT 19160.9 4983.75 19286.9 4988.36 ;
      RECT 19160.9 5001.58 19286.9 5006.19 ;
      RECT 19160.9 5055.75 19286.9 5060.36 ;
      RECT 19160.9 5073.58 19286.9 5078.19 ;
      RECT 19160.9 5127.75 19286.9 5132.36 ;
      RECT 19160.9 5145.58 19286.9 5150.19 ;
      RECT 19160.9 5199.75 19286.9 5204.36 ;
      RECT 19160.9 5217.58 19286.9 5222.19 ;
      RECT 19160.9 5271.75 19286.9 5276.36 ;
      RECT 19160.9 5289.58 19286.9 5294.19 ;
      RECT 19160.9 5343.75 19286.9 5348.36 ;
      RECT 19160.9 5361.58 19286.9 5366.19 ;
      RECT 19160.9 5415.75 19286.9 5420.36 ;
      RECT 19160.9 5433.58 19286.9 5438.19 ;
      RECT 19160.9 5487.75 19286.9 5492.36 ;
      RECT 19160.9 5505.58 19286.9 5510.19 ;
      RECT 19160.9 5559.75 19286.9 5564.36 ;
      RECT 19160.9 5577.58 19286.9 5582.19 ;
      RECT 19160.9 5631.75 19286.9 5636.36 ;
      RECT 19160.9 5649.58 19286.9 5654.19 ;
      RECT 19160.9 5703.75 19286.9 5708.36 ;
      RECT 19160.9 5721.58 19286.9 5726.19 ;
      RECT 19160.9 5775.75 19286.9 5780.36 ;
      RECT 19160.9 5793.58 19286.9 5798.19 ;
      RECT 19160.9 5847.75 19286.9 5852.36 ;
      RECT 19160.9 5865.58 19286.9 5870.19 ;
      RECT 19160.9 5919.75 19286.9 5924.36 ;
      RECT 19160.9 5937.58 19286.9 5942.19 ;
      RECT 19160.9 5991.75 19286.9 5996.36 ;
      RECT 19160.9 6009.58 19286.9 6014.19 ;
      RECT 19160.9 6063.75 19286.9 6068.36 ;
      RECT 19160.9 6081.58 19286.9 6086.19 ;
      RECT 19160.9 6135.75 19286.9 6140.36 ;
      RECT 19160.9 6153.58 19286.9 6158.19 ;
      RECT 19160.9 6207.75 19286.9 6212.36 ;
      RECT 19160.9 6225.58 19286.9 6230.19 ;
      RECT 19160.9 6279.75 19286.9 6284.36 ;
      RECT 19160.9 6297.58 19286.9 6302.19 ;
      RECT 19160.9 6351.75 19286.9 6356.36 ;
      RECT 19160.9 6369.58 19286.9 6374.19 ;
      RECT 19160.9 6423.75 19286.9 6428.36 ;
      RECT 19160.9 6441.58 19286.9 6446.19 ;
      RECT 19160.9 6495.75 19286.9 6500.36 ;
      RECT 19160.9 6513.58 19286.9 6518.19 ;
      RECT 19160.9 6567.75 19286.9 6572.36 ;
      RECT 19160.9 6585.58 19286.9 6590.19 ;
      RECT 19160.9 6639.75 19286.9 6644.36 ;
      RECT 19160.9 6657.58 19286.9 6662.19 ;
      RECT 19160.9 6711.75 19286.9 6716.36 ;
      RECT 19160.9 6729.58 19286.9 6734.19 ;
      RECT 19160.9 6783.75 19286.9 6788.36 ;
      RECT 19160.9 6801.58 19286.9 6806.19 ;
      RECT 19160.9 6855.75 19286.9 6860.36 ;
      RECT 19160.9 6873.58 19286.9 6878.19 ;
      RECT 19160.9 6927.75 19286.9 6932.36 ;
      RECT 19160.9 6945.58 19286.9 6950.19 ;
      RECT 19160.9 6999.75 19286.9 7004.36 ;
      RECT 19160.9 7017.58 19286.9 7022.19 ;
      RECT 19160.9 7071.75 19286.9 7076.36 ;
      RECT 19160.9 7089.58 19286.9 7094.19 ;
      RECT 19160.9 7143.75 19286.9 7148.36 ;
      RECT 19160.9 7161.58 19286.9 7166.19 ;
      RECT 19160.9 7215.75 19286.9 7220.36 ;
      RECT 19160.9 7233.58 19286.9 7238.19 ;
      RECT 19160.9 7287.75 19286.9 7292.36 ;
      RECT 19160.9 7305.58 19286.9 7310.19 ;
      RECT 19160.9 7359.75 19286.9 7364.36 ;
      RECT 19160.9 7377.58 19286.9 7382.19 ;
      RECT 19160.9 7431.75 19286.9 7436.36 ;
      RECT 19160.9 7449.58 19286.9 7454.19 ;
      RECT 19160.9 7503.75 19286.9 7508.36 ;
      RECT 19160.9 7521.58 19286.9 7526.19 ;
      RECT 19160.9 7575.75 19286.9 7580.36 ;
      RECT 19160.9 7593.58 19286.9 7598.19 ;
      RECT 19160.9 7647.75 19286.9 7652.36 ;
      RECT 19160.9 7665.58 19286.9 7670.19 ;
      RECT 19160.9 7719.75 19286.9 7724.36 ;
      RECT 19160.9 7737.58 19286.9 7742.19 ;
      RECT 19160.9 7791.75 19286.9 7796.36 ;
      RECT 19160.9 7809.58 19286.9 7814.19 ;
      RECT 19160.9 7863.75 19286.9 7868.36 ;
      RECT 19160.9 7881.58 19286.9 7886.19 ;
      RECT 19160.9 7935.75 19286.9 7940.36 ;
      RECT 19160.9 7953.58 19286.9 7958.19 ;
      RECT 19160.9 8007.75 19286.9 8012.36 ;
      RECT 19160.9 8025.58 19286.9 8030.19 ;
      RECT 19160.9 8079.75 19286.9 8084.36 ;
      RECT 19160.9 8097.58 19286.9 8102.19 ;
      RECT 19160.9 8151.75 19286.9 8156.36 ;
      RECT 19160.9 8169.58 19286.9 8174.19 ;
      RECT 19160.9 8223.75 19286.9 8228.36 ;
      RECT 19160.9 8241.58 19286.9 8246.19 ;
      RECT 19160.9 8295.75 19286.9 8300.36 ;
      RECT 19160.9 8313.58 19286.9 8318.19 ;
      RECT 19160.9 8367.75 19286.9 8372.36 ;
      RECT 19160.9 8385.58 19286.9 8390.19 ;
      RECT 19160.9 8439.75 19286.9 8444.36 ;
      RECT 19160.9 8457.58 19286.9 8462.19 ;
      RECT 19160.9 8511.75 19286.9 8516.36 ;
      RECT 19160.9 8529.58 19286.9 8534.19 ;
      RECT 19160.9 8583.75 19286.9 8588.36 ;
      RECT 19160.9 8601.58 19286.9 8606.19 ;
      RECT 19160.9 8655.75 19286.9 8660.36 ;
      RECT 19160.9 8673.58 19286.9 8678.19 ;
      RECT 19160.9 8727.75 19286.9 8732.36 ;
      RECT 19160.9 8745.58 19286.9 8750.19 ;
      RECT 19160.9 8799.75 19286.9 8804.36 ;
      RECT 19160.9 8817.58 19286.9 8822.19 ;
      RECT 19160.9 8871.75 19286.9 8876.36 ;
      RECT 19160.9 8889.58 19286.9 8894.19 ;
      RECT 19160.9 8943.75 19286.9 8948.36 ;
      RECT 19160.9 8961.58 19286.9 8966.19 ;
      RECT 19160.9 9015.75 19286.9 9020.36 ;
      RECT 19160.9 9033.58 19286.9 9038.19 ;
      RECT 19160.9 9087.75 19286.9 9092.36 ;
      RECT 19160.9 9105.58 19286.9 9110.19 ;
      RECT 19160.9 9159.75 19286.9 9164.36 ;
      RECT 19160.9 9177.58 19286.9 9182.19 ;
      RECT 19160.9 9231.75 19286.9 9236.36 ;
      RECT 19160.9 9249.58 19286.9 9254.19 ;
      RECT 19160.9 9303.75 19286.9 9308.36 ;
      RECT 19160.9 9321.58 19286.9 9326.19 ;
      RECT 19160.9 9375.75 19286.9 9380.36 ;
      RECT 19160.9 9393.58 19286.9 9398.19 ;
      RECT 19160.9 9447.75 19286.9 9452.36 ;
      RECT 19160.9 1072.24 19246.9 1086.27 ;
      RECT 19160.9 1089.24 19246.9 1117.27 ;
      RECT 19160.9 1151.24 19246.9 1165.27 ;
      RECT 19040 1198.55 19246.9 1231.55 ;
      RECT 19160.9 1425.2 19246.9 1436.74 ;
      RECT 19160.9 1497.2 19246.9 1508.74 ;
      RECT 19160.9 1569.2 19246.9 1580.74 ;
      RECT 19160.9 1641.2 19246.9 1652.74 ;
      RECT 19160.9 1713.2 19246.9 1724.74 ;
      RECT 19160.9 1785.2 19246.9 1796.74 ;
      RECT 19160.9 1857.2 19246.9 1868.74 ;
      RECT 19160.9 1929.2 19246.9 1940.74 ;
      RECT 19160.9 2001.2 19246.9 2012.74 ;
      RECT 19160.9 2073.2 19246.9 2084.74 ;
      RECT 19160.9 2145.2 19246.9 2156.74 ;
      RECT 19160.9 2217.2 19246.9 2228.74 ;
      RECT 19160.9 2289.2 19246.9 2300.74 ;
      RECT 19160.9 2361.2 19246.9 2372.74 ;
      RECT 19160.9 2433.2 19246.9 2444.74 ;
      RECT 19160.9 2505.2 19246.9 2516.74 ;
      RECT 19160.9 2577.2 19246.9 2588.74 ;
      RECT 19160.9 2649.2 19246.9 2660.74 ;
      RECT 19160.9 2721.2 19246.9 2732.74 ;
      RECT 19160.9 2793.2 19246.9 2804.74 ;
      RECT 19160.9 2865.2 19246.9 2876.74 ;
      RECT 19160.9 2937.2 19246.9 2948.74 ;
      RECT 19160.9 3009.2 19246.9 3020.74 ;
      RECT 19160.9 3081.2 19246.9 3092.74 ;
      RECT 19160.9 3153.2 19246.9 3164.74 ;
      RECT 19160.9 3225.2 19246.9 3236.74 ;
      RECT 19160.9 3297.2 19246.9 3308.74 ;
      RECT 19160.9 3369.2 19246.9 3380.74 ;
      RECT 19160.9 3441.2 19246.9 3452.74 ;
      RECT 19160.9 3513.2 19246.9 3524.74 ;
      RECT 19160.9 3585.2 19246.9 3596.74 ;
      RECT 19160.9 3657.2 19246.9 3668.74 ;
      RECT 19160.9 3729.2 19246.9 3740.74 ;
      RECT 19160.9 3801.2 19246.9 3812.74 ;
      RECT 19160.9 3873.2 19246.9 3884.74 ;
      RECT 19160.9 3945.2 19246.9 3956.74 ;
      RECT 19160.9 4017.2 19246.9 4028.74 ;
      RECT 19160.9 4089.2 19246.9 4100.74 ;
      RECT 19160.9 4161.2 19246.9 4172.74 ;
      RECT 19160.9 4233.2 19246.9 4244.74 ;
      RECT 19160.9 4305.2 19246.9 4316.74 ;
      RECT 19160.9 4377.2 19246.9 4388.74 ;
      RECT 19160.9 4449.2 19246.9 4460.74 ;
      RECT 19160.9 4521.2 19246.9 4532.74 ;
      RECT 19160.9 4593.2 19246.9 4604.74 ;
      RECT 19160.9 4665.2 19246.9 4676.74 ;
      RECT 19160.9 4737.2 19246.9 4748.74 ;
      RECT 19160.9 4809.2 19246.9 4820.74 ;
      RECT 19160.9 4881.2 19246.9 4892.74 ;
      RECT 19160.9 4953.2 19246.9 4964.74 ;
      RECT 19160.9 5025.2 19246.9 5036.74 ;
      RECT 19160.9 5097.2 19246.9 5108.74 ;
      RECT 19160.9 5169.2 19246.9 5180.74 ;
      RECT 19160.9 5241.2 19246.9 5252.74 ;
      RECT 19160.9 5313.2 19246.9 5324.74 ;
      RECT 19160.9 5385.2 19246.9 5396.74 ;
      RECT 19160.9 5457.2 19246.9 5468.74 ;
      RECT 19160.9 5529.2 19246.9 5540.74 ;
      RECT 19160.9 5601.2 19246.9 5612.74 ;
      RECT 19160.9 5673.2 19246.9 5684.74 ;
      RECT 19160.9 5745.2 19246.9 5756.74 ;
      RECT 19160.9 5817.2 19246.9 5828.74 ;
      RECT 19160.9 5889.2 19246.9 5900.74 ;
      RECT 19160.9 5961.2 19246.9 5972.74 ;
      RECT 19160.9 6033.2 19246.9 6044.74 ;
      RECT 19160.9 6105.2 19246.9 6116.74 ;
      RECT 19160.9 6177.2 19246.9 6188.74 ;
      RECT 19160.9 6249.2 19246.9 6260.74 ;
      RECT 19160.9 6321.2 19246.9 6332.74 ;
      RECT 19160.9 6393.2 19246.9 6404.74 ;
      RECT 19160.9 6465.2 19246.9 6476.74 ;
      RECT 19160.9 6537.2 19246.9 6548.74 ;
      RECT 19160.9 6609.2 19246.9 6620.74 ;
      RECT 19160.9 6681.2 19246.9 6692.74 ;
      RECT 19160.9 6753.2 19246.9 6764.74 ;
      RECT 19160.9 6825.2 19246.9 6836.74 ;
      RECT 19160.9 6897.2 19246.9 6908.74 ;
      RECT 19160.9 6969.2 19246.9 6980.74 ;
      RECT 19160.9 7041.2 19246.9 7052.74 ;
      RECT 19160.9 7113.2 19246.9 7124.74 ;
      RECT 19160.9 7185.2 19246.9 7196.74 ;
      RECT 19160.9 7257.2 19246.9 7268.74 ;
      RECT 19160.9 7329.2 19246.9 7340.74 ;
      RECT 19160.9 7401.2 19246.9 7412.74 ;
      RECT 19160.9 7473.2 19246.9 7484.74 ;
      RECT 19160.9 7545.2 19246.9 7556.74 ;
      RECT 19160.9 7617.2 19246.9 7628.74 ;
      RECT 19160.9 7689.2 19246.9 7700.74 ;
      RECT 19160.9 7761.2 19246.9 7772.74 ;
      RECT 19160.9 7833.2 19246.9 7844.74 ;
      RECT 19160.9 7905.2 19246.9 7916.74 ;
      RECT 19160.9 7977.2 19246.9 7988.74 ;
      RECT 19160.9 8049.2 19246.9 8060.74 ;
      RECT 19160.9 8121.2 19246.9 8132.74 ;
      RECT 19160.9 8193.2 19246.9 8204.74 ;
      RECT 19160.9 8265.2 19246.9 8276.74 ;
      RECT 19160.9 8337.2 19246.9 8348.74 ;
      RECT 19160.9 8409.2 19246.9 8420.74 ;
      RECT 19160.9 8481.2 19246.9 8492.74 ;
      RECT 19160.9 8553.2 19246.9 8564.74 ;
      RECT 19160.9 8625.2 19246.9 8636.74 ;
      RECT 19160.9 8697.2 19246.9 8708.74 ;
      RECT 19160.9 8769.2 19246.9 8780.74 ;
      RECT 19160.9 8841.2 19246.9 8852.74 ;
      RECT 19160.9 8913.2 19246.9 8924.74 ;
      RECT 19160.9 8985.2 19246.9 8996.74 ;
      RECT 19160.9 9057.2 19246.9 9068.74 ;
      RECT 19160.9 9129.2 19246.9 9140.74 ;
      RECT 19160.9 9201.2 19246.9 9212.74 ;
      RECT 19160.9 9273.2 19246.9 9284.74 ;
      RECT 19160.9 9345.2 19246.9 9356.74 ;
      RECT 19160.9 9417.2 19246.9 9428.74 ;
      RECT 19160.9 1417.43 19206.9 1423.2 ;
      RECT 19160.9 1438.74 19206.9 1444.51 ;
      RECT 19160.9 1489.43 19206.9 1495.2 ;
      RECT 19160.9 1510.74 19206.9 1516.51 ;
      RECT 19160.9 1561.43 19206.9 1567.2 ;
      RECT 19160.9 1582.74 19206.9 1588.51 ;
      RECT 19160.9 1633.43 19206.9 1639.2 ;
      RECT 19160.9 1654.74 19206.9 1660.51 ;
      RECT 19160.9 1705.43 19206.9 1711.2 ;
      RECT 19160.9 1726.74 19206.9 1732.51 ;
      RECT 19160.9 1777.43 19206.9 1783.2 ;
      RECT 19160.9 1798.74 19206.9 1804.51 ;
      RECT 19160.9 1849.43 19206.9 1855.2 ;
      RECT 19160.9 1870.74 19206.9 1876.51 ;
      RECT 19160.9 1921.43 19206.9 1927.2 ;
      RECT 19160.9 1942.74 19206.9 1948.51 ;
      RECT 19160.9 1993.43 19206.9 1999.2 ;
      RECT 19160.9 2014.74 19206.9 2020.51 ;
      RECT 19160.9 2065.43 19206.9 2071.2 ;
      RECT 19160.9 2086.74 19206.9 2092.51 ;
      RECT 19160.9 2137.43 19206.9 2143.2 ;
      RECT 19160.9 2158.74 19206.9 2164.51 ;
      RECT 19160.9 2209.43 19206.9 2215.2 ;
      RECT 19160.9 2230.74 19206.9 2236.51 ;
      RECT 19160.9 2281.43 19206.9 2287.2 ;
      RECT 19160.9 2302.74 19206.9 2308.51 ;
      RECT 19160.9 2353.43 19206.9 2359.2 ;
      RECT 19160.9 2374.74 19206.9 2380.51 ;
      RECT 19160.9 2425.43 19206.9 2431.2 ;
      RECT 19160.9 2446.74 19206.9 2452.51 ;
      RECT 19160.9 2497.43 19206.9 2503.2 ;
      RECT 19160.9 2518.74 19206.9 2524.51 ;
      RECT 19160.9 2569.43 19206.9 2575.2 ;
      RECT 19160.9 2590.74 19206.9 2596.51 ;
      RECT 19160.9 2641.43 19206.9 2647.2 ;
      RECT 19160.9 2662.74 19206.9 2668.51 ;
      RECT 19160.9 2713.43 19206.9 2719.2 ;
      RECT 19160.9 2734.74 19206.9 2740.51 ;
      RECT 19160.9 2785.43 19206.9 2791.2 ;
      RECT 19160.9 2806.74 19206.9 2812.51 ;
      RECT 19160.9 2857.43 19206.9 2863.2 ;
      RECT 19160.9 2878.74 19206.9 2884.51 ;
      RECT 19160.9 2929.43 19206.9 2935.2 ;
      RECT 19160.9 2950.74 19206.9 2956.51 ;
      RECT 19160.9 3001.43 19206.9 3007.2 ;
      RECT 19160.9 3022.74 19206.9 3028.51 ;
      RECT 19160.9 3073.43 19206.9 3079.2 ;
      RECT 19160.9 3094.74 19206.9 3100.51 ;
      RECT 19160.9 3145.43 19206.9 3151.2 ;
      RECT 19160.9 3166.74 19206.9 3172.51 ;
      RECT 19160.9 3217.43 19206.9 3223.2 ;
      RECT 19160.9 3238.74 19206.9 3244.51 ;
      RECT 19160.9 3289.43 19206.9 3295.2 ;
      RECT 19160.9 3310.74 19206.9 3316.51 ;
      RECT 19160.9 3361.43 19206.9 3367.2 ;
      RECT 19160.9 3382.74 19206.9 3388.51 ;
      RECT 19160.9 3433.43 19206.9 3439.2 ;
      RECT 19160.9 3454.74 19206.9 3460.51 ;
      RECT 19160.9 3505.43 19206.9 3511.2 ;
      RECT 19160.9 3526.74 19206.9 3532.51 ;
      RECT 19160.9 3577.43 19206.9 3583.2 ;
      RECT 19160.9 3598.74 19206.9 3604.51 ;
      RECT 19160.9 3649.43 19206.9 3655.2 ;
      RECT 19160.9 3670.74 19206.9 3676.51 ;
      RECT 19160.9 3721.43 19206.9 3727.2 ;
      RECT 19160.9 3742.74 19206.9 3748.51 ;
      RECT 19160.9 3793.43 19206.9 3799.2 ;
      RECT 19160.9 3814.74 19206.9 3820.51 ;
      RECT 19160.9 3865.43 19206.9 3871.2 ;
      RECT 19160.9 3886.74 19206.9 3892.51 ;
      RECT 19160.9 3937.43 19206.9 3943.2 ;
      RECT 19160.9 3958.74 19206.9 3964.51 ;
      RECT 19160.9 4009.43 19206.9 4015.2 ;
      RECT 19160.9 4030.74 19206.9 4036.51 ;
      RECT 19160.9 4081.43 19206.9 4087.2 ;
      RECT 19160.9 4102.74 19206.9 4108.51 ;
      RECT 19160.9 4153.43 19206.9 4159.2 ;
      RECT 19160.9 4174.74 19206.9 4180.51 ;
      RECT 19160.9 4225.43 19206.9 4231.2 ;
      RECT 19160.9 4246.74 19206.9 4252.51 ;
      RECT 19160.9 4297.43 19206.9 4303.2 ;
      RECT 19160.9 4318.74 19206.9 4324.51 ;
      RECT 19160.9 4369.43 19206.9 4375.2 ;
      RECT 19160.9 4390.74 19206.9 4396.51 ;
      RECT 19160.9 4441.43 19206.9 4447.2 ;
      RECT 19160.9 4462.74 19206.9 4468.51 ;
      RECT 19160.9 4513.43 19206.9 4519.2 ;
      RECT 19160.9 4534.74 19206.9 4540.51 ;
      RECT 19160.9 4585.43 19206.9 4591.2 ;
      RECT 19160.9 4606.74 19206.9 4612.51 ;
      RECT 19160.9 4657.43 19206.9 4663.2 ;
      RECT 19160.9 4678.74 19206.9 4684.51 ;
      RECT 19160.9 4729.43 19206.9 4735.2 ;
      RECT 19160.9 4750.74 19206.9 4756.51 ;
      RECT 19160.9 4801.43 19206.9 4807.2 ;
      RECT 19160.9 4822.74 19206.9 4828.51 ;
      RECT 19160.9 4873.43 19206.9 4879.2 ;
      RECT 19160.9 4894.74 19206.9 4900.51 ;
      RECT 19160.9 4945.43 19206.9 4951.2 ;
      RECT 19160.9 4966.74 19206.9 4972.51 ;
      RECT 19160.9 5017.43 19206.9 5023.2 ;
      RECT 19160.9 5038.74 19206.9 5044.51 ;
      RECT 19160.9 5089.43 19206.9 5095.2 ;
      RECT 19160.9 5110.74 19206.9 5116.51 ;
      RECT 19160.9 5161.43 19206.9 5167.2 ;
      RECT 19160.9 5182.74 19206.9 5188.51 ;
      RECT 19160.9 5233.43 19206.9 5239.2 ;
      RECT 19160.9 5254.74 19206.9 5260.51 ;
      RECT 19160.9 5305.43 19206.9 5311.2 ;
      RECT 19160.9 5326.74 19206.9 5332.51 ;
      RECT 19160.9 5377.43 19206.9 5383.2 ;
      RECT 19160.9 5398.74 19206.9 5404.51 ;
      RECT 19160.9 5449.43 19206.9 5455.2 ;
      RECT 19160.9 5470.74 19206.9 5476.51 ;
      RECT 19160.9 5521.43 19206.9 5527.2 ;
      RECT 19160.9 5542.74 19206.9 5548.51 ;
      RECT 19160.9 5593.43 19206.9 5599.2 ;
      RECT 19160.9 5614.74 19206.9 5620.51 ;
      RECT 19160.9 5665.43 19206.9 5671.2 ;
      RECT 19160.9 5686.74 19206.9 5692.51 ;
      RECT 19160.9 5737.43 19206.9 5743.2 ;
      RECT 19160.9 5758.74 19206.9 5764.51 ;
      RECT 19160.9 5809.43 19206.9 5815.2 ;
      RECT 19160.9 5830.74 19206.9 5836.51 ;
      RECT 19160.9 5881.43 19206.9 5887.2 ;
      RECT 19160.9 5902.74 19206.9 5908.51 ;
      RECT 19160.9 5953.43 19206.9 5959.2 ;
      RECT 19160.9 5974.74 19206.9 5980.51 ;
      RECT 19160.9 6025.43 19206.9 6031.2 ;
      RECT 19160.9 6046.74 19206.9 6052.51 ;
      RECT 19160.9 6097.43 19206.9 6103.2 ;
      RECT 19160.9 6118.74 19206.9 6124.51 ;
      RECT 19160.9 6169.43 19206.9 6175.2 ;
      RECT 19160.9 6190.74 19206.9 6196.51 ;
      RECT 19160.9 6241.43 19206.9 6247.2 ;
      RECT 19160.9 6262.74 19206.9 6268.51 ;
      RECT 19160.9 6313.43 19206.9 6319.2 ;
      RECT 19160.9 6334.74 19206.9 6340.51 ;
      RECT 19160.9 6385.43 19206.9 6391.2 ;
      RECT 19160.9 6406.74 19206.9 6412.51 ;
      RECT 19160.9 6457.43 19206.9 6463.2 ;
      RECT 19160.9 6478.74 19206.9 6484.51 ;
      RECT 19160.9 6529.43 19206.9 6535.2 ;
      RECT 19160.9 6550.74 19206.9 6556.51 ;
      RECT 19160.9 6601.43 19206.9 6607.2 ;
      RECT 19160.9 6622.74 19206.9 6628.51 ;
      RECT 19160.9 6673.43 19206.9 6679.2 ;
      RECT 19160.9 6694.74 19206.9 6700.51 ;
      RECT 19160.9 6745.43 19206.9 6751.2 ;
      RECT 19160.9 6766.74 19206.9 6772.51 ;
      RECT 19160.9 6817.43 19206.9 6823.2 ;
      RECT 19160.9 6838.74 19206.9 6844.51 ;
      RECT 19160.9 6889.43 19206.9 6895.2 ;
      RECT 19160.9 6910.74 19206.9 6916.51 ;
      RECT 19160.9 6961.43 19206.9 6967.2 ;
      RECT 19160.9 6982.74 19206.9 6988.51 ;
      RECT 19160.9 7033.43 19206.9 7039.2 ;
      RECT 19160.9 7054.74 19206.9 7060.51 ;
      RECT 19160.9 7105.43 19206.9 7111.2 ;
      RECT 19160.9 7126.74 19206.9 7132.51 ;
      RECT 19160.9 7177.43 19206.9 7183.2 ;
      RECT 19160.9 7198.74 19206.9 7204.51 ;
      RECT 19160.9 7249.43 19206.9 7255.2 ;
      RECT 19160.9 7270.74 19206.9 7276.51 ;
      RECT 19160.9 7321.43 19206.9 7327.2 ;
      RECT 19160.9 7342.74 19206.9 7348.51 ;
      RECT 19160.9 7393.43 19206.9 7399.2 ;
      RECT 19160.9 7414.74 19206.9 7420.51 ;
      RECT 19160.9 7465.43 19206.9 7471.2 ;
      RECT 19160.9 7486.74 19206.9 7492.51 ;
      RECT 19160.9 7537.43 19206.9 7543.2 ;
      RECT 19160.9 7558.74 19206.9 7564.51 ;
      RECT 19160.9 7609.43 19206.9 7615.2 ;
      RECT 19160.9 7630.74 19206.9 7636.51 ;
      RECT 19160.9 7681.43 19206.9 7687.2 ;
      RECT 19160.9 7702.74 19206.9 7708.51 ;
      RECT 19160.9 7753.43 19206.9 7759.2 ;
      RECT 19160.9 7774.74 19206.9 7780.51 ;
      RECT 19160.9 7825.43 19206.9 7831.2 ;
      RECT 19160.9 7846.74 19206.9 7852.51 ;
      RECT 19160.9 7897.43 19206.9 7903.2 ;
      RECT 19160.9 7918.74 19206.9 7924.51 ;
      RECT 19160.9 7969.43 19206.9 7975.2 ;
      RECT 19160.9 7990.74 19206.9 7996.51 ;
      RECT 19160.9 8041.43 19206.9 8047.2 ;
      RECT 19160.9 8062.74 19206.9 8068.51 ;
      RECT 19160.9 8113.43 19206.9 8119.2 ;
      RECT 19160.9 8134.74 19206.9 8140.51 ;
      RECT 19160.9 8185.43 19206.9 8191.2 ;
      RECT 19160.9 8206.74 19206.9 8212.51 ;
      RECT 19160.9 8257.43 19206.9 8263.2 ;
      RECT 19160.9 8278.74 19206.9 8284.51 ;
      RECT 19160.9 8329.43 19206.9 8335.2 ;
      RECT 19160.9 8350.74 19206.9 8356.51 ;
      RECT 19160.9 8401.43 19206.9 8407.2 ;
      RECT 19160.9 8422.74 19206.9 8428.51 ;
      RECT 19160.9 8473.43 19206.9 8479.2 ;
      RECT 19160.9 8494.74 19206.9 8500.51 ;
      RECT 19160.9 8545.43 19206.9 8551.2 ;
      RECT 19160.9 8566.74 19206.9 8572.51 ;
      RECT 19160.9 8617.43 19206.9 8623.2 ;
      RECT 19160.9 8638.74 19206.9 8644.51 ;
      RECT 19160.9 8689.43 19206.9 8695.2 ;
      RECT 19160.9 8710.74 19206.9 8716.51 ;
      RECT 19160.9 8761.43 19206.9 8767.2 ;
      RECT 19160.9 8782.74 19206.9 8788.51 ;
      RECT 19160.9 8833.43 19206.9 8839.2 ;
      RECT 19160.9 8854.74 19206.9 8860.51 ;
      RECT 19160.9 8905.43 19206.9 8911.2 ;
      RECT 19160.9 8926.74 19206.9 8932.51 ;
      RECT 19160.9 8977.43 19206.9 8983.2 ;
      RECT 19160.9 8998.74 19206.9 9004.51 ;
      RECT 19160.9 9049.43 19206.9 9055.2 ;
      RECT 19160.9 9070.74 19206.9 9076.51 ;
      RECT 19160.9 9121.43 19206.9 9127.2 ;
      RECT 19160.9 9142.74 19206.9 9148.51 ;
      RECT 19160.9 9193.43 19206.9 9199.2 ;
      RECT 19160.9 9214.74 19206.9 9220.51 ;
      RECT 19160.9 9265.43 19206.9 9271.2 ;
      RECT 19160.9 9286.74 19206.9 9292.51 ;
      RECT 19160.9 9337.43 19206.9 9343.2 ;
      RECT 19160.9 9358.74 19206.9 9364.51 ;
      RECT 19160.9 9409.43 19206.9 9415.2 ;
      RECT 19160.9 9430.74 19206.9 9436.51 ;
      RECT 913.1 1198.55 1120 1231.55 ;
      RECT 913.1 1327.55 1120 1355.26 ;
      RECT 753.1 1050.27 999.1 1052.27 ;
      RECT 833.1 1055.24 999.1 1069.27 ;
      RECT 913.1 1072.24 999.1 1086.27 ;
      RECT 913.1 1089.24 999.1 1117.27 ;
      RECT 833.1 1120.24 999.1 1148.27 ;
      RECT 913.1 1151.24 999.1 1165.27 ;
      RECT 833.1 1168.24 999.1 1182.27 ;
      RECT 873.1 1359.26 999.1 1369.26 ;
      RECT 753.1 1371.26 999.1 1373.26 ;
      RECT 833.1 1394.97 999.1 1399.58 ;
      RECT 873.1 1401.58 999.1 1406.19 ;
      RECT 793.1 1408.19 999.1 1409.31 ;
      RECT 953.1 1417.43 999.1 1423.2 ;
      RECT 913.1 1425.2 999.1 1436.74 ;
      RECT 953.1 1438.74 999.1 1444.51 ;
      RECT 793.1 1452.63 999.1 1453.75 ;
      RECT 873.1 1455.75 999.1 1460.36 ;
      RECT 833.1 1462.36 999.1 1471.58 ;
      RECT 873.1 1473.58 999.1 1478.19 ;
      RECT 793.1 1480.19 999.1 1481.31 ;
      RECT 953.1 1489.43 999.1 1495.2 ;
      RECT 913.1 1497.2 999.1 1508.74 ;
      RECT 953.1 1510.74 999.1 1516.51 ;
      RECT 793.1 1524.63 999.1 1525.75 ;
      RECT 873.1 1527.75 999.1 1532.36 ;
      RECT 833.1 1534.36 999.1 1543.58 ;
      RECT 873.1 1545.58 999.1 1550.19 ;
      RECT 793.1 1552.19 999.1 1553.31 ;
      RECT 953.1 1561.43 999.1 1567.2 ;
      RECT 913.1 1569.2 999.1 1580.74 ;
      RECT 953.1 1582.74 999.1 1588.51 ;
      RECT 793.1 1596.63 999.1 1597.75 ;
      RECT 873.1 1599.75 999.1 1604.36 ;
      RECT 833.1 1606.36 999.1 1615.58 ;
      RECT 873.1 1617.58 999.1 1622.19 ;
      RECT 793.1 1624.19 999.1 1625.31 ;
      RECT 953.1 1633.43 999.1 1639.2 ;
      RECT 913.1 1641.2 999.1 1652.74 ;
      RECT 953.1 1654.74 999.1 1660.51 ;
      RECT 793.1 1668.63 999.1 1669.75 ;
      RECT 873.1 1671.75 999.1 1676.36 ;
      RECT 833.1 1678.36 999.1 1687.58 ;
      RECT 873.1 1689.58 999.1 1694.19 ;
      RECT 793.1 1696.19 999.1 1697.31 ;
      RECT 953.1 1705.43 999.1 1711.2 ;
      RECT 913.1 1713.2 999.1 1724.74 ;
      RECT 953.1 1726.74 999.1 1732.51 ;
      RECT 793.1 1740.63 999.1 1741.75 ;
      RECT 873.1 1743.75 999.1 1748.36 ;
      RECT 833.1 1750.36 999.1 1759.58 ;
      RECT 873.1 1761.58 999.1 1766.19 ;
      RECT 793.1 1768.19 999.1 1769.31 ;
      RECT 953.1 1777.43 999.1 1783.2 ;
      RECT 913.1 1785.2 999.1 1796.74 ;
      RECT 953.1 1798.74 999.1 1804.51 ;
      RECT 793.1 1812.63 999.1 1813.75 ;
      RECT 873.1 1815.75 999.1 1820.36 ;
      RECT 833.1 1822.36 999.1 1831.58 ;
      RECT 873.1 1833.58 999.1 1838.19 ;
      RECT 793.1 1840.19 999.1 1841.31 ;
      RECT 953.1 1849.43 999.1 1855.2 ;
      RECT 913.1 1857.2 999.1 1868.74 ;
      RECT 953.1 1870.74 999.1 1876.51 ;
      RECT 793.1 1884.63 999.1 1885.75 ;
      RECT 873.1 1887.75 999.1 1892.36 ;
      RECT 833.1 1894.36 999.1 1903.58 ;
      RECT 873.1 1905.58 999.1 1910.19 ;
      RECT 793.1 1912.19 999.1 1913.31 ;
      RECT 953.1 1921.43 999.1 1927.2 ;
      RECT 913.1 1929.2 999.1 1940.74 ;
      RECT 953.1 1942.74 999.1 1948.51 ;
      RECT 793.1 1956.63 999.1 1957.75 ;
      RECT 873.1 1959.75 999.1 1964.36 ;
      RECT 833.1 1966.36 999.1 1975.58 ;
      RECT 873.1 1977.58 999.1 1982.19 ;
      RECT 793.1 1984.19 999.1 1985.31 ;
      RECT 953.1 1993.43 999.1 1999.2 ;
      RECT 913.1 2001.2 999.1 2012.74 ;
      RECT 953.1 2014.74 999.1 2020.51 ;
      RECT 793.1 2028.63 999.1 2029.75 ;
      RECT 873.1 2031.75 999.1 2036.36 ;
      RECT 833.1 2038.36 999.1 2047.58 ;
      RECT 873.1 2049.58 999.1 2054.19 ;
      RECT 793.1 2056.19 999.1 2057.31 ;
      RECT 953.1 2065.43 999.1 2071.2 ;
      RECT 913.1 2073.2 999.1 2084.74 ;
      RECT 953.1 2086.74 999.1 2092.51 ;
      RECT 793.1 2100.63 999.1 2101.75 ;
      RECT 873.1 2103.75 999.1 2108.36 ;
      RECT 833.1 2110.36 999.1 2119.58 ;
      RECT 873.1 2121.58 999.1 2126.19 ;
      RECT 793.1 2128.19 999.1 2129.31 ;
      RECT 953.1 2137.43 999.1 2143.2 ;
      RECT 913.1 2145.2 999.1 2156.74 ;
      RECT 953.1 2158.74 999.1 2164.51 ;
      RECT 793.1 2172.63 999.1 2173.75 ;
      RECT 873.1 2175.75 999.1 2180.36 ;
      RECT 833.1 2182.36 999.1 2191.58 ;
      RECT 873.1 2193.58 999.1 2198.19 ;
      RECT 793.1 2200.19 999.1 2201.31 ;
      RECT 953.1 2209.43 999.1 2215.2 ;
      RECT 913.1 2217.2 999.1 2228.74 ;
      RECT 953.1 2230.74 999.1 2236.51 ;
      RECT 793.1 2244.63 999.1 2245.75 ;
      RECT 873.1 2247.75 999.1 2252.36 ;
      RECT 833.1 2254.36 999.1 2263.58 ;
      RECT 873.1 2265.58 999.1 2270.19 ;
      RECT 793.1 2272.19 999.1 2273.31 ;
      RECT 953.1 2281.43 999.1 2287.2 ;
      RECT 913.1 2289.2 999.1 2300.74 ;
      RECT 953.1 2302.74 999.1 2308.51 ;
      RECT 793.1 2316.63 999.1 2317.75 ;
      RECT 873.1 2319.75 999.1 2324.36 ;
      RECT 833.1 2326.36 999.1 2335.58 ;
      RECT 873.1 2337.58 999.1 2342.19 ;
      RECT 793.1 2344.19 999.1 2345.31 ;
      RECT 953.1 2353.43 999.1 2359.2 ;
      RECT 913.1 2361.2 999.1 2372.74 ;
      RECT 953.1 2374.74 999.1 2380.51 ;
      RECT 793.1 2388.63 999.1 2389.75 ;
      RECT 873.1 2391.75 999.1 2396.36 ;
      RECT 833.1 2398.36 999.1 2407.58 ;
      RECT 873.1 2409.58 999.1 2414.19 ;
      RECT 793.1 2416.19 999.1 2417.31 ;
      RECT 953.1 2425.43 999.1 2431.2 ;
      RECT 913.1 2433.2 999.1 2444.74 ;
      RECT 953.1 2446.74 999.1 2452.51 ;
      RECT 793.1 2460.63 999.1 2461.75 ;
      RECT 873.1 2463.75 999.1 2468.36 ;
      RECT 833.1 2470.36 999.1 2479.58 ;
      RECT 873.1 2481.58 999.1 2486.19 ;
      RECT 793.1 2488.19 999.1 2489.31 ;
      RECT 953.1 2497.43 999.1 2503.2 ;
      RECT 913.1 2505.2 999.1 2516.74 ;
      RECT 953.1 2518.74 999.1 2524.51 ;
      RECT 793.1 2532.63 999.1 2533.75 ;
      RECT 873.1 2535.75 999.1 2540.36 ;
      RECT 833.1 2542.36 999.1 2551.58 ;
      RECT 873.1 2553.58 999.1 2558.19 ;
      RECT 793.1 2560.19 999.1 2561.31 ;
      RECT 953.1 2569.43 999.1 2575.2 ;
      RECT 913.1 2577.2 999.1 2588.74 ;
      RECT 953.1 2590.74 999.1 2596.51 ;
      RECT 793.1 2604.63 999.1 2605.75 ;
      RECT 873.1 2607.75 999.1 2612.36 ;
      RECT 833.1 2614.36 999.1 2623.58 ;
      RECT 873.1 2625.58 999.1 2630.19 ;
      RECT 793.1 2632.19 999.1 2633.31 ;
      RECT 953.1 2641.43 999.1 2647.2 ;
      RECT 913.1 2649.2 999.1 2660.74 ;
      RECT 953.1 2662.74 999.1 2668.51 ;
      RECT 793.1 2676.63 999.1 2677.75 ;
      RECT 873.1 2679.75 999.1 2684.36 ;
      RECT 833.1 2686.36 999.1 2695.58 ;
      RECT 873.1 2697.58 999.1 2702.19 ;
      RECT 793.1 2704.19 999.1 2705.31 ;
      RECT 953.1 2713.43 999.1 2719.2 ;
      RECT 913.1 2721.2 999.1 2732.74 ;
      RECT 953.1 2734.74 999.1 2740.51 ;
      RECT 793.1 2748.63 999.1 2749.75 ;
      RECT 873.1 2751.75 999.1 2756.36 ;
      RECT 833.1 2758.36 999.1 2767.58 ;
      RECT 873.1 2769.58 999.1 2774.19 ;
      RECT 793.1 2776.19 999.1 2777.31 ;
      RECT 953.1 2785.43 999.1 2791.2 ;
      RECT 913.1 2793.2 999.1 2804.74 ;
      RECT 953.1 2806.74 999.1 2812.51 ;
      RECT 793.1 2820.63 999.1 2821.75 ;
      RECT 873.1 2823.75 999.1 2828.36 ;
      RECT 833.1 2830.36 999.1 2839.58 ;
      RECT 873.1 2841.58 999.1 2846.19 ;
      RECT 793.1 2848.19 999.1 2849.31 ;
      RECT 953.1 2857.43 999.1 2863.2 ;
      RECT 913.1 2865.2 999.1 2876.74 ;
      RECT 953.1 2878.74 999.1 2884.51 ;
      RECT 793.1 2892.63 999.1 2893.75 ;
      RECT 873.1 2895.75 999.1 2900.36 ;
      RECT 833.1 2902.36 999.1 2911.58 ;
      RECT 873.1 2913.58 999.1 2918.19 ;
      RECT 793.1 2920.19 999.1 2921.31 ;
      RECT 953.1 2929.43 999.1 2935.2 ;
      RECT 913.1 2937.2 999.1 2948.74 ;
      RECT 953.1 2950.74 999.1 2956.51 ;
      RECT 793.1 2964.63 999.1 2965.75 ;
      RECT 873.1 2967.75 999.1 2972.36 ;
      RECT 833.1 2974.36 999.1 2983.58 ;
      RECT 873.1 2985.58 999.1 2990.19 ;
      RECT 793.1 2992.19 999.1 2993.31 ;
      RECT 953.1 3001.43 999.1 3007.2 ;
      RECT 913.1 3009.2 999.1 3020.74 ;
      RECT 953.1 3022.74 999.1 3028.51 ;
      RECT 793.1 3036.63 999.1 3037.75 ;
      RECT 873.1 3039.75 999.1 3044.36 ;
      RECT 833.1 3046.36 999.1 3055.58 ;
      RECT 873.1 3057.58 999.1 3062.19 ;
      RECT 793.1 3064.19 999.1 3065.31 ;
      RECT 953.1 3073.43 999.1 3079.2 ;
      RECT 913.1 3081.2 999.1 3092.74 ;
      RECT 953.1 3094.74 999.1 3100.51 ;
      RECT 793.1 3108.63 999.1 3109.75 ;
      RECT 873.1 3111.75 999.1 3116.36 ;
      RECT 833.1 3118.36 999.1 3127.58 ;
      RECT 873.1 3129.58 999.1 3134.19 ;
      RECT 793.1 3136.19 999.1 3137.31 ;
      RECT 953.1 3145.43 999.1 3151.2 ;
      RECT 913.1 3153.2 999.1 3164.74 ;
      RECT 953.1 3166.74 999.1 3172.51 ;
      RECT 793.1 3180.63 999.1 3181.75 ;
      RECT 873.1 3183.75 999.1 3188.36 ;
      RECT 833.1 3190.36 999.1 3199.58 ;
      RECT 873.1 3201.58 999.1 3206.19 ;
      RECT 793.1 3208.19 999.1 3209.31 ;
      RECT 953.1 3217.43 999.1 3223.2 ;
      RECT 913.1 3225.2 999.1 3236.74 ;
      RECT 953.1 3238.74 999.1 3244.51 ;
      RECT 793.1 3252.63 999.1 3253.75 ;
      RECT 873.1 3255.75 999.1 3260.36 ;
      RECT 833.1 3262.36 999.1 3271.58 ;
      RECT 873.1 3273.58 999.1 3278.19 ;
      RECT 793.1 3280.19 999.1 3281.31 ;
      RECT 953.1 3289.43 999.1 3295.2 ;
      RECT 913.1 3297.2 999.1 3308.74 ;
      RECT 953.1 3310.74 999.1 3316.51 ;
      RECT 793.1 3324.63 999.1 3325.75 ;
      RECT 873.1 3327.75 999.1 3332.36 ;
      RECT 833.1 3334.36 999.1 3343.58 ;
      RECT 873.1 3345.58 999.1 3350.19 ;
      RECT 793.1 3352.19 999.1 3353.31 ;
      RECT 953.1 3361.43 999.1 3367.2 ;
      RECT 913.1 3369.2 999.1 3380.74 ;
      RECT 953.1 3382.74 999.1 3388.51 ;
      RECT 793.1 3396.63 999.1 3397.75 ;
      RECT 873.1 3399.75 999.1 3404.36 ;
      RECT 833.1 3406.36 999.1 3415.58 ;
      RECT 873.1 3417.58 999.1 3422.19 ;
      RECT 793.1 3424.19 999.1 3425.31 ;
      RECT 953.1 3433.43 999.1 3439.2 ;
      RECT 913.1 3441.2 999.1 3452.74 ;
      RECT 953.1 3454.74 999.1 3460.51 ;
      RECT 793.1 3468.63 999.1 3469.75 ;
      RECT 873.1 3471.75 999.1 3476.36 ;
      RECT 833.1 3478.36 999.1 3487.58 ;
      RECT 873.1 3489.58 999.1 3494.19 ;
      RECT 793.1 3496.19 999.1 3497.31 ;
      RECT 953.1 3505.43 999.1 3511.2 ;
      RECT 913.1 3513.2 999.1 3524.74 ;
      RECT 953.1 3526.74 999.1 3532.51 ;
      RECT 793.1 3540.63 999.1 3541.75 ;
      RECT 873.1 3543.75 999.1 3548.36 ;
      RECT 833.1 3550.36 999.1 3559.58 ;
      RECT 873.1 3561.58 999.1 3566.19 ;
      RECT 793.1 3568.19 999.1 3569.31 ;
      RECT 953.1 3577.43 999.1 3583.2 ;
      RECT 913.1 3585.2 999.1 3596.74 ;
      RECT 953.1 3598.74 999.1 3604.51 ;
      RECT 793.1 3612.63 999.1 3613.75 ;
      RECT 873.1 3615.75 999.1 3620.36 ;
      RECT 833.1 3622.36 999.1 3631.58 ;
      RECT 873.1 3633.58 999.1 3638.19 ;
      RECT 793.1 3640.19 999.1 3641.31 ;
      RECT 953.1 3649.43 999.1 3655.2 ;
      RECT 913.1 3657.2 999.1 3668.74 ;
      RECT 953.1 3670.74 999.1 3676.51 ;
      RECT 793.1 3684.63 999.1 3685.75 ;
      RECT 873.1 3687.75 999.1 3692.36 ;
      RECT 833.1 3694.36 999.1 3703.58 ;
      RECT 873.1 3705.58 999.1 3710.19 ;
      RECT 793.1 3712.19 999.1 3713.31 ;
      RECT 953.1 3721.43 999.1 3727.2 ;
      RECT 913.1 3729.2 999.1 3740.74 ;
      RECT 953.1 3742.74 999.1 3748.51 ;
      RECT 793.1 3756.63 999.1 3757.75 ;
      RECT 873.1 3759.75 999.1 3764.36 ;
      RECT 833.1 3766.36 999.1 3775.58 ;
      RECT 873.1 3777.58 999.1 3782.19 ;
      RECT 793.1 3784.19 999.1 3785.31 ;
      RECT 953.1 3793.43 999.1 3799.2 ;
      RECT 913.1 3801.2 999.1 3812.74 ;
      RECT 953.1 3814.74 999.1 3820.51 ;
      RECT 793.1 3828.63 999.1 3829.75 ;
      RECT 873.1 3831.75 999.1 3836.36 ;
      RECT 833.1 3838.36 999.1 3847.58 ;
      RECT 873.1 3849.58 999.1 3854.19 ;
      RECT 793.1 3856.19 999.1 3857.31 ;
      RECT 953.1 3865.43 999.1 3871.2 ;
      RECT 913.1 3873.2 999.1 3884.74 ;
      RECT 953.1 3886.74 999.1 3892.51 ;
      RECT 793.1 3900.63 999.1 3901.75 ;
      RECT 873.1 3903.75 999.1 3908.36 ;
      RECT 833.1 3910.36 999.1 3919.58 ;
      RECT 873.1 3921.58 999.1 3926.19 ;
      RECT 793.1 3928.19 999.1 3929.31 ;
      RECT 953.1 3937.43 999.1 3943.2 ;
      RECT 913.1 3945.2 999.1 3956.74 ;
      RECT 953.1 3958.74 999.1 3964.51 ;
      RECT 793.1 3972.63 999.1 3973.75 ;
      RECT 873.1 3975.75 999.1 3980.36 ;
      RECT 833.1 3982.36 999.1 3991.58 ;
      RECT 873.1 3993.58 999.1 3998.19 ;
      RECT 793.1 4000.19 999.1 4001.31 ;
      RECT 953.1 4009.43 999.1 4015.2 ;
      RECT 913.1 4017.2 999.1 4028.74 ;
      RECT 953.1 4030.74 999.1 4036.51 ;
      RECT 793.1 4044.63 999.1 4045.75 ;
      RECT 873.1 4047.75 999.1 4052.36 ;
      RECT 833.1 4054.36 999.1 4063.58 ;
      RECT 873.1 4065.58 999.1 4070.19 ;
      RECT 793.1 4072.19 999.1 4073.31 ;
      RECT 953.1 4081.43 999.1 4087.2 ;
      RECT 913.1 4089.2 999.1 4100.74 ;
      RECT 953.1 4102.74 999.1 4108.51 ;
      RECT 793.1 4116.63 999.1 4117.75 ;
      RECT 873.1 4119.75 999.1 4124.36 ;
      RECT 833.1 4126.36 999.1 4135.58 ;
      RECT 873.1 4137.58 999.1 4142.19 ;
      RECT 793.1 4144.19 999.1 4145.31 ;
      RECT 953.1 4153.43 999.1 4159.2 ;
      RECT 913.1 4161.2 999.1 4172.74 ;
      RECT 953.1 4174.74 999.1 4180.51 ;
      RECT 793.1 4188.63 999.1 4189.75 ;
      RECT 873.1 4191.75 999.1 4196.36 ;
      RECT 833.1 4198.36 999.1 4207.58 ;
      RECT 873.1 4209.58 999.1 4214.19 ;
      RECT 793.1 4216.19 999.1 4217.31 ;
      RECT 953.1 4225.43 999.1 4231.2 ;
      RECT 913.1 4233.2 999.1 4244.74 ;
      RECT 953.1 4246.74 999.1 4252.51 ;
      RECT 793.1 4260.63 999.1 4261.75 ;
      RECT 873.1 4263.75 999.1 4268.36 ;
      RECT 833.1 4270.36 999.1 4279.58 ;
      RECT 873.1 4281.58 999.1 4286.19 ;
      RECT 793.1 4288.19 999.1 4289.31 ;
      RECT 953.1 4297.43 999.1 4303.2 ;
      RECT 913.1 4305.2 999.1 4316.74 ;
      RECT 953.1 4318.74 999.1 4324.51 ;
      RECT 793.1 4332.63 999.1 4333.75 ;
      RECT 873.1 4335.75 999.1 4340.36 ;
      RECT 833.1 4342.36 999.1 4351.58 ;
      RECT 873.1 4353.58 999.1 4358.19 ;
      RECT 793.1 4360.19 999.1 4361.31 ;
      RECT 953.1 4369.43 999.1 4375.2 ;
      RECT 913.1 4377.2 999.1 4388.74 ;
      RECT 953.1 4390.74 999.1 4396.51 ;
      RECT 793.1 4404.63 999.1 4405.75 ;
      RECT 873.1 4407.75 999.1 4412.36 ;
      RECT 833.1 4414.36 999.1 4423.58 ;
      RECT 873.1 4425.58 999.1 4430.19 ;
      RECT 793.1 4432.19 999.1 4433.31 ;
      RECT 953.1 4441.43 999.1 4447.2 ;
      RECT 913.1 4449.2 999.1 4460.74 ;
      RECT 953.1 4462.74 999.1 4468.51 ;
      RECT 793.1 4476.63 999.1 4477.75 ;
      RECT 873.1 4479.75 999.1 4484.36 ;
      RECT 833.1 4486.36 999.1 4495.58 ;
      RECT 873.1 4497.58 999.1 4502.19 ;
      RECT 793.1 4504.19 999.1 4505.31 ;
      RECT 953.1 4513.43 999.1 4519.2 ;
      RECT 913.1 4521.2 999.1 4532.74 ;
      RECT 953.1 4534.74 999.1 4540.51 ;
      RECT 793.1 4548.63 999.1 4549.75 ;
      RECT 873.1 4551.75 999.1 4556.36 ;
      RECT 833.1 4558.36 999.1 4567.58 ;
      RECT 873.1 4569.58 999.1 4574.19 ;
      RECT 793.1 4576.19 999.1 4577.31 ;
      RECT 953.1 4585.43 999.1 4591.2 ;
      RECT 913.1 4593.2 999.1 4604.74 ;
      RECT 953.1 4606.74 999.1 4612.51 ;
      RECT 793.1 4620.63 999.1 4621.75 ;
      RECT 873.1 4623.75 999.1 4628.36 ;
      RECT 833.1 4630.36 999.1 4639.58 ;
      RECT 873.1 4641.58 999.1 4646.19 ;
      RECT 793.1 4648.19 999.1 4649.31 ;
      RECT 953.1 4657.43 999.1 4663.2 ;
      RECT 913.1 4665.2 999.1 4676.74 ;
      RECT 953.1 4678.74 999.1 4684.51 ;
      RECT 793.1 4692.63 999.1 4693.75 ;
      RECT 873.1 4695.75 999.1 4700.36 ;
      RECT 833.1 4702.36 999.1 4711.58 ;
      RECT 873.1 4713.58 999.1 4718.19 ;
      RECT 793.1 4720.19 999.1 4721.31 ;
      RECT 953.1 4729.43 999.1 4735.2 ;
      RECT 913.1 4737.2 999.1 4748.74 ;
      RECT 953.1 4750.74 999.1 4756.51 ;
      RECT 793.1 4764.63 999.1 4765.75 ;
      RECT 873.1 4767.75 999.1 4772.36 ;
      RECT 833.1 4774.36 999.1 4783.58 ;
      RECT 873.1 4785.58 999.1 4790.19 ;
      RECT 793.1 4792.19 999.1 4793.31 ;
      RECT 953.1 4801.43 999.1 4807.2 ;
      RECT 913.1 4809.2 999.1 4820.74 ;
      RECT 953.1 4822.74 999.1 4828.51 ;
      RECT 793.1 4836.63 999.1 4837.75 ;
      RECT 873.1 4839.75 999.1 4844.36 ;
      RECT 833.1 4846.36 999.1 4855.58 ;
      RECT 873.1 4857.58 999.1 4862.19 ;
      RECT 793.1 4864.19 999.1 4865.31 ;
      RECT 953.1 4873.43 999.1 4879.2 ;
      RECT 913.1 4881.2 999.1 4892.74 ;
      RECT 953.1 4894.74 999.1 4900.51 ;
      RECT 793.1 4908.63 999.1 4909.75 ;
      RECT 873.1 4911.75 999.1 4916.36 ;
      RECT 833.1 4918.36 999.1 4927.58 ;
      RECT 873.1 4929.58 999.1 4934.19 ;
      RECT 793.1 4936.19 999.1 4937.31 ;
      RECT 953.1 4945.43 999.1 4951.2 ;
      RECT 913.1 4953.2 999.1 4964.74 ;
      RECT 953.1 4966.74 999.1 4972.51 ;
      RECT 793.1 4980.63 999.1 4981.75 ;
      RECT 873.1 4983.75 999.1 4988.36 ;
      RECT 833.1 4990.36 999.1 4999.58 ;
      RECT 873.1 5001.58 999.1 5006.19 ;
      RECT 793.1 5008.19 999.1 5009.31 ;
      RECT 953.1 5017.43 999.1 5023.2 ;
      RECT 913.1 5025.2 999.1 5036.74 ;
      RECT 953.1 5038.74 999.1 5044.51 ;
      RECT 793.1 5052.63 999.1 5053.75 ;
      RECT 873.1 5055.75 999.1 5060.36 ;
      RECT 833.1 5062.36 999.1 5071.58 ;
      RECT 873.1 5073.58 999.1 5078.19 ;
      RECT 793.1 5080.19 999.1 5081.31 ;
      RECT 953.1 5089.43 999.1 5095.2 ;
      RECT 913.1 5097.2 999.1 5108.74 ;
      RECT 953.1 5110.74 999.1 5116.51 ;
      RECT 793.1 5124.63 999.1 5125.75 ;
      RECT 873.1 5127.75 999.1 5132.36 ;
      RECT 833.1 5134.36 999.1 5143.58 ;
      RECT 873.1 5145.58 999.1 5150.19 ;
      RECT 793.1 5152.19 999.1 5153.31 ;
      RECT 953.1 5161.43 999.1 5167.2 ;
      RECT 913.1 5169.2 999.1 5180.74 ;
      RECT 953.1 5182.74 999.1 5188.51 ;
      RECT 793.1 5196.63 999.1 5197.75 ;
      RECT 873.1 5199.75 999.1 5204.36 ;
      RECT 833.1 5206.36 999.1 5215.58 ;
      RECT 873.1 5217.58 999.1 5222.19 ;
      RECT 793.1 5224.19 999.1 5225.31 ;
      RECT 953.1 5233.43 999.1 5239.2 ;
      RECT 913.1 5241.2 999.1 5252.74 ;
      RECT 953.1 5254.74 999.1 5260.51 ;
      RECT 793.1 5268.63 999.1 5269.75 ;
      RECT 873.1 5271.75 999.1 5276.36 ;
      RECT 833.1 5278.36 999.1 5287.58 ;
      RECT 873.1 5289.58 999.1 5294.19 ;
      RECT 793.1 5296.19 999.1 5297.31 ;
      RECT 953.1 5305.43 999.1 5311.2 ;
      RECT 913.1 5313.2 999.1 5324.74 ;
      RECT 953.1 5326.74 999.1 5332.51 ;
      RECT 793.1 5340.63 999.1 5341.75 ;
      RECT 873.1 5343.75 999.1 5348.36 ;
      RECT 833.1 5350.36 999.1 5359.58 ;
      RECT 873.1 5361.58 999.1 5366.19 ;
      RECT 793.1 5368.19 999.1 5369.31 ;
      RECT 953.1 5377.43 999.1 5383.2 ;
      RECT 913.1 5385.2 999.1 5396.74 ;
      RECT 953.1 5398.74 999.1 5404.51 ;
      RECT 793.1 5412.63 999.1 5413.75 ;
      RECT 873.1 5415.75 999.1 5420.36 ;
      RECT 833.1 5422.36 999.1 5431.58 ;
      RECT 873.1 5433.58 999.1 5438.19 ;
      RECT 793.1 5440.19 999.1 5441.31 ;
      RECT 953.1 5449.43 999.1 5455.2 ;
      RECT 913.1 5457.2 999.1 5468.74 ;
      RECT 953.1 5470.74 999.1 5476.51 ;
      RECT 793.1 5484.63 999.1 5485.75 ;
      RECT 873.1 5487.75 999.1 5492.36 ;
      RECT 833.1 5494.36 999.1 5503.58 ;
      RECT 873.1 5505.58 999.1 5510.19 ;
      RECT 793.1 5512.19 999.1 5513.31 ;
      RECT 953.1 5521.43 999.1 5527.2 ;
      RECT 913.1 5529.2 999.1 5540.74 ;
      RECT 953.1 5542.74 999.1 5548.51 ;
      RECT 793.1 5556.63 999.1 5557.75 ;
      RECT 873.1 5559.75 999.1 5564.36 ;
      RECT 833.1 5566.36 999.1 5575.58 ;
      RECT 873.1 5577.58 999.1 5582.19 ;
      RECT 793.1 5584.19 999.1 5585.31 ;
      RECT 953.1 5593.43 999.1 5599.2 ;
      RECT 913.1 5601.2 999.1 5612.74 ;
      RECT 953.1 5614.74 999.1 5620.51 ;
      RECT 793.1 5628.63 999.1 5629.75 ;
      RECT 873.1 5631.75 999.1 5636.36 ;
      RECT 833.1 5638.36 999.1 5647.58 ;
      RECT 873.1 5649.58 999.1 5654.19 ;
      RECT 793.1 5656.19 999.1 5657.31 ;
      RECT 953.1 5665.43 999.1 5671.2 ;
      RECT 913.1 5673.2 999.1 5684.74 ;
      RECT 953.1 5686.74 999.1 5692.51 ;
      RECT 793.1 5700.63 999.1 5701.75 ;
      RECT 873.1 5703.75 999.1 5708.36 ;
      RECT 833.1 5710.36 999.1 5719.58 ;
      RECT 873.1 5721.58 999.1 5726.19 ;
      RECT 793.1 5728.19 999.1 5729.31 ;
      RECT 953.1 5737.43 999.1 5743.2 ;
      RECT 913.1 5745.2 999.1 5756.74 ;
      RECT 953.1 5758.74 999.1 5764.51 ;
      RECT 793.1 5772.63 999.1 5773.75 ;
      RECT 873.1 5775.75 999.1 5780.36 ;
      RECT 833.1 5782.36 999.1 5791.58 ;
      RECT 873.1 5793.58 999.1 5798.19 ;
      RECT 793.1 5800.19 999.1 5801.31 ;
      RECT 953.1 5809.43 999.1 5815.2 ;
      RECT 913.1 5817.2 999.1 5828.74 ;
      RECT 953.1 5830.74 999.1 5836.51 ;
      RECT 793.1 5844.63 999.1 5845.75 ;
      RECT 873.1 5847.75 999.1 5852.36 ;
      RECT 833.1 5854.36 999.1 5863.58 ;
      RECT 873.1 5865.58 999.1 5870.19 ;
      RECT 793.1 5872.19 999.1 5873.31 ;
      RECT 953.1 5881.43 999.1 5887.2 ;
      RECT 913.1 5889.2 999.1 5900.74 ;
      RECT 953.1 5902.74 999.1 5908.51 ;
      RECT 793.1 5916.63 999.1 5917.75 ;
      RECT 873.1 5919.75 999.1 5924.36 ;
      RECT 833.1 5926.36 999.1 5935.58 ;
      RECT 873.1 5937.58 999.1 5942.19 ;
      RECT 793.1 5944.19 999.1 5945.31 ;
      RECT 953.1 5953.43 999.1 5959.2 ;
      RECT 913.1 5961.2 999.1 5972.74 ;
      RECT 953.1 5974.74 999.1 5980.51 ;
      RECT 793.1 5988.63 999.1 5989.75 ;
      RECT 873.1 5991.75 999.1 5996.36 ;
      RECT 833.1 5998.36 999.1 6007.58 ;
      RECT 873.1 6009.58 999.1 6014.19 ;
      RECT 793.1 6016.19 999.1 6017.31 ;
      RECT 953.1 6025.43 999.1 6031.2 ;
      RECT 913.1 6033.2 999.1 6044.74 ;
      RECT 953.1 6046.74 999.1 6052.51 ;
      RECT 793.1 6060.63 999.1 6061.75 ;
      RECT 873.1 6063.75 999.1 6068.36 ;
      RECT 833.1 6070.36 999.1 6079.58 ;
      RECT 873.1 6081.58 999.1 6086.19 ;
      RECT 793.1 6088.19 999.1 6089.31 ;
      RECT 953.1 6097.43 999.1 6103.2 ;
      RECT 913.1 6105.2 999.1 6116.74 ;
      RECT 953.1 6118.74 999.1 6124.51 ;
      RECT 793.1 6132.63 999.1 6133.75 ;
      RECT 873.1 6135.75 999.1 6140.36 ;
      RECT 833.1 6142.36 999.1 6151.58 ;
      RECT 873.1 6153.58 999.1 6158.19 ;
      RECT 793.1 6160.19 999.1 6161.31 ;
      RECT 953.1 6169.43 999.1 6175.2 ;
      RECT 913.1 6177.2 999.1 6188.74 ;
      RECT 953.1 6190.74 999.1 6196.51 ;
      RECT 793.1 6204.63 999.1 6205.75 ;
      RECT 873.1 6207.75 999.1 6212.36 ;
      RECT 833.1 6214.36 999.1 6223.58 ;
      RECT 873.1 6225.58 999.1 6230.19 ;
      RECT 793.1 6232.19 999.1 6233.31 ;
      RECT 953.1 6241.43 999.1 6247.2 ;
      RECT 913.1 6249.2 999.1 6260.74 ;
      RECT 953.1 6262.74 999.1 6268.51 ;
      RECT 793.1 6276.63 999.1 6277.75 ;
      RECT 873.1 6279.75 999.1 6284.36 ;
      RECT 833.1 6286.36 999.1 6295.58 ;
      RECT 873.1 6297.58 999.1 6302.19 ;
      RECT 793.1 6304.19 999.1 6305.31 ;
      RECT 953.1 6313.43 999.1 6319.2 ;
      RECT 913.1 6321.2 999.1 6332.74 ;
      RECT 953.1 6334.74 999.1 6340.51 ;
      RECT 793.1 6348.63 999.1 6349.75 ;
      RECT 873.1 6351.75 999.1 6356.36 ;
      RECT 833.1 6358.36 999.1 6367.58 ;
      RECT 873.1 6369.58 999.1 6374.19 ;
      RECT 793.1 6376.19 999.1 6377.31 ;
      RECT 953.1 6385.43 999.1 6391.2 ;
      RECT 913.1 6393.2 999.1 6404.74 ;
      RECT 953.1 6406.74 999.1 6412.51 ;
      RECT 793.1 6420.63 999.1 6421.75 ;
      RECT 873.1 6423.75 999.1 6428.36 ;
      RECT 833.1 6430.36 999.1 6439.58 ;
      RECT 873.1 6441.58 999.1 6446.19 ;
      RECT 793.1 6448.19 999.1 6449.31 ;
      RECT 953.1 6457.43 999.1 6463.2 ;
      RECT 913.1 6465.2 999.1 6476.74 ;
      RECT 953.1 6478.74 999.1 6484.51 ;
      RECT 793.1 6492.63 999.1 6493.75 ;
      RECT 873.1 6495.75 999.1 6500.36 ;
      RECT 833.1 6502.36 999.1 6511.58 ;
      RECT 873.1 6513.58 999.1 6518.19 ;
      RECT 793.1 6520.19 999.1 6521.31 ;
      RECT 953.1 6529.43 999.1 6535.2 ;
      RECT 913.1 6537.2 999.1 6548.74 ;
      RECT 953.1 6550.74 999.1 6556.51 ;
      RECT 793.1 6564.63 999.1 6565.75 ;
      RECT 873.1 6567.75 999.1 6572.36 ;
      RECT 833.1 6574.36 999.1 6583.58 ;
      RECT 873.1 6585.58 999.1 6590.19 ;
      RECT 793.1 6592.19 999.1 6593.31 ;
      RECT 953.1 6601.43 999.1 6607.2 ;
      RECT 913.1 6609.2 999.1 6620.74 ;
      RECT 953.1 6622.74 999.1 6628.51 ;
      RECT 793.1 6636.63 999.1 6637.75 ;
      RECT 873.1 6639.75 999.1 6644.36 ;
      RECT 833.1 6646.36 999.1 6655.58 ;
      RECT 873.1 6657.58 999.1 6662.19 ;
      RECT 793.1 6664.19 999.1 6665.31 ;
      RECT 953.1 6673.43 999.1 6679.2 ;
      RECT 913.1 6681.2 999.1 6692.74 ;
      RECT 953.1 6694.74 999.1 6700.51 ;
      RECT 793.1 6708.63 999.1 6709.75 ;
      RECT 873.1 6711.75 999.1 6716.36 ;
      RECT 833.1 6718.36 999.1 6727.58 ;
      RECT 873.1 6729.58 999.1 6734.19 ;
      RECT 793.1 6736.19 999.1 6737.31 ;
      RECT 953.1 6745.43 999.1 6751.2 ;
      RECT 913.1 6753.2 999.1 6764.74 ;
      RECT 953.1 6766.74 999.1 6772.51 ;
      RECT 793.1 6780.63 999.1 6781.75 ;
      RECT 873.1 6783.75 999.1 6788.36 ;
      RECT 833.1 6790.36 999.1 6799.58 ;
      RECT 873.1 6801.58 999.1 6806.19 ;
      RECT 793.1 6808.19 999.1 6809.31 ;
      RECT 953.1 6817.43 999.1 6823.2 ;
      RECT 913.1 6825.2 999.1 6836.74 ;
      RECT 953.1 6838.74 999.1 6844.51 ;
      RECT 793.1 6852.63 999.1 6853.75 ;
      RECT 873.1 6855.75 999.1 6860.36 ;
      RECT 833.1 6862.36 999.1 6871.58 ;
      RECT 873.1 6873.58 999.1 6878.19 ;
      RECT 793.1 6880.19 999.1 6881.31 ;
      RECT 953.1 6889.43 999.1 6895.2 ;
      RECT 913.1 6897.2 999.1 6908.74 ;
      RECT 953.1 6910.74 999.1 6916.51 ;
      RECT 793.1 6924.63 999.1 6925.75 ;
      RECT 873.1 6927.75 999.1 6932.36 ;
      RECT 833.1 6934.36 999.1 6943.58 ;
      RECT 873.1 6945.58 999.1 6950.19 ;
      RECT 793.1 6952.19 999.1 6953.31 ;
      RECT 953.1 6961.43 999.1 6967.2 ;
      RECT 913.1 6969.2 999.1 6980.74 ;
      RECT 953.1 6982.74 999.1 6988.51 ;
      RECT 793.1 6996.63 999.1 6997.75 ;
      RECT 873.1 6999.75 999.1 7004.36 ;
      RECT 833.1 7006.36 999.1 7015.58 ;
      RECT 873.1 7017.58 999.1 7022.19 ;
      RECT 793.1 7024.19 999.1 7025.31 ;
      RECT 953.1 7033.43 999.1 7039.2 ;
      RECT 913.1 7041.2 999.1 7052.74 ;
      RECT 953.1 7054.74 999.1 7060.51 ;
      RECT 793.1 7068.63 999.1 7069.75 ;
      RECT 873.1 7071.75 999.1 7076.36 ;
      RECT 833.1 7078.36 999.1 7087.58 ;
      RECT 873.1 7089.58 999.1 7094.19 ;
      RECT 793.1 7096.19 999.1 7097.31 ;
      RECT 953.1 7105.43 999.1 7111.2 ;
      RECT 913.1 7113.2 999.1 7124.74 ;
      RECT 953.1 7126.74 999.1 7132.51 ;
      RECT 793.1 7140.63 999.1 7141.75 ;
      RECT 873.1 7143.75 999.1 7148.36 ;
      RECT 833.1 7150.36 999.1 7159.58 ;
      RECT 873.1 7161.58 999.1 7166.19 ;
      RECT 793.1 7168.19 999.1 7169.31 ;
      RECT 953.1 7177.43 999.1 7183.2 ;
      RECT 913.1 7185.2 999.1 7196.74 ;
      RECT 953.1 7198.74 999.1 7204.51 ;
      RECT 793.1 7212.63 999.1 7213.75 ;
      RECT 873.1 7215.75 999.1 7220.36 ;
      RECT 833.1 7222.36 999.1 7231.58 ;
      RECT 873.1 7233.58 999.1 7238.19 ;
      RECT 793.1 7240.19 999.1 7241.31 ;
      RECT 953.1 7249.43 999.1 7255.2 ;
      RECT 913.1 7257.2 999.1 7268.74 ;
      RECT 953.1 7270.74 999.1 7276.51 ;
      RECT 793.1 7284.63 999.1 7285.75 ;
      RECT 873.1 7287.75 999.1 7292.36 ;
      RECT 833.1 7294.36 999.1 7303.58 ;
      RECT 873.1 7305.58 999.1 7310.19 ;
      RECT 793.1 7312.19 999.1 7313.31 ;
      RECT 953.1 7321.43 999.1 7327.2 ;
      RECT 913.1 7329.2 999.1 7340.74 ;
      RECT 953.1 7342.74 999.1 7348.51 ;
      RECT 793.1 7356.63 999.1 7357.75 ;
      RECT 873.1 7359.75 999.1 7364.36 ;
      RECT 833.1 7366.36 999.1 7375.58 ;
      RECT 873.1 7377.58 999.1 7382.19 ;
      RECT 793.1 7384.19 999.1 7385.31 ;
      RECT 953.1 7393.43 999.1 7399.2 ;
      RECT 913.1 7401.2 999.1 7412.74 ;
      RECT 953.1 7414.74 999.1 7420.51 ;
      RECT 793.1 7428.63 999.1 7429.75 ;
      RECT 873.1 7431.75 999.1 7436.36 ;
      RECT 833.1 7438.36 999.1 7447.58 ;
      RECT 873.1 7449.58 999.1 7454.19 ;
      RECT 793.1 7456.19 999.1 7457.31 ;
      RECT 953.1 7465.43 999.1 7471.2 ;
      RECT 913.1 7473.2 999.1 7484.74 ;
      RECT 953.1 7486.74 999.1 7492.51 ;
      RECT 793.1 7500.63 999.1 7501.75 ;
      RECT 873.1 7503.75 999.1 7508.36 ;
      RECT 833.1 7510.36 999.1 7519.58 ;
      RECT 873.1 7521.58 999.1 7526.19 ;
      RECT 793.1 7528.19 999.1 7529.31 ;
      RECT 953.1 7537.43 999.1 7543.2 ;
      RECT 913.1 7545.2 999.1 7556.74 ;
      RECT 953.1 7558.74 999.1 7564.51 ;
      RECT 793.1 7572.63 999.1 7573.75 ;
      RECT 873.1 7575.75 999.1 7580.36 ;
      RECT 833.1 7582.36 999.1 7591.58 ;
      RECT 873.1 7593.58 999.1 7598.19 ;
      RECT 793.1 7600.19 999.1 7601.31 ;
      RECT 953.1 7609.43 999.1 7615.2 ;
      RECT 913.1 7617.2 999.1 7628.74 ;
      RECT 953.1 7630.74 999.1 7636.51 ;
      RECT 793.1 7644.63 999.1 7645.75 ;
      RECT 873.1 7647.75 999.1 7652.36 ;
      RECT 833.1 7654.36 999.1 7663.58 ;
      RECT 873.1 7665.58 999.1 7670.19 ;
      RECT 793.1 7672.19 999.1 7673.31 ;
      RECT 953.1 7681.43 999.1 7687.2 ;
      RECT 913.1 7689.2 999.1 7700.74 ;
      RECT 953.1 7702.74 999.1 7708.51 ;
      RECT 793.1 7716.63 999.1 7717.75 ;
      RECT 873.1 7719.75 999.1 7724.36 ;
      RECT 833.1 7726.36 999.1 7735.58 ;
      RECT 873.1 7737.58 999.1 7742.19 ;
      RECT 793.1 7744.19 999.1 7745.31 ;
      RECT 953.1 7753.43 999.1 7759.2 ;
      RECT 913.1 7761.2 999.1 7772.74 ;
      RECT 953.1 7774.74 999.1 7780.51 ;
      RECT 793.1 7788.63 999.1 7789.75 ;
      RECT 873.1 7791.75 999.1 7796.36 ;
      RECT 833.1 7798.36 999.1 7807.58 ;
      RECT 873.1 7809.58 999.1 7814.19 ;
      RECT 793.1 7816.19 999.1 7817.31 ;
      RECT 953.1 7825.43 999.1 7831.2 ;
      RECT 913.1 7833.2 999.1 7844.74 ;
      RECT 953.1 7846.74 999.1 7852.51 ;
      RECT 793.1 7860.63 999.1 7861.75 ;
      RECT 873.1 7863.75 999.1 7868.36 ;
      RECT 833.1 7870.36 999.1 7879.58 ;
      RECT 873.1 7881.58 999.1 7886.19 ;
      RECT 793.1 7888.19 999.1 7889.31 ;
      RECT 953.1 7897.43 999.1 7903.2 ;
      RECT 913.1 7905.2 999.1 7916.74 ;
      RECT 953.1 7918.74 999.1 7924.51 ;
      RECT 793.1 7932.63 999.1 7933.75 ;
      RECT 873.1 7935.75 999.1 7940.36 ;
      RECT 833.1 7942.36 999.1 7951.58 ;
      RECT 873.1 7953.58 999.1 7958.19 ;
      RECT 793.1 7960.19 999.1 7961.31 ;
      RECT 953.1 7969.43 999.1 7975.2 ;
      RECT 913.1 7977.2 999.1 7988.74 ;
      RECT 953.1 7990.74 999.1 7996.51 ;
      RECT 793.1 8004.63 999.1 8005.75 ;
      RECT 873.1 8007.75 999.1 8012.36 ;
      RECT 833.1 8014.36 999.1 8023.58 ;
      RECT 873.1 8025.58 999.1 8030.19 ;
      RECT 793.1 8032.19 999.1 8033.31 ;
      RECT 953.1 8041.43 999.1 8047.2 ;
      RECT 913.1 8049.2 999.1 8060.74 ;
      RECT 953.1 8062.74 999.1 8068.51 ;
      RECT 793.1 8076.63 999.1 8077.75 ;
      RECT 873.1 8079.75 999.1 8084.36 ;
      RECT 833.1 8086.36 999.1 8095.58 ;
      RECT 873.1 8097.58 999.1 8102.19 ;
      RECT 793.1 8104.19 999.1 8105.31 ;
      RECT 953.1 8113.43 999.1 8119.2 ;
      RECT 913.1 8121.2 999.1 8132.74 ;
      RECT 953.1 8134.74 999.1 8140.51 ;
      RECT 793.1 8148.63 999.1 8149.75 ;
      RECT 873.1 8151.75 999.1 8156.36 ;
      RECT 833.1 8158.36 999.1 8167.58 ;
      RECT 873.1 8169.58 999.1 8174.19 ;
      RECT 793.1 8176.19 999.1 8177.31 ;
      RECT 953.1 8185.43 999.1 8191.2 ;
      RECT 913.1 8193.2 999.1 8204.74 ;
      RECT 953.1 8206.74 999.1 8212.51 ;
      RECT 793.1 8220.63 999.1 8221.75 ;
      RECT 873.1 8223.75 999.1 8228.36 ;
      RECT 833.1 8230.36 999.1 8239.58 ;
      RECT 873.1 8241.58 999.1 8246.19 ;
      RECT 793.1 8248.19 999.1 8249.31 ;
      RECT 953.1 8257.43 999.1 8263.2 ;
      RECT 913.1 8265.2 999.1 8276.74 ;
      RECT 953.1 8278.74 999.1 8284.51 ;
      RECT 793.1 8292.63 999.1 8293.75 ;
      RECT 873.1 8295.75 999.1 8300.36 ;
      RECT 833.1 8302.36 999.1 8311.58 ;
      RECT 873.1 8313.58 999.1 8318.19 ;
      RECT 793.1 8320.19 999.1 8321.31 ;
      RECT 953.1 8329.43 999.1 8335.2 ;
      RECT 913.1 8337.2 999.1 8348.74 ;
      RECT 953.1 8350.74 999.1 8356.51 ;
      RECT 793.1 8364.63 999.1 8365.75 ;
      RECT 873.1 8367.75 999.1 8372.36 ;
      RECT 833.1 8374.36 999.1 8383.58 ;
      RECT 873.1 8385.58 999.1 8390.19 ;
      RECT 793.1 8392.19 999.1 8393.31 ;
      RECT 953.1 8401.43 999.1 8407.2 ;
      RECT 913.1 8409.2 999.1 8420.74 ;
      RECT 953.1 8422.74 999.1 8428.51 ;
      RECT 793.1 8436.63 999.1 8437.75 ;
      RECT 873.1 8439.75 999.1 8444.36 ;
      RECT 833.1 8446.36 999.1 8455.58 ;
      RECT 873.1 8457.58 999.1 8462.19 ;
      RECT 793.1 8464.19 999.1 8465.31 ;
      RECT 953.1 8473.43 999.1 8479.2 ;
      RECT 913.1 8481.2 999.1 8492.74 ;
      RECT 953.1 8494.74 999.1 8500.51 ;
      RECT 793.1 8508.63 999.1 8509.75 ;
      RECT 873.1 8511.75 999.1 8516.36 ;
      RECT 833.1 8518.36 999.1 8527.58 ;
      RECT 873.1 8529.58 999.1 8534.19 ;
      RECT 793.1 8536.19 999.1 8537.31 ;
      RECT 953.1 8545.43 999.1 8551.2 ;
      RECT 913.1 8553.2 999.1 8564.74 ;
      RECT 953.1 8566.74 999.1 8572.51 ;
      RECT 793.1 8580.63 999.1 8581.75 ;
      RECT 873.1 8583.75 999.1 8588.36 ;
      RECT 833.1 8590.36 999.1 8599.58 ;
      RECT 873.1 8601.58 999.1 8606.19 ;
      RECT 793.1 8608.19 999.1 8609.31 ;
      RECT 953.1 8617.43 999.1 8623.2 ;
      RECT 913.1 8625.2 999.1 8636.74 ;
      RECT 953.1 8638.74 999.1 8644.51 ;
      RECT 793.1 8652.63 999.1 8653.75 ;
      RECT 873.1 8655.75 999.1 8660.36 ;
      RECT 833.1 8662.36 999.1 8671.58 ;
      RECT 873.1 8673.58 999.1 8678.19 ;
      RECT 793.1 8680.19 999.1 8681.31 ;
      RECT 953.1 8689.43 999.1 8695.2 ;
      RECT 913.1 8697.2 999.1 8708.74 ;
      RECT 953.1 8710.74 999.1 8716.51 ;
      RECT 793.1 8724.63 999.1 8725.75 ;
      RECT 873.1 8727.75 999.1 8732.36 ;
      RECT 833.1 8734.36 999.1 8743.58 ;
      RECT 873.1 8745.58 999.1 8750.19 ;
      RECT 793.1 8752.19 999.1 8753.31 ;
      RECT 953.1 8761.43 999.1 8767.2 ;
      RECT 913.1 8769.2 999.1 8780.74 ;
      RECT 953.1 8782.74 999.1 8788.51 ;
      RECT 793.1 8796.63 999.1 8797.75 ;
      RECT 873.1 8799.75 999.1 8804.36 ;
      RECT 833.1 8806.36 999.1 8815.58 ;
      RECT 873.1 8817.58 999.1 8822.19 ;
      RECT 793.1 8824.19 999.1 8825.31 ;
      RECT 953.1 8833.43 999.1 8839.2 ;
      RECT 913.1 8841.2 999.1 8852.74 ;
      RECT 953.1 8854.74 999.1 8860.51 ;
      RECT 793.1 8868.63 999.1 8869.75 ;
      RECT 873.1 8871.75 999.1 8876.36 ;
      RECT 833.1 8878.36 999.1 8887.58 ;
      RECT 873.1 8889.58 999.1 8894.19 ;
      RECT 793.1 8896.19 999.1 8897.31 ;
      RECT 953.1 8905.43 999.1 8911.2 ;
      RECT 913.1 8913.2 999.1 8924.74 ;
      RECT 953.1 8926.74 999.1 8932.51 ;
      RECT 793.1 8940.63 999.1 8941.75 ;
      RECT 873.1 8943.75 999.1 8948.36 ;
      RECT 833.1 8950.36 999.1 8959.58 ;
      RECT 873.1 8961.58 999.1 8966.19 ;
      RECT 793.1 8968.19 999.1 8969.31 ;
      RECT 953.1 8977.43 999.1 8983.2 ;
      RECT 913.1 8985.2 999.1 8996.74 ;
      RECT 953.1 8998.74 999.1 9004.51 ;
      RECT 793.1 9012.63 999.1 9013.75 ;
      RECT 873.1 9015.75 999.1 9020.36 ;
      RECT 833.1 9022.36 999.1 9031.58 ;
      RECT 873.1 9033.58 999.1 9038.19 ;
      RECT 793.1 9040.19 999.1 9041.31 ;
      RECT 953.1 9049.43 999.1 9055.2 ;
      RECT 913.1 9057.2 999.1 9068.74 ;
      RECT 953.1 9070.74 999.1 9076.51 ;
      RECT 793.1 9084.63 999.1 9085.75 ;
      RECT 873.1 9087.75 999.1 9092.36 ;
      RECT 833.1 9094.36 999.1 9103.58 ;
      RECT 873.1 9105.58 999.1 9110.19 ;
      RECT 793.1 9112.19 999.1 9113.31 ;
      RECT 953.1 9121.43 999.1 9127.2 ;
      RECT 913.1 9129.2 999.1 9140.74 ;
      RECT 953.1 9142.74 999.1 9148.51 ;
      RECT 793.1 9156.63 999.1 9157.75 ;
      RECT 873.1 9159.75 999.1 9164.36 ;
      RECT 833.1 9166.36 999.1 9175.58 ;
      RECT 873.1 9177.58 999.1 9182.19 ;
      RECT 793.1 9184.19 999.1 9185.31 ;
      RECT 953.1 9193.43 999.1 9199.2 ;
      RECT 913.1 9201.2 999.1 9212.74 ;
      RECT 953.1 9214.74 999.1 9220.51 ;
      RECT 793.1 9228.63 999.1 9229.75 ;
      RECT 873.1 9231.75 999.1 9236.36 ;
      RECT 833.1 9238.36 999.1 9247.58 ;
      RECT 873.1 9249.58 999.1 9254.19 ;
      RECT 793.1 9256.19 999.1 9257.31 ;
      RECT 953.1 9265.43 999.1 9271.2 ;
      RECT 913.1 9273.2 999.1 9284.74 ;
      RECT 953.1 9286.74 999.1 9292.51 ;
      RECT 793.1 9300.63 999.1 9301.75 ;
      RECT 873.1 9303.75 999.1 9308.36 ;
      RECT 833.1 9310.36 999.1 9319.58 ;
      RECT 873.1 9321.58 999.1 9326.19 ;
      RECT 793.1 9328.19 999.1 9329.31 ;
      RECT 953.1 9337.43 999.1 9343.2 ;
      RECT 913.1 9345.2 999.1 9356.74 ;
      RECT 953.1 9358.74 999.1 9364.51 ;
      RECT 793.1 9372.63 999.1 9373.75 ;
      RECT 873.1 9375.75 999.1 9380.36 ;
      RECT 833.1 9382.36 999.1 9391.58 ;
      RECT 873.1 9393.58 999.1 9398.19 ;
      RECT 793.1 9400.19 999.1 9401.31 ;
      RECT 953.1 9409.43 999.1 9415.2 ;
      RECT 913.1 9417.2 999.1 9428.74 ;
      RECT 953.1 9430.74 999.1 9436.51 ;
      RECT 793.1 9444.63 999.1 9445.75 ;
      RECT 873.1 9447.75 999.1 9452.36 ;
      RECT 833.1 9454.36 999.1 9458.97 ;
    LAYER TOP_M SPACING 0.46 ;
      RECT 998.1 1048.165 19161.9 10000 ;
      RECT 19047.23 1046.435 19161.9 10000 ;
      RECT 963.1 1238.18 19196.9 1292.55 ;
      RECT 724.1 1288.91 19475.9 1290.55 ;
      RECT 19454.63 1238.18 19475.9 1290.55 ;
      RECT 748.83 1265.55 19451.17 1290.55 ;
      RECT 724.1 1238.18 745.37 1290.55 ;
      RECT 19454.63 1238.18 19567.9 1288.18 ;
      RECT 632.1 1238.18 745.37 1288.18 ;
      RECT 748.83 1238.18 19451.17 1263.55 ;
      RECT 19030.25 1046.435 19032.77 10000 ;
      RECT 19014.73 1046.435 19015.79 10000 ;
      RECT 18984.21 1046.435 18985.27 10000 ;
      RECT 18967.23 1046.435 18969.75 10000 ;
      RECT 18950.25 1046.435 18952.77 10000 ;
      RECT 18934.73 1046.435 18935.79 10000 ;
      RECT 18904.21 1046.435 18905.27 10000 ;
      RECT 18887.23 1046.435 18889.75 10000 ;
      RECT 18870.25 1046.435 18872.77 10000 ;
      RECT 18854.73 1046.435 18855.79 10000 ;
      RECT 18824.21 1046.435 18825.27 10000 ;
      RECT 18807.23 1046.435 18809.75 10000 ;
      RECT 18790.25 1046.435 18792.77 10000 ;
      RECT 18774.73 1046.435 18775.79 10000 ;
      RECT 18744.21 1046.435 18745.27 10000 ;
      RECT 18727.23 1046.435 18729.75 10000 ;
      RECT 18710.25 1046.435 18712.77 10000 ;
      RECT 18694.73 1046.435 18695.79 10000 ;
      RECT 18664.21 1046.435 18665.27 10000 ;
      RECT 18647.23 1046.435 18649.75 10000 ;
      RECT 18630.25 1046.435 18632.77 10000 ;
      RECT 18614.73 1046.435 18615.79 10000 ;
      RECT 18584.21 1046.435 18585.27 10000 ;
      RECT 18567.23 1046.435 18569.75 10000 ;
      RECT 18550.25 1046.435 18552.77 10000 ;
      RECT 18534.73 1046.435 18535.79 10000 ;
      RECT 18504.21 1046.435 18505.27 10000 ;
      RECT 18487.23 1046.435 18489.75 10000 ;
      RECT 18470.25 1046.435 18472.77 10000 ;
      RECT 18454.73 1046.435 18455.79 10000 ;
      RECT 18424.21 1046.435 18425.27 10000 ;
      RECT 18407.23 1046.435 18409.75 10000 ;
      RECT 18390.25 1046.435 18392.77 10000 ;
      RECT 18374.73 1046.435 18375.79 10000 ;
      RECT 18344.21 1046.435 18345.27 10000 ;
      RECT 18327.23 1046.435 18329.75 10000 ;
      RECT 18310.25 1046.435 18312.77 10000 ;
      RECT 18294.73 1046.435 18295.79 10000 ;
      RECT 18264.21 1046.435 18265.27 10000 ;
      RECT 18247.23 1046.435 18249.75 10000 ;
      RECT 18230.25 1046.435 18232.77 10000 ;
      RECT 18214.73 1046.435 18215.79 10000 ;
      RECT 18184.21 1046.435 18185.27 10000 ;
      RECT 18167.23 1046.435 18169.75 10000 ;
      RECT 18150.25 1046.435 18152.77 10000 ;
      RECT 18134.73 1046.435 18135.79 10000 ;
      RECT 18104.21 1046.435 18105.27 10000 ;
      RECT 18087.23 1046.435 18089.75 10000 ;
      RECT 18070.25 1046.435 18072.77 10000 ;
      RECT 18054.73 1046.435 18055.79 10000 ;
      RECT 18024.21 1046.435 18025.27 10000 ;
      RECT 18007.23 1046.435 18009.75 10000 ;
      RECT 17990.25 1046.435 17992.77 10000 ;
      RECT 17974.73 1046.435 17975.79 10000 ;
      RECT 17944.21 1046.435 17945.27 10000 ;
      RECT 17927.23 1046.435 17929.75 10000 ;
      RECT 17910.25 1046.435 17912.77 10000 ;
      RECT 17894.73 1046.435 17895.79 10000 ;
      RECT 17864.21 1046.435 17865.27 10000 ;
      RECT 17847.23 1046.435 17849.75 10000 ;
      RECT 17830.25 1046.435 17832.77 10000 ;
      RECT 17814.73 1046.435 17815.79 10000 ;
      RECT 17784.21 1046.435 17785.27 10000 ;
      RECT 17767.23 1046.435 17769.75 10000 ;
      RECT 17750.25 1046.435 17752.77 10000 ;
      RECT 17734.73 1046.435 17735.79 10000 ;
      RECT 17704.21 1046.435 17705.27 10000 ;
      RECT 17687.23 1046.435 17689.75 10000 ;
      RECT 17670.25 1046.435 17672.77 10000 ;
      RECT 17654.73 1046.435 17655.79 10000 ;
      RECT 17624.21 1046.435 17625.27 10000 ;
      RECT 17607.23 1046.435 17609.75 10000 ;
      RECT 17590.25 1046.435 17592.77 10000 ;
      RECT 17574.73 1046.435 17575.79 10000 ;
      RECT 17544.21 1046.435 17545.27 10000 ;
      RECT 17527.23 1046.435 17529.75 10000 ;
      RECT 17510.25 1046.435 17512.77 10000 ;
      RECT 17494.73 1046.435 17495.79 10000 ;
      RECT 17464.21 1046.435 17465.27 10000 ;
      RECT 17447.23 1046.435 17449.75 10000 ;
      RECT 17430.25 1046.435 17432.77 10000 ;
      RECT 17414.73 1046.435 17415.79 10000 ;
      RECT 17384.21 1046.435 17385.27 10000 ;
      RECT 17367.23 1046.435 17369.75 10000 ;
      RECT 17350.25 1046.435 17352.77 10000 ;
      RECT 17334.73 1046.435 17335.79 10000 ;
      RECT 17304.21 1046.435 17305.27 10000 ;
      RECT 17287.23 1046.435 17289.75 10000 ;
      RECT 17270.25 1046.435 17272.77 10000 ;
      RECT 17254.73 1046.435 17255.79 10000 ;
      RECT 17224.21 1046.435 17225.27 10000 ;
      RECT 17207.23 1046.435 17209.75 10000 ;
      RECT 17190.25 1046.435 17192.77 10000 ;
      RECT 17174.73 1046.435 17175.79 10000 ;
      RECT 17144.21 1046.435 17145.27 10000 ;
      RECT 17127.23 1046.435 17129.75 10000 ;
      RECT 17110.25 1046.435 17112.77 10000 ;
      RECT 17094.73 1046.435 17095.79 10000 ;
      RECT 17064.21 1046.435 17065.27 10000 ;
      RECT 17047.23 1046.435 17049.75 10000 ;
      RECT 17030.25 1046.435 17032.77 10000 ;
      RECT 17014.73 1046.435 17015.79 10000 ;
      RECT 16984.21 1046.435 16985.27 10000 ;
      RECT 16967.23 1046.435 16969.75 10000 ;
      RECT 16950.25 1046.435 16952.77 10000 ;
      RECT 16934.73 1046.435 16935.79 10000 ;
      RECT 16904.21 1046.435 16905.27 10000 ;
      RECT 16887.23 1046.435 16889.75 10000 ;
      RECT 16870.25 1046.435 16872.77 10000 ;
      RECT 16854.73 1046.435 16855.79 10000 ;
      RECT 16824.21 1046.435 16825.27 10000 ;
      RECT 16807.23 1046.435 16809.75 10000 ;
      RECT 16790.25 1046.435 16792.77 10000 ;
      RECT 16774.73 1046.435 16775.79 10000 ;
      RECT 16744.21 1046.435 16745.27 10000 ;
      RECT 16727.23 1046.435 16729.75 10000 ;
      RECT 16710.25 1046.435 16712.77 10000 ;
      RECT 16694.73 1046.435 16695.79 10000 ;
      RECT 16664.21 1046.435 16665.27 10000 ;
      RECT 16647.23 1046.435 16649.75 10000 ;
      RECT 16630.25 1046.435 16632.77 10000 ;
      RECT 16614.73 1046.435 16615.79 10000 ;
      RECT 16584.21 1046.435 16585.27 10000 ;
      RECT 16567.23 1046.435 16569.75 10000 ;
      RECT 16550.25 1046.435 16552.77 10000 ;
      RECT 16534.73 1046.435 16535.79 10000 ;
      RECT 16504.21 1046.435 16505.27 10000 ;
      RECT 16487.23 1046.435 16489.75 10000 ;
      RECT 16470.25 1046.435 16472.77 10000 ;
      RECT 16454.73 1046.435 16455.79 10000 ;
      RECT 16424.21 1046.435 16425.27 10000 ;
      RECT 16407.23 1046.435 16409.75 10000 ;
      RECT 16390.25 1046.435 16392.77 10000 ;
      RECT 16374.73 1046.435 16375.79 10000 ;
      RECT 16344.21 1046.435 16345.27 10000 ;
      RECT 16327.23 1046.435 16329.75 10000 ;
      RECT 16310.25 1046.435 16312.77 10000 ;
      RECT 16294.73 1046.435 16295.79 10000 ;
      RECT 16264.21 1046.435 16265.27 10000 ;
      RECT 16247.23 1046.435 16249.75 10000 ;
      RECT 16230.25 1046.435 16232.77 10000 ;
      RECT 16214.73 1046.435 16215.79 10000 ;
      RECT 16184.21 1046.435 16185.27 10000 ;
      RECT 16167.23 1046.435 16169.75 10000 ;
      RECT 16150.25 1046.435 16152.77 10000 ;
      RECT 16134.73 1046.435 16135.79 10000 ;
      RECT 16104.21 1046.435 16105.27 10000 ;
      RECT 16087.23 1046.435 16089.75 10000 ;
      RECT 16070.25 1046.435 16072.77 10000 ;
      RECT 16054.73 1046.435 16055.79 10000 ;
      RECT 16024.21 1046.435 16025.27 10000 ;
      RECT 16007.23 1046.435 16009.75 10000 ;
      RECT 15990.25 1046.435 15992.77 10000 ;
      RECT 15974.73 1046.435 15975.79 10000 ;
      RECT 15944.21 1046.435 15945.27 10000 ;
      RECT 15927.23 1046.435 15929.75 10000 ;
      RECT 15910.25 1046.435 15912.77 10000 ;
      RECT 15894.73 1046.435 15895.79 10000 ;
      RECT 15864.21 1046.435 15865.27 10000 ;
      RECT 15847.23 1046.435 15849.75 10000 ;
      RECT 15830.25 1046.435 15832.77 10000 ;
      RECT 15814.73 1046.435 15815.79 10000 ;
      RECT 15784.21 1046.435 15785.27 10000 ;
      RECT 15767.23 1046.435 15769.75 10000 ;
      RECT 15750.25 1046.435 15752.77 10000 ;
      RECT 15734.73 1046.435 15735.79 10000 ;
      RECT 15704.21 1046.435 15705.27 10000 ;
      RECT 15687.23 1046.435 15689.75 10000 ;
      RECT 15670.25 1046.435 15672.77 10000 ;
      RECT 15654.73 1046.435 15655.79 10000 ;
      RECT 15624.21 1046.435 15625.27 10000 ;
      RECT 15607.23 1046.435 15609.75 10000 ;
      RECT 15590.25 1046.435 15592.77 10000 ;
      RECT 15574.73 1046.435 15575.79 10000 ;
      RECT 15544.21 1046.435 15545.27 10000 ;
      RECT 15527.23 1046.435 15529.75 10000 ;
      RECT 15510.25 1046.435 15512.77 10000 ;
      RECT 15494.73 1046.435 15495.79 10000 ;
      RECT 15464.21 1046.435 15465.27 10000 ;
      RECT 15447.23 1046.435 15449.75 10000 ;
      RECT 15430.25 1046.435 15432.77 10000 ;
      RECT 15414.73 1046.435 15415.79 10000 ;
      RECT 15384.21 1046.435 15385.27 10000 ;
      RECT 15367.23 1046.435 15369.75 10000 ;
      RECT 15350.25 1046.435 15352.77 10000 ;
      RECT 15334.73 1046.435 15335.79 10000 ;
      RECT 15304.21 1046.435 15305.27 10000 ;
      RECT 15287.23 1046.435 15289.75 10000 ;
      RECT 15270.25 1046.435 15272.77 10000 ;
      RECT 15254.73 1046.435 15255.79 10000 ;
      RECT 15224.21 1046.435 15225.27 10000 ;
      RECT 15207.23 1046.435 15209.75 10000 ;
      RECT 15190.25 1046.435 15192.77 10000 ;
      RECT 15174.73 1046.435 15175.79 10000 ;
      RECT 15144.21 1046.435 15145.27 10000 ;
      RECT 15127.23 1046.435 15129.75 10000 ;
      RECT 15110.25 1046.435 15112.77 10000 ;
      RECT 15094.73 1046.435 15095.79 10000 ;
      RECT 15064.21 1046.435 15065.27 10000 ;
      RECT 15047.23 1046.435 15049.75 10000 ;
      RECT 15030.25 1046.435 15032.77 10000 ;
      RECT 15014.73 1046.435 15015.79 10000 ;
      RECT 14984.21 1046.435 14985.27 10000 ;
      RECT 14967.23 1046.435 14969.75 10000 ;
      RECT 14950.25 1046.435 14952.77 10000 ;
      RECT 14934.73 1046.435 14935.79 10000 ;
      RECT 14904.21 1046.435 14905.27 10000 ;
      RECT 14887.23 1046.435 14889.75 10000 ;
      RECT 14870.25 1046.435 14872.77 10000 ;
      RECT 14854.73 1046.435 14855.79 10000 ;
      RECT 14824.21 1046.435 14825.27 10000 ;
      RECT 14807.23 1046.435 14809.75 10000 ;
      RECT 14790.25 1046.435 14792.77 10000 ;
      RECT 14774.73 1046.435 14775.79 10000 ;
      RECT 14744.21 1046.435 14745.27 10000 ;
      RECT 14727.23 1046.435 14729.75 10000 ;
      RECT 14710.25 1046.435 14712.77 10000 ;
      RECT 14694.73 1046.435 14695.79 10000 ;
      RECT 14664.21 1046.435 14665.27 10000 ;
      RECT 14647.23 1046.435 14649.75 10000 ;
      RECT 14630.25 1046.435 14632.77 10000 ;
      RECT 14614.73 1046.435 14615.79 10000 ;
      RECT 14584.21 1046.435 14585.27 10000 ;
      RECT 14567.23 1046.435 14569.75 10000 ;
      RECT 14550.25 1046.435 14552.77 10000 ;
      RECT 14534.73 1046.435 14535.79 10000 ;
      RECT 14504.21 1046.435 14505.27 10000 ;
      RECT 14487.23 1046.435 14489.75 10000 ;
      RECT 14470.25 1046.435 14472.77 10000 ;
      RECT 14454.73 1046.435 14455.79 10000 ;
      RECT 14424.21 1046.435 14425.27 10000 ;
      RECT 14407.23 1046.435 14409.75 10000 ;
      RECT 14390.25 1046.435 14392.77 10000 ;
      RECT 14374.73 1046.435 14375.79 10000 ;
      RECT 14344.21 1046.435 14345.27 10000 ;
      RECT 14327.23 1046.435 14329.75 10000 ;
      RECT 14310.25 1046.435 14312.77 10000 ;
      RECT 14294.73 1046.435 14295.79 10000 ;
      RECT 14264.21 1046.435 14265.27 10000 ;
      RECT 14247.23 1046.435 14249.75 10000 ;
      RECT 14230.25 1046.435 14232.77 10000 ;
      RECT 14214.73 1046.435 14215.79 10000 ;
      RECT 14184.21 1046.435 14185.27 10000 ;
      RECT 14167.23 1046.435 14169.75 10000 ;
      RECT 14150.25 1046.435 14152.77 10000 ;
      RECT 14134.73 1046.435 14135.79 10000 ;
      RECT 14104.21 1046.435 14105.27 10000 ;
      RECT 14087.23 1046.435 14089.75 10000 ;
      RECT 14070.25 1046.435 14072.77 10000 ;
      RECT 14054.73 1046.435 14055.79 10000 ;
      RECT 14024.21 1046.435 14025.27 10000 ;
      RECT 14007.23 1046.435 14009.75 10000 ;
      RECT 13990.25 1046.435 13992.77 10000 ;
      RECT 13974.73 1046.435 13975.79 10000 ;
      RECT 13944.21 1046.435 13945.27 10000 ;
      RECT 13927.23 1046.435 13929.75 10000 ;
      RECT 13910.25 1046.435 13912.77 10000 ;
      RECT 13894.73 1046.435 13895.79 10000 ;
      RECT 13864.21 1046.435 13865.27 10000 ;
      RECT 13847.23 1046.435 13849.75 10000 ;
      RECT 13830.25 1046.435 13832.77 10000 ;
      RECT 13814.73 1046.435 13815.79 10000 ;
      RECT 13784.21 1046.435 13785.27 10000 ;
      RECT 13767.23 1046.435 13769.75 10000 ;
      RECT 13750.25 1046.435 13752.77 10000 ;
      RECT 13734.73 1046.435 13735.79 10000 ;
      RECT 13704.21 1046.435 13705.27 10000 ;
      RECT 13687.23 1046.435 13689.75 10000 ;
      RECT 13670.25 1046.435 13672.77 10000 ;
      RECT 13654.73 1046.435 13655.79 10000 ;
      RECT 13624.21 1046.435 13625.27 10000 ;
      RECT 13607.23 1046.435 13609.75 10000 ;
      RECT 13590.25 1046.435 13592.77 10000 ;
      RECT 13574.73 1046.435 13575.79 10000 ;
      RECT 13544.21 1046.435 13545.27 10000 ;
      RECT 13527.23 1046.435 13529.75 10000 ;
      RECT 13510.25 1046.435 13512.77 10000 ;
      RECT 13494.73 1046.435 13495.79 10000 ;
      RECT 13464.21 1046.435 13465.27 10000 ;
      RECT 13447.23 1046.435 13449.75 10000 ;
      RECT 13430.25 1046.435 13432.77 10000 ;
      RECT 13414.73 1046.435 13415.79 10000 ;
      RECT 13384.21 1046.435 13385.27 10000 ;
      RECT 13367.23 1046.435 13369.75 10000 ;
      RECT 13350.25 1046.435 13352.77 10000 ;
      RECT 13334.73 1046.435 13335.79 10000 ;
      RECT 13304.21 1046.435 13305.27 10000 ;
      RECT 13287.23 1046.435 13289.75 10000 ;
      RECT 13270.25 1046.435 13272.77 10000 ;
      RECT 13254.73 1046.435 13255.79 10000 ;
      RECT 13224.21 1046.435 13225.27 10000 ;
      RECT 13207.23 1046.435 13209.75 10000 ;
      RECT 13190.25 1046.435 13192.77 10000 ;
      RECT 13174.73 1046.435 13175.79 10000 ;
      RECT 13144.21 1046.435 13145.27 10000 ;
      RECT 13127.23 1046.435 13129.75 10000 ;
      RECT 13110.25 1046.435 13112.77 10000 ;
      RECT 13094.73 1046.435 13095.79 10000 ;
      RECT 13064.21 1046.435 13065.27 10000 ;
      RECT 13047.23 1046.435 13049.75 10000 ;
      RECT 13030.25 1046.435 13032.77 10000 ;
      RECT 13014.73 1046.435 13015.79 10000 ;
      RECT 12984.21 1046.435 12985.27 10000 ;
      RECT 12967.23 1046.435 12969.75 10000 ;
      RECT 12950.25 1046.435 12952.77 10000 ;
      RECT 12934.73 1046.435 12935.79 10000 ;
      RECT 12904.21 1046.435 12905.27 10000 ;
      RECT 12887.23 1046.435 12889.75 10000 ;
      RECT 12870.25 1046.435 12872.77 10000 ;
      RECT 12854.73 1046.435 12855.79 10000 ;
      RECT 12824.21 1046.435 12825.27 10000 ;
      RECT 12807.23 1046.435 12809.75 10000 ;
      RECT 12790.25 1046.435 12792.77 10000 ;
      RECT 12774.73 1046.435 12775.79 10000 ;
      RECT 12744.21 1046.435 12745.27 10000 ;
      RECT 12727.23 1046.435 12729.75 10000 ;
      RECT 12710.25 1046.435 12712.77 10000 ;
      RECT 12694.73 1046.435 12695.79 10000 ;
      RECT 12664.21 1046.435 12665.27 10000 ;
      RECT 12647.23 1046.435 12649.75 10000 ;
      RECT 12630.25 1046.435 12632.77 10000 ;
      RECT 12614.73 1046.435 12615.79 10000 ;
      RECT 12584.21 1046.435 12585.27 10000 ;
      RECT 12567.23 1046.435 12569.75 10000 ;
      RECT 12550.25 1046.435 12552.77 10000 ;
      RECT 12534.73 1046.435 12535.79 10000 ;
      RECT 12504.21 1046.435 12505.27 10000 ;
      RECT 12487.23 1046.435 12489.75 10000 ;
      RECT 12470.25 1046.435 12472.77 10000 ;
      RECT 12454.73 1046.435 12455.79 10000 ;
      RECT 12424.21 1046.435 12425.27 10000 ;
      RECT 12407.23 1046.435 12409.75 10000 ;
      RECT 12390.25 1046.435 12392.77 10000 ;
      RECT 12374.73 1046.435 12375.79 10000 ;
      RECT 12344.21 1046.435 12345.27 10000 ;
      RECT 12327.23 1046.435 12329.75 10000 ;
      RECT 12310.25 1046.435 12312.77 10000 ;
      RECT 12294.73 1046.435 12295.79 10000 ;
      RECT 12264.21 1046.435 12265.27 10000 ;
      RECT 12247.23 1046.435 12249.75 10000 ;
      RECT 12230.25 1046.435 12232.77 10000 ;
      RECT 12214.73 1046.435 12215.79 10000 ;
      RECT 12184.21 1046.435 12185.27 10000 ;
      RECT 12167.23 1046.435 12169.75 10000 ;
      RECT 12150.25 1046.435 12152.77 10000 ;
      RECT 12134.73 1046.435 12135.79 10000 ;
      RECT 12104.21 1046.435 12105.27 10000 ;
      RECT 12087.23 1046.435 12089.75 10000 ;
      RECT 12070.25 1046.435 12072.77 10000 ;
      RECT 12054.73 1046.435 12055.79 10000 ;
      RECT 12024.21 1046.435 12025.27 10000 ;
      RECT 12007.23 1046.435 12009.75 10000 ;
      RECT 11990.25 1046.435 11992.77 10000 ;
      RECT 11974.73 1046.435 11975.79 10000 ;
      RECT 11944.21 1046.435 11945.27 10000 ;
      RECT 11927.23 1046.435 11929.75 10000 ;
      RECT 11910.25 1046.435 11912.77 10000 ;
      RECT 11894.73 1046.435 11895.79 10000 ;
      RECT 11864.21 1046.435 11865.27 10000 ;
      RECT 11847.23 1046.435 11849.75 10000 ;
      RECT 11830.25 1046.435 11832.77 10000 ;
      RECT 11814.73 1046.435 11815.79 10000 ;
      RECT 11784.21 1046.435 11785.27 10000 ;
      RECT 11767.23 1046.435 11769.75 10000 ;
      RECT 11750.25 1046.435 11752.77 10000 ;
      RECT 11734.73 1046.435 11735.79 10000 ;
      RECT 11704.21 1046.435 11705.27 10000 ;
      RECT 11687.23 1046.435 11689.75 10000 ;
      RECT 11670.25 1046.435 11672.77 10000 ;
      RECT 11654.73 1046.435 11655.79 10000 ;
      RECT 11624.21 1046.435 11625.27 10000 ;
      RECT 11607.23 1046.435 11609.75 10000 ;
      RECT 11590.25 1046.435 11592.77 10000 ;
      RECT 11574.73 1046.435 11575.79 10000 ;
      RECT 11544.21 1046.435 11545.27 10000 ;
      RECT 11527.23 1046.435 11529.75 10000 ;
      RECT 11510.25 1046.435 11512.77 10000 ;
      RECT 11494.73 1046.435 11495.79 10000 ;
      RECT 11464.21 1046.435 11465.27 10000 ;
      RECT 11447.23 1046.435 11449.75 10000 ;
      RECT 11430.25 1046.435 11432.77 10000 ;
      RECT 11414.73 1046.435 11415.79 10000 ;
      RECT 11384.21 1046.435 11385.27 10000 ;
      RECT 11367.23 1046.435 11369.75 10000 ;
      RECT 11350.25 1046.435 11352.77 10000 ;
      RECT 11334.73 1046.435 11335.79 10000 ;
      RECT 11304.21 1046.435 11305.27 10000 ;
      RECT 11287.23 1046.435 11289.75 10000 ;
      RECT 11270.25 1046.435 11272.77 10000 ;
      RECT 11254.73 1046.435 11255.79 10000 ;
      RECT 11224.21 1046.435 11225.27 10000 ;
      RECT 11207.23 1046.435 11209.75 10000 ;
      RECT 11190.25 1046.435 11192.77 10000 ;
      RECT 11174.73 1046.435 11175.79 10000 ;
      RECT 11144.21 1046.435 11145.27 10000 ;
      RECT 11127.23 1046.435 11129.75 10000 ;
      RECT 11110.25 1046.435 11112.77 10000 ;
      RECT 11094.73 1046.435 11095.79 10000 ;
      RECT 11064.21 1046.435 11065.27 10000 ;
      RECT 11047.23 1046.435 11049.75 10000 ;
      RECT 11030.25 1046.435 11032.77 10000 ;
      RECT 11014.73 1046.435 11015.79 10000 ;
      RECT 10984.21 1046.435 10985.27 10000 ;
      RECT 10967.23 1046.435 10969.75 10000 ;
      RECT 10950.25 1046.435 10952.77 10000 ;
      RECT 10934.73 1046.435 10935.79 10000 ;
      RECT 10904.21 1046.435 10905.27 10000 ;
      RECT 10887.23 1046.435 10889.75 10000 ;
      RECT 10870.25 1046.435 10872.77 10000 ;
      RECT 10854.73 1046.435 10855.79 10000 ;
      RECT 10824.21 1046.435 10825.27 10000 ;
      RECT 10807.23 1046.435 10809.75 10000 ;
      RECT 10790.25 1046.435 10792.77 10000 ;
      RECT 10774.73 1046.435 10775.79 10000 ;
      RECT 10744.21 1046.435 10745.27 10000 ;
      RECT 10727.23 1046.435 10729.75 10000 ;
      RECT 10710.25 1046.435 10712.77 10000 ;
      RECT 10694.73 1046.435 10695.79 10000 ;
      RECT 10664.21 1046.435 10665.27 10000 ;
      RECT 10647.23 1046.435 10649.75 10000 ;
      RECT 10630.25 1046.435 10632.77 10000 ;
      RECT 10614.73 1046.435 10615.79 10000 ;
      RECT 10584.21 1046.435 10585.27 10000 ;
      RECT 10567.23 1046.435 10569.75 10000 ;
      RECT 10550.25 1046.435 10552.77 10000 ;
      RECT 10534.73 1046.435 10535.79 10000 ;
      RECT 10504.21 1046.435 10505.27 10000 ;
      RECT 10487.23 1046.435 10489.75 10000 ;
      RECT 10470.25 1046.435 10472.77 10000 ;
      RECT 10454.73 1046.435 10455.79 10000 ;
      RECT 10424.21 1046.435 10425.27 10000 ;
      RECT 10407.23 1046.435 10409.75 10000 ;
      RECT 10390.25 1046.435 10392.77 10000 ;
      RECT 10374.73 1046.435 10375.79 10000 ;
      RECT 10344.21 1046.435 10345.27 10000 ;
      RECT 10327.23 1046.435 10329.75 10000 ;
      RECT 10310.25 1046.435 10312.77 10000 ;
      RECT 10294.73 1046.435 10295.79 10000 ;
      RECT 10264.21 1046.435 10265.27 10000 ;
      RECT 10247.23 1046.435 10249.75 10000 ;
      RECT 10230.25 1046.435 10232.77 10000 ;
      RECT 10214.73 1046.435 10215.79 10000 ;
      RECT 10184.21 1046.435 10185.27 10000 ;
      RECT 10167.23 1046.435 10169.75 10000 ;
      RECT 10150.25 1046.435 10152.77 10000 ;
      RECT 10134.73 1046.435 10135.79 10000 ;
      RECT 10104.21 1046.435 10105.27 10000 ;
      RECT 10087.23 1046.435 10089.75 10000 ;
      RECT 10070.25 1046.435 10072.77 10000 ;
      RECT 10054.73 1046.435 10055.79 10000 ;
      RECT 10024.21 1046.435 10025.27 10000 ;
      RECT 10007.23 1046.435 10009.75 10000 ;
      RECT 9990.25 1046.435 9992.77 10000 ;
      RECT 9974.73 1046.435 9975.79 10000 ;
      RECT 9944.21 1046.435 9945.27 10000 ;
      RECT 9927.23 1046.435 9929.75 10000 ;
      RECT 9910.25 1046.435 9912.77 10000 ;
      RECT 9894.73 1046.435 9895.79 10000 ;
      RECT 9864.21 1046.435 9865.27 10000 ;
      RECT 9847.23 1046.435 9849.75 10000 ;
      RECT 9830.25 1046.435 9832.77 10000 ;
      RECT 9814.73 1046.435 9815.79 10000 ;
      RECT 9784.21 1046.435 9785.27 10000 ;
      RECT 9767.23 1046.435 9769.75 10000 ;
      RECT 9750.25 1046.435 9752.77 10000 ;
      RECT 9734.73 1046.435 9735.79 10000 ;
      RECT 9704.21 1046.435 9705.27 10000 ;
      RECT 9687.23 1046.435 9689.75 10000 ;
      RECT 9670.25 1046.435 9672.77 10000 ;
      RECT 9654.73 1046.435 9655.79 10000 ;
      RECT 9624.21 1046.435 9625.27 10000 ;
      RECT 9607.23 1046.435 9609.75 10000 ;
      RECT 9590.25 1046.435 9592.77 10000 ;
      RECT 9574.73 1046.435 9575.79 10000 ;
      RECT 9544.21 1046.435 9545.27 10000 ;
      RECT 9527.23 1046.435 9529.75 10000 ;
      RECT 9510.25 1046.435 9512.77 10000 ;
      RECT 9494.73 1046.435 9495.79 10000 ;
      RECT 9464.21 1046.435 9465.27 10000 ;
      RECT 9447.23 1046.435 9449.75 10000 ;
      RECT 9430.25 1046.435 9432.77 10000 ;
      RECT 9414.73 1046.435 9415.79 10000 ;
      RECT 9384.21 1046.435 9385.27 10000 ;
      RECT 9367.23 1046.435 9369.75 10000 ;
      RECT 9350.25 1046.435 9352.77 10000 ;
      RECT 9334.73 1046.435 9335.79 10000 ;
      RECT 9304.21 1046.435 9305.27 10000 ;
      RECT 9287.23 1046.435 9289.75 10000 ;
      RECT 9270.25 1046.435 9272.77 10000 ;
      RECT 9254.73 1046.435 9255.79 10000 ;
      RECT 9224.21 1046.435 9225.27 10000 ;
      RECT 9207.23 1046.435 9209.75 10000 ;
      RECT 9190.25 1046.435 9192.77 10000 ;
      RECT 9174.73 1046.435 9175.79 10000 ;
      RECT 9144.21 1046.435 9145.27 10000 ;
      RECT 9127.23 1046.435 9129.75 10000 ;
      RECT 9110.25 1046.435 9112.77 10000 ;
      RECT 9094.73 1046.435 9095.79 10000 ;
      RECT 9064.21 1046.435 9065.27 10000 ;
      RECT 9047.23 1046.435 9049.75 10000 ;
      RECT 9030.25 1046.435 9032.77 10000 ;
      RECT 9014.73 1046.435 9015.79 10000 ;
      RECT 8984.21 1046.435 8985.27 10000 ;
      RECT 8967.23 1046.435 8969.75 10000 ;
      RECT 8950.25 1046.435 8952.77 10000 ;
      RECT 8934.73 1046.435 8935.79 10000 ;
      RECT 8904.21 1046.435 8905.27 10000 ;
      RECT 8887.23 1046.435 8889.75 10000 ;
      RECT 8870.25 1046.435 8872.77 10000 ;
      RECT 8854.73 1046.435 8855.79 10000 ;
      RECT 8824.21 1046.435 8825.27 10000 ;
      RECT 8807.23 1046.435 8809.75 10000 ;
      RECT 8790.25 1046.435 8792.77 10000 ;
      RECT 8774.73 1046.435 8775.79 10000 ;
      RECT 8744.21 1046.435 8745.27 10000 ;
      RECT 8727.23 1046.435 8729.75 10000 ;
      RECT 8710.25 1046.435 8712.77 10000 ;
      RECT 8694.73 1046.435 8695.79 10000 ;
      RECT 8664.21 1046.435 8665.27 10000 ;
      RECT 8647.23 1046.435 8649.75 10000 ;
      RECT 8630.25 1046.435 8632.77 10000 ;
      RECT 8614.73 1046.435 8615.79 10000 ;
      RECT 8584.21 1046.435 8585.27 10000 ;
      RECT 8567.23 1046.435 8569.75 10000 ;
      RECT 8550.25 1046.435 8552.77 10000 ;
      RECT 8534.73 1046.435 8535.79 10000 ;
      RECT 8504.21 1046.435 8505.27 10000 ;
      RECT 8487.23 1046.435 8489.75 10000 ;
      RECT 8470.25 1046.435 8472.77 10000 ;
      RECT 8454.73 1046.435 8455.79 10000 ;
      RECT 8424.21 1046.435 8425.27 10000 ;
      RECT 8407.23 1046.435 8409.75 10000 ;
      RECT 8390.25 1046.435 8392.77 10000 ;
      RECT 8374.73 1046.435 8375.79 10000 ;
      RECT 8344.21 1046.435 8345.27 10000 ;
      RECT 8327.23 1046.435 8329.75 10000 ;
      RECT 8310.25 1046.435 8312.77 10000 ;
      RECT 8294.73 1046.435 8295.79 10000 ;
      RECT 8264.21 1046.435 8265.27 10000 ;
      RECT 8247.23 1046.435 8249.75 10000 ;
      RECT 8230.25 1046.435 8232.77 10000 ;
      RECT 8214.73 1046.435 8215.79 10000 ;
      RECT 8184.21 1046.435 8185.27 10000 ;
      RECT 8167.23 1046.435 8169.75 10000 ;
      RECT 8150.25 1046.435 8152.77 10000 ;
      RECT 8134.73 1046.435 8135.79 10000 ;
      RECT 8104.21 1046.435 8105.27 10000 ;
      RECT 8087.23 1046.435 8089.75 10000 ;
      RECT 8070.25 1046.435 8072.77 10000 ;
      RECT 8054.73 1046.435 8055.79 10000 ;
      RECT 8024.21 1046.435 8025.27 10000 ;
      RECT 8007.23 1046.435 8009.75 10000 ;
      RECT 7990.25 1046.435 7992.77 10000 ;
      RECT 7974.73 1046.435 7975.79 10000 ;
      RECT 7944.21 1046.435 7945.27 10000 ;
      RECT 7927.23 1046.435 7929.75 10000 ;
      RECT 7910.25 1046.435 7912.77 10000 ;
      RECT 7894.73 1046.435 7895.79 10000 ;
      RECT 7864.21 1046.435 7865.27 10000 ;
      RECT 7847.23 1046.435 7849.75 10000 ;
      RECT 7830.25 1046.435 7832.77 10000 ;
      RECT 7814.73 1046.435 7815.79 10000 ;
      RECT 7784.21 1046.435 7785.27 10000 ;
      RECT 7767.23 1046.435 7769.75 10000 ;
      RECT 7750.25 1046.435 7752.77 10000 ;
      RECT 7734.73 1046.435 7735.79 10000 ;
      RECT 7704.21 1046.435 7705.27 10000 ;
      RECT 7687.23 1046.435 7689.75 10000 ;
      RECT 7670.25 1046.435 7672.77 10000 ;
      RECT 7654.73 1046.435 7655.79 10000 ;
      RECT 7624.21 1046.435 7625.27 10000 ;
      RECT 7607.23 1046.435 7609.75 10000 ;
      RECT 7590.25 1046.435 7592.77 10000 ;
      RECT 7574.73 1046.435 7575.79 10000 ;
      RECT 7544.21 1046.435 7545.27 10000 ;
      RECT 7527.23 1046.435 7529.75 10000 ;
      RECT 7510.25 1046.435 7512.77 10000 ;
      RECT 7494.73 1046.435 7495.79 10000 ;
      RECT 7464.21 1046.435 7465.27 10000 ;
      RECT 7447.23 1046.435 7449.75 10000 ;
      RECT 7430.25 1046.435 7432.77 10000 ;
      RECT 7414.73 1046.435 7415.79 10000 ;
      RECT 7384.21 1046.435 7385.27 10000 ;
      RECT 7367.23 1046.435 7369.75 10000 ;
      RECT 7350.25 1046.435 7352.77 10000 ;
      RECT 7334.73 1046.435 7335.79 10000 ;
      RECT 7304.21 1046.435 7305.27 10000 ;
      RECT 7287.23 1046.435 7289.75 10000 ;
      RECT 7270.25 1046.435 7272.77 10000 ;
      RECT 7254.73 1046.435 7255.79 10000 ;
      RECT 7224.21 1046.435 7225.27 10000 ;
      RECT 7207.23 1046.435 7209.75 10000 ;
      RECT 7190.25 1046.435 7192.77 10000 ;
      RECT 7174.73 1046.435 7175.79 10000 ;
      RECT 7144.21 1046.435 7145.27 10000 ;
      RECT 7127.23 1046.435 7129.75 10000 ;
      RECT 7110.25 1046.435 7112.77 10000 ;
      RECT 7094.73 1046.435 7095.79 10000 ;
      RECT 7064.21 1046.435 7065.27 10000 ;
      RECT 7047.23 1046.435 7049.75 10000 ;
      RECT 7030.25 1046.435 7032.77 10000 ;
      RECT 7014.73 1046.435 7015.79 10000 ;
      RECT 6984.21 1046.435 6985.27 10000 ;
      RECT 6967.23 1046.435 6969.75 10000 ;
      RECT 6950.25 1046.435 6952.77 10000 ;
      RECT 6934.73 1046.435 6935.79 10000 ;
      RECT 6904.21 1046.435 6905.27 10000 ;
      RECT 6887.23 1046.435 6889.75 10000 ;
      RECT 6870.25 1046.435 6872.77 10000 ;
      RECT 6854.73 1046.435 6855.79 10000 ;
      RECT 6824.21 1046.435 6825.27 10000 ;
      RECT 6807.23 1046.435 6809.75 10000 ;
      RECT 6790.25 1046.435 6792.77 10000 ;
      RECT 6774.73 1046.435 6775.79 10000 ;
      RECT 6744.21 1046.435 6745.27 10000 ;
      RECT 6727.23 1046.435 6729.75 10000 ;
      RECT 6710.25 1046.435 6712.77 10000 ;
      RECT 6694.73 1046.435 6695.79 10000 ;
      RECT 6664.21 1046.435 6665.27 10000 ;
      RECT 6647.23 1046.435 6649.75 10000 ;
      RECT 6630.25 1046.435 6632.77 10000 ;
      RECT 6614.73 1046.435 6615.79 10000 ;
      RECT 6584.21 1046.435 6585.27 10000 ;
      RECT 6567.23 1046.435 6569.75 10000 ;
      RECT 6550.25 1046.435 6552.77 10000 ;
      RECT 6534.73 1046.435 6535.79 10000 ;
      RECT 6504.21 1046.435 6505.27 10000 ;
      RECT 6487.23 1046.435 6489.75 10000 ;
      RECT 6470.25 1046.435 6472.77 10000 ;
      RECT 6454.73 1046.435 6455.79 10000 ;
      RECT 6424.21 1046.435 6425.27 10000 ;
      RECT 6407.23 1046.435 6409.75 10000 ;
      RECT 6390.25 1046.435 6392.77 10000 ;
      RECT 6374.73 1046.435 6375.79 10000 ;
      RECT 6344.21 1046.435 6345.27 10000 ;
      RECT 6327.23 1046.435 6329.75 10000 ;
      RECT 6310.25 1046.435 6312.77 10000 ;
      RECT 6294.73 1046.435 6295.79 10000 ;
      RECT 6264.21 1046.435 6265.27 10000 ;
      RECT 6247.23 1046.435 6249.75 10000 ;
      RECT 6230.25 1046.435 6232.77 10000 ;
      RECT 6214.73 1046.435 6215.79 10000 ;
      RECT 6184.21 1046.435 6185.27 10000 ;
      RECT 6167.23 1046.435 6169.75 10000 ;
      RECT 6150.25 1046.435 6152.77 10000 ;
      RECT 6134.73 1046.435 6135.79 10000 ;
      RECT 6104.21 1046.435 6105.27 10000 ;
      RECT 6087.23 1046.435 6089.75 10000 ;
      RECT 6070.25 1046.435 6072.77 10000 ;
      RECT 6054.73 1046.435 6055.79 10000 ;
      RECT 6024.21 1046.435 6025.27 10000 ;
      RECT 6007.23 1046.435 6009.75 10000 ;
      RECT 5990.25 1046.435 5992.77 10000 ;
      RECT 5974.73 1046.435 5975.79 10000 ;
      RECT 5944.21 1046.435 5945.27 10000 ;
      RECT 5927.23 1046.435 5929.75 10000 ;
      RECT 5910.25 1046.435 5912.77 10000 ;
      RECT 5894.73 1046.435 5895.79 10000 ;
      RECT 5864.21 1046.435 5865.27 10000 ;
      RECT 5847.23 1046.435 5849.75 10000 ;
      RECT 5830.25 1046.435 5832.77 10000 ;
      RECT 5814.73 1046.435 5815.79 10000 ;
      RECT 5784.21 1046.435 5785.27 10000 ;
      RECT 5767.23 1046.435 5769.75 10000 ;
      RECT 5750.25 1046.435 5752.77 10000 ;
      RECT 5734.73 1046.435 5735.79 10000 ;
      RECT 5704.21 1046.435 5705.27 10000 ;
      RECT 5687.23 1046.435 5689.75 10000 ;
      RECT 5670.25 1046.435 5672.77 10000 ;
      RECT 5654.73 1046.435 5655.79 10000 ;
      RECT 5624.21 1046.435 5625.27 10000 ;
      RECT 5607.23 1046.435 5609.75 10000 ;
      RECT 5590.25 1046.435 5592.77 10000 ;
      RECT 5574.73 1046.435 5575.79 10000 ;
      RECT 5544.21 1046.435 5545.27 10000 ;
      RECT 5527.23 1046.435 5529.75 10000 ;
      RECT 5510.25 1046.435 5512.77 10000 ;
      RECT 5494.73 1046.435 5495.79 10000 ;
      RECT 5464.21 1046.435 5465.27 10000 ;
      RECT 5447.23 1046.435 5449.75 10000 ;
      RECT 5430.25 1046.435 5432.77 10000 ;
      RECT 5414.73 1046.435 5415.79 10000 ;
      RECT 5384.21 1046.435 5385.27 10000 ;
      RECT 5367.23 1046.435 5369.75 10000 ;
      RECT 5350.25 1046.435 5352.77 10000 ;
      RECT 5334.73 1046.435 5335.79 10000 ;
      RECT 5304.21 1046.435 5305.27 10000 ;
      RECT 5287.23 1046.435 5289.75 10000 ;
      RECT 5270.25 1046.435 5272.77 10000 ;
      RECT 5254.73 1046.435 5255.79 10000 ;
      RECT 5224.21 1046.435 5225.27 10000 ;
      RECT 5207.23 1046.435 5209.75 10000 ;
      RECT 5190.25 1046.435 5192.77 10000 ;
      RECT 5174.73 1046.435 5175.79 10000 ;
      RECT 5144.21 1046.435 5145.27 10000 ;
      RECT 5127.23 1046.435 5129.75 10000 ;
      RECT 5110.25 1046.435 5112.77 10000 ;
      RECT 5094.73 1046.435 5095.79 10000 ;
      RECT 5064.21 1046.435 5065.27 10000 ;
      RECT 5047.23 1046.435 5049.75 10000 ;
      RECT 5030.25 1046.435 5032.77 10000 ;
      RECT 5014.73 1046.435 5015.79 10000 ;
      RECT 4984.21 1046.435 4985.27 10000 ;
      RECT 4967.23 1046.435 4969.75 10000 ;
      RECT 4950.25 1046.435 4952.77 10000 ;
      RECT 4934.73 1046.435 4935.79 10000 ;
      RECT 4904.21 1046.435 4905.27 10000 ;
      RECT 4887.23 1046.435 4889.75 10000 ;
      RECT 4870.25 1046.435 4872.77 10000 ;
      RECT 4854.73 1046.435 4855.79 10000 ;
      RECT 4824.21 1046.435 4825.27 10000 ;
      RECT 4807.23 1046.435 4809.75 10000 ;
      RECT 4790.25 1046.435 4792.77 10000 ;
      RECT 4774.73 1046.435 4775.79 10000 ;
      RECT 4744.21 1046.435 4745.27 10000 ;
      RECT 4727.23 1046.435 4729.75 10000 ;
      RECT 4710.25 1046.435 4712.77 10000 ;
      RECT 4694.73 1046.435 4695.79 10000 ;
      RECT 4664.21 1046.435 4665.27 10000 ;
      RECT 4647.23 1046.435 4649.75 10000 ;
      RECT 4630.25 1046.435 4632.77 10000 ;
      RECT 4614.73 1046.435 4615.79 10000 ;
      RECT 4584.21 1046.435 4585.27 10000 ;
      RECT 4567.23 1046.435 4569.75 10000 ;
      RECT 4550.25 1046.435 4552.77 10000 ;
      RECT 4534.73 1046.435 4535.79 10000 ;
      RECT 4504.21 1046.435 4505.27 10000 ;
      RECT 4487.23 1046.435 4489.75 10000 ;
      RECT 4470.25 1046.435 4472.77 10000 ;
      RECT 4454.73 1046.435 4455.79 10000 ;
      RECT 4424.21 1046.435 4425.27 10000 ;
      RECT 4407.23 1046.435 4409.75 10000 ;
      RECT 4390.25 1046.435 4392.77 10000 ;
      RECT 4374.73 1046.435 4375.79 10000 ;
      RECT 4344.21 1046.435 4345.27 10000 ;
      RECT 4327.23 1046.435 4329.75 10000 ;
      RECT 4310.25 1046.435 4312.77 10000 ;
      RECT 4294.73 1046.435 4295.79 10000 ;
      RECT 4264.21 1046.435 4265.27 10000 ;
      RECT 4247.23 1046.435 4249.75 10000 ;
      RECT 4230.25 1046.435 4232.77 10000 ;
      RECT 4214.73 1046.435 4215.79 10000 ;
      RECT 4184.21 1046.435 4185.27 10000 ;
      RECT 4167.23 1046.435 4169.75 10000 ;
      RECT 4150.25 1046.435 4152.77 10000 ;
      RECT 4134.73 1046.435 4135.79 10000 ;
      RECT 4104.21 1046.435 4105.27 10000 ;
      RECT 4087.23 1046.435 4089.75 10000 ;
      RECT 4070.25 1046.435 4072.77 10000 ;
      RECT 4054.73 1046.435 4055.79 10000 ;
      RECT 4024.21 1046.435 4025.27 10000 ;
      RECT 4007.23 1046.435 4009.75 10000 ;
      RECT 3990.25 1046.435 3992.77 10000 ;
      RECT 3974.73 1046.435 3975.79 10000 ;
      RECT 3944.21 1046.435 3945.27 10000 ;
      RECT 3927.23 1046.435 3929.75 10000 ;
      RECT 3910.25 1046.435 3912.77 10000 ;
      RECT 3894.73 1046.435 3895.79 10000 ;
      RECT 3864.21 1046.435 3865.27 10000 ;
      RECT 3847.23 1046.435 3849.75 10000 ;
      RECT 3830.25 1046.435 3832.77 10000 ;
      RECT 3814.73 1046.435 3815.79 10000 ;
      RECT 3784.21 1046.435 3785.27 10000 ;
      RECT 3767.23 1046.435 3769.75 10000 ;
      RECT 3750.25 1046.435 3752.77 10000 ;
      RECT 3734.73 1046.435 3735.79 10000 ;
      RECT 3704.21 1046.435 3705.27 10000 ;
      RECT 3687.23 1046.435 3689.75 10000 ;
      RECT 3670.25 1046.435 3672.77 10000 ;
      RECT 3654.73 1046.435 3655.79 10000 ;
      RECT 3624.21 1046.435 3625.27 10000 ;
      RECT 3607.23 1046.435 3609.75 10000 ;
      RECT 3590.25 1046.435 3592.77 10000 ;
      RECT 3574.73 1046.435 3575.79 10000 ;
      RECT 3544.21 1046.435 3545.27 10000 ;
      RECT 3527.23 1046.435 3529.75 10000 ;
      RECT 3510.25 1046.435 3512.77 10000 ;
      RECT 3494.73 1046.435 3495.79 10000 ;
      RECT 3464.21 1046.435 3465.27 10000 ;
      RECT 3447.23 1046.435 3449.75 10000 ;
      RECT 3430.25 1046.435 3432.77 10000 ;
      RECT 3414.73 1046.435 3415.79 10000 ;
      RECT 3384.21 1046.435 3385.27 10000 ;
      RECT 3367.23 1046.435 3369.75 10000 ;
      RECT 3350.25 1046.435 3352.77 10000 ;
      RECT 3334.73 1046.435 3335.79 10000 ;
      RECT 3304.21 1046.435 3305.27 10000 ;
      RECT 3287.23 1046.435 3289.75 10000 ;
      RECT 3270.25 1046.435 3272.77 10000 ;
      RECT 3254.73 1046.435 3255.79 10000 ;
      RECT 3224.21 1046.435 3225.27 10000 ;
      RECT 3207.23 1046.435 3209.75 10000 ;
      RECT 3190.25 1046.435 3192.77 10000 ;
      RECT 3174.73 1046.435 3175.79 10000 ;
      RECT 3144.21 1046.435 3145.27 10000 ;
      RECT 3127.23 1046.435 3129.75 10000 ;
      RECT 3110.25 1046.435 3112.77 10000 ;
      RECT 3094.73 1046.435 3095.79 10000 ;
      RECT 3064.21 1046.435 3065.27 10000 ;
      RECT 3047.23 1046.435 3049.75 10000 ;
      RECT 3030.25 1046.435 3032.77 10000 ;
      RECT 3014.73 1046.435 3015.79 10000 ;
      RECT 2984.21 1046.435 2985.27 10000 ;
      RECT 2967.23 1046.435 2969.75 10000 ;
      RECT 2950.25 1046.435 2952.77 10000 ;
      RECT 2934.73 1046.435 2935.79 10000 ;
      RECT 2904.21 1046.435 2905.27 10000 ;
      RECT 2887.23 1046.435 2889.75 10000 ;
      RECT 2870.25 1046.435 2872.77 10000 ;
      RECT 2854.73 1046.435 2855.79 10000 ;
      RECT 2824.21 1046.435 2825.27 10000 ;
      RECT 2807.23 1046.435 2809.75 10000 ;
      RECT 2790.25 1046.435 2792.77 10000 ;
      RECT 2774.73 1046.435 2775.79 10000 ;
      RECT 2744.21 1046.435 2745.27 10000 ;
      RECT 2727.23 1046.435 2729.75 10000 ;
      RECT 2710.25 1046.435 2712.77 10000 ;
      RECT 2694.73 1046.435 2695.79 10000 ;
      RECT 2664.21 1046.435 2665.27 10000 ;
      RECT 2647.23 1046.435 2649.75 10000 ;
      RECT 2630.25 1046.435 2632.77 10000 ;
      RECT 2614.73 1046.435 2615.79 10000 ;
      RECT 2584.21 1046.435 2585.27 10000 ;
      RECT 2567.23 1046.435 2569.75 10000 ;
      RECT 2550.25 1046.435 2552.77 10000 ;
      RECT 2534.73 1046.435 2535.79 10000 ;
      RECT 2504.21 1046.435 2505.27 10000 ;
      RECT 2487.23 1046.435 2489.75 10000 ;
      RECT 2470.25 1046.435 2472.77 10000 ;
      RECT 2454.73 1046.435 2455.79 10000 ;
      RECT 2424.21 1046.435 2425.27 10000 ;
      RECT 2407.23 1046.435 2409.75 10000 ;
      RECT 2390.25 1046.435 2392.77 10000 ;
      RECT 2374.73 1046.435 2375.79 10000 ;
      RECT 2344.21 1046.435 2345.27 10000 ;
      RECT 2327.23 1046.435 2329.75 10000 ;
      RECT 2310.25 1046.435 2312.77 10000 ;
      RECT 2294.73 1046.435 2295.79 10000 ;
      RECT 2264.21 1046.435 2265.27 10000 ;
      RECT 2247.23 1046.435 2249.75 10000 ;
      RECT 2230.25 1046.435 2232.77 10000 ;
      RECT 2214.73 1046.435 2215.79 10000 ;
      RECT 2184.21 1046.435 2185.27 10000 ;
      RECT 2167.23 1046.435 2169.75 10000 ;
      RECT 2150.25 1046.435 2152.77 10000 ;
      RECT 2134.73 1046.435 2135.79 10000 ;
      RECT 2104.21 1046.435 2105.27 10000 ;
      RECT 2087.23 1046.435 2089.75 10000 ;
      RECT 2070.25 1046.435 2072.77 10000 ;
      RECT 2054.73 1046.435 2055.79 10000 ;
      RECT 2024.21 1046.435 2025.27 10000 ;
      RECT 2007.23 1046.435 2009.75 10000 ;
      RECT 1990.25 1046.435 1992.77 10000 ;
      RECT 1974.73 1046.435 1975.79 10000 ;
      RECT 1944.21 1046.435 1945.27 10000 ;
      RECT 1927.23 1046.435 1929.75 10000 ;
      RECT 1910.25 1046.435 1912.77 10000 ;
      RECT 1894.73 1046.435 1895.79 10000 ;
      RECT 1864.21 1046.435 1865.27 10000 ;
      RECT 1847.23 1046.435 1849.75 10000 ;
      RECT 1830.25 1046.435 1832.77 10000 ;
      RECT 1814.73 1046.435 1815.79 10000 ;
      RECT 1784.21 1046.435 1785.27 10000 ;
      RECT 1767.23 1046.435 1769.75 10000 ;
      RECT 1750.25 1046.435 1752.77 10000 ;
      RECT 1734.73 1046.435 1735.79 10000 ;
      RECT 1704.21 1046.435 1705.27 10000 ;
      RECT 1687.23 1046.435 1689.75 10000 ;
      RECT 1670.25 1046.435 1672.77 10000 ;
      RECT 1654.73 1046.435 1655.79 10000 ;
      RECT 1624.21 1046.435 1625.27 10000 ;
      RECT 1607.23 1046.435 1609.75 10000 ;
      RECT 1590.25 1046.435 1592.77 10000 ;
      RECT 1574.73 1046.435 1575.79 10000 ;
      RECT 1544.21 1046.435 1545.27 10000 ;
      RECT 1527.23 1046.435 1529.75 10000 ;
      RECT 1510.25 1046.435 1512.77 10000 ;
      RECT 1494.73 1046.435 1495.79 10000 ;
      RECT 1464.21 1046.435 1465.27 10000 ;
      RECT 1447.23 1046.435 1449.75 10000 ;
      RECT 1430.25 1046.435 1432.77 10000 ;
      RECT 1414.73 1046.435 1415.79 10000 ;
      RECT 1384.21 1046.435 1385.27 10000 ;
      RECT 1367.23 1046.435 1369.75 10000 ;
      RECT 1350.25 1046.435 1352.77 10000 ;
      RECT 1334.73 1046.435 1335.79 10000 ;
      RECT 1304.21 1046.435 1305.27 10000 ;
      RECT 1287.23 1046.435 1289.75 10000 ;
      RECT 1270.25 1046.435 1272.77 10000 ;
      RECT 1254.73 1046.435 1255.79 10000 ;
      RECT 1224.21 1046.435 1225.27 10000 ;
      RECT 1207.23 1046.435 1209.75 10000 ;
      RECT 1190.25 1046.435 1192.77 10000 ;
      RECT 1174.73 1046.435 1175.79 10000 ;
      RECT 1144.21 1046.435 1145.27 10000 ;
      RECT 998.1 1046.435 1129.75 10000 ;
      RECT 19584.63 680.155 19623.26 715.155 ;
      RECT 19584.63 800.155 19623.26 835.155 ;
      RECT 19584.63 920.155 19623.26 955.155 ;
      RECT 19584.63 1040.155 19623.26 1075.155 ;
      RECT 19584.63 1280.155 19623.26 1315.155 ;
      RECT 19584.63 1400.155 19623.26 1435.155 ;
      RECT 19584.63 8720.155 19623.26 8755.155 ;
      RECT 19584.63 8840.155 19623.26 8875.155 ;
      RECT 19584.63 8960.155 19623.26 8995.155 ;
      RECT 19584.63 9080.155 19623.26 9115.155 ;
      RECT 19584.63 9200.155 19623.26 9235.155 ;
      RECT 19584.63 9320.155 19623.26 9355.155 ;
      RECT 19454.63 638.18 19567.9 688.18 ;
      RECT 19454.63 758.18 19567.9 808.18 ;
      RECT 19454.63 878.18 19567.9 928.18 ;
      RECT 19454.63 998.18 19567.9 1048.18 ;
      RECT 19454.63 1118.18 19567.9 1168.18 ;
      RECT 19454.63 1358.18 19567.9 1408.18 ;
      RECT 19454.63 1478.18 19567.9 1528.18 ;
      RECT 19454.63 1598.18 19567.9 1648.18 ;
      RECT 19454.63 1718.18 19567.9 1768.18 ;
      RECT 19454.63 1838.18 19567.9 1888.18 ;
      RECT 19454.63 1958.18 19567.9 2008.18 ;
      RECT 19454.63 2078.18 19567.9 2128.18 ;
      RECT 19454.63 2198.18 19567.9 2248.18 ;
      RECT 19454.63 2318.18 19567.9 2368.18 ;
      RECT 19454.63 2438.18 19567.9 2488.18 ;
      RECT 19454.63 2558.18 19567.9 2608.18 ;
      RECT 19454.63 2678.18 19567.9 2728.18 ;
      RECT 19454.63 2798.18 19567.9 2848.18 ;
      RECT 19454.63 2918.18 19567.9 2968.18 ;
      RECT 19454.63 3038.18 19567.9 3088.18 ;
      RECT 19454.63 3158.18 19567.9 3208.18 ;
      RECT 19454.63 3278.18 19567.9 3328.18 ;
      RECT 19454.63 3398.18 19567.9 3448.18 ;
      RECT 19454.63 3518.18 19567.9 3568.18 ;
      RECT 19454.63 3638.18 19567.9 3688.18 ;
      RECT 19454.63 3758.18 19567.9 3808.18 ;
      RECT 19454.63 3878.18 19567.9 3928.18 ;
      RECT 19454.63 3998.18 19567.9 4048.18 ;
      RECT 19454.63 4118.18 19567.9 4168.18 ;
      RECT 19454.63 4238.18 19567.9 4288.18 ;
      RECT 19454.63 4358.18 19567.9 4408.18 ;
      RECT 19454.63 4478.18 19567.9 4528.18 ;
      RECT 19454.63 4598.18 19567.9 4648.18 ;
      RECT 19454.63 4718.18 19567.9 4768.18 ;
      RECT 19454.63 4838.18 19567.9 4888.18 ;
      RECT 19454.63 4958.18 19567.9 5008.18 ;
      RECT 19454.63 5078.18 19567.9 5128.18 ;
      RECT 19454.63 5198.18 19567.9 5248.18 ;
      RECT 19454.63 5318.18 19567.9 5368.18 ;
      RECT 19454.63 5438.18 19567.9 5488.18 ;
      RECT 19454.63 5558.18 19567.9 5608.18 ;
      RECT 19454.63 5678.18 19567.9 5728.18 ;
      RECT 19454.63 5798.18 19567.9 5848.18 ;
      RECT 19454.63 5918.18 19567.9 5968.18 ;
      RECT 19454.63 6038.18 19567.9 6088.18 ;
      RECT 19454.63 6158.18 19567.9 6208.18 ;
      RECT 19454.63 6278.18 19567.9 6328.18 ;
      RECT 19454.63 6398.18 19567.9 6448.18 ;
      RECT 19454.63 6518.18 19567.9 6568.18 ;
      RECT 19454.63 6638.18 19567.9 6688.18 ;
      RECT 19454.63 6758.18 19567.9 6808.18 ;
      RECT 19454.63 6878.18 19567.9 6928.18 ;
      RECT 19454.63 6998.18 19567.9 7048.18 ;
      RECT 19454.63 7118.18 19567.9 7168.18 ;
      RECT 19454.63 7238.18 19567.9 7288.18 ;
      RECT 19454.63 7358.18 19567.9 7408.18 ;
      RECT 19454.63 7478.18 19567.9 7528.18 ;
      RECT 19454.63 7598.18 19567.9 7648.18 ;
      RECT 19454.63 7718.18 19567.9 7768.18 ;
      RECT 19454.63 7838.18 19567.9 7888.18 ;
      RECT 19454.63 7958.18 19567.9 8008.18 ;
      RECT 19454.63 8078.18 19567.9 8128.18 ;
      RECT 19454.63 8198.18 19567.9 8248.18 ;
      RECT 19454.63 8318.18 19567.9 8368.18 ;
      RECT 19454.63 8438.18 19567.9 8488.18 ;
      RECT 19454.63 8558.18 19567.9 8608.18 ;
      RECT 19454.63 8678.18 19567.9 8728.18 ;
      RECT 19454.63 8798.18 19567.9 8848.18 ;
      RECT 19454.63 8918.18 19567.9 8968.18 ;
      RECT 19454.63 9038.18 19567.9 9088.18 ;
      RECT 19454.63 9158.18 19567.9 9208.18 ;
      RECT 19454.63 9278.18 19567.9 9328.18 ;
      RECT 19454.63 9398.18 19567.9 9448.18 ;
      RECT 632.1 638.18 745.37 688.18 ;
      RECT 632.1 758.18 745.37 808.18 ;
      RECT 632.1 878.18 745.37 928.18 ;
      RECT 632.1 998.18 745.37 1048.18 ;
      RECT 632.1 1118.18 745.37 1168.18 ;
      RECT 632.1 1358.18 745.37 1408.18 ;
      RECT 632.1 1478.18 745.37 1528.18 ;
      RECT 632.1 1598.18 745.37 1648.18 ;
      RECT 632.1 1718.18 745.37 1768.18 ;
      RECT 632.1 1838.18 745.37 1888.18 ;
      RECT 632.1 1958.18 745.37 2008.18 ;
      RECT 632.1 2078.18 745.37 2128.18 ;
      RECT 632.1 2198.18 745.37 2248.18 ;
      RECT 632.1 2318.18 745.37 2368.18 ;
      RECT 632.1 2438.18 745.37 2488.18 ;
      RECT 632.1 2558.18 745.37 2608.18 ;
      RECT 632.1 2678.18 745.37 2728.18 ;
      RECT 632.1 2798.18 745.37 2848.18 ;
      RECT 632.1 2918.18 745.37 2968.18 ;
      RECT 632.1 3038.18 745.37 3088.18 ;
      RECT 632.1 3158.18 745.37 3208.18 ;
      RECT 632.1 3278.18 745.37 3328.18 ;
      RECT 632.1 3398.18 745.37 3448.18 ;
      RECT 632.1 3518.18 745.37 3568.18 ;
      RECT 632.1 3638.18 745.37 3688.18 ;
      RECT 632.1 3758.18 745.37 3808.18 ;
      RECT 632.1 3878.18 745.37 3928.18 ;
      RECT 632.1 3998.18 745.37 4048.18 ;
      RECT 632.1 4118.18 745.37 4168.18 ;
      RECT 632.1 4238.18 745.37 4288.18 ;
      RECT 632.1 4358.18 745.37 4408.18 ;
      RECT 632.1 4478.18 745.37 4528.18 ;
      RECT 632.1 4598.18 745.37 4648.18 ;
      RECT 632.1 4718.18 745.37 4768.18 ;
      RECT 632.1 4838.18 745.37 4888.18 ;
      RECT 632.1 4958.18 745.37 5008.18 ;
      RECT 632.1 5078.18 745.37 5128.18 ;
      RECT 632.1 5198.18 745.37 5248.18 ;
      RECT 632.1 5318.18 745.37 5368.18 ;
      RECT 632.1 5438.18 745.37 5488.18 ;
      RECT 632.1 5558.18 745.37 5608.18 ;
      RECT 632.1 5678.18 745.37 5728.18 ;
      RECT 632.1 5798.18 745.37 5848.18 ;
      RECT 632.1 5918.18 745.37 5968.18 ;
      RECT 632.1 6038.18 745.37 6088.18 ;
      RECT 632.1 6158.18 745.37 6208.18 ;
      RECT 632.1 6278.18 745.37 6328.18 ;
      RECT 632.1 6398.18 745.37 6448.18 ;
      RECT 632.1 6518.18 745.37 6568.18 ;
      RECT 632.1 6638.18 745.37 6688.18 ;
      RECT 632.1 6758.18 745.37 6808.18 ;
      RECT 632.1 6878.18 745.37 6928.18 ;
      RECT 632.1 6998.18 745.37 7048.18 ;
      RECT 632.1 7118.18 745.37 7168.18 ;
      RECT 632.1 7238.18 745.37 7288.18 ;
      RECT 632.1 7358.18 745.37 7408.18 ;
      RECT 632.1 7478.18 745.37 7528.18 ;
      RECT 632.1 7598.18 745.37 7648.18 ;
      RECT 632.1 7718.18 745.37 7768.18 ;
      RECT 632.1 7838.18 745.37 7888.18 ;
      RECT 632.1 7958.18 745.37 8008.18 ;
      RECT 632.1 8078.18 745.37 8128.18 ;
      RECT 632.1 8198.18 745.37 8248.18 ;
      RECT 632.1 8318.18 745.37 8368.18 ;
      RECT 632.1 8438.18 745.37 8488.18 ;
      RECT 632.1 8558.18 745.37 8608.18 ;
      RECT 632.1 8678.18 745.37 8728.18 ;
      RECT 632.1 8798.18 745.37 8848.18 ;
      RECT 632.1 8918.18 745.37 8968.18 ;
      RECT 632.1 9038.18 745.37 9088.18 ;
      RECT 632.1 9158.18 745.37 9208.18 ;
      RECT 632.1 9278.18 745.37 9328.18 ;
      RECT 632.1 9398.18 745.37 9448.18 ;
      RECT 576.74 680.155 615.37 715.155 ;
      RECT 576.74 800.155 615.37 835.155 ;
      RECT 576.74 920.155 615.37 955.155 ;
      RECT 576.74 1040.155 615.37 1075.155 ;
      RECT 576.74 1160.155 615.37 1195.155 ;
      RECT 502.1 1298.18 615.37 1348.18 ;
      RECT 576.74 8720.155 615.37 8755.155 ;
      RECT 576.74 8840.155 615.37 8875.155 ;
      RECT 576.74 8960.155 615.37 8995.155 ;
      RECT 576.74 9080.155 615.37 9115.155 ;
      RECT 576.74 9200.155 615.37 9235.155 ;
      RECT 576.74 9320.155 615.37 9355.155 ;
    LAYER M1 ;
      POLYGON 19148.125 1036.14 19146.625 1036.14 19146.625 661.71 1013.375 661.71 1013.375 1034.64 19146.625 1034.64 19146.625 1036.14 1011.875 1036.14 1011.875 660.21 19148.125 660.21 ;
  END
END MONOPIX_TOP

END LIBRARY
