VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO digital_ring
  CLASS BLOCK ;
  ORIGIN -12.895 -16.205 ;
  FOREIGN digital_ring 12.895 16.205 ;
  SIZE 18163.8 BY 400.56 ;
  SYMMETRY X Y R90 ;
  PIN PSUB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 18171.195 20.725 18172.195 419.145 ;
        RECT 17.395 20.725 18172.195 21.725 ;
        RECT 17.395 20.725 18.395 419.145 ;
    END
  END PSUB
  PIN VDDP
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 26.67 404.43 18162.92 405.93 ;
        RECT 18161.42 30 18162.92 405.93 ;
        RECT 26.67 30 18162.92 31.5 ;
        RECT 26.67 30 28.17 405.93 ;
    END
  END VDDP
END digital_ring

END LIBRARY
